magic
tech sky130A
magscale 1 2
timestamp 1671334348
<< error_p >>
rect -125 322 -67 328
rect 67 322 125 328
rect -125 288 -113 322
rect 67 288 79 322
rect -125 282 -67 288
rect 67 282 125 288
rect -221 -288 -163 -282
rect -29 -288 29 -282
rect 163 -288 221 -282
rect -221 -322 -209 -288
rect -29 -322 -17 -288
rect 163 -322 175 -288
rect -221 -328 -163 -322
rect -29 -328 29 -322
rect 163 -328 221 -322
<< pwell >>
rect -407 -460 407 460
<< nmos >>
rect -207 -250 -177 250
rect -111 -250 -81 250
rect -15 -250 15 250
rect 81 -250 111 250
rect 177 -250 207 250
<< ndiff >>
rect -269 238 -207 250
rect -269 -238 -257 238
rect -223 -238 -207 238
rect -269 -250 -207 -238
rect -177 238 -111 250
rect -177 -238 -161 238
rect -127 -238 -111 238
rect -177 -250 -111 -238
rect -81 238 -15 250
rect -81 -238 -65 238
rect -31 -238 -15 238
rect -81 -250 -15 -238
rect 15 238 81 250
rect 15 -238 31 238
rect 65 -238 81 238
rect 15 -250 81 -238
rect 111 238 177 250
rect 111 -238 127 238
rect 161 -238 177 238
rect 111 -250 177 -238
rect 207 238 269 250
rect 207 -238 223 238
rect 257 -238 269 238
rect 207 -250 269 -238
<< ndiffc >>
rect -257 -238 -223 238
rect -161 -238 -127 238
rect -65 -238 -31 238
rect 31 -238 65 238
rect 127 -238 161 238
rect 223 -238 257 238
<< psubdiff >>
rect -371 390 -275 424
rect 275 390 371 424
rect -371 328 -337 390
rect 337 328 371 390
rect -371 -390 -337 -328
rect 337 -390 371 -328
rect -371 -424 -275 -390
rect 275 -424 371 -390
<< psubdiffcont >>
rect -275 390 275 424
rect -371 -328 -337 328
rect 337 -328 371 328
rect -275 -424 275 -390
<< poly >>
rect -129 322 -63 338
rect -129 288 -113 322
rect -79 288 -63 322
rect -207 250 -177 276
rect -129 272 -63 288
rect 63 322 129 338
rect 63 288 79 322
rect 113 288 129 322
rect -111 250 -81 272
rect -15 250 15 276
rect 63 272 129 288
rect 81 250 111 272
rect 177 250 207 276
rect -207 -272 -177 -250
rect -225 -288 -159 -272
rect -111 -276 -81 -250
rect -15 -272 15 -250
rect -225 -322 -209 -288
rect -175 -322 -159 -288
rect -225 -338 -159 -322
rect -33 -288 33 -272
rect 81 -276 111 -250
rect 177 -272 207 -250
rect -33 -322 -17 -288
rect 17 -322 33 -288
rect -33 -338 33 -322
rect 159 -288 225 -272
rect 159 -322 175 -288
rect 209 -322 225 -288
rect 159 -338 225 -322
<< polycont >>
rect -113 288 -79 322
rect 79 288 113 322
rect -209 -322 -175 -288
rect -17 -322 17 -288
rect 175 -322 209 -288
<< locali >>
rect -371 390 -275 424
rect 275 390 371 424
rect -371 328 -337 390
rect 337 328 371 390
rect -129 288 -113 322
rect -79 288 -63 322
rect 63 288 79 322
rect 113 288 129 322
rect -257 238 -223 254
rect -257 -254 -223 -238
rect -161 238 -127 254
rect -161 -254 -127 -238
rect -65 238 -31 254
rect -65 -254 -31 -238
rect 31 238 65 254
rect 31 -254 65 -238
rect 127 238 161 254
rect 127 -254 161 -238
rect 223 238 257 254
rect 223 -254 257 -238
rect -225 -322 -209 -288
rect -175 -322 -159 -288
rect -33 -322 -17 -288
rect 17 -322 33 -288
rect 159 -322 175 -288
rect 209 -322 225 -288
rect -371 -390 -337 -328
rect 337 -390 371 -328
rect -371 -424 -275 -390
rect 275 -424 371 -390
<< viali >>
rect -113 288 -79 322
rect 79 288 113 322
rect -257 -238 -223 238
rect -161 -238 -127 238
rect -65 -238 -31 238
rect 31 -238 65 238
rect 127 -238 161 238
rect 223 -238 257 238
rect -209 -322 -175 -288
rect -17 -322 17 -288
rect 175 -322 209 -288
<< metal1 >>
rect -125 322 -67 328
rect -125 288 -113 322
rect -79 288 -67 322
rect -125 282 -67 288
rect 67 322 125 328
rect 67 288 79 322
rect 113 288 125 322
rect 67 282 125 288
rect -263 238 -217 250
rect -263 -238 -257 238
rect -223 -238 -217 238
rect -263 -250 -217 -238
rect -167 238 -121 250
rect -167 -238 -161 238
rect -127 -238 -121 238
rect -167 -250 -121 -238
rect -71 238 -25 250
rect -71 -238 -65 238
rect -31 -238 -25 238
rect -71 -250 -25 -238
rect 25 238 71 250
rect 25 -238 31 238
rect 65 -238 71 238
rect 25 -250 71 -238
rect 121 238 167 250
rect 121 -238 127 238
rect 161 -238 167 238
rect 121 -250 167 -238
rect 217 238 263 250
rect 217 -238 223 238
rect 257 -238 263 238
rect 217 -250 263 -238
rect -221 -288 -163 -282
rect -221 -322 -209 -288
rect -175 -322 -163 -288
rect -221 -328 -163 -322
rect -29 -288 29 -282
rect -29 -322 -17 -288
rect 17 -322 29 -288
rect -29 -328 29 -322
rect 163 -288 221 -282
rect 163 -322 175 -288
rect 209 -322 221 -288
rect 163 -328 221 -322
<< properties >>
string FIXED_BBOX -354 -407 354 407
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2.5 l 0.150 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
