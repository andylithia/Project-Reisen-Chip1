* NGSPICE file created from swcap_array_1.ext - technology: sky130A

X0 tcap_200f_60/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X1 tcap_200f_60/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X3 tcap_200f_50/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X4 tcap_200f_50/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5 C tcap_200f_50/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X6 tcap_200f_61/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X7 tcap_200f_61/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8 C tcap_200f_61/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X9 tcap_200f_40/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X10 tcap_200f_40/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11 C tcap_200f_40/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X12 tcap_200f_51/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X13 tcap_200f_51/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14 C tcap_200f_51/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X15 tcap_200f_62/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X16 tcap_200f_62/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X17 C tcap_200f_62/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X18 tcap_200f_30/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X19 tcap_200f_30/a_173_157# B6 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X20 C tcap_200f_30/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X21 tcap_200f_41/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X22 tcap_200f_41/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X23 C tcap_200f_41/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X24 tcap_200f_52/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X25 tcap_200f_52/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X26 C tcap_200f_52/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X27 tcap_200f_63/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X28 tcap_200f_63/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X29 C tcap_200f_63/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X30 tcap_50f_0/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=7.85e+06u
X31 tcap_50f_0/a_173_157# B0 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X32 C tcap_50f_0/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=7.85e+06u
X33 tcap_200f_31/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X34 tcap_200f_31/a_173_157# B6 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X35 C tcap_200f_31/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X36 tcap_200f_42/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X37 tcap_200f_42/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X38 C tcap_200f_42/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X39 tcap_200f_20/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X40 tcap_200f_20/a_173_157# B6 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X41 C tcap_200f_20/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X42 tcap_200f_53/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X43 tcap_200f_53/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X44 C tcap_200f_53/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X45 tcap_200f_64/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X46 tcap_200f_64/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X47 C tcap_200f_64/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X48 tcap_200f_32/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X49 tcap_200f_32/a_173_157# B6 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X50 C tcap_200f_32/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X51 tcap_200f_33/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X52 tcap_200f_33/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X53 C tcap_200f_33/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X54 tcap_200f_43/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X55 tcap_200f_43/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X56 C tcap_200f_43/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X57 tcap_200f_22/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X58 tcap_200f_22/a_173_157# B6 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X59 C tcap_200f_22/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X60 tcap_200f_44/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X61 tcap_200f_44/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X62 C tcap_200f_44/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X63 tcap_200f_21/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X64 tcap_200f_21/a_173_157# B6 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X65 C tcap_200f_21/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X66 tcap_200f_10/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X67 tcap_200f_10/a_173_157# B5 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X68 C tcap_200f_10/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X69 tcap_200f_54/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X70 tcap_200f_54/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X71 C tcap_200f_54/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X72 tcap_200f_11/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X73 tcap_200f_11/a_173_157# B5 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X74 C tcap_200f_11/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X75 tcap_200f_55/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X76 tcap_200f_55/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X77 C tcap_200f_55/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X78 tcap_200f_65/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X79 tcap_200f_65/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X80 C tcap_200f_65/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X81 tcap_200f_34/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X82 tcap_200f_34/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X83 C tcap_200f_34/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X84 tcap_200f_23/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X85 tcap_200f_23/a_173_157# B6 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X86 C tcap_200f_23/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X87 tcap_200f_45/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X88 tcap_200f_45/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X89 C tcap_200f_45/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X90 tcap_200f_12/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X91 tcap_200f_12/a_173_157# B5 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X92 C tcap_200f_12/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X93 tcap_200f_0/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X94 tcap_200f_0/a_173_157# B5 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X95 C tcap_200f_0/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X96 tcap_200f_56/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X97 tcap_200f_56/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X98 C tcap_200f_56/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X99 tcap_200f_35/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X100 tcap_200f_35/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X101 C tcap_200f_35/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X102 tcap_200f_24/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X103 tcap_200f_24/a_173_157# B6 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X104 C tcap_200f_24/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X105 tcap_200f_46/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X106 tcap_200f_46/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X107 C tcap_200f_46/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X108 tcap_200f_13/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X109 tcap_200f_13/a_173_157# B5 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X110 C tcap_200f_13/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X111 tcap_200f_57/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X112 tcap_200f_57/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X113 C tcap_200f_57/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X114 tcap_200f_36/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X115 tcap_200f_36/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X116 C tcap_200f_36/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X117 tcap_200f_25/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X118 tcap_200f_25/a_173_157# B6 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X119 C tcap_200f_25/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X120 tcap_200f_47/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X121 tcap_200f_47/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X122 C tcap_200f_47/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X123 tcap_200f_14/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X124 tcap_200f_14/a_173_157# B5 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X125 C tcap_200f_14/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X126 tcap_200f_58/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X127 tcap_200f_58/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X128 C tcap_200f_58/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X129 tcap_200f_37/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X130 tcap_200f_37/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X131 C tcap_200f_37/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X132 tcap_200f_26/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X133 tcap_200f_26/a_173_157# B6 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X134 C tcap_200f_26/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X135 tcap_200f_15/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X136 tcap_200f_15/a_173_157# B6 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X137 C tcap_200f_15/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X138 tcap_200f_48/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X139 tcap_200f_48/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X140 C tcap_200f_48/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X141 tcap_200f_59/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X142 tcap_200f_59/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X143 C tcap_200f_59/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X144 tcap_200f_3/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X145 tcap_200f_3/a_173_157# B2 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X146 C tcap_200f_3/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X147 tcap_200f_38/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X148 tcap_200f_38/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X149 C tcap_200f_38/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X150 tcap_200f_27/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X151 tcap_200f_27/a_173_157# B6 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X152 C tcap_200f_27/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X153 tcap_200f_16/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X154 tcap_200f_16/a_173_157# B5 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X155 C tcap_200f_16/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X156 tcap_200f_49/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X157 tcap_200f_49/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X158 C tcap_200f_49/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X159 tcap_200f_4/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X160 tcap_200f_4/a_173_157# B3 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X161 C tcap_200f_4/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X162 tcap_200f_28/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X163 tcap_200f_28/a_173_157# B6 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X164 C tcap_200f_28/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X165 tcap_200f_39/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X166 tcap_200f_39/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X167 C tcap_200f_39/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X168 tcap_200f_17/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X169 tcap_200f_17/a_173_157# B5 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X170 C tcap_200f_17/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X171 tcap_200f_5/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X172 tcap_200f_5/a_173_157# B3 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X173 C tcap_200f_5/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X174 tcap_200f_29/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X175 tcap_200f_29/a_173_157# B6 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X176 C tcap_200f_29/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X177 tcap_200f_18/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X178 tcap_200f_18/a_173_157# B6 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X179 C tcap_200f_18/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X180 tcap_200f_6/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X181 tcap_200f_6/a_173_157# B4 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X182 C tcap_200f_6/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X183 tcap_200f_19/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X184 tcap_200f_19/a_173_157# B6 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X185 C tcap_200f_19/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X186 tcap_200f_8/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X187 tcap_200f_8/a_173_157# B4 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X188 C tcap_200f_8/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X189 tcap_200f_7/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X190 tcap_200f_7/a_173_157# B4 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X191 C tcap_200f_7/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X192 tcap_200f_9/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X193 tcap_200f_9/a_173_157# B4 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X194 C tcap_200f_9/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X195 tcap_100f_0/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=1.57e+07u
X196 tcap_100f_0/a_173_157# B1 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X197 C tcap_100f_0/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=1.57e+07u
C0 C tcap_100f_0/a_173_157# 5.85fF
C1 tcap_200f_36/a_173_157# tcap_200f_37/a_173_157# 4.48fF
C2 tcap_200f_38/a_173_157# tcap_200f_37/a_173_157# 4.48fF
C3 tcap_200f_28/a_173_157# tcap_200f_31/a_173_157# 4.47fF
C4 tcap_200f_10/a_173_157# tcap_200f_13/a_173_157# 4.47fF
C5 tcap_200f_45/a_173_157# C 12.05fF
C6 tcap_200f_44/a_173_157# C 12.05fF
C7 tcap_200f_16/a_173_157# tcap_200f_14/a_173_157# 4.47fF
C8 C tcap_200f_52/a_173_157# 12.05fF
C9 tcap_200f_57/a_173_157# tcap_200f_58/a_173_157# 4.48fF
C10 tcap_200f_17/a_173_157# tcap_200f_16/a_173_157# 4.47fF
C11 tcap_200f_18/a_173_157# C 12.05fF
C12 tcap_200f_12/a_173_157# C 12.05fF
C13 tcap_200f_47/a_173_157# tcap_200f_46/a_173_157# 4.48fF
C14 tcap_200f_49/a_173_157# tcap_200f_50/a_173_157# 4.48fF
C15 tcap_200f_56/a_173_157# C 12.05fF
C16 tcap_200f_54/a_173_157# tcap_200f_53/a_173_157# 4.48fF
C17 tcap_200f_41/a_173_157# tcap_200f_40/a_173_157# 4.48fF
C18 tcap_200f_15/a_173_157# C 12.05fF
C19 C tcap_200f_7/a_173_157# 12.05fF
C20 tcap_200f_15/a_173_157# tcap_200f_25/a_173_157# 4.47fF
C21 tcap_200f_36/a_173_157# C 12.05fF
C22 tcap_200f_38/a_173_157# C 12.05fF
C23 tcap_200f_5/a_173_157# C 12.05fF
C24 tcap_200f_22/a_173_157# C 12.05fF
C25 tcap_200f_42/a_173_157# C 12.05fF
C26 tcap_200f_48/a_173_157# tcap_200f_47/a_173_157# 4.48fF
C27 tcap_200f_34/a_173_157# C 11.79fF
C28 tcap_200f_52/a_173_157# tcap_200f_53/a_173_157# 4.48fF
C29 C tcap_200f_6/a_173_157# 12.05fF
C30 tcap_200f_44/a_173_157# tcap_200f_43/a_173_157# 4.48fF
C31 tcap_200f_31/a_173_157# tcap_200f_30/a_173_157# 4.47fF
C32 tcap_200f_36/a_173_157# tcap_200f_35/a_173_157# 4.48fF
C33 tcap_200f_39/a_173_157# C 12.05fF
C34 tcap_200f_45/a_173_157# tcap_200f_46/a_173_157# 4.48fF
C35 tcap_200f_4/a_173_157# tcap_200f_3/a_173_157# 4.47fF
C36 tcap_200f_16/a_173_157# C 12.05fF
C37 tcap_200f_59/a_173_157# C 12.05fF
C38 tcap_200f_14/a_173_157# C 12.05fF
C39 tcap_200f_23/a_173_157# tcap_200f_22/a_173_157# 4.47fF
C40 tcap_200f_34/a_173_157# tcap_200f_35/a_173_157# 4.48fF
C41 tcap_200f_61/a_173_157# tcap_200f_62/a_173_157# 4.48fF
C42 tcap_200f_55/a_173_157# tcap_200f_54/a_173_157# 4.48fF
C43 C tcap_200f_37/a_173_157# 12.05fF
C44 tcap_200f_15/a_173_157# tcap_200f_27/a_173_157# 4.47fF
C45 tcap_200f_51/a_173_157# tcap_200f_50/a_173_157# 4.48fF
C46 tcap_200f_63/a_173_157# tcap_200f_62/a_173_157# 4.48fF
C47 tcap_200f_57/a_173_157# tcap_200f_56/a_173_157# 4.48fF
C48 tcap_200f_17/a_173_157# C 12.05fF
C49 tcap_200f_11/a_173_157# tcap_200f_0/a_173_157# 4.47fF
C50 tcap_50f_0/a_173_157# C 3.01fF
C51 tcap_200f_8/a_173_157# tcap_200f_7/a_173_157# 4.47fF
C52 tcap_200f_11/a_173_157# C 12.05fF
C53 tcap_200f_42/a_173_157# tcap_200f_43/a_173_157# 4.48fF
C54 tcap_200f_60/a_173_157# tcap_200f_61/a_173_157# 4.48fF
C55 tcap_200f_3/a_173_157# tcap_100f_0/a_173_157# 2.53fF
C56 tcap_200f_21/a_173_157# tcap_200f_22/a_173_157# 4.47fF
C57 tcap_200f_0/a_173_157# C 12.05fF
C58 tcap_200f_24/a_173_157# C 12.05fF
C59 tcap_200f_52/a_173_157# tcap_200f_51/a_173_157# 4.48fF
C60 tcap_200f_55/a_173_157# tcap_200f_56/a_173_157# 4.48fF
C61 tcap_200f_24/a_173_157# tcap_200f_25/a_173_157# 4.47fF
C62 tcap_200f_64/a_173_157# C 11.71fF
C63 tcap_200f_29/a_173_157# C 12.05fF
C64 B4 B5 3.35fF
C65 tcap_200f_20/a_173_157# C 12.05fF
C66 tcap_200f_42/a_173_157# tcap_200f_41/a_173_157# 4.48fF
C67 tcap_200f_25/a_173_157# C 12.05fF
C68 tcap_200f_18/a_173_157# tcap_200f_19/a_173_157# 4.47fF
C69 tcap_200f_23/a_173_157# tcap_200f_24/a_173_157# 4.47fF
C70 tcap_200f_10/a_173_157# tcap_200f_11/a_173_157# 4.47fF
C71 tcap_200f_12/a_173_157# tcap_200f_13/a_173_157# 4.47fF
C72 C tcap_200f_35/a_173_157# 12.05fF
C73 tcap_200f_5/a_173_157# tcap_200f_4/a_173_157# 4.47fF
C74 B5 B6 6.53fF
C75 tcap_200f_29/a_173_157# tcap_200f_28/a_173_157# 4.47fF
C76 tcap_200f_23/a_173_157# C 12.05fF
C77 tcap_200f_26/a_173_157# tcap_200f_29/a_173_157# 4.47fF
C78 tcap_200f_28/a_173_157# C 12.05fF
C79 tcap_200f_44/a_173_157# tcap_200f_45/a_173_157# 4.48fF
C80 tcap_200f_26/a_173_157# C 12.05fF
C81 tcap_200f_9/a_173_157# tcap_200f_0/a_173_157# 4.47fF
C82 tcap_200f_32/a_173_157# C 11.60fF
C83 tcap_200f_10/a_173_157# C 12.05fF
C84 tcap_200f_27/a_173_157# C 12.05fF
C85 tcap_200f_39/a_173_157# tcap_200f_40/a_173_157# 4.48fF
C86 tcap_200f_34/a_173_157# tcap_200f_33/a_173_157# 4.48fF
C87 C tcap_200f_53/a_173_157# 12.05fF
C88 tcap_200f_57/a_173_157# C 12.05fF
C89 tcap_200f_43/a_173_157# C 12.05fF
C90 tcap_200f_9/a_173_157# C 12.05fF
C91 tcap_200f_49/a_173_157# C 12.05fF
C92 C tcap_200f_8/a_173_157# 12.05fF
C93 C tcap_200f_46/a_173_157# 12.05fF
C94 tcap_200f_21/a_173_157# C 12.05fF
C95 tcap_200f_21/a_173_157# tcap_200f_20/a_173_157# 4.47fF
C96 tcap_200f_59/a_173_157# tcap_200f_58/a_173_157# 4.48fF
C97 tcap_200f_64/a_173_157# tcap_200f_65/a_173_157# 4.48fF
C98 C tcap_200f_65/a_173_157# 10.91fF
C99 tcap_200f_41/a_173_157# C 12.05fF
C100 tcap_200f_26/a_173_157# tcap_200f_27/a_173_157# 4.47fF
C101 tcap_200f_48/a_173_157# C 12.05fF
C102 tcap_200f_55/a_173_157# C 12.05fF
C103 tcap_200f_59/a_173_157# tcap_200f_60/a_173_157# 4.48fF
C104 C tcap_200f_30/a_173_157# 11.79fF
C105 tcap_200f_4/a_173_157# C 11.89fF
C106 B7 B6 9.55fF
C107 C tcap_200f_62/a_173_157# 12.05fF
C108 C tcap_200f_51/a_173_157# 12.05fF
C109 tcap_200f_19/a_173_157# C 12.05fF
C110 tcap_200f_19/a_173_157# tcap_200f_20/a_173_157# 4.47fF
C111 tcap_200f_9/a_173_157# tcap_200f_8/a_173_157# 4.47fF
C112 C tcap_200f_40/a_173_157# 12.05fF
C113 C tcap_200f_13/a_173_157# 12.05fF
C114 tcap_200f_6/a_173_157# tcap_200f_7/a_173_157# 4.47fF
C115 C tcap_200f_3/a_173_157# 11.41fF
C116 tcap_200f_33/a_173_157# C 11.60fF
C117 tcap_200f_61/a_173_157# C 12.05fF
C118 tcap_200f_14/a_173_157# tcap_200f_12/a_173_157# 4.47fF
C119 tcap_200f_47/a_173_157# C 12.05fF
C120 tcap_200f_58/a_173_157# C 12.05fF
C121 C tcap_200f_31/a_173_157# 12.05fF
C122 tcap_200f_64/a_173_157# tcap_200f_63/a_173_157# 4.48fF
C123 tcap_200f_5/a_173_157# tcap_200f_6/a_173_157# 4.47fF
C124 tcap_200f_32/a_173_157# tcap_200f_30/a_173_157# 4.47fF
C125 C tcap_200f_50/a_173_157# 12.05fF
C126 tcap_200f_39/a_173_157# tcap_200f_38/a_173_157# 4.48fF
C127 C tcap_200f_63/a_173_157# 12.04fF
C128 tcap_200f_18/a_173_157# tcap_200f_17/a_173_157# 4.47fF
C129 tcap_200f_48/a_173_157# tcap_200f_49/a_173_157# 4.48fF
C130 tcap_200f_60/a_173_157# C 12.05fF
C131 tcap_200f_54/a_173_157# C 12.05fF
C132 tcap_100f_0/a_173_157# VSUB 4.99fF $ **FLOATING
C133 tcap_200f_9/a_173_157# VSUB 7.94fF $ **FLOATING
C134 tcap_200f_7/a_173_157# VSUB 7.94fF $ **FLOATING
C135 tcap_200f_8/a_173_157# VSUB 7.94fF $ **FLOATING
C136 tcap_200f_19/a_173_157# VSUB 7.94fF $ **FLOATING
C137 tcap_200f_6/a_173_157# VSUB 7.94fF $ **FLOATING
C138 B4 VSUB 5.01fF $ **FLOATING
C139 tcap_200f_18/a_173_157# VSUB 7.94fF $ **FLOATING
C140 B6 VSUB 22.15fF $ **FLOATING
C141 tcap_200f_29/a_173_157# VSUB 7.94fF $ **FLOATING
C142 tcap_200f_5/a_173_157# VSUB 7.94fF $ **FLOATING
C143 tcap_200f_17/a_173_157# VSUB 7.94fF $ **FLOATING
C144 tcap_200f_39/a_173_157# VSUB 7.96fF $ **FLOATING
C145 tcap_200f_28/a_173_157# VSUB 7.94fF $ **FLOATING
C146 tcap_200f_4/a_173_157# VSUB 7.94fF $ **FLOATING
C147 B3 VSUB 2.41fF $ **FLOATING
C148 tcap_200f_49/a_173_157# VSUB 7.96fF $ **FLOATING
C149 tcap_200f_16/a_173_157# VSUB 7.94fF $ **FLOATING
C150 tcap_200f_27/a_173_157# VSUB 7.94fF $ **FLOATING
C151 tcap_200f_38/a_173_157# VSUB 7.96fF $ **FLOATING
C152 tcap_200f_3/a_173_157# VSUB 7.94fF $ **FLOATING
C153 tcap_200f_59/a_173_157# VSUB 7.95fF $ **FLOATING
C154 tcap_200f_48/a_173_157# VSUB 7.96fF $ **FLOATING
C155 tcap_200f_15/a_173_157# VSUB 7.94fF $ **FLOATING
C156 tcap_200f_26/a_173_157# VSUB 7.94fF $ **FLOATING
C157 tcap_200f_37/a_173_157# VSUB 7.96fF $ **FLOATING
C158 tcap_200f_58/a_173_157# VSUB 7.95fF $ **FLOATING
C159 tcap_200f_14/a_173_157# VSUB 7.94fF $ **FLOATING
C160 tcap_200f_47/a_173_157# VSUB 7.96fF $ **FLOATING
C161 tcap_200f_25/a_173_157# VSUB 7.94fF $ **FLOATING
C162 tcap_200f_36/a_173_157# VSUB 7.96fF $ **FLOATING
C163 tcap_200f_57/a_173_157# VSUB 7.95fF $ **FLOATING
C164 tcap_200f_13/a_173_157# VSUB 7.94fF $ **FLOATING
C165 tcap_200f_46/a_173_157# VSUB 7.96fF $ **FLOATING
C166 tcap_200f_24/a_173_157# VSUB 7.94fF $ **FLOATING
C167 tcap_200f_35/a_173_157# VSUB 7.96fF $ **FLOATING
C168 tcap_200f_56/a_173_157# VSUB 7.95fF $ **FLOATING
C169 tcap_200f_0/a_173_157# VSUB 7.94fF $ **FLOATING
C170 B5 VSUB 10.51fF $ **FLOATING
C171 tcap_200f_12/a_173_157# VSUB 7.94fF $ **FLOATING
C172 tcap_200f_45/a_173_157# VSUB 7.96fF $ **FLOATING
C173 tcap_200f_23/a_173_157# VSUB 7.94fF $ **FLOATING
C174 tcap_200f_34/a_173_157# VSUB 7.95fF $ **FLOATING
C175 C VSUB 71.74fF $ **FLOATING
C176 tcap_200f_65/a_173_157# VSUB 7.92fF $ **FLOATING
C177 B7 VSUB 28.92fF $ **FLOATING
C178 tcap_200f_55/a_173_157# VSUB 7.95fF $ **FLOATING
C179 tcap_200f_11/a_173_157# VSUB 7.94fF $ **FLOATING
C180 tcap_200f_54/a_173_157# VSUB 7.95fF $ **FLOATING
C181 tcap_200f_10/a_173_157# VSUB 7.94fF $ **FLOATING
C182 tcap_200f_21/a_173_157# VSUB 7.94fF $ **FLOATING
C183 tcap_200f_44/a_173_157# VSUB 7.96fF $ **FLOATING
C184 tcap_200f_22/a_173_157# VSUB 7.94fF $ **FLOATING
C185 tcap_200f_43/a_173_157# VSUB 7.96fF $ **FLOATING
C186 tcap_200f_33/a_173_157# VSUB 7.96fF $ **FLOATING
C187 tcap_200f_32/a_173_157# VSUB 7.96fF $ **FLOATING
C188 tcap_200f_64/a_173_157# VSUB 7.93fF $ **FLOATING
C189 tcap_200f_53/a_173_157# VSUB 7.95fF $ **FLOATING
C190 tcap_200f_20/a_173_157# VSUB 7.94fF $ **FLOATING
C191 tcap_200f_42/a_173_157# VSUB 7.96fF $ **FLOATING
C192 tcap_200f_31/a_173_157# VSUB 7.94fF $ **FLOATING
C193 tcap_50f_0/a_173_157# VSUB 3.60fF $ **FLOATING
C194 tcap_200f_63/a_173_157# VSUB 7.94fF $ **FLOATING
C195 tcap_200f_52/a_173_157# VSUB 7.95fF $ **FLOATING
C196 tcap_200f_41/a_173_157# VSUB 7.96fF $ **FLOATING
C197 tcap_200f_30/a_173_157# VSUB 7.94fF $ **FLOATING
C198 tcap_200f_62/a_173_157# VSUB 7.94fF $ **FLOATING
C199 tcap_200f_51/a_173_157# VSUB 7.95fF $ **FLOATING
C200 tcap_200f_40/a_173_157# VSUB 7.96fF $ **FLOATING
C201 tcap_200f_61/a_173_157# VSUB 7.95fF $ **FLOATING
C202 tcap_200f_50/a_173_157# VSUB 7.95fF $ **FLOATING
C203 tcap_200f_60/a_173_157# VSUB 7.95fF $ **FLOATING
