magic
tech sky130A
magscale 1 2
timestamp 1671388962
<< nwell >>
rect -2918 1664 4934 2036
rect -2918 628 4934 1000
rect -1766 332 4934 628
<< pwell >>
rect -1888 3552 -1466 3682
rect -1888 3499 -1708 3552
rect -1654 3499 -1466 3552
rect -1888 2838 -1466 3499
rect -1888 2785 -1708 2838
rect -1654 2785 -1466 2838
rect -1888 2148 -1466 2785
rect -1106 3552 -684 3682
rect -1106 3499 -918 3552
rect -864 3499 -684 3552
rect -1106 2838 -684 3499
rect -1106 2785 -918 2838
rect -864 2785 -684 2838
rect -1106 2148 -684 2785
rect -2805 1381 -2595 1580
rect -1436 1381 -1162 1580
rect -1136 1381 -519 1527
rect 5 1381 187 1587
rect 208 1381 825 1527
rect 880 1381 1497 1527
rect 1552 1381 2169 1527
rect 2224 1381 2841 1527
rect 2896 1381 3513 1527
rect 3568 1381 4185 1527
rect 4240 1381 4602 1527
rect -2880 1283 4896 1381
rect -2805 1084 -2595 1283
rect -1436 1084 -1162 1283
rect -1151 1084 -291 1283
rect -284 1084 -2 1283
rect 5 1077 187 1283
rect 198 1140 3839 1283
rect 198 1114 2265 1140
rect 198 1103 2170 1114
rect 854 1097 2170 1103
rect 854 1060 1218 1097
rect 1639 1071 2170 1097
rect 2538 1084 3839 1140
rect 3841 1084 4031 1283
rect 4033 1084 4895 1283
rect 2935 1042 3123 1084
rect -1653 49 -1443 248
rect -284 49 -10 248
rect 5 49 187 255
rect 854 235 1218 272
rect 1639 235 2170 261
rect 2935 248 3123 290
rect 854 229 2170 235
rect 198 218 2170 229
rect 198 192 2265 218
rect 2538 192 3839 248
rect 198 49 3839 192
rect 3841 49 4031 248
rect 4033 49 4895 273
rect -1728 0 4896 49
rect -1539 -218 -1117 -88
rect -1539 -271 -1351 -218
rect -1297 -271 -1117 -218
rect -1539 -932 -1117 -271
rect -1539 -985 -1351 -932
rect -1297 -985 -1117 -932
rect -1539 -1622 -1117 -985
<< nmos >>
rect -1692 3072 -1662 3472
rect -1692 2358 -1662 2758
rect -910 3072 -880 3472
rect -910 2358 -880 2758
rect -1343 -698 -1313 -298
rect -1343 -1412 -1313 -1012
<< scpmos >>
rect -2710 1700 -2680 1924
rect -1356 1700 -1326 1924
rect -1266 1700 -1236 1924
rect -1070 1724 -870 1924
rect -815 1724 -615 1924
rect 274 1724 474 1924
rect 529 1724 729 1924
rect 946 1724 1146 1924
rect 1201 1724 1401 1924
rect 1618 1724 1818 1924
rect 1873 1724 2073 1924
rect 2290 1724 2490 1924
rect 2545 1724 2745 1924
rect 2962 1724 3162 1924
rect 3217 1724 3417 1924
rect 3634 1724 3834 1924
rect 3889 1724 4089 1924
rect 4306 1724 4506 1924
rect -2710 740 -2680 964
rect -1356 740 -1326 964
rect -1266 740 -1236 964
rect -1066 796 -1036 964
rect -959 764 -929 964
rect -766 764 -736 964
rect -658 764 -628 964
rect -544 764 -514 964
rect -420 740 -390 964
rect -204 740 -174 964
rect -114 740 -84 964
rect 278 740 308 868
rect 368 740 398 868
rect 446 740 476 868
rect 536 740 566 868
rect 738 740 768 868
rect 940 740 970 964
rect 1030 740 1060 964
rect 1232 784 1262 868
rect 1316 784 1346 868
rect 1423 740 1453 868
rect 1754 740 1784 908
rect 1838 740 1868 908
rect 1946 740 1976 908
rect 2148 740 2178 908
rect 2226 740 2256 908
rect 2333 740 2363 824
rect 2411 740 2441 824
rect 2616 740 2646 940
rect 2718 740 2748 940
rect 2802 740 2832 940
rect 3004 805 3034 933
rect 3240 740 3270 964
rect 3330 740 3360 964
rect 3529 748 3559 948
rect 3634 740 3664 964
rect 3724 740 3754 964
rect 4119 740 4149 964
rect 4371 740 4401 964
rect 4471 740 4501 964
rect 4770 740 4800 964
rect -1558 368 -1528 592
rect -204 368 -174 592
rect -114 368 -84 592
rect 278 464 308 592
rect 368 464 398 592
rect 446 464 476 592
rect 536 464 566 592
rect 738 464 768 592
rect 940 368 970 592
rect 1030 368 1060 592
rect 1232 464 1262 548
rect 1316 464 1346 548
rect 1423 464 1453 592
rect 1754 424 1784 592
rect 1838 424 1868 592
rect 1946 424 1976 592
rect 2148 424 2178 592
rect 2226 424 2256 592
rect 2333 508 2363 592
rect 2411 508 2441 592
rect 2616 392 2646 592
rect 2718 392 2748 592
rect 2802 392 2832 592
rect 3004 399 3034 527
rect 3240 368 3270 592
rect 3330 368 3360 592
rect 3529 384 3559 584
rect 3634 368 3664 592
rect 3724 368 3754 592
rect 4119 409 4149 577
rect 4209 409 4239 577
rect 4304 409 4334 577
rect 4399 409 4429 577
rect 4506 368 4536 592
rect 4600 368 4630 592
rect 4690 368 4720 592
rect 4780 368 4810 592
<< nmoslvt >>
rect -2708 1406 -2678 1554
rect -1353 1406 -1323 1554
rect -1275 1406 -1245 1554
rect -1057 1417 -857 1501
rect -801 1417 -601 1501
rect 287 1417 487 1501
rect 543 1417 743 1501
rect 959 1417 1159 1501
rect 1215 1417 1415 1501
rect 1631 1417 1831 1501
rect 1887 1417 2087 1501
rect 2303 1417 2503 1501
rect 2559 1417 2759 1501
rect 2975 1417 3175 1501
rect 3231 1417 3431 1501
rect 3647 1417 3847 1501
rect 3903 1417 4103 1501
rect 4319 1417 4519 1501
rect -2708 1110 -2678 1258
rect -1353 1110 -1323 1258
rect -1275 1110 -1245 1258
rect -1068 1110 -1038 1220
rect -956 1110 -926 1258
rect -878 1110 -848 1258
rect -739 1110 -709 1258
rect -547 1110 -517 1258
rect -404 1110 -374 1258
rect -201 1110 -171 1258
rect -115 1110 -85 1258
rect 281 1129 311 1213
rect 359 1129 389 1213
rect 525 1129 555 1213
rect 603 1129 633 1213
rect 739 1129 769 1213
rect 937 1086 967 1234
rect 1105 1086 1135 1234
rect 1347 1123 1377 1207
rect 1419 1123 1449 1207
rect 1510 1123 1540 1207
rect 1757 1097 1787 1207
rect 1843 1097 1873 1207
rect 1964 1097 1994 1207
rect 2064 1097 2094 1207
rect 2159 1140 2189 1250
rect 2409 1166 2439 1250
rect 2487 1166 2517 1250
rect 2614 1110 2644 1258
rect 2718 1110 2748 1258
rect 2804 1110 2834 1258
rect 3017 1068 3047 1152
rect 3223 1110 3253 1258
rect 3309 1110 3339 1258
rect 3521 1110 3551 1238
rect 3641 1110 3671 1258
rect 3727 1110 3757 1258
rect 4116 1110 4146 1258
rect 4202 1110 4232 1258
rect 4288 1110 4318 1258
rect 4374 1110 4404 1258
rect 4468 1110 4498 1258
rect 4560 1110 4590 1258
rect 4660 1110 4690 1258
rect 4773 1110 4803 1258
rect -1556 74 -1526 222
rect -201 74 -171 222
rect -123 74 -93 222
rect 281 119 311 203
rect 359 119 389 203
rect 525 119 555 203
rect 603 119 633 203
rect 739 119 769 203
rect 937 98 967 246
rect 1105 98 1135 246
rect 1347 125 1377 209
rect 1419 125 1449 209
rect 1510 125 1540 209
rect 1757 125 1787 235
rect 1843 125 1873 235
rect 1964 125 1994 235
rect 2064 125 2094 235
rect 2159 82 2189 192
rect 2409 82 2439 166
rect 2487 82 2517 166
rect 2614 74 2644 222
rect 2718 74 2748 222
rect 2804 74 2834 222
rect 3017 180 3047 264
rect 3223 74 3253 222
rect 3309 74 3339 222
rect 3521 94 3551 222
rect 3641 74 3671 222
rect 3727 74 3757 222
rect 4116 119 4146 247
rect 4206 119 4236 247
rect 4301 119 4331 247
rect 4392 119 4422 247
rect 4494 99 4524 247
rect 4610 99 4640 247
rect 4696 99 4726 247
rect 4782 99 4812 247
<< ndiff >>
rect -1750 3460 -1692 3472
rect -1750 3084 -1738 3460
rect -1704 3084 -1692 3460
rect -1750 3072 -1692 3084
rect -1662 3460 -1604 3472
rect -1662 3084 -1650 3460
rect -1616 3084 -1604 3460
rect -1662 3072 -1604 3084
rect -1750 2746 -1692 2758
rect -1750 2370 -1738 2746
rect -1704 2370 -1692 2746
rect -1750 2358 -1692 2370
rect -1662 2746 -1604 2758
rect -1662 2370 -1650 2746
rect -1616 2370 -1604 2746
rect -1662 2358 -1604 2370
rect -968 3460 -910 3472
rect -968 3084 -956 3460
rect -922 3084 -910 3460
rect -968 3072 -910 3084
rect -880 3460 -822 3472
rect -880 3084 -868 3460
rect -834 3084 -822 3460
rect -880 3072 -822 3084
rect -968 2746 -910 2758
rect -968 2370 -956 2746
rect -922 2370 -910 2746
rect -968 2358 -910 2370
rect -880 2746 -822 2758
rect -880 2370 -868 2746
rect -834 2370 -822 2746
rect -880 2358 -822 2370
rect -2779 1542 -2708 1554
rect -2779 1508 -2767 1542
rect -2733 1508 -2708 1542
rect -2779 1452 -2708 1508
rect -2779 1418 -2767 1452
rect -2733 1418 -2708 1452
rect -2779 1406 -2708 1418
rect -2678 1542 -2621 1554
rect -2678 1508 -2667 1542
rect -2633 1508 -2621 1542
rect -2678 1452 -2621 1508
rect -1410 1534 -1353 1554
rect -1410 1500 -1398 1534
rect -1364 1500 -1353 1534
rect -2678 1418 -2667 1452
rect -2633 1418 -2621 1452
rect -2678 1406 -2621 1418
rect -1410 1452 -1353 1500
rect -1410 1418 -1398 1452
rect -1364 1418 -1353 1452
rect -1410 1406 -1353 1418
rect -1323 1406 -1275 1554
rect -1245 1534 -1188 1554
rect -1245 1500 -1234 1534
rect -1200 1500 -1188 1534
rect -1245 1452 -1188 1500
rect -1245 1418 -1234 1452
rect -1200 1418 -1188 1452
rect -1245 1406 -1188 1418
rect -1110 1477 -1057 1501
rect -1110 1443 -1102 1477
rect -1068 1443 -1057 1477
rect -1110 1417 -1057 1443
rect -857 1477 -801 1501
rect -857 1443 -846 1477
rect -812 1443 -801 1477
rect -857 1417 -801 1443
rect -601 1477 -545 1501
rect -601 1443 -590 1477
rect -556 1443 -545 1477
rect -601 1417 -545 1443
rect 234 1477 287 1501
rect 234 1443 242 1477
rect 276 1443 287 1477
rect 234 1417 287 1443
rect 487 1477 543 1501
rect 487 1443 498 1477
rect 532 1443 543 1477
rect 487 1417 543 1443
rect 743 1477 799 1501
rect 743 1443 754 1477
rect 788 1443 799 1477
rect 743 1417 799 1443
rect 906 1477 959 1501
rect 906 1443 914 1477
rect 948 1443 959 1477
rect 906 1417 959 1443
rect 1159 1477 1215 1501
rect 1159 1443 1170 1477
rect 1204 1443 1215 1477
rect 1159 1417 1215 1443
rect 1415 1477 1471 1501
rect 1415 1443 1426 1477
rect 1460 1443 1471 1477
rect 1415 1417 1471 1443
rect 1578 1477 1631 1501
rect 1578 1443 1586 1477
rect 1620 1443 1631 1477
rect 1578 1417 1631 1443
rect 1831 1477 1887 1501
rect 1831 1443 1842 1477
rect 1876 1443 1887 1477
rect 1831 1417 1887 1443
rect 2087 1477 2143 1501
rect 2087 1443 2098 1477
rect 2132 1443 2143 1477
rect 2087 1417 2143 1443
rect 2250 1477 2303 1501
rect 2250 1443 2258 1477
rect 2292 1443 2303 1477
rect 2250 1417 2303 1443
rect 2503 1477 2559 1501
rect 2503 1443 2514 1477
rect 2548 1443 2559 1477
rect 2503 1417 2559 1443
rect 2759 1477 2815 1501
rect 2759 1443 2770 1477
rect 2804 1443 2815 1477
rect 2759 1417 2815 1443
rect 2922 1477 2975 1501
rect 2922 1443 2930 1477
rect 2964 1443 2975 1477
rect 2922 1417 2975 1443
rect 3175 1477 3231 1501
rect 3175 1443 3186 1477
rect 3220 1443 3231 1477
rect 3175 1417 3231 1443
rect 3431 1477 3487 1501
rect 3431 1443 3442 1477
rect 3476 1443 3487 1477
rect 3431 1417 3487 1443
rect 3594 1477 3647 1501
rect 3594 1443 3602 1477
rect 3636 1443 3647 1477
rect 3594 1417 3647 1443
rect 3847 1477 3903 1501
rect 3847 1443 3858 1477
rect 3892 1443 3903 1477
rect 3847 1417 3903 1443
rect 4103 1477 4159 1501
rect 4103 1443 4114 1477
rect 4148 1443 4159 1477
rect 4103 1417 4159 1443
rect 4266 1477 4319 1501
rect 4266 1443 4274 1477
rect 4308 1443 4319 1477
rect 4266 1417 4319 1443
rect 4519 1477 4576 1501
rect 4519 1443 4530 1477
rect 4564 1443 4576 1477
rect 4519 1417 4576 1443
rect -2779 1246 -2708 1258
rect -2779 1212 -2767 1246
rect -2733 1212 -2708 1246
rect -2779 1156 -2708 1212
rect -2779 1122 -2767 1156
rect -2733 1122 -2708 1156
rect -2779 1110 -2708 1122
rect -2678 1246 -2621 1258
rect -2678 1212 -2667 1246
rect -2633 1212 -2621 1246
rect -2678 1156 -2621 1212
rect -1410 1246 -1353 1258
rect -1410 1212 -1398 1246
rect -1364 1212 -1353 1246
rect -2678 1122 -2667 1156
rect -2633 1122 -2621 1156
rect -2678 1110 -2621 1122
rect -1410 1164 -1353 1212
rect -1410 1130 -1398 1164
rect -1364 1130 -1353 1164
rect -1410 1110 -1353 1130
rect -1323 1110 -1275 1258
rect -1245 1246 -1188 1258
rect -1023 1246 -956 1258
rect -1245 1212 -1234 1246
rect -1200 1212 -1188 1246
rect -1023 1220 -1006 1246
rect -1245 1164 -1188 1212
rect -1245 1130 -1234 1164
rect -1200 1130 -1188 1164
rect -1245 1110 -1188 1130
rect -1125 1182 -1068 1220
rect -1125 1148 -1113 1182
rect -1079 1148 -1068 1182
rect -1125 1110 -1068 1148
rect -1038 1212 -1006 1220
rect -972 1212 -956 1246
rect -1038 1156 -956 1212
rect -1038 1122 -1024 1156
rect -990 1122 -956 1156
rect -1038 1110 -956 1122
rect -926 1110 -878 1258
rect -848 1238 -739 1258
rect -848 1204 -811 1238
rect -777 1204 -739 1238
rect -848 1110 -739 1204
rect -709 1110 -547 1258
rect -517 1220 -404 1258
rect -517 1186 -477 1220
rect -443 1186 -404 1220
rect -517 1110 -404 1186
rect -374 1246 -317 1258
rect -374 1212 -363 1246
rect -329 1212 -317 1246
rect -374 1156 -317 1212
rect -374 1122 -363 1156
rect -329 1122 -317 1156
rect -374 1110 -317 1122
rect -258 1246 -201 1258
rect -258 1212 -246 1246
rect -212 1212 -201 1246
rect -258 1156 -201 1212
rect -258 1122 -246 1156
rect -212 1122 -201 1156
rect -258 1110 -201 1122
rect -171 1246 -115 1258
rect -171 1212 -160 1246
rect -126 1212 -115 1246
rect -171 1156 -115 1212
rect -171 1122 -160 1156
rect -126 1122 -115 1156
rect -171 1110 -115 1122
rect -85 1246 -28 1258
rect -85 1212 -74 1246
rect -40 1212 -28 1246
rect -85 1156 -28 1212
rect -85 1122 -74 1156
rect -40 1122 -28 1156
rect -85 1110 -28 1122
rect 982 1284 1040 1296
rect 982 1250 994 1284
rect 1028 1250 1040 1284
rect 982 1234 1040 1250
rect 1270 1248 1332 1260
rect 224 1196 281 1213
rect 224 1162 236 1196
rect 270 1162 281 1196
rect 224 1129 281 1162
rect 311 1129 359 1213
rect 389 1191 525 1213
rect 389 1157 400 1191
rect 434 1157 480 1191
rect 514 1157 525 1191
rect 389 1129 525 1157
rect 555 1129 603 1213
rect 633 1197 739 1213
rect 633 1163 644 1197
rect 678 1163 739 1197
rect 633 1129 739 1163
rect 769 1186 826 1213
rect 769 1152 780 1186
rect 814 1152 826 1186
rect 769 1129 826 1152
rect 880 1132 937 1234
rect 880 1098 892 1132
rect 926 1098 937 1132
rect 880 1086 937 1098
rect 967 1086 1105 1234
rect 1135 1197 1192 1234
rect 1135 1163 1146 1197
rect 1180 1163 1192 1197
rect 1135 1129 1192 1163
rect 1135 1095 1146 1129
rect 1180 1095 1192 1129
rect 1270 1214 1284 1248
rect 1318 1214 1332 1248
rect 1270 1207 1332 1214
rect 1665 1247 1742 1259
rect 2532 1280 2599 1292
rect 2532 1250 2548 1280
rect 1665 1213 1686 1247
rect 1720 1213 1742 1247
rect 1665 1207 1742 1213
rect 2109 1207 2159 1250
rect 1270 1123 1347 1207
rect 1377 1123 1419 1207
rect 1449 1182 1510 1207
rect 1449 1148 1465 1182
rect 1499 1148 1510 1182
rect 1449 1123 1510 1148
rect 1540 1187 1611 1207
rect 1540 1153 1565 1187
rect 1599 1153 1611 1187
rect 1540 1123 1611 1153
rect 1135 1086 1192 1095
rect 1665 1097 1757 1207
rect 1787 1177 1843 1207
rect 1787 1143 1798 1177
rect 1832 1143 1843 1177
rect 1787 1097 1843 1143
rect 1873 1195 1964 1207
rect 1873 1161 1908 1195
rect 1942 1161 1964 1195
rect 1873 1097 1964 1161
rect 1994 1195 2064 1207
rect 1994 1161 2019 1195
rect 2053 1161 2064 1195
rect 1994 1097 2064 1161
rect 2094 1140 2159 1207
rect 2189 1212 2409 1250
rect 2189 1178 2200 1212
rect 2234 1178 2282 1212
rect 2316 1178 2364 1212
rect 2398 1178 2409 1212
rect 2189 1166 2409 1178
rect 2439 1166 2487 1250
rect 2517 1246 2548 1250
rect 2582 1258 2599 1280
rect 2849 1267 2907 1279
rect 2849 1258 2861 1267
rect 2582 1246 2614 1258
rect 2517 1166 2614 1246
rect 2189 1140 2239 1166
rect 2094 1097 2144 1140
rect 2564 1110 2614 1166
rect 2644 1246 2718 1258
rect 2644 1212 2664 1246
rect 2698 1212 2718 1246
rect 2644 1110 2718 1212
rect 2748 1194 2804 1258
rect 2748 1160 2759 1194
rect 2793 1160 2804 1194
rect 2748 1110 2804 1160
rect 2834 1233 2861 1258
rect 2895 1233 2907 1267
rect 2834 1110 2907 1233
rect 3170 1246 3223 1258
rect 3170 1212 3178 1246
rect 3212 1212 3223 1246
rect 3170 1156 3223 1212
rect 3170 1152 3178 1156
rect 2961 1115 3017 1152
rect 2961 1081 2972 1115
rect 3006 1081 3017 1115
rect 2961 1068 3017 1081
rect 3047 1122 3178 1152
rect 3212 1122 3223 1156
rect 3047 1110 3223 1122
rect 3253 1246 3309 1258
rect 3253 1212 3264 1246
rect 3298 1212 3309 1246
rect 3253 1156 3309 1212
rect 3253 1122 3264 1156
rect 3298 1122 3309 1156
rect 3253 1110 3309 1122
rect 3339 1246 3401 1258
rect 3339 1212 3350 1246
rect 3384 1212 3401 1246
rect 3570 1246 3641 1258
rect 3570 1238 3582 1246
rect 3339 1156 3401 1212
rect 3339 1122 3350 1156
rect 3384 1122 3401 1156
rect 3339 1110 3401 1122
rect 3464 1220 3521 1238
rect 3464 1186 3476 1220
rect 3510 1186 3521 1220
rect 3464 1152 3521 1186
rect 3464 1118 3476 1152
rect 3510 1118 3521 1152
rect 3464 1110 3521 1118
rect 3551 1212 3582 1238
rect 3616 1212 3641 1246
rect 3551 1172 3641 1212
rect 3551 1138 3582 1172
rect 3616 1138 3641 1172
rect 3551 1110 3641 1138
rect 3671 1246 3727 1258
rect 3671 1212 3682 1246
rect 3716 1212 3727 1246
rect 3671 1172 3727 1212
rect 3671 1138 3682 1172
rect 3716 1138 3727 1172
rect 3671 1110 3727 1138
rect 3757 1246 3813 1258
rect 3757 1212 3768 1246
rect 3802 1212 3813 1246
rect 3757 1156 3813 1212
rect 3757 1122 3768 1156
rect 3802 1122 3813 1156
rect 3757 1110 3813 1122
rect 3867 1250 4005 1258
rect 3867 1216 3883 1250
rect 3917 1216 3955 1250
rect 3989 1216 4005 1250
rect 3867 1110 4005 1216
rect 4059 1246 4116 1258
rect 4059 1212 4071 1246
rect 4105 1212 4116 1246
rect 4059 1156 4116 1212
rect 4059 1122 4071 1156
rect 4105 1122 4116 1156
rect 4059 1110 4116 1122
rect 4146 1224 4202 1258
rect 4146 1190 4157 1224
rect 4191 1190 4202 1224
rect 4146 1110 4202 1190
rect 4232 1246 4288 1258
rect 4232 1212 4243 1246
rect 4277 1212 4288 1246
rect 4232 1156 4288 1212
rect 4232 1122 4243 1156
rect 4277 1122 4288 1156
rect 4232 1110 4288 1122
rect 4318 1224 4374 1258
rect 4318 1190 4329 1224
rect 4363 1190 4374 1224
rect 4318 1110 4374 1190
rect 4404 1246 4468 1258
rect 4404 1212 4415 1246
rect 4449 1212 4468 1246
rect 4404 1156 4468 1212
rect 4404 1122 4415 1156
rect 4449 1122 4468 1156
rect 4404 1110 4468 1122
rect 4498 1192 4560 1258
rect 4498 1158 4515 1192
rect 4549 1158 4560 1192
rect 4498 1110 4560 1158
rect 4590 1224 4660 1258
rect 4590 1190 4615 1224
rect 4649 1190 4660 1224
rect 4590 1110 4660 1190
rect 4690 1192 4773 1258
rect 4690 1158 4719 1192
rect 4753 1158 4773 1192
rect 4690 1110 4773 1158
rect 4803 1224 4869 1258
rect 4803 1190 4823 1224
rect 4857 1190 4869 1224
rect 4803 1110 4869 1190
rect 3047 1068 3097 1110
rect -1627 210 -1556 222
rect -1627 176 -1615 210
rect -1581 176 -1556 210
rect -1627 120 -1556 176
rect -1627 86 -1615 120
rect -1581 86 -1556 120
rect -1627 74 -1556 86
rect -1526 210 -1469 222
rect -1526 176 -1515 210
rect -1481 176 -1469 210
rect -1526 120 -1469 176
rect -258 202 -201 222
rect -258 168 -246 202
rect -212 168 -201 202
rect -1526 86 -1515 120
rect -1481 86 -1469 120
rect -1526 74 -1469 86
rect -258 120 -201 168
rect -258 86 -246 120
rect -212 86 -201 120
rect -258 74 -201 86
rect -171 74 -123 222
rect -93 202 -36 222
rect -93 168 -82 202
rect -48 168 -36 202
rect -93 120 -36 168
rect -93 86 -82 120
rect -48 86 -36 120
rect -93 74 -36 86
rect 880 234 937 246
rect 224 170 281 203
rect 224 136 236 170
rect 270 136 281 170
rect 224 119 281 136
rect 311 119 359 203
rect 389 175 525 203
rect 389 141 400 175
rect 434 141 480 175
rect 514 141 525 175
rect 389 119 525 141
rect 555 119 603 203
rect 633 169 739 203
rect 633 135 644 169
rect 678 135 739 169
rect 633 119 739 135
rect 769 180 826 203
rect 769 146 780 180
rect 814 146 826 180
rect 769 119 826 146
rect 880 200 892 234
rect 926 200 937 234
rect 880 98 937 200
rect 967 98 1105 246
rect 1135 237 1192 246
rect 1135 203 1146 237
rect 1180 203 1192 237
rect 1135 169 1192 203
rect 1135 135 1146 169
rect 1180 135 1192 169
rect 1135 98 1192 135
rect 1270 125 1347 209
rect 1377 125 1419 209
rect 1449 184 1510 209
rect 1449 150 1465 184
rect 1499 150 1510 184
rect 1449 125 1510 150
rect 1540 179 1611 209
rect 1540 145 1565 179
rect 1599 145 1611 179
rect 1540 125 1611 145
rect 1665 125 1757 235
rect 1787 189 1843 235
rect 1787 155 1798 189
rect 1832 155 1843 189
rect 1787 125 1843 155
rect 1873 171 1964 235
rect 1873 137 1908 171
rect 1942 137 1964 171
rect 1873 125 1964 137
rect 1994 171 2064 235
rect 1994 137 2019 171
rect 2053 137 2064 171
rect 1994 125 2064 137
rect 2094 192 2144 235
rect 2094 125 2159 192
rect 1270 118 1332 125
rect 982 82 1040 98
rect 982 48 994 82
rect 1028 48 1040 82
rect 982 36 1040 48
rect 1270 84 1284 118
rect 1318 84 1332 118
rect 1270 72 1332 84
rect 1665 119 1742 125
rect 1665 85 1686 119
rect 1720 85 1742 119
rect 1665 73 1742 85
rect 2109 82 2159 125
rect 2189 166 2239 192
rect 2961 251 3017 264
rect 2564 166 2614 222
rect 2189 154 2409 166
rect 2189 120 2200 154
rect 2234 120 2282 154
rect 2316 120 2364 154
rect 2398 120 2409 154
rect 2189 82 2409 120
rect 2439 82 2487 166
rect 2517 86 2614 166
rect 2517 82 2548 86
rect 2532 52 2548 82
rect 2582 74 2614 86
rect 2644 120 2718 222
rect 2644 86 2664 120
rect 2698 86 2718 120
rect 2644 74 2718 86
rect 2748 172 2804 222
rect 2748 138 2759 172
rect 2793 138 2804 172
rect 2748 74 2804 138
rect 2834 99 2907 222
rect 2961 217 2972 251
rect 3006 217 3017 251
rect 2961 180 3017 217
rect 3047 222 3097 264
rect 4059 235 4116 247
rect 3047 210 3223 222
rect 3047 180 3178 210
rect 3170 176 3178 180
rect 3212 176 3223 210
rect 2834 74 2861 99
rect 2582 52 2599 74
rect 2532 40 2599 52
rect 2849 65 2861 74
rect 2895 65 2907 99
rect 3170 120 3223 176
rect 3170 86 3178 120
rect 3212 86 3223 120
rect 3170 74 3223 86
rect 3253 210 3309 222
rect 3253 176 3264 210
rect 3298 176 3309 210
rect 3253 120 3309 176
rect 3253 86 3264 120
rect 3298 86 3309 120
rect 3253 74 3309 86
rect 3339 210 3401 222
rect 3339 176 3350 210
rect 3384 176 3401 210
rect 3339 120 3401 176
rect 3339 86 3350 120
rect 3384 86 3401 120
rect 3464 214 3521 222
rect 3464 180 3476 214
rect 3510 180 3521 214
rect 3464 146 3521 180
rect 3464 112 3476 146
rect 3510 112 3521 146
rect 3464 94 3521 112
rect 3551 194 3641 222
rect 3551 160 3582 194
rect 3616 160 3641 194
rect 3551 120 3641 160
rect 3551 94 3582 120
rect 3339 74 3401 86
rect 2849 53 2907 65
rect 3570 86 3582 94
rect 3616 86 3641 120
rect 3570 74 3641 86
rect 3671 194 3727 222
rect 3671 160 3682 194
rect 3716 160 3727 194
rect 3671 120 3727 160
rect 3671 86 3682 120
rect 3716 86 3727 120
rect 3671 74 3727 86
rect 3757 210 3813 222
rect 3757 176 3768 210
rect 3802 176 3813 210
rect 3757 120 3813 176
rect 3757 86 3768 120
rect 3802 86 3813 120
rect 3757 74 3813 86
rect 3867 116 4005 222
rect 4059 201 4071 235
rect 4105 201 4116 235
rect 4059 165 4116 201
rect 4059 131 4071 165
rect 4105 131 4116 165
rect 4059 119 4116 131
rect 4146 168 4206 247
rect 4146 134 4161 168
rect 4195 134 4206 168
rect 4146 119 4206 134
rect 4236 239 4301 247
rect 4236 205 4247 239
rect 4281 205 4301 239
rect 4236 161 4301 205
rect 4236 127 4247 161
rect 4281 127 4301 161
rect 4236 119 4301 127
rect 4331 229 4392 247
rect 4331 195 4347 229
rect 4381 195 4392 229
rect 4331 161 4392 195
rect 4331 127 4347 161
rect 4381 127 4392 161
rect 4331 119 4392 127
rect 4422 235 4494 247
rect 4422 201 4449 235
rect 4483 201 4494 235
rect 4422 157 4494 201
rect 4422 123 4449 157
rect 4483 123 4494 157
rect 4422 119 4494 123
rect 3867 82 3883 116
rect 3917 82 3955 116
rect 3989 82 4005 116
rect 3867 74 4005 82
rect 4437 99 4494 119
rect 4524 219 4610 247
rect 4524 185 4551 219
rect 4585 185 4610 219
rect 4524 145 4610 185
rect 4524 111 4551 145
rect 4585 111 4610 145
rect 4524 99 4610 111
rect 4640 151 4696 247
rect 4640 117 4651 151
rect 4685 117 4696 151
rect 4640 99 4696 117
rect 4726 235 4782 247
rect 4726 201 4737 235
rect 4771 201 4782 235
rect 4726 145 4782 201
rect 4726 111 4737 145
rect 4771 111 4782 145
rect 4726 99 4782 111
rect 4812 235 4869 247
rect 4812 201 4823 235
rect 4857 201 4869 235
rect 4812 145 4869 201
rect 4812 111 4823 145
rect 4857 111 4869 145
rect 4812 99 4869 111
rect -1401 -310 -1343 -298
rect -1401 -686 -1389 -310
rect -1355 -686 -1343 -310
rect -1401 -698 -1343 -686
rect -1313 -310 -1255 -298
rect -1313 -686 -1301 -310
rect -1267 -686 -1255 -310
rect -1313 -698 -1255 -686
rect -1401 -1024 -1343 -1012
rect -1401 -1400 -1389 -1024
rect -1355 -1400 -1343 -1024
rect -1401 -1412 -1343 -1400
rect -1313 -1024 -1255 -1012
rect -1313 -1400 -1301 -1024
rect -1267 -1400 -1255 -1024
rect -1313 -1412 -1255 -1400
<< pdiff >>
rect -2779 1912 -2710 1924
rect -2779 1878 -2767 1912
rect -2733 1878 -2710 1912
rect -2779 1842 -2710 1878
rect -2779 1808 -2767 1842
rect -2733 1808 -2710 1842
rect -2779 1772 -2710 1808
rect -2779 1738 -2767 1772
rect -2733 1738 -2710 1772
rect -2779 1700 -2710 1738
rect -2680 1912 -2621 1924
rect -2680 1878 -2667 1912
rect -2633 1878 -2621 1912
rect -2680 1829 -2621 1878
rect -2680 1795 -2667 1829
rect -2633 1795 -2621 1829
rect -2680 1746 -2621 1795
rect -1413 1912 -1356 1924
rect -1413 1878 -1403 1912
rect -1369 1878 -1356 1912
rect -1413 1829 -1356 1878
rect -1413 1795 -1403 1829
rect -1369 1795 -1356 1829
rect -2680 1712 -2667 1746
rect -2633 1712 -2621 1746
rect -2680 1700 -2621 1712
rect -1413 1746 -1356 1795
rect -1413 1712 -1403 1746
rect -1369 1712 -1356 1746
rect -1413 1700 -1356 1712
rect -1326 1912 -1266 1924
rect -1326 1878 -1313 1912
rect -1279 1878 -1266 1912
rect -1326 1829 -1266 1878
rect -1326 1795 -1313 1829
rect -1279 1795 -1266 1829
rect -1326 1746 -1266 1795
rect -1326 1712 -1313 1746
rect -1279 1712 -1266 1746
rect -1326 1700 -1266 1712
rect -1236 1912 -1179 1924
rect -1236 1878 -1223 1912
rect -1189 1878 -1179 1912
rect -1236 1829 -1179 1878
rect -1236 1795 -1223 1829
rect -1189 1795 -1179 1829
rect -1236 1746 -1179 1795
rect -1236 1712 -1223 1746
rect -1189 1712 -1179 1746
rect -1125 1912 -1070 1924
rect -1125 1878 -1117 1912
rect -1083 1878 -1070 1912
rect -1125 1841 -1070 1878
rect -1125 1807 -1117 1841
rect -1083 1807 -1070 1841
rect -1125 1770 -1070 1807
rect -1125 1736 -1117 1770
rect -1083 1736 -1070 1770
rect -1125 1724 -1070 1736
rect -870 1912 -815 1924
rect -870 1878 -859 1912
rect -825 1878 -815 1912
rect -870 1841 -815 1878
rect -870 1807 -859 1841
rect -825 1807 -815 1841
rect -870 1770 -815 1807
rect -870 1736 -859 1770
rect -825 1736 -815 1770
rect -870 1724 -815 1736
rect -615 1912 -558 1924
rect -615 1878 -604 1912
rect -570 1878 -558 1912
rect -615 1841 -558 1878
rect -615 1807 -604 1841
rect -570 1807 -558 1841
rect -615 1770 -558 1807
rect -615 1736 -604 1770
rect -570 1736 -558 1770
rect 219 1912 274 1924
rect 219 1878 227 1912
rect 261 1878 274 1912
rect 219 1841 274 1878
rect 219 1807 227 1841
rect 261 1807 274 1841
rect 219 1770 274 1807
rect -615 1724 -558 1736
rect 219 1736 227 1770
rect 261 1736 274 1770
rect 219 1724 274 1736
rect 474 1912 529 1924
rect 474 1878 485 1912
rect 519 1878 529 1912
rect 474 1841 529 1878
rect 474 1807 485 1841
rect 519 1807 529 1841
rect 474 1770 529 1807
rect 474 1736 485 1770
rect 519 1736 529 1770
rect 474 1724 529 1736
rect 729 1912 786 1924
rect 729 1878 740 1912
rect 774 1878 786 1912
rect 729 1841 786 1878
rect 729 1807 740 1841
rect 774 1807 786 1841
rect 729 1770 786 1807
rect 729 1736 740 1770
rect 774 1736 786 1770
rect 729 1724 786 1736
rect 891 1912 946 1924
rect 891 1878 899 1912
rect 933 1878 946 1912
rect 891 1841 946 1878
rect 891 1807 899 1841
rect 933 1807 946 1841
rect 891 1770 946 1807
rect 891 1736 899 1770
rect 933 1736 946 1770
rect 891 1724 946 1736
rect 1146 1912 1201 1924
rect 1146 1878 1157 1912
rect 1191 1878 1201 1912
rect 1146 1841 1201 1878
rect 1146 1807 1157 1841
rect 1191 1807 1201 1841
rect 1146 1770 1201 1807
rect 1146 1736 1157 1770
rect 1191 1736 1201 1770
rect 1146 1724 1201 1736
rect 1401 1912 1458 1924
rect 1401 1878 1412 1912
rect 1446 1878 1458 1912
rect 1401 1841 1458 1878
rect 1401 1807 1412 1841
rect 1446 1807 1458 1841
rect 1401 1770 1458 1807
rect 1401 1736 1412 1770
rect 1446 1736 1458 1770
rect 1401 1724 1458 1736
rect 1563 1912 1618 1924
rect 1563 1878 1571 1912
rect 1605 1878 1618 1912
rect 1563 1841 1618 1878
rect 1563 1807 1571 1841
rect 1605 1807 1618 1841
rect 1563 1770 1618 1807
rect 1563 1736 1571 1770
rect 1605 1736 1618 1770
rect 1563 1724 1618 1736
rect 1818 1912 1873 1924
rect 1818 1878 1829 1912
rect 1863 1878 1873 1912
rect 1818 1841 1873 1878
rect 1818 1807 1829 1841
rect 1863 1807 1873 1841
rect 1818 1770 1873 1807
rect 1818 1736 1829 1770
rect 1863 1736 1873 1770
rect 1818 1724 1873 1736
rect 2073 1912 2130 1924
rect 2073 1878 2084 1912
rect 2118 1878 2130 1912
rect 2073 1841 2130 1878
rect 2073 1807 2084 1841
rect 2118 1807 2130 1841
rect 2073 1770 2130 1807
rect 2073 1736 2084 1770
rect 2118 1736 2130 1770
rect 2073 1724 2130 1736
rect 2235 1912 2290 1924
rect 2235 1878 2243 1912
rect 2277 1878 2290 1912
rect 2235 1841 2290 1878
rect 2235 1807 2243 1841
rect 2277 1807 2290 1841
rect 2235 1770 2290 1807
rect 2235 1736 2243 1770
rect 2277 1736 2290 1770
rect 2235 1724 2290 1736
rect 2490 1912 2545 1924
rect 2490 1878 2501 1912
rect 2535 1878 2545 1912
rect 2490 1841 2545 1878
rect 2490 1807 2501 1841
rect 2535 1807 2545 1841
rect 2490 1770 2545 1807
rect 2490 1736 2501 1770
rect 2535 1736 2545 1770
rect 2490 1724 2545 1736
rect 2745 1912 2802 1924
rect 2745 1878 2756 1912
rect 2790 1878 2802 1912
rect 2745 1841 2802 1878
rect 2745 1807 2756 1841
rect 2790 1807 2802 1841
rect 2745 1770 2802 1807
rect 2745 1736 2756 1770
rect 2790 1736 2802 1770
rect 2745 1724 2802 1736
rect 2907 1912 2962 1924
rect 2907 1878 2915 1912
rect 2949 1878 2962 1912
rect 2907 1841 2962 1878
rect 2907 1807 2915 1841
rect 2949 1807 2962 1841
rect 2907 1770 2962 1807
rect 2907 1736 2915 1770
rect 2949 1736 2962 1770
rect 2907 1724 2962 1736
rect 3162 1912 3217 1924
rect 3162 1878 3173 1912
rect 3207 1878 3217 1912
rect 3162 1841 3217 1878
rect 3162 1807 3173 1841
rect 3207 1807 3217 1841
rect 3162 1770 3217 1807
rect 3162 1736 3173 1770
rect 3207 1736 3217 1770
rect 3162 1724 3217 1736
rect 3417 1912 3474 1924
rect 3417 1878 3428 1912
rect 3462 1878 3474 1912
rect 3417 1841 3474 1878
rect 3417 1807 3428 1841
rect 3462 1807 3474 1841
rect 3417 1770 3474 1807
rect 3417 1736 3428 1770
rect 3462 1736 3474 1770
rect 3417 1724 3474 1736
rect 3579 1912 3634 1924
rect 3579 1878 3587 1912
rect 3621 1878 3634 1912
rect 3579 1841 3634 1878
rect 3579 1807 3587 1841
rect 3621 1807 3634 1841
rect 3579 1770 3634 1807
rect 3579 1736 3587 1770
rect 3621 1736 3634 1770
rect 3579 1724 3634 1736
rect 3834 1912 3889 1924
rect 3834 1878 3845 1912
rect 3879 1878 3889 1912
rect 3834 1841 3889 1878
rect 3834 1807 3845 1841
rect 3879 1807 3889 1841
rect 3834 1770 3889 1807
rect 3834 1736 3845 1770
rect 3879 1736 3889 1770
rect 3834 1724 3889 1736
rect 4089 1912 4146 1924
rect 4089 1878 4100 1912
rect 4134 1878 4146 1912
rect 4089 1841 4146 1878
rect 4089 1807 4100 1841
rect 4134 1807 4146 1841
rect 4089 1770 4146 1807
rect 4089 1736 4100 1770
rect 4134 1736 4146 1770
rect 4089 1724 4146 1736
rect 4251 1912 4306 1924
rect 4251 1878 4259 1912
rect 4293 1878 4306 1912
rect 4251 1841 4306 1878
rect 4251 1807 4259 1841
rect 4293 1807 4306 1841
rect 4251 1770 4306 1807
rect 4251 1736 4259 1770
rect 4293 1736 4306 1770
rect 4251 1724 4306 1736
rect 4506 1912 4563 1924
rect 4506 1878 4517 1912
rect 4551 1878 4563 1912
rect 4506 1841 4563 1878
rect 4506 1807 4517 1841
rect 4551 1807 4563 1841
rect 4506 1770 4563 1807
rect 4506 1736 4517 1770
rect 4551 1736 4563 1770
rect 4506 1724 4563 1736
rect -1236 1700 -1179 1712
rect -2779 926 -2710 964
rect -2779 892 -2767 926
rect -2733 892 -2710 926
rect -2779 856 -2710 892
rect -2779 822 -2767 856
rect -2733 822 -2710 856
rect -2779 786 -2710 822
rect -2779 752 -2767 786
rect -2733 752 -2710 786
rect -2779 740 -2710 752
rect -2680 952 -2621 964
rect -2680 918 -2667 952
rect -2633 918 -2621 952
rect -2680 869 -2621 918
rect -1413 952 -1356 964
rect -1413 918 -1403 952
rect -1369 918 -1356 952
rect -2680 835 -2667 869
rect -2633 835 -2621 869
rect -2680 786 -2621 835
rect -2680 752 -2667 786
rect -2633 752 -2621 786
rect -2680 740 -2621 752
rect -1413 869 -1356 918
rect -1413 835 -1403 869
rect -1369 835 -1356 869
rect -1413 786 -1356 835
rect -1413 752 -1403 786
rect -1369 752 -1356 786
rect -1413 740 -1356 752
rect -1326 952 -1266 964
rect -1326 918 -1313 952
rect -1279 918 -1266 952
rect -1326 869 -1266 918
rect -1326 835 -1313 869
rect -1279 835 -1266 869
rect -1326 786 -1266 835
rect -1326 752 -1313 786
rect -1279 752 -1266 786
rect -1326 740 -1266 752
rect -1236 952 -1179 964
rect -1236 918 -1223 952
rect -1189 918 -1179 952
rect -1236 869 -1179 918
rect -1236 835 -1223 869
rect -1189 835 -1179 869
rect -1236 786 -1179 835
rect -1125 937 -1066 964
rect -1125 903 -1113 937
rect -1079 903 -1066 937
rect -1125 842 -1066 903
rect -1125 808 -1113 842
rect -1079 808 -1066 842
rect -1125 796 -1066 808
rect -1036 847 -959 964
rect -1036 813 -1006 847
rect -972 813 -959 847
rect -1036 796 -959 813
rect -1236 752 -1223 786
rect -1189 752 -1179 786
rect -1018 764 -959 796
rect -929 764 -766 964
rect -736 952 -658 964
rect -736 918 -723 952
rect -689 918 -658 952
rect -736 835 -658 918
rect -736 801 -723 835
rect -689 801 -658 835
rect -736 764 -658 801
rect -628 764 -544 964
rect -514 952 -420 964
rect -514 918 -477 952
rect -443 918 -420 952
rect -514 869 -420 918
rect -514 835 -477 869
rect -443 835 -420 869
rect -514 786 -420 835
rect -514 764 -477 786
rect -1236 740 -1179 752
rect -489 752 -477 764
rect -443 752 -420 786
rect -489 740 -420 752
rect -390 952 -331 964
rect -390 918 -377 952
rect -343 918 -331 952
rect -390 869 -331 918
rect -390 835 -377 869
rect -343 835 -331 869
rect -390 786 -331 835
rect -390 752 -377 786
rect -343 752 -331 786
rect -390 740 -331 752
rect -261 926 -204 964
rect -261 892 -251 926
rect -217 892 -204 926
rect -261 856 -204 892
rect -261 822 -251 856
rect -217 822 -204 856
rect -261 786 -204 822
rect -261 752 -251 786
rect -217 752 -204 786
rect -261 740 -204 752
rect -174 952 -114 964
rect -174 918 -161 952
rect -127 918 -114 952
rect -174 869 -114 918
rect -174 835 -161 869
rect -127 835 -114 869
rect -174 786 -114 835
rect -174 752 -161 786
rect -127 752 -114 786
rect -174 740 -114 752
rect -84 952 -27 964
rect -84 918 -71 952
rect -37 918 -27 952
rect -84 869 -27 918
rect -84 835 -71 869
rect -37 835 -27 869
rect -84 786 -27 835
rect -84 752 -71 786
rect -37 752 -27 786
rect -84 740 -27 752
rect 881 926 940 964
rect 881 892 893 926
rect 927 892 940 926
rect 219 855 278 868
rect 219 821 231 855
rect 265 821 278 855
rect 219 786 278 821
rect 219 752 231 786
rect 265 752 278 786
rect 219 740 278 752
rect 308 787 368 868
rect 308 753 321 787
rect 355 753 368 787
rect 308 740 368 753
rect 398 740 446 868
rect 476 846 536 868
rect 476 812 489 846
rect 523 812 536 846
rect 476 740 536 812
rect 566 856 625 868
rect 566 822 579 856
rect 613 822 625 856
rect 566 786 625 822
rect 566 752 579 786
rect 613 752 625 786
rect 566 740 625 752
rect 679 856 738 868
rect 679 822 691 856
rect 725 822 738 856
rect 679 786 738 822
rect 679 752 691 786
rect 725 752 738 786
rect 679 740 738 752
rect 768 856 827 868
rect 768 822 781 856
rect 815 822 827 856
rect 768 786 827 822
rect 768 752 781 786
rect 815 752 827 786
rect 768 740 827 752
rect 881 856 940 892
rect 881 822 893 856
rect 927 822 940 856
rect 881 786 940 822
rect 881 752 893 786
rect 927 752 940 786
rect 881 740 940 752
rect 970 864 1030 964
rect 970 830 983 864
rect 1017 830 1030 864
rect 970 786 1030 830
rect 970 752 983 786
rect 1017 752 1030 786
rect 970 740 1030 752
rect 1060 948 1119 964
rect 1060 914 1073 948
rect 1107 914 1119 948
rect 1060 867 1119 914
rect 1060 833 1073 867
rect 1107 833 1119 867
rect 1060 786 1119 833
rect 1060 752 1073 786
rect 1107 752 1119 786
rect 1173 838 1232 868
rect 1173 804 1185 838
rect 1219 804 1232 838
rect 1173 784 1232 804
rect 1262 784 1316 868
rect 1346 846 1423 868
rect 1346 812 1376 846
rect 1410 812 1423 846
rect 1346 784 1423 812
rect 1060 740 1119 752
rect 1364 740 1423 784
rect 1453 846 1522 868
rect 1453 812 1476 846
rect 1510 812 1522 846
rect 1453 740 1522 812
rect 1576 786 1754 908
rect 1576 752 1588 786
rect 1622 752 1707 786
rect 1741 752 1754 786
rect 1576 740 1754 752
rect 1784 740 1838 908
rect 1868 823 1946 908
rect 1868 789 1881 823
rect 1915 789 1946 823
rect 1868 740 1946 789
rect 1976 896 2035 908
rect 1976 862 1989 896
rect 2023 862 2035 896
rect 1976 786 2035 862
rect 1976 752 1989 786
rect 2023 752 2035 786
rect 1976 740 2035 752
rect 2089 858 2148 908
rect 2089 824 2101 858
rect 2135 824 2148 858
rect 2089 786 2148 824
rect 2089 752 2101 786
rect 2135 752 2148 786
rect 2089 740 2148 752
rect 2178 740 2226 908
rect 2256 896 2315 908
rect 2256 862 2269 896
rect 2303 862 2315 896
rect 2256 824 2315 862
rect 2557 864 2616 940
rect 2557 830 2569 864
rect 2603 830 2616 864
rect 2256 786 2333 824
rect 2256 752 2269 786
rect 2303 752 2333 786
rect 2256 740 2333 752
rect 2363 740 2411 824
rect 2441 791 2500 824
rect 2441 757 2454 791
rect 2488 757 2500 791
rect 2441 740 2500 757
rect 2557 786 2616 830
rect 2557 752 2569 786
rect 2603 752 2616 786
rect 2557 740 2616 752
rect 2646 791 2718 940
rect 2646 757 2669 791
rect 2703 757 2718 791
rect 2646 740 2718 757
rect 2748 740 2802 940
rect 2832 904 2891 940
rect 3187 933 3240 964
rect 2832 870 2845 904
rect 2879 870 2891 904
rect 2832 786 2891 870
rect 2945 915 3004 933
rect 2945 881 2957 915
rect 2991 881 3004 915
rect 2945 805 3004 881
rect 3034 919 3240 933
rect 3034 885 3176 919
rect 3210 885 3240 919
rect 3034 837 3240 885
rect 3034 805 3176 837
rect 2832 752 2845 786
rect 2879 752 2891 786
rect 3052 803 3176 805
rect 3210 803 3240 837
rect 2832 740 2891 752
rect 3052 747 3240 803
rect 3052 713 3064 747
rect 3098 713 3176 747
rect 3210 740 3240 747
rect 3270 952 3330 964
rect 3270 918 3283 952
rect 3317 918 3330 952
rect 3270 869 3330 918
rect 3270 835 3283 869
rect 3317 835 3330 869
rect 3270 786 3330 835
rect 3270 752 3283 786
rect 3317 752 3330 786
rect 3270 740 3330 752
rect 3360 926 3417 964
rect 3581 948 3634 964
rect 3360 892 3373 926
rect 3407 892 3417 926
rect 3360 856 3417 892
rect 3360 822 3373 856
rect 3407 822 3417 856
rect 3360 786 3417 822
rect 3360 752 3373 786
rect 3407 752 3417 786
rect 3360 740 3417 752
rect 3471 936 3529 948
rect 3471 902 3482 936
rect 3516 902 3529 936
rect 3471 865 3529 902
rect 3471 831 3482 865
rect 3516 831 3529 865
rect 3471 794 3529 831
rect 3471 760 3482 794
rect 3516 760 3529 794
rect 3471 748 3529 760
rect 3559 940 3634 948
rect 3559 906 3587 940
rect 3621 906 3634 940
rect 3559 868 3634 906
rect 3559 834 3587 868
rect 3621 834 3634 868
rect 3559 790 3634 834
rect 3559 756 3587 790
rect 3621 756 3634 790
rect 3559 748 3634 756
rect 3210 713 3222 740
rect 3577 740 3634 748
rect 3664 952 3724 964
rect 3664 918 3677 952
rect 3711 918 3724 952
rect 3664 869 3724 918
rect 3664 835 3677 869
rect 3711 835 3724 869
rect 3664 786 3724 835
rect 3664 752 3677 786
rect 3711 752 3724 786
rect 3664 740 3724 752
rect 3754 952 3813 964
rect 3754 918 3767 952
rect 3801 918 3813 952
rect 3754 869 3813 918
rect 3754 835 3767 869
rect 3801 835 3813 869
rect 3754 786 3813 835
rect 3754 752 3767 786
rect 3801 752 3813 786
rect 3754 740 3813 752
rect 3867 782 4005 964
rect 3867 748 3883 782
rect 3917 748 3955 782
rect 3989 748 4005 782
rect 3867 740 4005 748
rect 4059 946 4119 964
rect 4059 912 4071 946
rect 4105 912 4119 946
rect 4059 866 4119 912
rect 4059 832 4071 866
rect 4105 832 4119 866
rect 4059 786 4119 832
rect 4059 752 4071 786
rect 4105 752 4119 786
rect 4059 740 4119 752
rect 4149 926 4371 964
rect 4149 892 4162 926
rect 4196 892 4242 926
rect 4276 892 4324 926
rect 4358 892 4371 926
rect 4149 855 4371 892
rect 4149 821 4162 855
rect 4196 821 4242 855
rect 4276 821 4324 855
rect 4358 821 4371 855
rect 4149 786 4371 821
rect 4149 752 4162 786
rect 4196 752 4242 786
rect 4276 752 4324 786
rect 4358 752 4371 786
rect 4149 740 4371 752
rect 4401 865 4471 964
rect 4401 831 4414 865
rect 4448 831 4471 865
rect 4401 786 4471 831
rect 4401 752 4414 786
rect 4448 752 4471 786
rect 4401 740 4471 752
rect 4501 926 4770 964
rect 4501 892 4514 926
rect 4548 892 4583 926
rect 4617 892 4654 926
rect 4688 892 4723 926
rect 4757 892 4770 926
rect 4501 855 4770 892
rect 4501 821 4514 855
rect 4548 821 4583 855
rect 4617 821 4654 855
rect 4688 821 4723 855
rect 4757 821 4770 855
rect 4501 786 4770 821
rect 4501 752 4514 786
rect 4548 752 4583 786
rect 4617 752 4654 786
rect 4688 752 4723 786
rect 4757 752 4770 786
rect 4501 740 4770 752
rect 4800 865 4869 964
rect 4800 831 4823 865
rect 4857 831 4869 865
rect 4800 786 4869 831
rect 4800 752 4823 786
rect 4857 752 4869 786
rect 4800 740 4869 752
rect 3052 701 3222 713
rect 3052 619 3222 631
rect -1627 580 -1558 592
rect -1627 546 -1615 580
rect -1581 546 -1558 580
rect -1627 510 -1558 546
rect -1627 476 -1615 510
rect -1581 476 -1558 510
rect -1627 440 -1558 476
rect -1627 406 -1615 440
rect -1581 406 -1558 440
rect -1627 368 -1558 406
rect -1528 580 -1469 592
rect -1528 546 -1515 580
rect -1481 546 -1469 580
rect -1528 497 -1469 546
rect -1528 463 -1515 497
rect -1481 463 -1469 497
rect -1528 414 -1469 463
rect -261 580 -204 592
rect -261 546 -251 580
rect -217 546 -204 580
rect -261 497 -204 546
rect -261 463 -251 497
rect -217 463 -204 497
rect -1528 380 -1515 414
rect -1481 380 -1469 414
rect -1528 368 -1469 380
rect -261 414 -204 463
rect -261 380 -251 414
rect -217 380 -204 414
rect -261 368 -204 380
rect -174 580 -114 592
rect -174 546 -161 580
rect -127 546 -114 580
rect -174 497 -114 546
rect -174 463 -161 497
rect -127 463 -114 497
rect -174 414 -114 463
rect -174 380 -161 414
rect -127 380 -114 414
rect -174 368 -114 380
rect -84 580 -27 592
rect -84 546 -71 580
rect -37 546 -27 580
rect -84 497 -27 546
rect -84 463 -71 497
rect -37 463 -27 497
rect -84 414 -27 463
rect 219 580 278 592
rect 219 546 231 580
rect 265 546 278 580
rect 219 511 278 546
rect 219 477 231 511
rect 265 477 278 511
rect 219 464 278 477
rect 308 579 368 592
rect 308 545 321 579
rect 355 545 368 579
rect 308 464 368 545
rect 398 464 446 592
rect 476 520 536 592
rect 476 486 489 520
rect 523 486 536 520
rect 476 464 536 486
rect 566 580 625 592
rect 566 546 579 580
rect 613 546 625 580
rect 566 510 625 546
rect 566 476 579 510
rect 613 476 625 510
rect 566 464 625 476
rect 679 580 738 592
rect 679 546 691 580
rect 725 546 738 580
rect 679 510 738 546
rect 679 476 691 510
rect 725 476 738 510
rect 679 464 738 476
rect 768 580 827 592
rect 768 546 781 580
rect 815 546 827 580
rect 768 510 827 546
rect 768 476 781 510
rect 815 476 827 510
rect 768 464 827 476
rect 881 580 940 592
rect 881 546 893 580
rect 927 546 940 580
rect 881 510 940 546
rect 881 476 893 510
rect 927 476 940 510
rect -84 380 -71 414
rect -37 380 -27 414
rect -84 368 -27 380
rect 881 440 940 476
rect 881 406 893 440
rect 927 406 940 440
rect 881 368 940 406
rect 970 580 1030 592
rect 970 546 983 580
rect 1017 546 1030 580
rect 970 502 1030 546
rect 970 468 983 502
rect 1017 468 1030 502
rect 970 368 1030 468
rect 1060 580 1119 592
rect 1060 546 1073 580
rect 1107 546 1119 580
rect 1364 548 1423 592
rect 1060 499 1119 546
rect 1060 465 1073 499
rect 1107 465 1119 499
rect 1060 418 1119 465
rect 1173 528 1232 548
rect 1173 494 1185 528
rect 1219 494 1232 528
rect 1173 464 1232 494
rect 1262 464 1316 548
rect 1346 520 1423 548
rect 1346 486 1376 520
rect 1410 486 1423 520
rect 1346 464 1423 486
rect 1453 520 1522 592
rect 1453 486 1476 520
rect 1510 486 1522 520
rect 1453 464 1522 486
rect 1576 580 1754 592
rect 1576 546 1588 580
rect 1622 546 1707 580
rect 1741 546 1754 580
rect 1060 384 1073 418
rect 1107 384 1119 418
rect 1060 368 1119 384
rect 1576 424 1754 546
rect 1784 424 1838 592
rect 1868 543 1946 592
rect 1868 509 1881 543
rect 1915 509 1946 543
rect 1868 424 1946 509
rect 1976 580 2035 592
rect 1976 546 1989 580
rect 2023 546 2035 580
rect 1976 470 2035 546
rect 1976 436 1989 470
rect 2023 436 2035 470
rect 1976 424 2035 436
rect 2089 580 2148 592
rect 2089 546 2101 580
rect 2135 546 2148 580
rect 2089 508 2148 546
rect 2089 474 2101 508
rect 2135 474 2148 508
rect 2089 424 2148 474
rect 2178 424 2226 592
rect 2256 580 2333 592
rect 2256 546 2269 580
rect 2303 546 2333 580
rect 2256 508 2333 546
rect 2363 508 2411 592
rect 2441 575 2500 592
rect 2441 541 2454 575
rect 2488 541 2500 575
rect 2441 508 2500 541
rect 2557 580 2616 592
rect 2557 546 2569 580
rect 2603 546 2616 580
rect 2256 470 2315 508
rect 2557 502 2616 546
rect 2256 436 2269 470
rect 2303 436 2315 470
rect 2256 424 2315 436
rect 2557 468 2569 502
rect 2603 468 2616 502
rect 2557 392 2616 468
rect 2646 575 2718 592
rect 2646 541 2669 575
rect 2703 541 2718 575
rect 2646 392 2718 541
rect 2748 392 2802 592
rect 2832 580 2891 592
rect 2832 546 2845 580
rect 2879 546 2891 580
rect 3052 585 3064 619
rect 3098 585 3176 619
rect 3210 592 3222 619
rect 3210 585 3240 592
rect 2832 462 2891 546
rect 3052 529 3240 585
rect 3052 527 3176 529
rect 2832 428 2845 462
rect 2879 428 2891 462
rect 2832 392 2891 428
rect 2945 451 3004 527
rect 2945 417 2957 451
rect 2991 417 3004 451
rect 2945 399 3004 417
rect 3034 495 3176 527
rect 3210 495 3240 529
rect 3034 447 3240 495
rect 3034 413 3176 447
rect 3210 413 3240 447
rect 3034 399 3240 413
rect 3187 368 3240 399
rect 3270 580 3330 592
rect 3270 546 3283 580
rect 3317 546 3330 580
rect 3270 497 3330 546
rect 3270 463 3283 497
rect 3317 463 3330 497
rect 3270 414 3330 463
rect 3270 380 3283 414
rect 3317 380 3330 414
rect 3270 368 3330 380
rect 3360 580 3417 592
rect 3577 584 3634 592
rect 3360 546 3373 580
rect 3407 546 3417 580
rect 3360 510 3417 546
rect 3360 476 3373 510
rect 3407 476 3417 510
rect 3360 440 3417 476
rect 3360 406 3373 440
rect 3407 406 3417 440
rect 3360 368 3417 406
rect 3471 572 3529 584
rect 3471 538 3482 572
rect 3516 538 3529 572
rect 3471 501 3529 538
rect 3471 467 3482 501
rect 3516 467 3529 501
rect 3471 430 3529 467
rect 3471 396 3482 430
rect 3516 396 3529 430
rect 3471 384 3529 396
rect 3559 576 3634 584
rect 3559 542 3587 576
rect 3621 542 3634 576
rect 3559 498 3634 542
rect 3559 464 3587 498
rect 3621 464 3634 498
rect 3559 426 3634 464
rect 3559 392 3587 426
rect 3621 392 3634 426
rect 3559 384 3634 392
rect 3581 368 3634 384
rect 3664 580 3724 592
rect 3664 546 3677 580
rect 3711 546 3724 580
rect 3664 497 3724 546
rect 3664 463 3677 497
rect 3711 463 3724 497
rect 3664 414 3724 463
rect 3664 380 3677 414
rect 3711 380 3724 414
rect 3664 368 3724 380
rect 3754 580 3813 592
rect 3754 546 3767 580
rect 3801 546 3813 580
rect 3754 497 3813 546
rect 3754 463 3767 497
rect 3801 463 3813 497
rect 3754 414 3813 463
rect 3754 380 3767 414
rect 3801 380 3813 414
rect 3754 368 3813 380
rect 3867 584 4005 592
rect 3867 550 3883 584
rect 3917 550 3955 584
rect 3989 550 4005 584
rect 4447 580 4506 592
rect 4447 577 4459 580
rect 3867 368 4005 550
rect 4060 565 4119 577
rect 4060 531 4072 565
rect 4106 531 4119 565
rect 4060 455 4119 531
rect 4060 421 4072 455
rect 4106 421 4119 455
rect 4060 409 4119 421
rect 4149 565 4209 577
rect 4149 531 4162 565
rect 4196 531 4209 565
rect 4149 455 4209 531
rect 4149 421 4162 455
rect 4196 421 4209 455
rect 4149 409 4209 421
rect 4239 568 4304 577
rect 4239 534 4252 568
rect 4286 534 4304 568
rect 4239 500 4304 534
rect 4239 466 4252 500
rect 4286 466 4304 500
rect 4239 409 4304 466
rect 4334 565 4399 577
rect 4334 531 4352 565
rect 4386 531 4399 565
rect 4334 455 4399 531
rect 4334 421 4352 455
rect 4386 421 4399 455
rect 4334 409 4399 421
rect 4429 546 4459 577
rect 4493 546 4506 580
rect 4429 508 4506 546
rect 4429 474 4459 508
rect 4493 474 4506 508
rect 4429 409 4506 474
rect 4453 368 4506 409
rect 4536 580 4600 592
rect 4536 546 4553 580
rect 4587 546 4600 580
rect 4536 499 4600 546
rect 4536 465 4553 499
rect 4587 465 4600 499
rect 4536 419 4600 465
rect 4536 385 4553 419
rect 4587 385 4600 419
rect 4536 368 4600 385
rect 4630 580 4690 592
rect 4630 546 4643 580
rect 4677 546 4690 580
rect 4630 487 4690 546
rect 4630 453 4643 487
rect 4677 453 4690 487
rect 4630 368 4690 453
rect 4720 580 4780 592
rect 4720 546 4733 580
rect 4767 546 4780 580
rect 4720 499 4780 546
rect 4720 465 4733 499
rect 4767 465 4780 499
rect 4720 419 4780 465
rect 4720 385 4733 419
rect 4767 385 4780 419
rect 4720 368 4780 385
rect 4810 580 4869 592
rect 4810 546 4823 580
rect 4857 546 4869 580
rect 4810 497 4869 546
rect 4810 463 4823 497
rect 4857 463 4869 497
rect 4810 414 4869 463
rect 4810 380 4823 414
rect 4857 380 4869 414
rect 4810 368 4869 380
<< ndiffc >>
rect -1738 3084 -1704 3460
rect -1650 3084 -1616 3460
rect -1738 2370 -1704 2746
rect -1650 2370 -1616 2746
rect -956 3084 -922 3460
rect -868 3084 -834 3460
rect -956 2370 -922 2746
rect -868 2370 -834 2746
rect -2767 1508 -2733 1542
rect -2767 1418 -2733 1452
rect -2667 1508 -2633 1542
rect -1398 1500 -1364 1534
rect -2667 1418 -2633 1452
rect -1398 1418 -1364 1452
rect -1234 1500 -1200 1534
rect -1234 1418 -1200 1452
rect -1102 1443 -1068 1477
rect -846 1443 -812 1477
rect -590 1443 -556 1477
rect 242 1443 276 1477
rect 498 1443 532 1477
rect 754 1443 788 1477
rect 914 1443 948 1477
rect 1170 1443 1204 1477
rect 1426 1443 1460 1477
rect 1586 1443 1620 1477
rect 1842 1443 1876 1477
rect 2098 1443 2132 1477
rect 2258 1443 2292 1477
rect 2514 1443 2548 1477
rect 2770 1443 2804 1477
rect 2930 1443 2964 1477
rect 3186 1443 3220 1477
rect 3442 1443 3476 1477
rect 3602 1443 3636 1477
rect 3858 1443 3892 1477
rect 4114 1443 4148 1477
rect 4274 1443 4308 1477
rect 4530 1443 4564 1477
rect -2767 1212 -2733 1246
rect -2767 1122 -2733 1156
rect -2667 1212 -2633 1246
rect -1398 1212 -1364 1246
rect -2667 1122 -2633 1156
rect -1398 1130 -1364 1164
rect -1234 1212 -1200 1246
rect -1234 1130 -1200 1164
rect -1113 1148 -1079 1182
rect -1006 1212 -972 1246
rect -1024 1122 -990 1156
rect -811 1204 -777 1238
rect -477 1186 -443 1220
rect -363 1212 -329 1246
rect -363 1122 -329 1156
rect -246 1212 -212 1246
rect -246 1122 -212 1156
rect -160 1212 -126 1246
rect -160 1122 -126 1156
rect -74 1212 -40 1246
rect -74 1122 -40 1156
rect 994 1250 1028 1284
rect 236 1162 270 1196
rect 400 1157 434 1191
rect 480 1157 514 1191
rect 644 1163 678 1197
rect 780 1152 814 1186
rect 892 1098 926 1132
rect 1146 1163 1180 1197
rect 1146 1095 1180 1129
rect 1284 1214 1318 1248
rect 1686 1213 1720 1247
rect 1465 1148 1499 1182
rect 1565 1153 1599 1187
rect 1798 1143 1832 1177
rect 1908 1161 1942 1195
rect 2019 1161 2053 1195
rect 2200 1178 2234 1212
rect 2282 1178 2316 1212
rect 2364 1178 2398 1212
rect 2548 1246 2582 1280
rect 2664 1212 2698 1246
rect 2759 1160 2793 1194
rect 2861 1233 2895 1267
rect 3178 1212 3212 1246
rect 2972 1081 3006 1115
rect 3178 1122 3212 1156
rect 3264 1212 3298 1246
rect 3264 1122 3298 1156
rect 3350 1212 3384 1246
rect 3350 1122 3384 1156
rect 3476 1186 3510 1220
rect 3476 1118 3510 1152
rect 3582 1212 3616 1246
rect 3582 1138 3616 1172
rect 3682 1212 3716 1246
rect 3682 1138 3716 1172
rect 3768 1212 3802 1246
rect 3768 1122 3802 1156
rect 3883 1216 3917 1250
rect 3955 1216 3989 1250
rect 4071 1212 4105 1246
rect 4071 1122 4105 1156
rect 4157 1190 4191 1224
rect 4243 1212 4277 1246
rect 4243 1122 4277 1156
rect 4329 1190 4363 1224
rect 4415 1212 4449 1246
rect 4415 1122 4449 1156
rect 4515 1158 4549 1192
rect 4615 1190 4649 1224
rect 4719 1158 4753 1192
rect 4823 1190 4857 1224
rect -1615 176 -1581 210
rect -1615 86 -1581 120
rect -1515 176 -1481 210
rect -246 168 -212 202
rect -1515 86 -1481 120
rect -246 86 -212 120
rect -82 168 -48 202
rect -82 86 -48 120
rect 236 136 270 170
rect 400 141 434 175
rect 480 141 514 175
rect 644 135 678 169
rect 780 146 814 180
rect 892 200 926 234
rect 1146 203 1180 237
rect 1146 135 1180 169
rect 1465 150 1499 184
rect 1565 145 1599 179
rect 1798 155 1832 189
rect 1908 137 1942 171
rect 2019 137 2053 171
rect 994 48 1028 82
rect 1284 84 1318 118
rect 1686 85 1720 119
rect 2200 120 2234 154
rect 2282 120 2316 154
rect 2364 120 2398 154
rect 2548 52 2582 86
rect 2664 86 2698 120
rect 2759 138 2793 172
rect 2972 217 3006 251
rect 3178 176 3212 210
rect 2861 65 2895 99
rect 3178 86 3212 120
rect 3264 176 3298 210
rect 3264 86 3298 120
rect 3350 176 3384 210
rect 3350 86 3384 120
rect 3476 180 3510 214
rect 3476 112 3510 146
rect 3582 160 3616 194
rect 3582 86 3616 120
rect 3682 160 3716 194
rect 3682 86 3716 120
rect 3768 176 3802 210
rect 3768 86 3802 120
rect 4071 201 4105 235
rect 4071 131 4105 165
rect 4161 134 4195 168
rect 4247 205 4281 239
rect 4247 127 4281 161
rect 4347 195 4381 229
rect 4347 127 4381 161
rect 4449 201 4483 235
rect 4449 123 4483 157
rect 3883 82 3917 116
rect 3955 82 3989 116
rect 4551 185 4585 219
rect 4551 111 4585 145
rect 4651 117 4685 151
rect 4737 201 4771 235
rect 4737 111 4771 145
rect 4823 201 4857 235
rect 4823 111 4857 145
rect -1389 -686 -1355 -310
rect -1301 -686 -1267 -310
rect -1389 -1400 -1355 -1024
rect -1301 -1400 -1267 -1024
<< pdiffc >>
rect -2767 1878 -2733 1912
rect -2767 1808 -2733 1842
rect -2767 1738 -2733 1772
rect -2667 1878 -2633 1912
rect -2667 1795 -2633 1829
rect -1403 1878 -1369 1912
rect -1403 1795 -1369 1829
rect -2667 1712 -2633 1746
rect -1403 1712 -1369 1746
rect -1313 1878 -1279 1912
rect -1313 1795 -1279 1829
rect -1313 1712 -1279 1746
rect -1223 1878 -1189 1912
rect -1223 1795 -1189 1829
rect -1223 1712 -1189 1746
rect -1117 1878 -1083 1912
rect -1117 1807 -1083 1841
rect -1117 1736 -1083 1770
rect -859 1878 -825 1912
rect -859 1807 -825 1841
rect -859 1736 -825 1770
rect -604 1878 -570 1912
rect -604 1807 -570 1841
rect -604 1736 -570 1770
rect 227 1878 261 1912
rect 227 1807 261 1841
rect 227 1736 261 1770
rect 485 1878 519 1912
rect 485 1807 519 1841
rect 485 1736 519 1770
rect 740 1878 774 1912
rect 740 1807 774 1841
rect 740 1736 774 1770
rect 899 1878 933 1912
rect 899 1807 933 1841
rect 899 1736 933 1770
rect 1157 1878 1191 1912
rect 1157 1807 1191 1841
rect 1157 1736 1191 1770
rect 1412 1878 1446 1912
rect 1412 1807 1446 1841
rect 1412 1736 1446 1770
rect 1571 1878 1605 1912
rect 1571 1807 1605 1841
rect 1571 1736 1605 1770
rect 1829 1878 1863 1912
rect 1829 1807 1863 1841
rect 1829 1736 1863 1770
rect 2084 1878 2118 1912
rect 2084 1807 2118 1841
rect 2084 1736 2118 1770
rect 2243 1878 2277 1912
rect 2243 1807 2277 1841
rect 2243 1736 2277 1770
rect 2501 1878 2535 1912
rect 2501 1807 2535 1841
rect 2501 1736 2535 1770
rect 2756 1878 2790 1912
rect 2756 1807 2790 1841
rect 2756 1736 2790 1770
rect 2915 1878 2949 1912
rect 2915 1807 2949 1841
rect 2915 1736 2949 1770
rect 3173 1878 3207 1912
rect 3173 1807 3207 1841
rect 3173 1736 3207 1770
rect 3428 1878 3462 1912
rect 3428 1807 3462 1841
rect 3428 1736 3462 1770
rect 3587 1878 3621 1912
rect 3587 1807 3621 1841
rect 3587 1736 3621 1770
rect 3845 1878 3879 1912
rect 3845 1807 3879 1841
rect 3845 1736 3879 1770
rect 4100 1878 4134 1912
rect 4100 1807 4134 1841
rect 4100 1736 4134 1770
rect 4259 1878 4293 1912
rect 4259 1807 4293 1841
rect 4259 1736 4293 1770
rect 4517 1878 4551 1912
rect 4517 1807 4551 1841
rect 4517 1736 4551 1770
rect -2767 892 -2733 926
rect -2767 822 -2733 856
rect -2767 752 -2733 786
rect -2667 918 -2633 952
rect -1403 918 -1369 952
rect -2667 835 -2633 869
rect -2667 752 -2633 786
rect -1403 835 -1369 869
rect -1403 752 -1369 786
rect -1313 918 -1279 952
rect -1313 835 -1279 869
rect -1313 752 -1279 786
rect -1223 918 -1189 952
rect -1223 835 -1189 869
rect -1113 903 -1079 937
rect -1113 808 -1079 842
rect -1006 813 -972 847
rect -1223 752 -1189 786
rect -723 918 -689 952
rect -723 801 -689 835
rect -477 918 -443 952
rect -477 835 -443 869
rect -477 752 -443 786
rect -377 918 -343 952
rect -377 835 -343 869
rect -377 752 -343 786
rect -251 892 -217 926
rect -251 822 -217 856
rect -251 752 -217 786
rect -161 918 -127 952
rect -161 835 -127 869
rect -161 752 -127 786
rect -71 918 -37 952
rect -71 835 -37 869
rect -71 752 -37 786
rect 893 892 927 926
rect 231 821 265 855
rect 231 752 265 786
rect 321 753 355 787
rect 489 812 523 846
rect 579 822 613 856
rect 579 752 613 786
rect 691 822 725 856
rect 691 752 725 786
rect 781 822 815 856
rect 781 752 815 786
rect 893 822 927 856
rect 893 752 927 786
rect 983 830 1017 864
rect 983 752 1017 786
rect 1073 914 1107 948
rect 1073 833 1107 867
rect 1073 752 1107 786
rect 1185 804 1219 838
rect 1376 812 1410 846
rect 1476 812 1510 846
rect 1588 752 1622 786
rect 1707 752 1741 786
rect 1881 789 1915 823
rect 1989 862 2023 896
rect 1989 752 2023 786
rect 2101 824 2135 858
rect 2101 752 2135 786
rect 2269 862 2303 896
rect 2569 830 2603 864
rect 2269 752 2303 786
rect 2454 757 2488 791
rect 2569 752 2603 786
rect 2669 757 2703 791
rect 2845 870 2879 904
rect 2957 881 2991 915
rect 3176 885 3210 919
rect 2845 752 2879 786
rect 3176 803 3210 837
rect 3064 713 3098 747
rect 3176 713 3210 747
rect 3283 918 3317 952
rect 3283 835 3317 869
rect 3283 752 3317 786
rect 3373 892 3407 926
rect 3373 822 3407 856
rect 3373 752 3407 786
rect 3482 902 3516 936
rect 3482 831 3516 865
rect 3482 760 3516 794
rect 3587 906 3621 940
rect 3587 834 3621 868
rect 3587 756 3621 790
rect 3677 918 3711 952
rect 3677 835 3711 869
rect 3677 752 3711 786
rect 3767 918 3801 952
rect 3767 835 3801 869
rect 3767 752 3801 786
rect 3883 748 3917 782
rect 3955 748 3989 782
rect 4071 912 4105 946
rect 4071 832 4105 866
rect 4071 752 4105 786
rect 4162 892 4196 926
rect 4242 892 4276 926
rect 4324 892 4358 926
rect 4162 821 4196 855
rect 4242 821 4276 855
rect 4324 821 4358 855
rect 4162 752 4196 786
rect 4242 752 4276 786
rect 4324 752 4358 786
rect 4414 831 4448 865
rect 4414 752 4448 786
rect 4514 892 4548 926
rect 4583 892 4617 926
rect 4654 892 4688 926
rect 4723 892 4757 926
rect 4514 821 4548 855
rect 4583 821 4617 855
rect 4654 821 4688 855
rect 4723 821 4757 855
rect 4514 752 4548 786
rect 4583 752 4617 786
rect 4654 752 4688 786
rect 4723 752 4757 786
rect 4823 831 4857 865
rect 4823 752 4857 786
rect -1615 546 -1581 580
rect -1615 476 -1581 510
rect -1615 406 -1581 440
rect -1515 546 -1481 580
rect -1515 463 -1481 497
rect -251 546 -217 580
rect -251 463 -217 497
rect -1515 380 -1481 414
rect -251 380 -217 414
rect -161 546 -127 580
rect -161 463 -127 497
rect -161 380 -127 414
rect -71 546 -37 580
rect -71 463 -37 497
rect 231 546 265 580
rect 231 477 265 511
rect 321 545 355 579
rect 489 486 523 520
rect 579 546 613 580
rect 579 476 613 510
rect 691 546 725 580
rect 691 476 725 510
rect 781 546 815 580
rect 781 476 815 510
rect 893 546 927 580
rect 893 476 927 510
rect -71 380 -37 414
rect 893 406 927 440
rect 983 546 1017 580
rect 983 468 1017 502
rect 1073 546 1107 580
rect 1073 465 1107 499
rect 1185 494 1219 528
rect 1376 486 1410 520
rect 1476 486 1510 520
rect 1588 546 1622 580
rect 1707 546 1741 580
rect 1073 384 1107 418
rect 1881 509 1915 543
rect 1989 546 2023 580
rect 1989 436 2023 470
rect 2101 546 2135 580
rect 2101 474 2135 508
rect 2269 546 2303 580
rect 2454 541 2488 575
rect 2569 546 2603 580
rect 2269 436 2303 470
rect 2569 468 2603 502
rect 2669 541 2703 575
rect 2845 546 2879 580
rect 3064 585 3098 619
rect 3176 585 3210 619
rect 2845 428 2879 462
rect 2957 417 2991 451
rect 3176 495 3210 529
rect 3176 413 3210 447
rect 3283 546 3317 580
rect 3283 463 3317 497
rect 3283 380 3317 414
rect 3373 546 3407 580
rect 3373 476 3407 510
rect 3373 406 3407 440
rect 3482 538 3516 572
rect 3482 467 3516 501
rect 3482 396 3516 430
rect 3587 542 3621 576
rect 3587 464 3621 498
rect 3587 392 3621 426
rect 3677 546 3711 580
rect 3677 463 3711 497
rect 3677 380 3711 414
rect 3767 546 3801 580
rect 3767 463 3801 497
rect 3767 380 3801 414
rect 3883 550 3917 584
rect 3955 550 3989 584
rect 4072 531 4106 565
rect 4072 421 4106 455
rect 4162 531 4196 565
rect 4162 421 4196 455
rect 4252 534 4286 568
rect 4252 466 4286 500
rect 4352 531 4386 565
rect 4352 421 4386 455
rect 4459 546 4493 580
rect 4459 474 4493 508
rect 4553 546 4587 580
rect 4553 465 4587 499
rect 4553 385 4587 419
rect 4643 546 4677 580
rect 4643 453 4677 487
rect 4733 546 4767 580
rect 4733 465 4767 499
rect 4733 385 4767 419
rect 4823 546 4857 580
rect 4823 463 4857 497
rect 4823 380 4857 414
<< psubdiff >>
rect -1852 3612 -1756 3646
rect -1598 3612 -1502 3646
rect -1852 3550 -1818 3612
rect -1536 3550 -1502 3612
rect -1852 2932 -1818 2994
rect -1536 2932 -1502 2994
rect -1852 2898 -1756 2932
rect -1598 2898 -1502 2932
rect -1852 2836 -1818 2898
rect -1536 2836 -1502 2898
rect -1852 2218 -1818 2280
rect -1536 2218 -1502 2280
rect -1852 2184 -1756 2218
rect -1598 2184 -1502 2218
rect -1070 3612 -974 3646
rect -816 3612 -720 3646
rect -1070 3550 -1036 3612
rect -754 3550 -720 3612
rect -1070 2932 -1036 2994
rect -754 2932 -720 2994
rect -1070 2898 -974 2932
rect -816 2898 -720 2932
rect -1070 2836 -1036 2898
rect -754 2836 -720 2898
rect -1070 2218 -1036 2280
rect -754 2218 -720 2280
rect -1070 2184 -974 2218
rect -816 2184 -720 2218
rect 31 1537 161 1561
rect 65 1503 127 1537
rect 31 1454 161 1503
rect 65 1420 127 1454
rect 31 1396 161 1420
rect 31 1244 161 1268
rect 65 1210 127 1244
rect 31 1161 161 1210
rect 65 1127 127 1161
rect 31 1103 161 1127
rect 31 205 161 229
rect 65 171 127 205
rect 31 122 161 171
rect 65 88 127 122
rect 31 64 161 88
rect -1503 -158 -1407 -124
rect -1249 -158 -1153 -124
rect -1503 -220 -1469 -158
rect -1187 -220 -1153 -158
rect -1503 -838 -1469 -776
rect -1187 -838 -1153 -776
rect -1503 -872 -1407 -838
rect -1249 -872 -1153 -838
rect -1503 -934 -1469 -872
rect -1187 -934 -1153 -872
rect -1503 -1552 -1469 -1490
rect -1187 -1552 -1153 -1490
rect -1503 -1586 -1407 -1552
rect -1249 -1586 -1153 -1552
<< nsubdiff >>
rect 31 1910 161 1934
rect 65 1876 127 1910
rect 31 1824 161 1876
rect 65 1790 127 1824
rect 31 1766 161 1790
rect 31 874 161 898
rect 65 840 127 874
rect 31 788 161 840
rect 65 754 127 788
rect 31 730 161 754
rect 31 578 161 602
rect 65 544 127 578
rect 31 492 161 544
rect 65 458 127 492
rect 31 434 161 458
<< psubdiffcont >>
rect -1756 3612 -1598 3646
rect -1852 2994 -1818 3550
rect -1536 2994 -1502 3550
rect -1756 2898 -1598 2932
rect -1852 2280 -1818 2836
rect -1536 2280 -1502 2836
rect -1756 2184 -1598 2218
rect -974 3612 -816 3646
rect -1070 2994 -1036 3550
rect -754 2994 -720 3550
rect -974 2898 -816 2932
rect -1070 2280 -1036 2836
rect -754 2280 -720 2836
rect -974 2184 -816 2218
rect 31 1503 65 1537
rect 127 1503 161 1537
rect 31 1420 65 1454
rect 127 1420 161 1454
rect 31 1210 65 1244
rect 127 1210 161 1244
rect 31 1127 65 1161
rect 127 1127 161 1161
rect 31 171 65 205
rect 127 171 161 205
rect 31 88 65 122
rect 127 88 161 122
rect -1407 -158 -1249 -124
rect -1503 -776 -1469 -220
rect -1187 -776 -1153 -220
rect -1407 -872 -1249 -838
rect -1503 -1490 -1469 -934
rect -1187 -1490 -1153 -934
rect -1407 -1586 -1249 -1552
<< nsubdiffcont >>
rect 31 1876 65 1910
rect 127 1876 161 1910
rect 31 1790 65 1824
rect 127 1790 161 1824
rect 31 840 65 874
rect 127 840 161 874
rect 31 754 65 788
rect 127 754 161 788
rect 31 544 65 578
rect 127 544 161 578
rect 31 458 65 492
rect 127 458 161 492
<< poly >>
rect -1710 3494 -1644 3560
rect -1692 3472 -1662 3494
rect -1692 3050 -1662 3072
rect -1710 3034 -1644 3050
rect -1710 3000 -1694 3034
rect -1660 3000 -1644 3034
rect -1710 2984 -1644 3000
rect -1710 2780 -1644 2846
rect -1692 2758 -1662 2780
rect -1692 2336 -1662 2358
rect -1710 2320 -1644 2336
rect -1710 2286 -1694 2320
rect -1660 2286 -1644 2320
rect -1710 2270 -1644 2286
rect -928 3494 -862 3560
rect -910 3472 -880 3494
rect -910 3050 -880 3072
rect -928 3034 -862 3050
rect -928 3000 -912 3034
rect -878 3000 -862 3034
rect -928 2984 -862 3000
rect -928 2780 -862 2846
rect -910 2758 -880 2780
rect -910 2336 -880 2358
rect -928 2320 -862 2336
rect -928 2286 -912 2320
rect -878 2286 -862 2320
rect -928 2270 -862 2286
rect -2710 1924 -2680 1950
rect -1356 1924 -1326 1950
rect -1266 1924 -1236 1950
rect -1070 1924 -870 1950
rect -815 1924 -615 1950
rect -2710 1685 -2680 1700
rect -2713 1658 -2677 1685
rect -2851 1651 -2677 1658
rect -2853 1642 -2677 1651
rect -2853 1608 -2835 1642
rect -2801 1608 -2767 1642
rect -2733 1608 -2677 1642
rect -2853 1599 -2677 1608
rect -2851 1592 -2677 1599
rect -2708 1554 -2678 1592
rect 274 1924 474 1950
rect 529 1924 729 1950
rect 946 1924 1146 1950
rect 1201 1924 1401 1950
rect 1618 1924 1818 1950
rect 1873 1924 2073 1950
rect 2290 1924 2490 1950
rect 2545 1924 2745 1950
rect 2962 1924 3162 1950
rect 3217 1924 3417 1950
rect 3634 1924 3834 1950
rect 3889 1924 4089 1950
rect 4306 1924 4506 1950
rect -1356 1685 -1326 1700
rect -1266 1685 -1236 1700
rect -1070 1698 -870 1724
rect -815 1698 -615 1724
rect -1359 1642 -1323 1685
rect -1269 1642 -1233 1685
rect -1419 1626 -1323 1642
rect -1419 1592 -1403 1626
rect -1369 1592 -1323 1626
rect -1419 1576 -1323 1592
rect -1353 1554 -1323 1576
rect -1275 1626 -1173 1642
rect -1275 1592 -1223 1626
rect -1189 1592 -1173 1626
rect -1275 1576 -1173 1592
rect -1070 1633 -1004 1698
rect -1070 1599 -1054 1633
rect -1020 1599 -1004 1633
rect -1070 1583 -1004 1599
rect -923 1632 -736 1648
rect -923 1598 -907 1632
rect -873 1598 -786 1632
rect -752 1598 -736 1632
rect -1275 1554 -1245 1576
rect -923 1570 -736 1598
rect -681 1633 -615 1698
rect -681 1599 -665 1633
rect -631 1599 -615 1633
rect -681 1583 -615 1599
rect 274 1698 474 1724
rect 529 1698 729 1724
rect 274 1633 340 1698
rect 274 1599 290 1633
rect 324 1599 340 1633
rect 274 1583 340 1599
rect 421 1632 608 1648
rect 421 1598 437 1632
rect 471 1598 558 1632
rect 592 1598 608 1632
rect -923 1541 -857 1570
rect -1057 1501 -857 1541
rect -801 1541 -736 1570
rect 421 1570 608 1598
rect 663 1633 729 1698
rect 663 1599 679 1633
rect 713 1599 729 1633
rect 663 1583 729 1599
rect 946 1698 1146 1724
rect 1201 1698 1401 1724
rect 946 1633 1012 1698
rect 946 1599 962 1633
rect 996 1599 1012 1633
rect 946 1583 1012 1599
rect 1093 1632 1280 1648
rect 1093 1598 1109 1632
rect 1143 1598 1230 1632
rect 1264 1598 1280 1632
rect -801 1501 -601 1541
rect 421 1541 487 1570
rect 287 1501 487 1541
rect 543 1541 608 1570
rect 1093 1570 1280 1598
rect 1335 1633 1401 1698
rect 1335 1599 1351 1633
rect 1385 1599 1401 1633
rect 1335 1583 1401 1599
rect 1618 1698 1818 1724
rect 1873 1698 2073 1724
rect 1618 1633 1684 1698
rect 1618 1599 1634 1633
rect 1668 1599 1684 1633
rect 1618 1583 1684 1599
rect 1765 1632 1952 1648
rect 1765 1598 1781 1632
rect 1815 1598 1902 1632
rect 1936 1598 1952 1632
rect 1093 1541 1159 1570
rect 543 1501 743 1541
rect 959 1501 1159 1541
rect 1215 1541 1280 1570
rect 1765 1570 1952 1598
rect 2007 1633 2073 1698
rect 2007 1599 2023 1633
rect 2057 1599 2073 1633
rect 2007 1583 2073 1599
rect 2290 1698 2490 1724
rect 2545 1698 2745 1724
rect 2290 1633 2356 1698
rect 2290 1599 2306 1633
rect 2340 1599 2356 1633
rect 2290 1583 2356 1599
rect 2437 1632 2624 1648
rect 2437 1598 2453 1632
rect 2487 1598 2574 1632
rect 2608 1598 2624 1632
rect 1765 1541 1831 1570
rect 1215 1501 1415 1541
rect 1631 1501 1831 1541
rect 1887 1541 1952 1570
rect 2437 1570 2624 1598
rect 2679 1633 2745 1698
rect 2679 1599 2695 1633
rect 2729 1599 2745 1633
rect 2679 1583 2745 1599
rect 2962 1698 3162 1724
rect 3217 1698 3417 1724
rect 2962 1633 3028 1698
rect 2962 1599 2978 1633
rect 3012 1599 3028 1633
rect 2962 1583 3028 1599
rect 3109 1632 3296 1648
rect 3109 1598 3125 1632
rect 3159 1598 3246 1632
rect 3280 1598 3296 1632
rect 2437 1541 2503 1570
rect 1887 1501 2087 1541
rect 2303 1501 2503 1541
rect 2559 1541 2624 1570
rect 3109 1570 3296 1598
rect 3351 1633 3417 1698
rect 3351 1599 3367 1633
rect 3401 1599 3417 1633
rect 3351 1583 3417 1599
rect 3634 1698 3834 1724
rect 3889 1698 4089 1724
rect 3634 1633 3700 1698
rect 3634 1599 3650 1633
rect 3684 1599 3700 1633
rect 3634 1583 3700 1599
rect 3781 1632 3968 1648
rect 3781 1598 3797 1632
rect 3831 1598 3918 1632
rect 3952 1598 3968 1632
rect 3109 1541 3175 1570
rect 2559 1501 2759 1541
rect 2975 1501 3175 1541
rect 3231 1541 3296 1570
rect 3781 1570 3968 1598
rect 4023 1633 4089 1698
rect 4023 1599 4039 1633
rect 4073 1599 4089 1633
rect 4023 1583 4089 1599
rect 4306 1698 4506 1724
rect 4306 1633 4372 1698
rect 4306 1599 4322 1633
rect 4356 1599 4372 1633
rect 4306 1583 4372 1599
rect 4453 1632 4519 1648
rect 4453 1598 4469 1632
rect 4503 1598 4519 1632
rect 3781 1541 3847 1570
rect 3231 1501 3431 1541
rect 3647 1501 3847 1541
rect 3903 1541 3968 1570
rect 4453 1541 4519 1598
rect 3903 1501 4103 1541
rect 4319 1501 4519 1541
rect -2708 1380 -2678 1406
rect -1353 1380 -1323 1406
rect -1275 1380 -1245 1406
rect -1057 1379 -857 1417
rect -801 1379 -601 1417
rect 287 1379 487 1417
rect 543 1379 743 1417
rect 959 1379 1159 1417
rect 1215 1379 1415 1417
rect 1631 1379 1831 1417
rect 1887 1379 2087 1417
rect 2303 1379 2503 1417
rect 2559 1379 2759 1417
rect 2975 1379 3175 1417
rect 3231 1379 3431 1417
rect 3647 1379 3847 1417
rect 3903 1379 4103 1417
rect 4319 1379 4519 1417
rect -2708 1258 -2678 1284
rect -1353 1258 -1323 1284
rect -1275 1258 -1245 1284
rect -956 1258 -926 1284
rect -878 1258 -848 1284
rect -739 1258 -709 1284
rect -547 1258 -517 1284
rect -404 1258 -374 1284
rect -201 1258 -171 1284
rect -115 1258 -85 1284
rect 359 1281 769 1311
rect -2708 1072 -2678 1110
rect -2851 1065 -2677 1072
rect -2853 1056 -2677 1065
rect -2853 1022 -2835 1056
rect -2801 1022 -2767 1056
rect -2733 1022 -2677 1056
rect -2853 1013 -2677 1022
rect -2851 1006 -2677 1013
rect -2713 979 -2677 1006
rect -2710 964 -2680 979
rect -1068 1220 -1038 1246
rect 281 1213 311 1239
rect 359 1213 389 1281
rect 525 1213 555 1239
rect 603 1213 633 1239
rect 739 1213 769 1281
rect 937 1234 967 1260
rect 1105 1281 2189 1311
rect 1105 1234 1135 1281
rect -1353 1088 -1323 1110
rect -1419 1072 -1323 1088
rect -1419 1038 -1403 1072
rect -1369 1038 -1323 1072
rect -1419 1022 -1323 1038
rect -1275 1088 -1245 1110
rect -1275 1072 -1173 1088
rect -1275 1038 -1223 1072
rect -1189 1038 -1173 1072
rect -1068 1062 -1038 1110
rect -956 1062 -926 1110
rect -878 1088 -848 1110
rect -739 1088 -709 1110
rect -1275 1022 -1173 1038
rect -1069 1046 -926 1062
rect -1359 979 -1323 1022
rect -1269 979 -1233 1022
rect -1069 1012 -1035 1046
rect -1001 1012 -926 1046
rect -883 1072 -817 1088
rect -883 1038 -867 1072
rect -833 1038 -817 1072
rect -883 1022 -817 1038
rect -775 1072 -709 1088
rect -775 1038 -759 1072
rect -725 1038 -709 1072
rect -775 1022 -709 1038
rect -661 1072 -595 1088
rect -661 1038 -645 1072
rect -611 1038 -595 1072
rect -661 1022 -595 1038
rect -547 1068 -517 1110
rect -404 1072 -374 1110
rect -201 1072 -171 1110
rect -115 1072 -85 1110
rect 281 1107 311 1129
rect 359 1107 389 1129
rect 236 1091 311 1107
rect -547 1052 -481 1068
rect -1069 996 -926 1012
rect -1069 979 -1033 996
rect -962 979 -926 996
rect -769 979 -733 1022
rect -661 979 -625 1022
rect -547 1018 -531 1052
rect -497 1018 -481 1052
rect -547 1002 -481 1018
rect -439 1056 -373 1072
rect -439 1022 -423 1056
rect -389 1022 -373 1056
rect -439 1006 -373 1022
rect -267 1056 -81 1072
rect -267 1022 -251 1056
rect -217 1042 -81 1056
rect -217 1022 -171 1042
rect -267 1006 -171 1022
rect -547 979 -511 1002
rect -423 979 -387 1006
rect -207 979 -171 1006
rect -117 979 -81 1042
rect 236 1057 252 1091
rect 286 1057 311 1091
rect 236 1023 311 1057
rect 236 989 252 1023
rect 286 989 311 1023
rect -1356 964 -1326 979
rect -1266 964 -1236 979
rect -1066 964 -1036 979
rect -959 964 -929 979
rect -766 964 -736 979
rect -658 964 -628 979
rect -544 964 -514 979
rect -420 964 -390 979
rect -204 964 -174 979
rect -114 964 -84 979
rect -1066 770 -1036 796
rect -2710 714 -2680 740
rect -1356 714 -1326 740
rect -1266 714 -1236 740
rect -959 738 -929 764
rect -766 738 -736 764
rect -658 738 -628 764
rect -544 738 -514 764
rect 236 955 311 989
rect 353 1091 419 1107
rect 353 1057 369 1091
rect 403 1057 419 1091
rect 353 1023 419 1057
rect 525 1040 555 1129
rect 353 989 369 1023
rect 403 989 419 1023
rect 353 973 419 989
rect 461 1024 555 1040
rect 461 990 505 1024
rect 539 990 555 1024
rect 461 974 555 990
rect 603 1000 633 1129
rect 739 1114 769 1129
rect 739 1084 857 1114
rect 1347 1207 1377 1233
rect 1419 1207 1449 1281
rect 2159 1250 2189 1281
rect 2409 1250 2439 1276
rect 2487 1250 2517 1276
rect 1510 1207 1540 1233
rect 1757 1207 1787 1233
rect 1843 1207 1873 1233
rect 1964 1207 1994 1233
rect 2064 1207 2094 1233
rect 1347 1108 1377 1123
rect 713 1020 779 1036
rect 713 1000 729 1020
rect 603 986 729 1000
rect 763 986 779 1020
rect 236 921 252 955
rect 286 921 311 955
rect 236 905 311 921
rect 275 883 311 905
rect 365 883 401 973
rect 461 925 491 974
rect 443 895 491 925
rect 603 970 779 986
rect 603 922 633 970
rect 827 922 857 1084
rect 937 1062 967 1086
rect 1105 1064 1135 1086
rect 905 1046 973 1062
rect 905 1012 921 1046
rect 955 1012 973 1046
rect 905 996 973 1012
rect 1015 1048 1135 1064
rect 1015 1014 1031 1048
rect 1065 1014 1135 1048
rect 1015 998 1135 1014
rect 1233 1078 1377 1108
rect 937 979 973 996
rect 1027 979 1063 998
rect 940 964 970 979
rect 1030 964 1060 979
rect 1233 966 1263 1078
rect 1311 1014 1377 1030
rect 1311 980 1327 1014
rect 1361 980 1377 1014
rect 443 883 479 895
rect 533 892 633 922
rect 735 892 857 922
rect 533 883 569 892
rect 735 883 771 892
rect 278 868 308 883
rect 368 868 398 883
rect 446 868 476 883
rect 536 868 566 883
rect 738 868 768 883
rect -420 714 -390 740
rect -204 714 -174 740
rect -114 714 -84 740
rect 1199 950 1265 966
rect 1311 964 1377 980
rect 1199 916 1215 950
rect 1249 916 1265 950
rect 1199 900 1265 916
rect 1229 883 1265 900
rect 1313 883 1349 964
rect 1419 913 1449 1123
rect 1510 1027 1540 1123
rect 2614 1258 2644 1284
rect 2718 1258 2748 1284
rect 2804 1258 2834 1284
rect 2159 1125 2189 1140
rect 1757 1075 1787 1097
rect 1843 1075 1873 1097
rect 1599 1059 1787 1075
rect 1491 1011 1557 1027
rect 1491 977 1507 1011
rect 1541 977 1557 1011
rect 1491 961 1557 977
rect 1599 1025 1615 1059
rect 1649 1045 1787 1059
rect 1649 1025 1665 1045
rect 1599 991 1665 1025
rect 1599 957 1615 991
rect 1649 957 1665 991
rect 1599 941 1665 957
rect 1751 923 1787 1045
rect 1835 1059 1901 1075
rect 1835 1025 1851 1059
rect 1885 1025 1901 1059
rect 1964 1042 1994 1097
rect 1835 991 1901 1025
rect 1835 957 1851 991
rect 1885 957 1901 991
rect 1835 941 1901 957
rect 1943 1026 2016 1042
rect 1943 992 1966 1026
rect 2000 992 2016 1026
rect 1943 976 2016 992
rect 2064 1016 2094 1097
rect 2159 1095 2361 1125
rect 2223 1031 2289 1047
rect 2064 1000 2181 1016
rect 1835 923 1871 941
rect 1943 923 1979 976
rect 2064 966 2131 1000
rect 2165 966 2181 1000
rect 2064 950 2181 966
rect 2145 923 2181 950
rect 2223 997 2239 1031
rect 2273 997 2289 1031
rect 2223 981 2289 997
rect 2223 923 2259 981
rect 2331 933 2361 1095
rect 2409 1079 2439 1166
rect 2487 1151 2517 1166
rect 2487 1121 2541 1151
rect 2403 1063 2469 1079
rect 2403 1029 2419 1063
rect 2453 1029 2469 1063
rect 2403 1013 2469 1029
rect 1419 883 1456 913
rect 1754 908 1784 923
rect 1838 908 1868 923
rect 1946 908 1976 923
rect 2148 908 2178 923
rect 2226 908 2256 923
rect 1232 868 1262 883
rect 1316 868 1346 883
rect 1423 868 1453 883
rect 1232 758 1262 784
rect 1316 758 1346 784
rect 2330 839 2366 933
rect 2511 922 2541 1121
rect 3223 1258 3253 1284
rect 3309 1258 3339 1284
rect 3017 1152 3047 1178
rect 2614 1088 2644 1110
rect 2718 1088 2748 1110
rect 2583 1072 2649 1088
rect 2583 1038 2599 1072
rect 2633 1038 2649 1072
rect 2583 1022 2649 1038
rect 2691 1072 2757 1088
rect 2691 1038 2707 1072
rect 2741 1038 2757 1072
rect 2804 1038 2834 1110
rect 3521 1238 3551 1264
rect 3641 1258 3671 1284
rect 3727 1258 3757 1284
rect 4116 1258 4146 1284
rect 4202 1258 4232 1284
rect 4288 1258 4318 1284
rect 4374 1258 4404 1284
rect 4468 1258 4498 1284
rect 4560 1258 4590 1284
rect 4660 1258 4690 1284
rect 4773 1258 4803 1284
rect 2691 1022 2757 1038
rect 2799 1022 2865 1038
rect 3017 1031 3047 1068
rect 3223 1062 3253 1110
rect 3309 1062 3339 1110
rect 3521 1062 3551 1110
rect 3641 1088 3671 1110
rect 3727 1088 3757 1110
rect 3599 1072 3757 1088
rect 3223 1046 3557 1062
rect 2613 955 2649 1022
rect 2715 955 2751 1022
rect 2799 988 2815 1022
rect 2849 988 2865 1022
rect 2799 972 2865 988
rect 2981 1015 3047 1031
rect 2981 981 2997 1015
rect 3031 981 3047 1015
rect 2799 955 2835 972
rect 2981 965 3047 981
rect 3089 1030 3557 1046
rect 3089 996 3105 1030
rect 3139 1003 3557 1030
rect 3599 1038 3615 1072
rect 3649 1038 3757 1072
rect 3599 1022 3757 1038
rect 3139 996 3155 1003
rect 3089 980 3155 996
rect 3237 979 3273 1003
rect 3327 979 3363 1003
rect 3526 1002 3557 1003
rect 2616 940 2646 955
rect 2718 940 2748 955
rect 2802 940 2832 955
rect 3001 948 3037 965
rect 3240 964 3270 979
rect 3330 964 3360 979
rect 2408 906 2541 922
rect 2408 872 2424 906
rect 2458 892 2541 906
rect 2458 872 2474 892
rect 2408 856 2474 872
rect 2408 839 2444 856
rect 2333 824 2363 839
rect 2411 824 2441 839
rect 3004 933 3034 948
rect 3004 779 3034 805
rect 278 714 308 740
rect 368 714 398 740
rect 446 714 476 740
rect 536 714 566 740
rect 738 714 768 740
rect 940 714 970 740
rect 1030 714 1060 740
rect 1423 714 1453 740
rect 1754 714 1784 740
rect 1838 714 1868 740
rect 1946 714 1976 740
rect 2148 714 2178 740
rect 2226 714 2256 740
rect 2333 714 2363 740
rect 2411 714 2441 740
rect 2616 714 2646 740
rect 2718 714 2748 740
rect 2802 714 2832 740
rect 3526 963 3562 1002
rect 3631 979 3667 1022
rect 3721 979 3757 1022
rect 4116 1062 4146 1110
rect 4202 1062 4232 1110
rect 4288 1062 4318 1110
rect 4374 1062 4404 1110
rect 4116 1046 4404 1062
rect 4116 1012 4150 1046
rect 4184 1012 4218 1046
rect 4252 1012 4286 1046
rect 4320 1012 4354 1046
rect 4388 1012 4404 1046
rect 4116 996 4404 1012
rect 4116 979 4152 996
rect 4368 979 4404 996
rect 4468 1062 4498 1110
rect 4560 1062 4590 1110
rect 4660 1062 4690 1110
rect 4773 1062 4803 1110
rect 4468 1046 4803 1062
rect 4468 1012 4537 1046
rect 4571 1012 4605 1046
rect 4639 1012 4673 1046
rect 4707 1012 4741 1046
rect 4775 1012 4803 1046
rect 4468 996 4803 1012
rect 4468 979 4504 996
rect 4767 979 4803 996
rect 3634 964 3664 979
rect 3724 964 3754 979
rect 4119 964 4149 979
rect 4371 964 4401 979
rect 4471 964 4501 979
rect 4770 964 4800 979
rect 3529 948 3559 963
rect 3240 714 3270 740
rect 3330 714 3360 740
rect 3529 722 3559 748
rect 3634 714 3664 740
rect 3724 714 3754 740
rect 4119 714 4149 740
rect 4371 714 4401 740
rect 4471 714 4501 740
rect 4770 714 4800 740
rect -1558 592 -1528 618
rect -204 592 -174 618
rect -114 592 -84 618
rect -1558 353 -1528 368
rect -1561 326 -1525 353
rect -1699 319 -1525 326
rect -1701 310 -1525 319
rect -1701 276 -1683 310
rect -1649 276 -1615 310
rect -1581 276 -1525 310
rect -1701 267 -1525 276
rect -1699 260 -1525 267
rect -1556 222 -1526 260
rect 278 592 308 618
rect 368 592 398 618
rect 446 592 476 618
rect 536 592 566 618
rect 738 592 768 618
rect 940 592 970 618
rect 1030 592 1060 618
rect 1423 592 1453 618
rect 1754 592 1784 618
rect 1838 592 1868 618
rect 1946 592 1976 618
rect 2148 592 2178 618
rect 2226 592 2256 618
rect 2333 592 2363 618
rect 2411 592 2441 618
rect 2616 592 2646 618
rect 2718 592 2748 618
rect 2802 592 2832 618
rect 278 449 308 464
rect 368 449 398 464
rect 446 449 476 464
rect 536 449 566 464
rect 738 449 768 464
rect 275 427 311 449
rect 236 411 311 427
rect 236 377 252 411
rect 286 377 311 411
rect -204 353 -174 368
rect -114 353 -84 368
rect -207 310 -171 353
rect -117 310 -81 353
rect 236 343 311 377
rect 365 359 401 449
rect 443 437 479 449
rect 533 440 569 449
rect 735 440 771 449
rect 443 407 491 437
rect 533 410 633 440
rect 735 410 857 440
rect -267 294 -171 310
rect -267 260 -251 294
rect -217 260 -171 294
rect -267 244 -171 260
rect -201 222 -171 244
rect -123 294 -21 310
rect -123 260 -71 294
rect -37 260 -21 294
rect -123 244 -21 260
rect 236 309 252 343
rect 286 309 311 343
rect 236 275 311 309
rect -123 222 -93 244
rect 236 241 252 275
rect 286 241 311 275
rect 236 225 311 241
rect 353 343 419 359
rect 353 309 369 343
rect 403 309 419 343
rect 353 275 419 309
rect 461 358 491 407
rect 603 362 633 410
rect 461 342 555 358
rect 461 308 505 342
rect 539 308 555 342
rect 461 292 555 308
rect 353 241 369 275
rect 403 241 419 275
rect 353 225 419 241
rect 281 203 311 225
rect 359 203 389 225
rect 525 203 555 292
rect 603 346 779 362
rect 603 332 729 346
rect 603 203 633 332
rect 713 312 729 332
rect 763 312 779 346
rect 713 296 779 312
rect 827 248 857 410
rect 1232 548 1262 574
rect 1316 548 1346 574
rect 1232 449 1262 464
rect 1316 449 1346 464
rect 1423 449 1453 464
rect 1229 432 1265 449
rect 1199 416 1265 432
rect 1199 382 1215 416
rect 1249 382 1265 416
rect 940 353 970 368
rect 1030 353 1060 368
rect 1199 366 1265 382
rect 1313 368 1349 449
rect 1419 419 1456 449
rect 2333 493 2363 508
rect 2411 493 2441 508
rect 937 336 973 353
rect 905 320 973 336
rect 1027 334 1063 353
rect 905 286 921 320
rect 955 286 973 320
rect 905 270 973 286
rect 1015 318 1135 334
rect 1015 284 1031 318
rect 1065 284 1135 318
rect 739 218 857 248
rect 937 246 967 270
rect 1015 268 1135 284
rect 1105 246 1135 268
rect 1233 254 1263 366
rect 1311 352 1377 368
rect 1311 318 1327 352
rect 1361 318 1377 352
rect 1311 302 1377 318
rect 739 203 769 218
rect 281 93 311 119
rect -1556 48 -1526 74
rect -201 48 -171 74
rect -123 48 -93 74
rect 359 51 389 119
rect 525 93 555 119
rect 603 93 633 119
rect 739 51 769 119
rect 1233 224 1377 254
rect 1347 209 1377 224
rect 1419 209 1449 419
rect 1754 409 1784 424
rect 1838 409 1868 424
rect 1946 409 1976 424
rect 2148 409 2178 424
rect 2226 409 2256 424
rect 1599 375 1665 391
rect 1491 355 1557 371
rect 1491 321 1507 355
rect 1541 321 1557 355
rect 1491 305 1557 321
rect 1599 341 1615 375
rect 1649 341 1665 375
rect 1599 307 1665 341
rect 1510 209 1540 305
rect 1599 273 1615 307
rect 1649 287 1665 307
rect 1751 287 1787 409
rect 1649 273 1787 287
rect 1599 257 1787 273
rect 1835 391 1871 409
rect 1835 375 1901 391
rect 1835 341 1851 375
rect 1885 341 1901 375
rect 1835 307 1901 341
rect 1835 273 1851 307
rect 1885 273 1901 307
rect 1943 356 1979 409
rect 2145 382 2181 409
rect 2064 366 2181 382
rect 1943 340 2016 356
rect 1943 306 1966 340
rect 2000 306 2016 340
rect 1943 290 2016 306
rect 2064 332 2131 366
rect 2165 332 2181 366
rect 2064 316 2181 332
rect 2223 351 2259 409
rect 2330 399 2366 493
rect 2408 476 2444 493
rect 2408 460 2474 476
rect 2408 426 2424 460
rect 2458 440 2474 460
rect 2458 426 2541 440
rect 2408 410 2541 426
rect 2223 335 2289 351
rect 1835 257 1901 273
rect 1757 235 1787 257
rect 1843 235 1873 257
rect 1964 235 1994 290
rect 2064 235 2094 316
rect 2223 301 2239 335
rect 2273 301 2289 335
rect 2223 285 2289 301
rect 2331 237 2361 399
rect 2403 303 2469 319
rect 2403 269 2419 303
rect 2453 269 2469 303
rect 2403 253 2469 269
rect 2159 207 2361 237
rect 2159 192 2189 207
rect 937 72 967 98
rect 359 21 769 51
rect 1105 51 1135 98
rect 1347 99 1377 125
rect 1419 51 1449 125
rect 1510 99 1540 125
rect 1757 99 1787 125
rect 1843 99 1873 125
rect 1964 99 1994 125
rect 2064 99 2094 125
rect 2409 166 2439 253
rect 2511 211 2541 410
rect 3240 592 3270 618
rect 3330 592 3360 618
rect 3004 527 3034 553
rect 2616 377 2646 392
rect 2718 377 2748 392
rect 2802 377 2832 392
rect 3004 384 3034 399
rect 2613 310 2649 377
rect 2715 310 2751 377
rect 2799 360 2835 377
rect 3001 367 3037 384
rect 3529 584 3559 610
rect 3634 592 3664 618
rect 3724 592 3754 618
rect 3529 369 3559 384
rect 2799 344 2865 360
rect 2799 310 2815 344
rect 2849 310 2865 344
rect 2583 294 2649 310
rect 2583 260 2599 294
rect 2633 260 2649 294
rect 2583 244 2649 260
rect 2691 294 2757 310
rect 2799 294 2865 310
rect 2981 351 3047 367
rect 3240 353 3270 368
rect 3330 353 3360 368
rect 2981 317 2997 351
rect 3031 317 3047 351
rect 2981 301 3047 317
rect 2691 260 2707 294
rect 2741 260 2757 294
rect 2691 244 2757 260
rect 2614 222 2644 244
rect 2718 222 2748 244
rect 2804 222 2834 294
rect 3017 264 3047 301
rect 3089 336 3155 352
rect 3089 302 3105 336
rect 3139 329 3155 336
rect 3237 329 3273 353
rect 3327 329 3363 353
rect 3526 330 3562 369
rect 4119 577 4149 603
rect 4209 577 4239 603
rect 4304 577 4334 603
rect 4399 577 4429 603
rect 4506 592 4536 618
rect 4600 592 4630 618
rect 4690 592 4720 618
rect 4780 592 4810 618
rect 4119 394 4149 409
rect 4209 394 4239 409
rect 4304 394 4334 409
rect 4399 394 4429 409
rect 3634 353 3664 368
rect 3724 353 3754 368
rect 3526 329 3557 330
rect 3139 302 3557 329
rect 3631 310 3667 353
rect 3721 310 3757 353
rect 3089 286 3557 302
rect 3223 270 3557 286
rect 3599 294 3757 310
rect 2487 181 2541 211
rect 2487 166 2517 181
rect 2159 51 2189 82
rect 2409 56 2439 82
rect 2487 56 2517 82
rect 1105 21 2189 51
rect 3223 222 3253 270
rect 3309 222 3339 270
rect 3521 222 3551 270
rect 3599 260 3615 294
rect 3649 260 3757 294
rect 3599 244 3757 260
rect 4116 262 4152 394
rect 4206 383 4242 394
rect 4301 383 4337 394
rect 4206 340 4337 383
rect 4206 306 4261 340
rect 4295 306 4337 340
rect 4396 335 4432 394
rect 4506 353 4536 368
rect 4600 353 4630 368
rect 4690 353 4720 368
rect 4780 353 4810 368
rect 4503 335 4539 353
rect 4597 335 4633 353
rect 4687 335 4723 353
rect 4777 335 4813 353
rect 4206 290 4337 306
rect 4379 319 4445 335
rect 4116 247 4146 262
rect 4206 247 4236 290
rect 4301 247 4331 290
rect 4379 285 4395 319
rect 4429 285 4445 319
rect 4379 269 4445 285
rect 4493 319 4813 335
rect 4493 285 4509 319
rect 4543 285 4577 319
rect 4611 285 4645 319
rect 4679 285 4813 319
rect 4493 269 4813 285
rect 4392 247 4422 269
rect 4494 247 4524 269
rect 4610 247 4640 269
rect 4696 247 4726 269
rect 4782 247 4812 269
rect 3641 222 3671 244
rect 3727 222 3757 244
rect 3017 154 3047 180
rect 2614 48 2644 74
rect 2718 48 2748 74
rect 2804 48 2834 74
rect 3223 48 3253 74
rect 3309 48 3339 74
rect 3521 68 3551 94
rect 3641 48 3671 74
rect 3727 48 3757 74
rect 4116 51 4146 119
rect 4206 93 4236 119
rect 4301 93 4331 119
rect 4392 51 4422 119
rect 4494 73 4524 99
rect 4610 73 4640 99
rect 4696 73 4726 99
rect 4782 73 4812 99
rect 4116 21 4422 51
rect -1361 -276 -1295 -210
rect -1343 -298 -1313 -276
rect -1343 -720 -1313 -698
rect -1361 -736 -1295 -720
rect -1361 -770 -1345 -736
rect -1311 -770 -1295 -736
rect -1361 -786 -1295 -770
rect -1361 -990 -1295 -924
rect -1343 -1012 -1313 -990
rect -1343 -1434 -1313 -1412
rect -1361 -1450 -1295 -1434
rect -1361 -1484 -1345 -1450
rect -1311 -1484 -1295 -1450
rect -1361 -1500 -1295 -1484
<< polycont >>
rect -1694 3000 -1660 3034
rect -1694 2286 -1660 2320
rect -912 3000 -878 3034
rect -912 2286 -878 2320
rect -2835 1608 -2801 1642
rect -2767 1608 -2733 1642
rect -1403 1592 -1369 1626
rect -1223 1592 -1189 1626
rect -1054 1599 -1020 1633
rect -907 1598 -873 1632
rect -786 1598 -752 1632
rect -665 1599 -631 1633
rect 290 1599 324 1633
rect 437 1598 471 1632
rect 558 1598 592 1632
rect 679 1599 713 1633
rect 962 1599 996 1633
rect 1109 1598 1143 1632
rect 1230 1598 1264 1632
rect 1351 1599 1385 1633
rect 1634 1599 1668 1633
rect 1781 1598 1815 1632
rect 1902 1598 1936 1632
rect 2023 1599 2057 1633
rect 2306 1599 2340 1633
rect 2453 1598 2487 1632
rect 2574 1598 2608 1632
rect 2695 1599 2729 1633
rect 2978 1599 3012 1633
rect 3125 1598 3159 1632
rect 3246 1598 3280 1632
rect 3367 1599 3401 1633
rect 3650 1599 3684 1633
rect 3797 1598 3831 1632
rect 3918 1598 3952 1632
rect 4039 1599 4073 1633
rect 4322 1599 4356 1633
rect 4469 1598 4503 1632
rect -2835 1022 -2801 1056
rect -2767 1022 -2733 1056
rect -1403 1038 -1369 1072
rect -1223 1038 -1189 1072
rect -1035 1012 -1001 1046
rect -867 1038 -833 1072
rect -759 1038 -725 1072
rect -645 1038 -611 1072
rect -531 1018 -497 1052
rect -423 1022 -389 1056
rect -251 1022 -217 1056
rect 252 1057 286 1091
rect 252 989 286 1023
rect 369 1057 403 1091
rect 369 989 403 1023
rect 505 990 539 1024
rect 729 986 763 1020
rect 252 921 286 955
rect 921 1012 955 1046
rect 1031 1014 1065 1048
rect 1327 980 1361 1014
rect 1215 916 1249 950
rect 1507 977 1541 1011
rect 1615 1025 1649 1059
rect 1615 957 1649 991
rect 1851 1025 1885 1059
rect 1851 957 1885 991
rect 1966 992 2000 1026
rect 2131 966 2165 1000
rect 2239 997 2273 1031
rect 2419 1029 2453 1063
rect 2599 1038 2633 1072
rect 2707 1038 2741 1072
rect 2815 988 2849 1022
rect 2997 981 3031 1015
rect 3105 996 3139 1030
rect 3615 1038 3649 1072
rect 2424 872 2458 906
rect 4150 1012 4184 1046
rect 4218 1012 4252 1046
rect 4286 1012 4320 1046
rect 4354 1012 4388 1046
rect 4537 1012 4571 1046
rect 4605 1012 4639 1046
rect 4673 1012 4707 1046
rect 4741 1012 4775 1046
rect -1683 276 -1649 310
rect -1615 276 -1581 310
rect 252 377 286 411
rect -251 260 -217 294
rect -71 260 -37 294
rect 252 309 286 343
rect 252 241 286 275
rect 369 309 403 343
rect 505 308 539 342
rect 369 241 403 275
rect 729 312 763 346
rect 1215 382 1249 416
rect 921 286 955 320
rect 1031 284 1065 318
rect 1327 318 1361 352
rect 1507 321 1541 355
rect 1615 341 1649 375
rect 1615 273 1649 307
rect 1851 341 1885 375
rect 1851 273 1885 307
rect 1966 306 2000 340
rect 2131 332 2165 366
rect 2424 426 2458 460
rect 2239 301 2273 335
rect 2419 269 2453 303
rect 2815 310 2849 344
rect 2599 260 2633 294
rect 2997 317 3031 351
rect 2707 260 2741 294
rect 3105 302 3139 336
rect 3615 260 3649 294
rect 4261 306 4295 340
rect 4395 285 4429 319
rect 4509 285 4543 319
rect 4577 285 4611 319
rect 4645 285 4679 319
rect -1345 -770 -1311 -736
rect -1345 -1484 -1311 -1450
<< xpolycontact >>
rect -2516 1467 -2084 1749
rect -1984 1467 -1552 1749
rect -2516 915 -2084 1197
rect -1984 915 -1552 1197
rect -1364 135 -932 417
rect -832 135 -400 417
<< xpolyres >>
rect -2084 1467 -1984 1749
rect -2084 915 -1984 1197
rect -932 135 -832 417
<< locali >>
rect -1852 3612 -1756 3646
rect -1598 3612 -1468 3646
rect -1852 3550 -1818 3612
rect -1536 3550 -1468 3612
rect -1738 3460 -1704 3476
rect -1738 3068 -1704 3084
rect -1650 3460 -1616 3476
rect -1650 3068 -1616 3084
rect -1710 3000 -1694 3034
rect -1660 3000 -1644 3034
rect -1852 2932 -1818 2994
rect -1502 2994 -1468 3550
rect -1536 2932 -1468 2994
rect -1852 2898 -1756 2932
rect -1598 2898 -1468 2932
rect -1852 2836 -1818 2898
rect -1536 2836 -1468 2898
rect -1738 2746 -1704 2762
rect -1738 2354 -1704 2370
rect -1650 2746 -1616 2762
rect -1650 2354 -1616 2370
rect -1710 2286 -1694 2320
rect -1660 2286 -1644 2320
rect -1852 2218 -1818 2280
rect -1502 2280 -1468 2836
rect -1536 2218 -1468 2280
rect -1852 2184 -1756 2218
rect -1598 2184 -1468 2218
rect -1104 3612 -974 3646
rect -816 3612 -720 3646
rect -1104 3550 -1036 3612
rect -1104 2994 -1070 3550
rect -754 3550 -720 3612
rect -956 3460 -922 3476
rect -956 3068 -922 3084
rect -868 3460 -834 3476
rect -868 3068 -834 3084
rect -928 3000 -912 3034
rect -878 3000 -862 3034
rect -1104 2932 -1036 2994
rect -754 2932 -720 2994
rect -1104 2898 -974 2932
rect -816 2898 -720 2932
rect -1104 2836 -1036 2898
rect -1104 2280 -1070 2836
rect -754 2836 -720 2898
rect -956 2746 -922 2762
rect -956 2354 -922 2370
rect -868 2746 -834 2762
rect -868 2354 -834 2370
rect -928 2286 -912 2320
rect -878 2286 -862 2320
rect -1104 2218 -1036 2280
rect -754 2218 -720 2280
rect -1104 2184 -974 2218
rect -816 2184 -720 2218
rect -2880 1981 -2849 2015
rect -2815 1981 -2753 2015
rect -2719 1981 -2657 2015
rect -2623 1981 -2561 2015
rect -2527 1981 -2465 2015
rect -2431 1981 -2369 2015
rect -2335 1981 -2273 2015
rect -2239 1981 -2177 2015
rect -2143 1981 -2081 2015
rect -2047 1981 -1985 2015
rect -1951 1981 -1889 2015
rect -1855 1981 -1793 2015
rect -1759 1981 -1697 2015
rect -1663 1981 -1601 2015
rect -1567 1981 -1505 2015
rect -1471 1981 -1409 2015
rect -1375 1981 -1313 2015
rect -1279 1981 -1217 2015
rect -1183 1981 -1121 2015
rect -1087 1981 -1025 2015
rect -991 1981 -929 2015
rect -895 1981 -833 2015
rect -799 1981 -737 2015
rect -703 1981 -641 2015
rect -607 1981 -545 2015
rect -511 1981 -449 2015
rect -415 1981 -353 2015
rect -319 1981 -257 2015
rect -223 1981 -161 2015
rect -127 1981 -65 2015
rect -31 1981 31 2015
rect 65 1981 127 2015
rect 161 1981 223 2015
rect 257 1981 319 2015
rect 353 1981 415 2015
rect 449 1981 511 2015
rect 545 1981 607 2015
rect 641 1981 703 2015
rect 737 1981 799 2015
rect 833 1981 895 2015
rect 929 1981 991 2015
rect 1025 1981 1087 2015
rect 1121 1981 1183 2015
rect 1217 1981 1279 2015
rect 1313 1981 1375 2015
rect 1409 1981 1471 2015
rect 1505 1981 1567 2015
rect 1601 1981 1663 2015
rect 1697 1981 1759 2015
rect 1793 1981 1855 2015
rect 1889 1981 1951 2015
rect 1985 1981 2047 2015
rect 2081 1981 2143 2015
rect 2177 1981 2239 2015
rect 2273 1981 2335 2015
rect 2369 1981 2431 2015
rect 2465 1981 2527 2015
rect 2561 1981 2623 2015
rect 2657 1981 2719 2015
rect 2753 1981 2815 2015
rect 2849 1981 2911 2015
rect 2945 1981 3007 2015
rect 3041 1981 3103 2015
rect 3137 1981 3199 2015
rect 3233 1981 3295 2015
rect 3329 1981 3391 2015
rect 3425 1981 3487 2015
rect 3521 1981 3583 2015
rect 3617 1981 3679 2015
rect 3713 1981 3775 2015
rect 3809 1981 3871 2015
rect 3905 1981 3967 2015
rect 4001 1981 4063 2015
rect 4097 1981 4159 2015
rect 4193 1981 4255 2015
rect 4289 1981 4351 2015
rect 4385 1981 4447 2015
rect 4481 1981 4543 2015
rect 4577 1981 4639 2015
rect 4673 1981 4735 2015
rect 4769 1981 4831 2015
rect 4865 1981 4896 2015
rect -2783 1912 -2717 1981
rect -2783 1878 -2767 1912
rect -2733 1878 -2717 1912
rect -2783 1842 -2717 1878
rect -2783 1808 -2767 1842
rect -2733 1808 -2717 1842
rect -2783 1772 -2717 1808
rect -2783 1738 -2767 1772
rect -2733 1738 -2717 1772
rect -2783 1722 -2717 1738
rect -2683 1912 -2617 1928
rect -2683 1878 -2667 1912
rect -2633 1878 -2617 1912
rect -2683 1829 -2617 1878
rect -2683 1795 -2667 1829
rect -2633 1795 -2617 1829
rect -2683 1746 -2617 1795
rect -1419 1912 -1353 1981
rect -1419 1878 -1403 1912
rect -1369 1878 -1353 1912
rect -1419 1829 -1353 1878
rect -1419 1795 -1403 1829
rect -1369 1795 -1353 1829
rect -2683 1712 -2667 1746
rect -2633 1712 -2617 1746
rect -2855 1642 -2717 1688
rect -2855 1608 -2839 1642
rect -2801 1608 -2767 1642
rect -2733 1608 -2717 1642
rect -2855 1592 -2717 1608
rect -2683 1659 -2617 1712
rect -2683 1600 -2516 1659
rect -2783 1542 -2717 1558
rect -2783 1508 -2767 1542
rect -2733 1508 -2717 1542
rect -2783 1452 -2717 1508
rect -2783 1418 -2767 1452
rect -2733 1418 -2717 1452
rect -2783 1349 -2717 1418
rect -2683 1542 -2617 1600
rect -2683 1508 -2667 1542
rect -2633 1508 -2617 1542
rect -2683 1452 -2617 1508
rect -1419 1746 -1353 1795
rect -1419 1712 -1403 1746
rect -1369 1712 -1353 1746
rect -1419 1696 -1353 1712
rect -1319 1912 -1273 1928
rect -1319 1878 -1313 1912
rect -1279 1878 -1273 1912
rect -1319 1829 -1273 1878
rect -1319 1795 -1313 1829
rect -1279 1795 -1273 1829
rect -1319 1746 -1273 1795
rect -1319 1712 -1313 1746
rect -1279 1712 -1273 1746
rect -1552 1626 -1353 1642
rect -1552 1592 -1403 1626
rect -1369 1592 -1353 1626
rect -1552 1576 -1353 1592
rect -1419 1568 -1353 1576
rect -1319 1568 -1273 1712
rect -1239 1912 -1173 1981
rect -1239 1878 -1223 1912
rect -1189 1878 -1173 1912
rect -1239 1829 -1173 1878
rect -1239 1795 -1223 1829
rect -1189 1795 -1173 1829
rect -1239 1746 -1173 1795
rect -1239 1712 -1223 1746
rect -1189 1712 -1173 1746
rect -1133 1912 -1067 1981
rect -1133 1878 -1117 1912
rect -1083 1878 -1067 1912
rect -1133 1841 -1067 1878
rect -1133 1807 -1117 1841
rect -1083 1807 -1067 1841
rect -1133 1770 -1067 1807
rect -1133 1736 -1117 1770
rect -1083 1736 -1067 1770
rect -1133 1718 -1067 1736
rect -923 1912 -736 1981
rect -923 1878 -859 1912
rect -825 1878 -736 1912
rect -923 1841 -736 1878
rect -923 1807 -859 1841
rect -825 1807 -736 1841
rect -923 1770 -736 1807
rect -923 1736 -859 1770
rect -825 1736 -736 1770
rect -1239 1696 -1173 1712
rect -1239 1626 -1173 1642
rect -1239 1592 -1223 1626
rect -1189 1592 -1173 1626
rect -1239 1568 -1173 1592
rect -1118 1633 -1004 1649
rect -1118 1599 -1054 1633
rect -1020 1599 -1004 1633
rect -1307 1534 -1273 1568
rect -1414 1500 -1398 1534
rect -1364 1500 -1348 1534
rect -1307 1500 -1234 1534
rect -1200 1500 -1184 1534
rect -2683 1418 -2667 1452
rect -2633 1418 -2617 1452
rect -2683 1402 -2617 1418
rect -1414 1452 -1348 1500
rect -1414 1418 -1398 1452
rect -1364 1418 -1348 1452
rect -1414 1349 -1348 1418
rect -1250 1458 -1184 1500
rect -1250 1452 -1233 1458
rect -1250 1418 -1234 1452
rect -1199 1424 -1184 1458
rect -1200 1418 -1184 1424
rect -1250 1402 -1184 1418
rect -1118 1477 -1004 1599
rect -923 1632 -736 1736
rect -620 1912 -554 1981
rect -620 1878 -604 1912
rect -570 1878 -554 1912
rect -620 1841 -554 1878
rect -620 1807 -604 1841
rect -570 1807 -554 1841
rect -620 1770 -554 1807
rect 18 1910 174 1945
rect 18 1876 31 1910
rect 65 1876 127 1910
rect 18 1870 127 1876
rect 161 1870 174 1910
rect 18 1824 174 1870
rect 18 1790 31 1824
rect 65 1790 127 1824
rect 161 1790 174 1824
rect 18 1774 174 1790
rect 211 1912 277 1981
rect 211 1878 227 1912
rect 261 1878 277 1912
rect 211 1841 277 1878
rect 211 1807 227 1841
rect 261 1807 277 1841
rect -620 1736 -604 1770
rect -570 1736 -554 1770
rect -620 1720 -554 1736
rect 211 1770 277 1807
rect 211 1736 227 1770
rect 261 1736 277 1770
rect 211 1718 277 1736
rect 421 1912 608 1981
rect 421 1878 485 1912
rect 519 1878 608 1912
rect 421 1841 608 1878
rect 421 1807 485 1841
rect 519 1807 608 1841
rect 421 1770 608 1807
rect 421 1736 485 1770
rect 519 1736 608 1770
rect -923 1598 -907 1632
rect -873 1598 -786 1632
rect -752 1598 -736 1632
rect -923 1582 -736 1598
rect -681 1633 -541 1648
rect -681 1599 -665 1633
rect -631 1599 -541 1633
rect -1118 1443 -1102 1477
rect -1068 1443 -1004 1477
rect -1118 1349 -1004 1443
rect -862 1477 -796 1493
rect -862 1443 -846 1477
rect -812 1443 -796 1477
rect -862 1349 -796 1443
rect -681 1477 -541 1599
rect 226 1633 340 1649
rect 226 1599 290 1633
rect 324 1599 340 1633
rect -681 1443 -590 1477
rect -556 1443 -541 1477
rect -681 1349 -541 1443
rect 18 1537 174 1553
rect 18 1503 31 1537
rect 65 1503 127 1537
rect 161 1503 174 1537
rect 18 1460 174 1503
rect 18 1420 31 1460
rect 65 1454 174 1460
rect 65 1420 127 1454
rect 161 1420 174 1454
rect 18 1385 174 1420
rect 226 1477 340 1599
rect 421 1632 608 1736
rect 724 1912 790 1981
rect 724 1878 740 1912
rect 774 1878 790 1912
rect 724 1841 790 1878
rect 724 1807 740 1841
rect 774 1807 790 1841
rect 724 1770 790 1807
rect 724 1736 740 1770
rect 774 1736 790 1770
rect 724 1720 790 1736
rect 883 1912 949 1981
rect 883 1878 899 1912
rect 933 1878 949 1912
rect 883 1841 949 1878
rect 883 1807 899 1841
rect 933 1807 949 1841
rect 883 1770 949 1807
rect 883 1736 899 1770
rect 933 1736 949 1770
rect 883 1718 949 1736
rect 1093 1912 1280 1981
rect 1093 1878 1157 1912
rect 1191 1878 1280 1912
rect 1093 1841 1280 1878
rect 1093 1807 1157 1841
rect 1191 1807 1280 1841
rect 1093 1770 1280 1807
rect 1093 1736 1157 1770
rect 1191 1736 1280 1770
rect 421 1598 437 1632
rect 471 1598 558 1632
rect 592 1598 608 1632
rect 421 1582 608 1598
rect 663 1633 803 1648
rect 663 1599 679 1633
rect 713 1599 803 1633
rect 226 1443 242 1477
rect 276 1443 340 1477
rect 226 1349 340 1443
rect 482 1477 548 1493
rect 482 1443 498 1477
rect 532 1443 548 1477
rect 482 1349 548 1443
rect 663 1477 803 1599
rect 663 1443 754 1477
rect 788 1443 803 1477
rect 663 1349 803 1443
rect 898 1633 1012 1649
rect 898 1599 962 1633
rect 996 1599 1012 1633
rect 898 1477 1012 1599
rect 1093 1632 1280 1736
rect 1396 1912 1462 1981
rect 1396 1878 1412 1912
rect 1446 1878 1462 1912
rect 1396 1841 1462 1878
rect 1396 1807 1412 1841
rect 1446 1807 1462 1841
rect 1396 1770 1462 1807
rect 1396 1736 1412 1770
rect 1446 1736 1462 1770
rect 1396 1720 1462 1736
rect 1555 1912 1621 1981
rect 1555 1878 1571 1912
rect 1605 1878 1621 1912
rect 1555 1841 1621 1878
rect 1555 1807 1571 1841
rect 1605 1807 1621 1841
rect 1555 1770 1621 1807
rect 1555 1736 1571 1770
rect 1605 1736 1621 1770
rect 1555 1718 1621 1736
rect 1765 1912 1952 1981
rect 1765 1878 1829 1912
rect 1863 1878 1952 1912
rect 1765 1841 1952 1878
rect 1765 1807 1829 1841
rect 1863 1807 1952 1841
rect 1765 1770 1952 1807
rect 1765 1736 1829 1770
rect 1863 1736 1952 1770
rect 1093 1598 1109 1632
rect 1143 1598 1230 1632
rect 1264 1598 1280 1632
rect 1093 1582 1280 1598
rect 1335 1633 1475 1648
rect 1335 1599 1351 1633
rect 1385 1599 1475 1633
rect 898 1443 914 1477
rect 948 1443 1012 1477
rect 898 1349 1012 1443
rect 1154 1477 1220 1493
rect 1154 1443 1170 1477
rect 1204 1443 1220 1477
rect 1154 1349 1220 1443
rect 1335 1477 1475 1599
rect 1335 1443 1426 1477
rect 1460 1443 1475 1477
rect 1335 1349 1475 1443
rect 1570 1633 1684 1649
rect 1570 1599 1634 1633
rect 1668 1599 1684 1633
rect 1570 1477 1684 1599
rect 1765 1632 1952 1736
rect 2068 1912 2134 1981
rect 2068 1878 2084 1912
rect 2118 1878 2134 1912
rect 2068 1841 2134 1878
rect 2068 1807 2084 1841
rect 2118 1807 2134 1841
rect 2068 1770 2134 1807
rect 2068 1736 2084 1770
rect 2118 1736 2134 1770
rect 2068 1720 2134 1736
rect 2227 1912 2293 1981
rect 2227 1878 2243 1912
rect 2277 1878 2293 1912
rect 2227 1841 2293 1878
rect 2227 1807 2243 1841
rect 2277 1807 2293 1841
rect 2227 1770 2293 1807
rect 2227 1736 2243 1770
rect 2277 1736 2293 1770
rect 2227 1718 2293 1736
rect 2437 1912 2624 1981
rect 2437 1878 2501 1912
rect 2535 1878 2624 1912
rect 2437 1841 2624 1878
rect 2437 1807 2501 1841
rect 2535 1807 2624 1841
rect 2437 1770 2624 1807
rect 2437 1736 2501 1770
rect 2535 1736 2624 1770
rect 1765 1598 1781 1632
rect 1815 1598 1902 1632
rect 1936 1598 1952 1632
rect 1765 1582 1952 1598
rect 2007 1633 2147 1648
rect 2007 1599 2023 1633
rect 2057 1599 2147 1633
rect 1570 1443 1586 1477
rect 1620 1443 1684 1477
rect 1570 1349 1684 1443
rect 1826 1477 1892 1493
rect 1826 1443 1842 1477
rect 1876 1443 1892 1477
rect 1826 1349 1892 1443
rect 2007 1477 2147 1599
rect 2007 1443 2098 1477
rect 2132 1443 2147 1477
rect 2007 1349 2147 1443
rect 2242 1633 2356 1649
rect 2242 1599 2306 1633
rect 2340 1599 2356 1633
rect 2242 1477 2356 1599
rect 2437 1632 2624 1736
rect 2740 1912 2806 1981
rect 2740 1878 2756 1912
rect 2790 1878 2806 1912
rect 2740 1841 2806 1878
rect 2740 1807 2756 1841
rect 2790 1807 2806 1841
rect 2740 1770 2806 1807
rect 2740 1736 2756 1770
rect 2790 1736 2806 1770
rect 2740 1720 2806 1736
rect 2899 1912 2965 1981
rect 2899 1878 2915 1912
rect 2949 1878 2965 1912
rect 2899 1841 2965 1878
rect 2899 1807 2915 1841
rect 2949 1807 2965 1841
rect 2899 1770 2965 1807
rect 2899 1736 2915 1770
rect 2949 1736 2965 1770
rect 2899 1718 2965 1736
rect 3109 1912 3296 1981
rect 3109 1878 3173 1912
rect 3207 1878 3296 1912
rect 3109 1841 3296 1878
rect 3109 1807 3173 1841
rect 3207 1807 3296 1841
rect 3109 1770 3296 1807
rect 3109 1736 3173 1770
rect 3207 1736 3296 1770
rect 2437 1598 2453 1632
rect 2487 1598 2574 1632
rect 2608 1598 2624 1632
rect 2437 1582 2624 1598
rect 2679 1633 2819 1648
rect 2679 1599 2695 1633
rect 2729 1599 2819 1633
rect 2242 1443 2258 1477
rect 2292 1443 2356 1477
rect 2242 1349 2356 1443
rect 2498 1477 2564 1493
rect 2498 1443 2514 1477
rect 2548 1443 2564 1477
rect 2498 1349 2564 1443
rect 2679 1477 2819 1599
rect 2679 1443 2770 1477
rect 2804 1443 2819 1477
rect 2679 1349 2819 1443
rect 2914 1633 3028 1649
rect 2914 1599 2978 1633
rect 3012 1599 3028 1633
rect 2914 1477 3028 1599
rect 3109 1632 3296 1736
rect 3412 1912 3478 1981
rect 3412 1878 3428 1912
rect 3462 1878 3478 1912
rect 3412 1841 3478 1878
rect 3412 1807 3428 1841
rect 3462 1807 3478 1841
rect 3412 1770 3478 1807
rect 3412 1736 3428 1770
rect 3462 1736 3478 1770
rect 3412 1720 3478 1736
rect 3571 1912 3637 1981
rect 3571 1878 3587 1912
rect 3621 1878 3637 1912
rect 3571 1841 3637 1878
rect 3571 1807 3587 1841
rect 3621 1807 3637 1841
rect 3571 1770 3637 1807
rect 3571 1736 3587 1770
rect 3621 1736 3637 1770
rect 3571 1718 3637 1736
rect 3781 1912 3968 1981
rect 3781 1878 3845 1912
rect 3879 1878 3968 1912
rect 3781 1841 3968 1878
rect 3781 1807 3845 1841
rect 3879 1807 3968 1841
rect 3781 1770 3968 1807
rect 3781 1736 3845 1770
rect 3879 1736 3968 1770
rect 3109 1598 3125 1632
rect 3159 1598 3246 1632
rect 3280 1598 3296 1632
rect 3109 1582 3296 1598
rect 3351 1633 3491 1648
rect 3351 1599 3367 1633
rect 3401 1599 3491 1633
rect 2914 1443 2930 1477
rect 2964 1443 3028 1477
rect 2914 1349 3028 1443
rect 3170 1477 3236 1493
rect 3170 1443 3186 1477
rect 3220 1443 3236 1477
rect 3170 1349 3236 1443
rect 3351 1477 3491 1599
rect 3351 1443 3442 1477
rect 3476 1443 3491 1477
rect 3351 1349 3491 1443
rect 3586 1633 3700 1649
rect 3586 1599 3650 1633
rect 3684 1599 3700 1633
rect 3586 1477 3700 1599
rect 3781 1632 3968 1736
rect 4084 1912 4150 1981
rect 4084 1878 4100 1912
rect 4134 1878 4150 1912
rect 4084 1841 4150 1878
rect 4084 1807 4100 1841
rect 4134 1807 4150 1841
rect 4084 1770 4150 1807
rect 4084 1736 4100 1770
rect 4134 1736 4150 1770
rect 4084 1720 4150 1736
rect 4243 1912 4309 1981
rect 4243 1878 4259 1912
rect 4293 1878 4309 1912
rect 4243 1841 4309 1878
rect 4243 1807 4259 1841
rect 4293 1807 4309 1841
rect 4243 1770 4309 1807
rect 4243 1736 4259 1770
rect 4293 1736 4309 1770
rect 4243 1718 4309 1736
rect 4453 1912 4567 1981
rect 4453 1878 4517 1912
rect 4551 1878 4567 1912
rect 4453 1841 4567 1878
rect 4453 1807 4517 1841
rect 4551 1807 4567 1841
rect 4453 1770 4567 1807
rect 4453 1736 4517 1770
rect 4551 1736 4567 1770
rect 3781 1598 3797 1632
rect 3831 1598 3918 1632
rect 3952 1598 3968 1632
rect 3781 1582 3968 1598
rect 4023 1633 4163 1648
rect 4023 1599 4039 1633
rect 4073 1599 4163 1633
rect 3586 1443 3602 1477
rect 3636 1443 3700 1477
rect 3586 1349 3700 1443
rect 3842 1477 3908 1493
rect 3842 1443 3858 1477
rect 3892 1443 3908 1477
rect 3842 1349 3908 1443
rect 4023 1477 4163 1599
rect 4023 1443 4114 1477
rect 4148 1443 4163 1477
rect 4023 1349 4163 1443
rect 4258 1633 4372 1649
rect 4258 1599 4322 1633
rect 4356 1599 4372 1633
rect 4258 1477 4372 1599
rect 4453 1632 4567 1736
rect 4453 1598 4469 1632
rect 4503 1598 4567 1632
rect 4453 1582 4567 1598
rect 4258 1443 4274 1477
rect 4308 1443 4372 1477
rect 4258 1349 4372 1443
rect 4514 1477 4580 1493
rect 4514 1443 4530 1477
rect 4564 1443 4580 1477
rect 4514 1349 4580 1443
rect -2880 1315 -2849 1349
rect -2815 1315 -2753 1349
rect -2719 1315 -2657 1349
rect -2623 1315 -2561 1349
rect -2527 1315 -2465 1349
rect -2431 1315 -2369 1349
rect -2335 1315 -2273 1349
rect -2239 1315 -2177 1349
rect -2143 1315 -2081 1349
rect -2047 1315 -1985 1349
rect -1951 1315 -1889 1349
rect -1855 1315 -1793 1349
rect -1759 1315 -1697 1349
rect -1663 1315 -1601 1349
rect -1567 1315 -1505 1349
rect -1471 1315 -1409 1349
rect -1375 1315 -1313 1349
rect -1279 1315 -1217 1349
rect -1183 1315 -1121 1349
rect -1087 1315 -1025 1349
rect -991 1315 -929 1349
rect -895 1315 -833 1349
rect -799 1315 -737 1349
rect -703 1315 -641 1349
rect -607 1315 -545 1349
rect -511 1315 -449 1349
rect -415 1315 -353 1349
rect -319 1315 -257 1349
rect -223 1315 -161 1349
rect -127 1315 -65 1349
rect -31 1315 31 1349
rect 65 1315 127 1349
rect 161 1315 223 1349
rect 257 1315 319 1349
rect 353 1315 415 1349
rect 449 1315 511 1349
rect 545 1315 607 1349
rect 641 1315 703 1349
rect 737 1315 799 1349
rect 833 1315 895 1349
rect 929 1315 991 1349
rect 1025 1315 1087 1349
rect 1121 1315 1183 1349
rect 1217 1315 1279 1349
rect 1313 1315 1375 1349
rect 1409 1315 1471 1349
rect 1505 1315 1567 1349
rect 1601 1315 1663 1349
rect 1697 1315 1759 1349
rect 1793 1315 1855 1349
rect 1889 1315 1951 1349
rect 1985 1315 2047 1349
rect 2081 1315 2143 1349
rect 2177 1315 2239 1349
rect 2273 1315 2335 1349
rect 2369 1315 2431 1349
rect 2465 1315 2527 1349
rect 2561 1315 2623 1349
rect 2657 1315 2719 1349
rect 2753 1315 2815 1349
rect 2849 1315 2911 1349
rect 2945 1315 3007 1349
rect 3041 1315 3103 1349
rect 3137 1315 3199 1349
rect 3233 1315 3295 1349
rect 3329 1315 3391 1349
rect 3425 1315 3487 1349
rect 3521 1315 3583 1349
rect 3617 1315 3679 1349
rect 3713 1315 3775 1349
rect 3809 1315 3871 1349
rect 3905 1315 3967 1349
rect 4001 1315 4063 1349
rect 4097 1315 4159 1349
rect 4193 1315 4255 1349
rect 4289 1315 4351 1349
rect 4385 1315 4447 1349
rect 4481 1315 4543 1349
rect 4577 1315 4639 1349
rect 4673 1315 4735 1349
rect 4769 1315 4831 1349
rect 4865 1315 4896 1349
rect -2783 1246 -2717 1315
rect -2783 1212 -2767 1246
rect -2733 1212 -2717 1246
rect -2783 1156 -2717 1212
rect -2783 1122 -2767 1156
rect -2733 1122 -2717 1156
rect -2783 1106 -2717 1122
rect -2683 1246 -2617 1262
rect -2683 1212 -2667 1246
rect -2633 1212 -2617 1246
rect -2683 1156 -2617 1212
rect -1414 1246 -1348 1315
rect -1414 1212 -1398 1246
rect -1364 1212 -1348 1246
rect -2683 1122 -2667 1156
rect -2633 1122 -2617 1156
rect -2855 1056 -2717 1072
rect -2855 1022 -2839 1056
rect -2801 1022 -2767 1056
rect -2733 1022 -2717 1056
rect -2855 976 -2717 1022
rect -2683 1064 -2617 1122
rect -2683 1005 -2516 1064
rect -2683 952 -2617 1005
rect -2783 926 -2717 942
rect -2783 892 -2767 926
rect -2733 892 -2717 926
rect -2783 856 -2717 892
rect -2783 822 -2767 856
rect -2733 822 -2717 856
rect -2783 786 -2717 822
rect -2783 752 -2767 786
rect -2733 752 -2717 786
rect -2783 683 -2717 752
rect -2683 918 -2667 952
rect -2633 918 -2617 952
rect -2683 869 -2617 918
rect -1414 1164 -1348 1212
rect -1250 1246 -1184 1262
rect -1250 1212 -1234 1246
rect -1200 1240 -1184 1246
rect -1250 1206 -1233 1212
rect -1199 1206 -1184 1240
rect -1027 1246 -951 1315
rect -1250 1164 -1184 1206
rect -1414 1130 -1398 1164
rect -1364 1130 -1348 1164
rect -1307 1130 -1234 1164
rect -1200 1130 -1184 1164
rect -1129 1182 -1063 1224
rect -1129 1148 -1113 1182
rect -1079 1148 -1063 1182
rect -1307 1096 -1273 1130
rect -1129 1106 -1063 1148
rect -1027 1212 -1006 1246
rect -972 1212 -951 1246
rect -1027 1196 -951 1212
rect -917 1238 -527 1254
rect -917 1204 -811 1238
rect -777 1204 -527 1238
rect -1027 1156 -985 1196
rect -917 1162 -883 1204
rect -1027 1122 -1024 1156
rect -990 1122 -985 1156
rect -1027 1106 -985 1122
rect -951 1128 -883 1162
rect -849 1136 -595 1170
rect -1419 1088 -1353 1096
rect -1552 1072 -1353 1088
rect -1552 1038 -1403 1072
rect -1369 1038 -1353 1072
rect -1552 1022 -1353 1038
rect -1419 952 -1353 968
rect -1419 918 -1403 952
rect -1369 918 -1353 952
rect -2683 835 -2667 869
rect -2633 835 -2617 869
rect -2683 786 -2617 835
rect -2683 752 -2667 786
rect -2633 752 -2617 786
rect -2683 736 -2617 752
rect -1419 869 -1353 918
rect -1419 835 -1403 869
rect -1369 835 -1353 869
rect -1419 786 -1353 835
rect -1419 752 -1403 786
rect -1369 752 -1353 786
rect -1419 683 -1353 752
rect -1319 952 -1273 1096
rect -1239 1072 -1173 1096
rect -1239 1038 -1223 1072
rect -1189 1038 -1173 1072
rect -1239 1022 -1173 1038
rect -1319 918 -1313 952
rect -1279 918 -1273 952
rect -1319 869 -1273 918
rect -1319 835 -1313 869
rect -1279 835 -1273 869
rect -1319 786 -1273 835
rect -1319 752 -1313 786
rect -1279 752 -1273 786
rect -1319 736 -1273 752
rect -1239 952 -1173 968
rect -1239 918 -1223 952
rect -1189 918 -1173 952
rect -1239 869 -1173 918
rect -1239 835 -1223 869
rect -1189 835 -1173 869
rect -1239 786 -1173 835
rect -1129 942 -1095 1106
rect -1051 1049 -985 1062
rect -1051 1015 -1036 1049
rect -1002 1046 -985 1049
rect -1051 1012 -1035 1015
rect -1001 1012 -985 1046
rect -1051 976 -985 1012
rect -951 988 -917 1128
rect -849 1088 -815 1136
rect -883 1072 -815 1088
rect -883 1038 -867 1072
rect -833 1038 -815 1072
rect -883 1022 -815 1038
rect -775 1072 -697 1096
rect -775 1038 -759 1072
rect -725 1038 -697 1072
rect -775 1022 -697 1038
rect -661 1074 -595 1136
rect -561 1136 -527 1204
rect -493 1220 -427 1315
rect -493 1186 -477 1220
rect -443 1186 -427 1220
rect -493 1170 -427 1186
rect -379 1246 -305 1262
rect -379 1212 -363 1246
rect -329 1212 -305 1246
rect -379 1156 -305 1212
rect -561 1102 -413 1136
rect -379 1122 -363 1156
rect -329 1122 -305 1156
rect -379 1106 -305 1122
rect -262 1246 -212 1315
rect -262 1212 -246 1246
rect -262 1156 -212 1212
rect -262 1122 -246 1156
rect -262 1106 -212 1122
rect -176 1246 -110 1262
rect -176 1212 -160 1246
rect -126 1212 -110 1246
rect -176 1156 -110 1212
rect -176 1122 -160 1156
rect -126 1122 -110 1156
rect -176 1106 -110 1122
rect -74 1246 -24 1315
rect -40 1212 -24 1246
rect -74 1156 -24 1212
rect -40 1122 -24 1156
rect -74 1106 -24 1122
rect 18 1244 174 1279
rect 18 1204 31 1244
rect 65 1210 127 1244
rect 161 1210 174 1244
rect 65 1204 174 1210
rect 18 1161 174 1204
rect 18 1127 31 1161
rect 65 1127 127 1161
rect 161 1127 174 1161
rect 18 1111 174 1127
rect 220 1196 286 1315
rect 220 1162 236 1196
rect 270 1162 286 1196
rect 220 1141 286 1162
rect 384 1191 530 1207
rect 384 1157 400 1191
rect 434 1157 480 1191
rect 514 1157 530 1191
rect 384 1141 530 1157
rect 628 1197 678 1315
rect 978 1284 1028 1315
rect 628 1163 644 1197
rect 628 1142 678 1163
rect 712 1247 899 1281
rect 220 1107 285 1141
rect 489 1108 530 1141
rect 712 1108 746 1247
rect -661 1038 -645 1074
rect -611 1038 -595 1074
rect -447 1072 -413 1102
rect -661 1022 -595 1038
rect -561 1052 -481 1068
rect -561 1018 -531 1052
rect -497 1018 -481 1052
rect -561 1002 -481 1018
rect -447 1056 -373 1072
rect -447 1022 -423 1056
rect -389 1022 -373 1056
rect -447 1006 -373 1022
rect -951 954 -673 988
rect -739 952 -673 954
rect -1129 937 -1063 942
rect -1129 903 -1113 937
rect -1079 920 -1063 937
rect -1079 903 -888 920
rect -1129 886 -888 903
rect -1129 842 -1063 886
rect -1129 808 -1113 842
rect -1079 808 -1063 842
rect -1129 792 -1063 808
rect -1022 847 -956 852
rect -1022 813 -1006 847
rect -972 813 -956 847
rect -1239 752 -1223 786
rect -1189 752 -1173 786
rect -1239 683 -1173 752
rect -1022 683 -956 813
rect -922 751 -888 886
rect -739 918 -723 952
rect -689 918 -673 952
rect -739 835 -673 918
rect -739 801 -723 835
rect -689 801 -673 835
rect -739 785 -673 801
rect -561 751 -527 1002
rect -339 968 -305 1106
rect -267 1061 -201 1072
rect -267 1027 -252 1061
rect -218 1056 -201 1061
rect -267 1022 -251 1027
rect -217 1022 -201 1056
rect -267 976 -201 1022
rect -922 717 -527 751
rect -493 952 -427 968
rect -493 918 -477 952
rect -443 918 -427 952
rect -493 869 -427 918
rect -493 835 -477 869
rect -443 835 -427 869
rect -493 786 -427 835
rect -493 752 -477 786
rect -443 752 -427 786
rect -493 683 -427 752
rect -393 952 -305 968
rect -393 918 -377 952
rect -343 918 -305 952
rect -167 952 -110 1106
rect 217 1091 455 1107
rect 217 1057 252 1091
rect 286 1057 369 1091
rect 403 1057 455 1091
rect 489 1074 746 1108
rect 780 1186 831 1213
rect 814 1152 831 1186
rect 865 1200 899 1247
rect 978 1250 994 1284
rect 978 1234 1028 1250
rect 1062 1247 1248 1281
rect 1062 1200 1096 1247
rect 865 1166 1096 1200
rect 1130 1197 1180 1213
rect 217 1040 455 1057
rect 217 1023 302 1040
rect 217 989 252 1023
rect 286 989 302 1023
rect -393 887 -305 918
rect -393 869 -360 887
rect -393 835 -377 869
rect -326 853 -305 887
rect -343 835 -305 853
rect -393 786 -305 835
rect -393 752 -377 786
rect -343 752 -305 786
rect -393 736 -305 752
rect -267 926 -201 942
rect -267 892 -251 926
rect -217 892 -201 926
rect -267 856 -201 892
rect -267 822 -251 856
rect -217 822 -201 856
rect -267 786 -201 822
rect -267 752 -251 786
rect -217 752 -201 786
rect -267 683 -201 752
rect -167 918 -161 952
rect -127 918 -110 952
rect -167 869 -110 918
rect -167 835 -161 869
rect -127 835 -110 869
rect -167 815 -110 835
rect -167 786 -158 815
rect -167 752 -161 786
rect -124 781 -110 815
rect -127 752 -110 781
rect -167 736 -110 752
rect -71 952 -21 968
rect -37 918 -21 952
rect -71 869 -21 918
rect 217 955 302 989
rect 353 1023 455 1040
rect 353 989 369 1023
rect 403 989 455 1023
rect 353 973 455 989
rect 489 1025 555 1040
rect 489 1024 509 1025
rect 489 990 505 1024
rect 543 991 555 1025
rect 539 990 555 991
rect 489 974 555 990
rect 217 921 252 955
rect 286 921 302 955
rect 589 940 623 1074
rect 780 1036 831 1152
rect 1130 1163 1146 1197
rect 876 1098 892 1132
rect 926 1098 1039 1132
rect 1005 1064 1039 1098
rect 1130 1129 1180 1163
rect 1214 1164 1248 1247
rect 1282 1248 1336 1315
rect 1282 1214 1284 1248
rect 1318 1214 1336 1248
rect 1282 1198 1336 1214
rect 1381 1245 1615 1279
rect 1381 1164 1415 1245
rect 1214 1130 1415 1164
rect 1449 1182 1515 1211
rect 1449 1148 1465 1182
rect 1499 1148 1515 1182
rect 1130 1096 1146 1129
rect 1115 1095 1146 1096
rect 1180 1095 1415 1096
rect 1115 1090 1415 1095
rect 713 1020 831 1036
rect 713 986 729 1020
rect 763 986 831 1020
rect 713 970 831 986
rect 889 1046 971 1062
rect 889 1012 917 1046
rect 955 1012 971 1046
rect 889 976 971 1012
rect 1005 1048 1081 1064
rect 1005 1014 1031 1048
rect 1065 1014 1081 1048
rect 1005 998 1081 1014
rect 1115 1062 1375 1090
rect 217 905 302 921
rect 489 906 623 940
rect -37 835 -21 869
rect -71 786 -21 835
rect -37 752 -21 786
rect -71 683 -21 752
rect 18 874 174 890
rect 18 840 31 874
rect 65 840 127 874
rect 161 840 174 874
rect 489 872 523 906
rect 18 794 174 840
rect 18 788 127 794
rect 18 754 31 788
rect 65 754 127 788
rect 161 754 174 794
rect 18 719 174 754
rect 215 855 439 871
rect 215 821 231 855
rect 265 837 439 855
rect 215 786 265 821
rect 215 752 231 786
rect 215 736 265 752
rect 305 787 371 803
rect 305 753 321 787
rect 355 753 371 787
rect 305 683 371 753
rect 405 751 439 837
rect 473 846 523 872
rect 473 812 489 846
rect 473 785 523 812
rect 563 856 629 872
rect 563 822 579 856
rect 613 822 629 856
rect 563 786 629 822
rect 563 752 579 786
rect 613 752 629 786
rect 563 751 629 752
rect 405 717 629 751
rect 675 856 741 872
rect 675 822 691 856
rect 725 822 741 856
rect 675 786 741 822
rect 675 752 691 786
rect 725 752 741 786
rect 675 683 741 752
rect 781 856 831 970
rect 1005 942 1039 998
rect 1115 964 1149 1062
rect 1311 1056 1375 1062
rect 1409 1056 1415 1090
rect 1449 1095 1515 1148
rect 1549 1187 1615 1245
rect 1661 1247 1916 1279
rect 1661 1213 1686 1247
rect 1720 1245 1916 1247
rect 1720 1213 1746 1245
rect 1661 1197 1746 1213
rect 1882 1211 1916 1245
rect 1549 1153 1565 1187
rect 1599 1163 1615 1187
rect 1782 1177 1848 1211
rect 1599 1153 1733 1163
rect 1549 1129 1733 1153
rect 1782 1143 1798 1177
rect 1832 1143 1848 1177
rect 1882 1195 1969 1211
rect 1882 1161 1908 1195
rect 1942 1161 1969 1195
rect 1882 1145 1969 1161
rect 2003 1195 2069 1315
rect 2528 1280 2603 1315
rect 2003 1161 2019 1195
rect 2053 1161 2069 1195
rect 2003 1144 2069 1161
rect 2103 1246 2494 1280
rect 2528 1246 2548 1280
rect 2582 1246 2603 1280
rect 2639 1267 2911 1281
rect 2639 1247 2861 1267
rect 2639 1246 2723 1247
rect 1449 1061 1665 1095
rect 1311 1027 1415 1056
rect 1599 1059 1665 1061
rect 1311 1014 1557 1027
rect 1311 980 1327 1014
rect 1361 1011 1557 1014
rect 1361 980 1507 1011
rect 1311 977 1507 980
rect 1541 977 1557 1011
rect 815 822 831 856
rect 781 786 831 822
rect 815 752 831 786
rect 781 736 831 752
rect 877 926 1039 942
rect 877 892 893 926
rect 927 908 1039 926
rect 1073 948 1149 964
rect 1107 914 1149 948
rect 877 856 927 892
rect 877 822 893 856
rect 877 786 927 822
rect 877 752 893 786
rect 877 736 927 752
rect 967 864 1033 874
rect 967 830 983 864
rect 1017 830 1033 864
rect 967 786 1033 830
rect 967 752 983 786
rect 1017 752 1033 786
rect 967 683 1033 752
rect 1073 867 1149 914
rect 1199 950 1265 966
rect 1311 964 1557 977
rect 1491 961 1557 964
rect 1599 1025 1615 1059
rect 1649 1025 1665 1059
rect 1599 991 1665 1025
rect 1199 916 1215 950
rect 1249 930 1265 950
rect 1599 957 1615 991
rect 1649 957 1665 991
rect 1249 916 1303 930
rect 1599 924 1665 957
rect 1199 896 1303 916
rect 1107 833 1149 867
rect 1073 786 1149 833
rect 1107 752 1149 786
rect 1073 736 1149 752
rect 1185 838 1235 862
rect 1219 804 1235 838
rect 1185 683 1235 804
rect 1269 751 1303 896
rect 1360 890 1665 924
rect 1360 846 1426 890
rect 1699 856 1733 1129
rect 1360 812 1376 846
rect 1410 812 1426 846
rect 1360 785 1426 812
rect 1460 846 1733 856
rect 1460 812 1476 846
rect 1510 822 1733 846
rect 1767 1109 1848 1143
rect 2103 1110 2137 1246
rect 2460 1212 2494 1246
rect 2639 1212 2664 1246
rect 2698 1212 2723 1246
rect 2845 1233 2861 1247
rect 2895 1233 2911 1267
rect 3157 1246 3214 1315
rect 2184 1178 2200 1212
rect 2234 1178 2282 1212
rect 2316 1178 2364 1212
rect 2398 1178 2414 1212
rect 2460 1178 2605 1212
rect 2759 1199 2809 1213
rect 3157 1212 3178 1246
rect 3212 1212 3214 1246
rect 2759 1194 3090 1199
rect 2184 1162 2414 1178
rect 2380 1144 2414 1162
rect 2571 1144 2725 1178
rect 2380 1110 2537 1144
rect 1767 907 1801 1109
rect 1882 1076 2137 1110
rect 2223 1090 2289 1096
rect 1882 1075 1916 1076
rect 1835 1059 1916 1075
rect 1835 1025 1851 1059
rect 1885 1025 1916 1059
rect 2223 1056 2239 1090
rect 2273 1076 2289 1090
rect 2273 1063 2469 1076
rect 2273 1056 2419 1063
rect 1835 991 1916 1025
rect 1835 957 1851 991
rect 1885 957 1916 991
rect 1950 1026 2081 1042
rect 1950 992 1966 1026
rect 2000 1016 2081 1026
rect 2223 1031 2419 1056
rect 2000 992 2047 1016
rect 1950 982 2047 992
rect 1950 976 2081 982
rect 2115 1000 2181 1016
rect 1835 941 1916 957
rect 2115 966 2131 1000
rect 2165 966 2181 1000
rect 2223 997 2239 1031
rect 2273 1029 2419 1031
rect 2453 1029 2469 1063
rect 2273 1016 2469 1029
rect 2273 997 2289 1016
rect 2223 981 2289 997
rect 2503 982 2537 1110
rect 2691 1106 2725 1144
rect 2793 1165 3090 1194
rect 2793 1160 2809 1165
rect 2759 1140 2809 1160
rect 3056 1131 3123 1165
rect 2913 1115 3022 1131
rect 2913 1106 2972 1115
rect 2583 1072 2657 1096
rect 2583 1038 2599 1072
rect 2633 1038 2657 1072
rect 2583 1016 2657 1038
rect 2691 1081 2972 1106
rect 3006 1081 3022 1115
rect 2691 1072 3022 1081
rect 2691 1038 2707 1072
rect 2741 1038 2757 1072
rect 2913 1065 3022 1072
rect 2691 1022 2757 1038
rect 2799 1022 2865 1038
rect 2583 982 2623 1016
rect 2799 988 2815 1022
rect 2849 988 2865 1022
rect 2115 942 2181 966
rect 1973 908 2181 942
rect 2340 948 2542 982
rect 2691 954 2865 988
rect 2691 948 2725 954
rect 2340 912 2374 948
rect 2508 914 2725 948
rect 2913 931 2947 1065
rect 3089 1046 3123 1131
rect 3157 1156 3214 1212
rect 3157 1122 3178 1156
rect 3212 1122 3214 1156
rect 3157 1106 3214 1122
rect 3248 1246 3314 1262
rect 3248 1212 3264 1246
rect 3298 1212 3314 1246
rect 3248 1156 3314 1212
rect 3248 1122 3264 1156
rect 3298 1122 3314 1156
rect 3248 1088 3314 1122
rect 3348 1246 3414 1315
rect 3348 1212 3350 1246
rect 3384 1212 3414 1246
rect 3566 1246 3632 1315
rect 3348 1156 3414 1212
rect 3348 1122 3350 1156
rect 3384 1122 3414 1156
rect 3348 1106 3414 1122
rect 3460 1220 3526 1224
rect 3460 1186 3476 1220
rect 3510 1186 3526 1220
rect 3460 1152 3526 1186
rect 3460 1118 3476 1152
rect 3510 1118 3526 1152
rect 3566 1212 3582 1246
rect 3616 1212 3632 1246
rect 3566 1172 3632 1212
rect 3566 1138 3582 1172
rect 3616 1138 3632 1172
rect 3566 1122 3632 1138
rect 3666 1246 3733 1262
rect 3666 1212 3682 1246
rect 3716 1212 3733 1246
rect 3666 1172 3733 1212
rect 3666 1138 3682 1172
rect 3716 1138 3733 1172
rect 3666 1122 3733 1138
rect 2981 1015 3047 1031
rect 2981 1014 2997 1015
rect 2981 980 2996 1014
rect 3031 981 3047 1015
rect 3030 980 3047 981
rect 2981 965 3047 980
rect 3089 1030 3155 1046
rect 3089 996 3105 1030
rect 3139 996 3155 1030
rect 3089 980 3155 996
rect 3267 1022 3314 1088
rect 3460 1088 3526 1118
rect 3460 1072 3665 1088
rect 3460 1038 3615 1072
rect 3649 1038 3665 1072
rect 3460 1022 3665 1038
rect 1973 907 2039 908
rect 1767 896 2039 907
rect 1767 873 1989 896
rect 1510 812 1526 822
rect 1460 785 1526 812
rect 1767 786 1801 873
rect 1973 862 1989 873
rect 2023 862 2039 896
rect 2253 896 2374 912
rect 1572 752 1588 786
rect 1622 752 1707 786
rect 1741 752 1801 786
rect 1865 823 1931 839
rect 1865 789 1881 823
rect 1915 789 1931 823
rect 1572 751 1757 752
rect 1269 717 1757 751
rect 1865 683 1931 789
rect 1973 786 2039 862
rect 1973 752 1989 786
rect 2023 752 2039 786
rect 1973 736 2039 752
rect 2085 858 2151 874
rect 2085 824 2101 858
rect 2135 824 2151 858
rect 2085 786 2151 824
rect 2085 752 2101 786
rect 2135 752 2151 786
rect 2085 683 2151 752
rect 2253 862 2269 896
rect 2303 878 2374 896
rect 2408 906 2474 914
rect 2303 862 2319 878
rect 2253 786 2319 862
rect 2408 872 2424 906
rect 2458 880 2474 906
rect 2829 904 2879 920
rect 2829 880 2845 904
rect 2458 872 2845 880
rect 2408 870 2845 872
rect 2408 864 2879 870
rect 2913 915 3007 931
rect 2913 881 2957 915
rect 2991 881 3007 915
rect 2913 865 3007 881
rect 2408 846 2569 864
rect 2553 830 2569 846
rect 2603 846 2879 864
rect 2603 830 2619 846
rect 2253 752 2269 786
rect 2303 752 2319 786
rect 2253 736 2319 752
rect 2438 791 2504 812
rect 2438 757 2454 791
rect 2488 757 2504 791
rect 2438 683 2504 757
rect 2553 786 2619 830
rect 2829 831 2879 846
rect 3089 831 3123 980
rect 3267 976 3335 1022
rect 3267 952 3317 976
rect 2553 752 2569 786
rect 2603 752 2619 786
rect 2553 736 2619 752
rect 2653 791 2719 812
rect 2653 757 2669 791
rect 2703 757 2719 791
rect 2653 683 2719 757
rect 2829 797 3123 831
rect 3157 919 3226 942
rect 3157 885 3176 919
rect 3210 885 3226 919
rect 3157 837 3226 885
rect 3157 803 3176 837
rect 3210 803 3226 837
rect 2829 786 2879 797
rect 2829 752 2845 786
rect 3157 763 3226 803
rect 2829 736 2879 752
rect 3048 747 3226 763
rect 3048 713 3064 747
rect 3098 713 3176 747
rect 3210 713 3226 747
rect 3267 918 3283 952
rect 3267 869 3317 918
rect 3267 835 3283 869
rect 3267 786 3317 835
rect 3267 752 3283 786
rect 3267 736 3317 752
rect 3357 926 3423 942
rect 3357 892 3373 926
rect 3407 892 3423 926
rect 3357 856 3423 892
rect 3357 822 3373 856
rect 3407 822 3423 856
rect 3357 786 3423 822
rect 3357 752 3373 786
rect 3407 752 3423 786
rect 3048 683 3226 713
rect 3357 683 3423 752
rect 3460 936 3532 1022
rect 3699 968 3733 1122
rect 3768 1246 3818 1315
rect 3802 1212 3818 1246
rect 3867 1250 4005 1315
rect 3867 1216 3883 1250
rect 3917 1216 3955 1250
rect 3989 1216 4005 1250
rect 4055 1246 4105 1262
rect 3768 1156 3818 1212
rect 3802 1122 3818 1156
rect 3768 1106 3818 1122
rect 4055 1212 4071 1246
rect 4055 1156 4105 1212
rect 4141 1224 4207 1315
rect 4141 1190 4157 1224
rect 4191 1190 4207 1224
rect 4141 1171 4207 1190
rect 4243 1246 4277 1262
rect 4055 1122 4071 1156
rect 4243 1156 4277 1212
rect 4313 1224 4379 1315
rect 4313 1190 4329 1224
rect 4363 1190 4379 1224
rect 4313 1171 4379 1190
rect 4415 1247 4873 1281
rect 4415 1246 4465 1247
rect 4449 1212 4465 1246
rect 4105 1122 4243 1130
rect 4415 1156 4465 1212
rect 4599 1224 4665 1247
rect 4277 1122 4415 1130
rect 4449 1122 4465 1156
rect 4055 1096 4465 1122
rect 4499 1192 4565 1210
rect 4499 1158 4515 1192
rect 4549 1158 4565 1192
rect 4599 1190 4615 1224
rect 4649 1190 4665 1224
rect 4807 1224 4873 1247
rect 4599 1171 4665 1190
rect 4699 1192 4773 1210
rect 4499 1130 4565 1158
rect 4699 1158 4719 1192
rect 4753 1158 4773 1192
rect 4807 1190 4823 1224
rect 4857 1190 4873 1224
rect 4807 1171 4873 1190
rect 4699 1130 4773 1158
rect 4499 1096 4871 1130
rect 4825 1080 4871 1096
rect 4134 1046 4487 1062
rect 4134 1012 4150 1046
rect 4184 1012 4218 1046
rect 4252 1012 4282 1046
rect 4320 1012 4354 1046
rect 4388 1012 4487 1046
rect 4134 996 4487 1012
rect 4249 976 4487 996
rect 4521 1046 4791 1062
rect 4521 1012 4537 1046
rect 4571 1012 4605 1046
rect 4639 1012 4669 1046
rect 4707 1012 4741 1046
rect 4775 1012 4791 1046
rect 4521 976 4791 1012
rect 4825 1000 4940 1080
rect 3460 902 3482 936
rect 3516 902 3532 936
rect 3460 865 3532 902
rect 3460 831 3482 865
rect 3516 831 3532 865
rect 3460 794 3532 831
rect 3460 760 3482 794
rect 3516 760 3532 794
rect 3460 744 3532 760
rect 3571 940 3637 968
rect 3571 906 3587 940
rect 3621 906 3637 940
rect 3571 868 3637 906
rect 3571 834 3587 868
rect 3621 834 3637 868
rect 3571 790 3637 834
rect 3571 756 3587 790
rect 3621 756 3637 790
rect 3571 683 3637 756
rect 3671 952 3733 968
rect 3671 918 3677 952
rect 3711 943 3733 952
rect 3671 909 3680 918
rect 3714 909 3733 943
rect 3671 871 3733 909
rect 3671 869 3680 871
rect 3671 835 3677 869
rect 3714 837 3733 871
rect 3711 835 3733 837
rect 3671 786 3733 835
rect 3671 752 3677 786
rect 3711 752 3733 786
rect 3671 736 3733 752
rect 3767 952 3817 968
rect 3801 918 3817 952
rect 3767 869 3817 918
rect 3801 835 3817 869
rect 3767 786 3817 835
rect 3801 752 3817 786
rect 4055 946 4121 962
rect 4055 912 4071 946
rect 4105 912 4121 946
rect 4825 942 4871 1000
rect 4055 866 4121 912
rect 4055 832 4071 866
rect 4105 832 4121 866
rect 4055 786 4121 832
rect 3767 683 3817 752
rect 3867 748 3883 782
rect 3917 748 3955 782
rect 3989 748 4005 782
rect 3867 683 4005 748
rect 4055 752 4071 786
rect 4105 752 4121 786
rect 4055 683 4121 752
rect 4155 926 4871 942
rect 4155 892 4162 926
rect 4196 892 4242 926
rect 4276 892 4324 926
rect 4358 908 4514 926
rect 4358 892 4364 908
rect 4155 855 4364 892
rect 4498 892 4514 908
rect 4548 892 4583 926
rect 4617 892 4654 926
rect 4688 892 4723 926
rect 4757 908 4871 926
rect 4757 892 4773 908
rect 4155 821 4162 855
rect 4196 821 4242 855
rect 4276 821 4324 855
rect 4358 821 4364 855
rect 4155 786 4364 821
rect 4155 752 4162 786
rect 4196 752 4242 786
rect 4276 752 4324 786
rect 4358 752 4364 786
rect 4155 736 4364 752
rect 4398 865 4464 874
rect 4398 831 4414 865
rect 4448 831 4464 865
rect 4398 786 4464 831
rect 4398 752 4414 786
rect 4448 752 4464 786
rect 4398 683 4464 752
rect 4498 855 4773 892
rect 4498 821 4514 855
rect 4548 821 4583 855
rect 4617 821 4654 855
rect 4688 821 4723 855
rect 4757 821 4773 855
rect 4498 786 4773 821
rect 4498 752 4514 786
rect 4548 752 4583 786
rect 4617 752 4654 786
rect 4688 752 4723 786
rect 4757 752 4773 786
rect 4498 736 4773 752
rect 4807 865 4873 874
rect 4807 831 4823 865
rect 4857 831 4873 865
rect 4807 786 4873 831
rect 4807 752 4823 786
rect 4857 752 4873 786
rect 4807 683 4873 752
rect -2880 649 -2849 683
rect -2815 649 -2753 683
rect -2719 649 -2657 683
rect -2623 649 -2561 683
rect -2527 649 -2465 683
rect -2431 649 -2369 683
rect -2335 649 -2273 683
rect -2239 649 -2177 683
rect -2143 649 -2081 683
rect -2047 649 -1985 683
rect -1951 649 -1889 683
rect -1855 649 -1793 683
rect -1759 649 -1697 683
rect -1663 649 -1601 683
rect -1567 649 -1505 683
rect -1471 649 -1409 683
rect -1375 649 -1313 683
rect -1279 649 -1217 683
rect -1183 649 -1121 683
rect -1087 649 -1025 683
rect -991 649 -929 683
rect -895 649 -833 683
rect -799 649 -737 683
rect -703 649 -641 683
rect -607 649 -545 683
rect -511 649 -449 683
rect -415 649 -353 683
rect -319 649 -257 683
rect -223 649 -161 683
rect -127 649 -65 683
rect -31 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 257 649 319 683
rect 353 649 415 683
rect 449 649 511 683
rect 545 649 607 683
rect 641 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1471 683
rect 1505 649 1567 683
rect 1601 649 1663 683
rect 1697 649 1759 683
rect 1793 649 1855 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 2657 649 2719 683
rect 2753 649 2815 683
rect 2849 649 2911 683
rect 2945 649 3007 683
rect 3041 649 3103 683
rect 3137 649 3199 683
rect 3233 649 3295 683
rect 3329 649 3391 683
rect 3425 649 3487 683
rect 3521 649 3583 683
rect 3617 649 3679 683
rect 3713 649 3775 683
rect 3809 649 3871 683
rect 3905 649 3967 683
rect 4001 649 4063 683
rect 4097 649 4159 683
rect 4193 649 4255 683
rect 4289 649 4351 683
rect 4385 649 4447 683
rect 4481 649 4543 683
rect 4577 649 4639 683
rect 4673 649 4735 683
rect 4769 649 4831 683
rect 4865 649 4896 683
rect -1631 580 -1565 649
rect -1631 546 -1615 580
rect -1581 546 -1565 580
rect -1631 510 -1565 546
rect -1631 476 -1615 510
rect -1581 476 -1565 510
rect -1631 440 -1565 476
rect -1631 406 -1615 440
rect -1581 406 -1565 440
rect -1631 390 -1565 406
rect -1531 580 -1465 596
rect -1531 546 -1515 580
rect -1481 546 -1465 580
rect -1531 497 -1465 546
rect -1531 463 -1515 497
rect -1481 463 -1465 497
rect -1531 414 -1465 463
rect -267 580 -201 649
rect -267 546 -251 580
rect -217 546 -201 580
rect -267 497 -201 546
rect -267 463 -251 497
rect -217 463 -201 497
rect -1531 380 -1515 414
rect -1481 380 -1465 414
rect -1703 310 -1565 356
rect -1703 276 -1687 310
rect -1649 276 -1615 310
rect -1581 276 -1565 310
rect -1703 260 -1565 276
rect -1531 327 -1465 380
rect -1531 268 -1364 327
rect -1631 210 -1565 226
rect -1631 176 -1615 210
rect -1581 176 -1565 210
rect -1631 120 -1565 176
rect -1631 86 -1615 120
rect -1581 86 -1565 120
rect -1631 17 -1565 86
rect -1531 210 -1465 268
rect -1531 176 -1515 210
rect -1481 176 -1465 210
rect -1531 120 -1465 176
rect -267 414 -201 463
rect -267 380 -251 414
rect -217 380 -201 414
rect -267 364 -201 380
rect -167 580 -121 596
rect -167 546 -161 580
rect -127 546 -121 580
rect -167 497 -121 546
rect -167 463 -161 497
rect -127 463 -121 497
rect -167 414 -121 463
rect -167 380 -161 414
rect -127 380 -121 414
rect -400 294 -201 310
rect -400 260 -251 294
rect -217 260 -201 294
rect -400 244 -201 260
rect -267 236 -201 244
rect -167 236 -121 380
rect -87 580 -21 649
rect -87 546 -71 580
rect -37 546 -21 580
rect -87 497 -21 546
rect -87 463 -71 497
rect -37 463 -21 497
rect -87 414 -21 463
rect 18 578 174 613
rect 18 544 31 578
rect 65 544 127 578
rect 18 538 127 544
rect 161 538 174 578
rect 18 492 174 538
rect 18 458 31 492
rect 65 458 127 492
rect 161 458 174 492
rect 215 580 265 596
rect 215 546 231 580
rect 215 511 265 546
rect 305 579 371 649
rect 305 545 321 579
rect 355 545 371 579
rect 305 529 371 545
rect 405 581 629 615
rect 215 477 231 511
rect 405 495 439 581
rect 563 580 629 581
rect 265 477 439 495
rect 215 461 439 477
rect 473 520 523 547
rect 473 486 489 520
rect 473 460 523 486
rect 563 546 579 580
rect 613 546 629 580
rect 563 510 629 546
rect 563 476 579 510
rect 613 476 629 510
rect 563 460 629 476
rect 675 580 741 649
rect 675 546 691 580
rect 725 546 741 580
rect 675 510 741 546
rect 675 476 691 510
rect 725 476 741 510
rect 675 460 741 476
rect 781 580 831 596
rect 815 546 831 580
rect 781 510 831 546
rect 815 476 831 510
rect 18 442 174 458
rect -87 380 -71 414
rect -37 380 -21 414
rect -87 364 -21 380
rect 217 411 302 427
rect 217 377 252 411
rect 286 377 302 411
rect 489 426 523 460
rect 489 392 623 426
rect 217 343 302 377
rect -87 294 -21 310
rect -87 260 -71 294
rect -37 260 -21 294
rect -87 236 -21 260
rect 217 309 252 343
rect 286 309 302 343
rect 217 292 302 309
rect 353 343 455 359
rect 353 309 369 343
rect 403 309 455 343
rect 353 292 455 309
rect 489 342 555 358
rect 489 308 505 342
rect 539 308 555 342
rect 489 292 555 308
rect 217 275 455 292
rect 217 241 252 275
rect 286 241 369 275
rect 403 241 455 275
rect 589 258 623 392
rect 781 362 831 476
rect 877 580 927 596
rect 877 546 893 580
rect 877 510 927 546
rect 877 476 893 510
rect 877 440 927 476
rect 967 580 1033 649
rect 967 546 983 580
rect 1017 546 1033 580
rect 967 502 1033 546
rect 967 468 983 502
rect 1017 468 1033 502
rect 967 458 1033 468
rect 1073 580 1149 596
rect 1107 546 1149 580
rect 1073 499 1149 546
rect 1107 465 1149 499
rect 1185 528 1235 649
rect 1219 494 1235 528
rect 1185 470 1235 494
rect 1269 581 1757 615
rect 877 406 893 440
rect 927 406 1039 424
rect 877 390 1039 406
rect 713 346 831 362
rect 713 312 729 346
rect 763 312 831 346
rect 713 296 831 312
rect -155 202 -121 236
rect 217 225 455 241
rect 18 205 174 221
rect -262 168 -246 202
rect -212 168 -196 202
rect -155 168 -82 202
rect -48 168 -32 202
rect -1531 86 -1515 120
rect -1481 86 -1465 120
rect -1531 70 -1465 86
rect -262 120 -196 168
rect -262 86 -246 120
rect -212 86 -196 120
rect -262 17 -196 86
rect -98 126 -32 168
rect -98 120 -81 126
rect -98 86 -82 120
rect -47 92 -32 126
rect -48 86 -32 92
rect -98 70 -32 86
rect 18 171 31 205
rect 65 171 127 205
rect 161 171 174 205
rect 18 128 174 171
rect 18 88 31 128
rect 65 122 174 128
rect 65 88 127 122
rect 161 88 174 122
rect 18 53 174 88
rect 220 170 286 225
rect 489 224 746 258
rect 489 191 530 224
rect 220 136 236 170
rect 270 136 286 170
rect 220 17 286 136
rect 384 175 530 191
rect 384 141 400 175
rect 434 141 480 175
rect 514 141 530 175
rect 384 125 530 141
rect 628 169 678 190
rect 628 135 644 169
rect 628 17 678 135
rect 712 85 746 224
rect 780 180 831 296
rect 889 320 971 356
rect 889 286 921 320
rect 955 286 971 320
rect 889 270 971 286
rect 1005 334 1039 390
rect 1073 418 1149 465
rect 1269 436 1303 581
rect 1572 580 1757 581
rect 1107 384 1149 418
rect 1073 368 1149 384
rect 1005 318 1081 334
rect 1005 284 1031 318
rect 1065 284 1081 318
rect 1005 268 1081 284
rect 1115 270 1149 368
rect 1199 416 1303 436
rect 1199 382 1215 416
rect 1249 402 1303 416
rect 1360 520 1426 547
rect 1360 486 1376 520
rect 1410 486 1426 520
rect 1360 442 1426 486
rect 1460 520 1526 547
rect 1572 546 1588 580
rect 1622 546 1707 580
rect 1741 546 1801 580
rect 1460 486 1476 520
rect 1510 510 1526 520
rect 1510 486 1733 510
rect 1460 476 1733 486
rect 1360 408 1665 442
rect 1249 382 1265 402
rect 1199 366 1265 382
rect 1599 375 1665 408
rect 1491 368 1557 371
rect 1311 355 1557 368
rect 1311 352 1507 355
rect 1311 318 1327 352
rect 1361 321 1507 352
rect 1541 321 1557 355
rect 1361 318 1557 321
rect 1311 305 1557 318
rect 1599 341 1615 375
rect 1649 341 1665 375
rect 1599 307 1665 341
rect 1311 276 1415 305
rect 1311 270 1375 276
rect 1005 234 1039 268
rect 1115 242 1375 270
rect 1409 242 1415 276
rect 1599 273 1615 307
rect 1649 273 1665 307
rect 1599 271 1665 273
rect 1115 237 1415 242
rect 1115 236 1146 237
rect 876 200 892 234
rect 926 200 1039 234
rect 1130 203 1146 236
rect 1180 236 1415 237
rect 1449 237 1665 271
rect 814 146 831 180
rect 1130 169 1180 203
rect 780 119 831 146
rect 865 132 1096 166
rect 865 85 899 132
rect 712 51 899 85
rect 978 82 1028 98
rect 978 48 994 82
rect 1062 85 1096 132
rect 1130 135 1146 169
rect 1130 119 1180 135
rect 1214 168 1415 202
rect 1214 85 1248 168
rect 1062 51 1248 85
rect 1282 118 1336 134
rect 1282 84 1284 118
rect 1318 84 1336 118
rect 978 17 1028 48
rect 1282 17 1336 84
rect 1381 87 1415 168
rect 1449 184 1515 237
rect 1699 203 1733 476
rect 1449 150 1465 184
rect 1499 150 1515 184
rect 1449 121 1515 150
rect 1549 179 1733 203
rect 1767 459 1801 546
rect 1865 543 1931 649
rect 1865 509 1881 543
rect 1915 509 1931 543
rect 1865 493 1931 509
rect 1973 580 2039 596
rect 1973 546 1989 580
rect 2023 546 2039 580
rect 1973 470 2039 546
rect 1973 459 1989 470
rect 1767 436 1989 459
rect 2023 436 2039 470
rect 2085 580 2151 649
rect 2085 546 2101 580
rect 2135 546 2151 580
rect 2085 508 2151 546
rect 2085 474 2101 508
rect 2135 474 2151 508
rect 2085 458 2151 474
rect 2253 580 2319 596
rect 2253 546 2269 580
rect 2303 546 2319 580
rect 2253 470 2319 546
rect 2438 575 2504 649
rect 2438 541 2454 575
rect 2488 541 2504 575
rect 2438 520 2504 541
rect 2553 580 2619 596
rect 2553 546 2569 580
rect 2603 546 2619 580
rect 2553 502 2619 546
rect 2653 575 2719 649
rect 3048 619 3226 649
rect 2653 541 2669 575
rect 2703 541 2719 575
rect 2653 520 2719 541
rect 2829 580 2879 596
rect 2829 546 2845 580
rect 3048 585 3064 619
rect 3098 585 3176 619
rect 3210 585 3226 619
rect 3048 569 3226 585
rect 2829 535 2879 546
rect 2553 486 2569 502
rect 1767 425 2039 436
rect 1767 223 1801 425
rect 1973 424 2039 425
rect 2253 436 2269 470
rect 2303 454 2319 470
rect 2408 468 2569 486
rect 2603 486 2619 502
rect 2829 501 3123 535
rect 2829 486 2879 501
rect 2603 468 2879 486
rect 2408 462 2879 468
rect 2408 460 2845 462
rect 2303 436 2374 454
rect 1835 375 1916 391
rect 1973 390 2181 424
rect 2253 420 2374 436
rect 1835 341 1851 375
rect 1885 341 1916 375
rect 2115 366 2181 390
rect 1835 307 1916 341
rect 1835 273 1851 307
rect 1885 273 1916 307
rect 1950 350 2081 356
rect 1950 340 2047 350
rect 1950 306 1966 340
rect 2000 316 2047 340
rect 2115 332 2131 366
rect 2165 332 2181 366
rect 2340 384 2374 420
rect 2408 426 2424 460
rect 2458 452 2845 460
rect 2458 426 2474 452
rect 2408 418 2474 426
rect 2829 428 2845 452
rect 2508 384 2725 418
rect 2829 412 2879 428
rect 2913 451 3007 467
rect 2913 417 2957 451
rect 2991 417 3007 451
rect 2115 316 2181 332
rect 2223 335 2289 351
rect 2340 350 2542 384
rect 2691 378 2725 384
rect 2913 401 3007 417
rect 2000 306 2081 316
rect 1950 290 2081 306
rect 2223 301 2239 335
rect 2273 316 2289 335
rect 2273 303 2469 316
rect 2273 301 2419 303
rect 1835 257 1916 273
rect 1882 256 1916 257
rect 2223 276 2419 301
rect 1767 189 1848 223
rect 1882 222 2137 256
rect 2223 242 2239 276
rect 2273 269 2419 276
rect 2453 269 2469 303
rect 2273 256 2469 269
rect 2273 242 2289 256
rect 2223 236 2289 242
rect 2503 222 2537 350
rect 2583 316 2623 350
rect 2691 344 2865 378
rect 2583 294 2657 316
rect 2799 310 2815 344
rect 2849 310 2865 344
rect 2583 260 2599 294
rect 2633 260 2657 294
rect 2583 236 2657 260
rect 2691 294 2757 310
rect 2799 294 2865 310
rect 2691 260 2707 294
rect 2741 260 2757 294
rect 2913 267 2947 401
rect 2981 353 3047 367
rect 2981 351 2998 353
rect 2981 317 2997 351
rect 3032 319 3047 353
rect 3031 317 3047 319
rect 2981 301 3047 317
rect 3089 352 3123 501
rect 3157 529 3226 569
rect 3157 495 3176 529
rect 3210 495 3226 529
rect 3267 580 3317 596
rect 3267 546 3283 580
rect 3267 505 3317 546
rect 3157 447 3226 495
rect 3157 413 3176 447
rect 3210 413 3226 447
rect 3157 390 3226 413
rect 3265 497 3317 505
rect 3265 490 3283 497
rect 3265 456 3274 490
rect 3308 456 3317 463
rect 3265 418 3317 456
rect 3265 384 3274 418
rect 3308 414 3317 418
rect 3357 580 3423 649
rect 3357 546 3373 580
rect 3407 546 3423 580
rect 3357 510 3423 546
rect 3357 476 3373 510
rect 3407 476 3423 510
rect 3357 440 3423 476
rect 3357 406 3373 440
rect 3407 406 3423 440
rect 3357 390 3423 406
rect 3460 572 3532 588
rect 3460 538 3482 572
rect 3516 538 3532 572
rect 3460 501 3532 538
rect 3460 467 3482 501
rect 3516 467 3532 501
rect 3460 430 3532 467
rect 3460 396 3482 430
rect 3516 396 3532 430
rect 3265 380 3283 384
rect 3265 369 3317 380
rect 3267 356 3317 369
rect 3089 336 3155 352
rect 3089 302 3105 336
rect 3139 302 3155 336
rect 3089 286 3155 302
rect 3267 310 3335 356
rect 3460 310 3532 396
rect 3571 576 3637 649
rect 3571 542 3587 576
rect 3621 542 3637 576
rect 3571 498 3637 542
rect 3571 464 3587 498
rect 3621 464 3637 498
rect 3571 426 3637 464
rect 3571 392 3587 426
rect 3621 392 3637 426
rect 3571 364 3637 392
rect 3671 580 3733 596
rect 3671 546 3677 580
rect 3711 546 3733 580
rect 3671 497 3733 546
rect 3671 463 3677 497
rect 3711 486 3733 497
rect 3671 452 3683 463
rect 3717 452 3733 486
rect 3671 414 3733 452
rect 3671 380 3677 414
rect 3717 380 3733 414
rect 3671 364 3733 380
rect 3767 580 3817 649
rect 3801 546 3817 580
rect 3867 584 4005 649
rect 3867 550 3883 584
rect 3917 550 3955 584
rect 3989 550 4005 584
rect 4056 565 4122 649
rect 3767 497 3817 546
rect 3801 463 3817 497
rect 3767 414 3817 463
rect 3801 380 3817 414
rect 4056 531 4072 565
rect 4106 531 4122 565
rect 4056 455 4122 531
rect 4056 421 4072 455
rect 4106 421 4122 455
rect 4056 405 4122 421
rect 4162 565 4196 581
rect 4162 455 4196 531
rect 4236 568 4302 649
rect 4236 534 4252 568
rect 4286 534 4302 568
rect 4236 500 4302 534
rect 4236 466 4252 500
rect 4286 466 4302 500
rect 4236 458 4302 466
rect 4336 565 4402 581
rect 4336 531 4352 565
rect 4386 531 4402 565
rect 4336 455 4402 531
rect 4443 580 4509 649
rect 4443 546 4459 580
rect 4493 546 4509 580
rect 4443 508 4509 546
rect 4443 474 4459 508
rect 4493 474 4509 508
rect 4443 458 4509 474
rect 4553 580 4603 596
rect 4587 546 4603 580
rect 4553 499 4603 546
rect 4587 465 4603 499
rect 4336 424 4352 455
rect 4196 421 4352 424
rect 4386 424 4402 455
rect 4386 421 4519 424
rect 3767 364 3817 380
rect 4162 390 4519 421
rect 2913 260 3022 267
rect 2691 251 3022 260
rect 1549 145 1565 179
rect 1599 169 1733 179
rect 1599 145 1615 169
rect 1549 87 1615 145
rect 1782 155 1798 189
rect 1832 155 1848 189
rect 1381 53 1615 87
rect 1661 119 1746 135
rect 1782 121 1848 155
rect 1882 171 1969 187
rect 1882 137 1908 171
rect 1942 137 1969 171
rect 1882 121 1969 137
rect 2003 171 2069 188
rect 2003 137 2019 171
rect 2053 137 2069 171
rect 1661 85 1686 119
rect 1720 87 1746 119
rect 1882 87 1916 121
rect 1720 85 1916 87
rect 1661 53 1916 85
rect 2003 17 2069 137
rect 2103 86 2137 222
rect 2380 188 2537 222
rect 2691 226 2972 251
rect 2691 188 2725 226
rect 2913 217 2972 226
rect 3006 217 3022 251
rect 2913 201 3022 217
rect 3089 201 3123 286
rect 3267 244 3314 310
rect 2380 170 2414 188
rect 2184 154 2414 170
rect 2571 154 2725 188
rect 2759 172 2809 192
rect 2184 120 2200 154
rect 2234 120 2282 154
rect 2316 120 2364 154
rect 2398 120 2414 154
rect 2460 120 2605 154
rect 2793 167 2809 172
rect 3056 167 3123 201
rect 3157 210 3214 226
rect 3157 176 3178 210
rect 3212 176 3214 210
rect 2793 138 3090 167
rect 2759 133 3090 138
rect 2460 86 2494 120
rect 2639 86 2664 120
rect 2698 86 2723 120
rect 2759 119 2809 133
rect 3157 120 3214 176
rect 2103 52 2494 86
rect 2528 52 2548 86
rect 2582 52 2603 86
rect 2528 17 2603 52
rect 2639 85 2723 86
rect 2845 85 2861 99
rect 2639 65 2861 85
rect 2895 65 2911 99
rect 2639 51 2911 65
rect 3157 86 3178 120
rect 3212 86 3214 120
rect 3157 17 3214 86
rect 3248 210 3314 244
rect 3460 294 3665 310
rect 3460 260 3615 294
rect 3649 260 3665 294
rect 3460 244 3665 260
rect 3248 176 3264 210
rect 3298 176 3314 210
rect 3248 120 3314 176
rect 3248 86 3264 120
rect 3298 86 3314 120
rect 3248 70 3314 86
rect 3348 210 3414 226
rect 3348 176 3350 210
rect 3384 176 3414 210
rect 3348 120 3414 176
rect 3348 86 3350 120
rect 3384 86 3414 120
rect 3460 214 3526 244
rect 3460 180 3476 214
rect 3510 180 3526 214
rect 3699 210 3733 364
rect 4162 256 4196 390
rect 4245 341 4311 356
rect 4245 340 4262 341
rect 4245 306 4261 340
rect 4296 307 4311 341
rect 4295 306 4311 307
rect 4245 290 4311 306
rect 4345 343 4445 356
rect 4345 334 4450 343
rect 4345 300 4387 334
rect 4421 319 4450 334
rect 4345 285 4395 300
rect 4429 291 4450 319
rect 4485 335 4519 390
rect 4553 419 4603 465
rect 4643 580 4693 649
rect 4677 546 4693 580
rect 4643 487 4693 546
rect 4677 453 4693 487
rect 4643 437 4693 453
rect 4733 580 4787 596
rect 4767 546 4787 580
rect 4733 499 4787 546
rect 4767 465 4787 499
rect 4587 403 4603 419
rect 4733 419 4787 465
rect 4587 385 4733 403
rect 4767 385 4787 419
rect 4553 369 4787 385
rect 4485 319 4695 335
rect 4429 285 4445 291
rect 4345 269 4445 285
rect 4485 285 4509 319
rect 4543 285 4577 319
rect 4611 285 4645 319
rect 4679 285 4695 319
rect 4729 327 4787 369
rect 4823 580 4873 649
rect 4857 546 4873 580
rect 4823 497 4873 546
rect 4857 463 4873 497
rect 4823 414 4873 463
rect 4857 380 4873 414
rect 4823 364 4873 380
rect 4916 327 4974 345
rect 4729 310 4974 327
rect 4485 269 4695 285
rect 4737 287 4974 310
rect 4055 235 4121 251
rect 3460 146 3526 180
rect 3460 112 3476 146
rect 3510 112 3526 146
rect 3460 108 3526 112
rect 3566 194 3632 210
rect 3566 160 3582 194
rect 3616 160 3632 194
rect 3566 120 3632 160
rect 3348 17 3414 86
rect 3566 86 3582 120
rect 3616 86 3632 120
rect 3566 17 3632 86
rect 3666 194 3733 210
rect 3666 160 3682 194
rect 3716 160 3733 194
rect 3666 120 3733 160
rect 3666 86 3682 120
rect 3716 86 3733 120
rect 3666 70 3733 86
rect 3768 210 3818 226
rect 3802 176 3818 210
rect 3768 120 3818 176
rect 3802 86 3818 120
rect 4055 201 4071 235
rect 4105 201 4121 235
rect 4162 239 4297 256
rect 4162 222 4247 239
rect 4055 165 4121 201
rect 4231 205 4247 222
rect 4281 205 4297 239
rect 4737 235 4787 287
rect 4916 265 4974 287
rect 4055 131 4071 165
rect 4105 131 4121 165
rect 3768 17 3818 86
rect 3867 82 3883 116
rect 3917 82 3955 116
rect 3989 82 4005 116
rect 3867 17 4005 82
rect 4055 17 4121 131
rect 4161 168 4195 188
rect 4161 85 4195 134
rect 4231 161 4297 205
rect 4231 127 4247 161
rect 4281 127 4297 161
rect 4231 119 4297 127
rect 4331 229 4397 235
rect 4331 195 4347 229
rect 4381 195 4397 229
rect 4331 161 4397 195
rect 4331 127 4347 161
rect 4381 127 4397 161
rect 4331 85 4397 127
rect 4161 51 4397 85
rect 4433 201 4449 235
rect 4483 201 4499 235
rect 4433 157 4499 201
rect 4433 123 4449 157
rect 4483 123 4499 157
rect 4433 17 4499 123
rect 4551 219 4737 235
rect 4585 201 4737 219
rect 4771 201 4787 235
rect 4585 185 4601 201
rect 4551 145 4601 185
rect 4585 111 4601 145
rect 4551 95 4601 111
rect 4635 151 4701 167
rect 4635 117 4651 151
rect 4685 117 4701 151
rect 4635 17 4701 117
rect 4737 145 4787 201
rect 4771 111 4787 145
rect 4737 95 4787 111
rect 4823 235 4873 251
rect 4857 201 4873 235
rect 4823 145 4873 201
rect 4857 111 4873 145
rect 4823 17 4873 111
rect -1728 -17 -1697 17
rect -1663 -17 -1601 17
rect -1567 -17 -1505 17
rect -1471 -17 -1409 17
rect -1375 -17 -1313 17
rect -1279 -17 -1217 17
rect -1183 -17 -1121 17
rect -1087 -17 -1025 17
rect -991 -17 -929 17
rect -895 -17 -833 17
rect -799 -17 -737 17
rect -703 -17 -641 17
rect -607 -17 -545 17
rect -511 -17 -449 17
rect -415 -17 -353 17
rect -319 -17 -257 17
rect -223 -17 -161 17
rect -127 -17 -65 17
rect -31 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3583 17
rect 3617 -17 3679 17
rect 3713 -17 3775 17
rect 3809 -17 3871 17
rect 3905 -17 3967 17
rect 4001 -17 4063 17
rect 4097 -17 4159 17
rect 4193 -17 4255 17
rect 4289 -17 4351 17
rect 4385 -17 4447 17
rect 4481 -17 4543 17
rect 4577 -17 4639 17
rect 4673 -17 4735 17
rect 4769 -17 4831 17
rect 4865 -17 4896 17
rect -1537 -158 -1407 -124
rect -1249 -158 -1153 -124
rect -1537 -220 -1469 -158
rect -1537 -776 -1503 -220
rect -1187 -220 -1153 -158
rect -1389 -310 -1355 -294
rect -1389 -702 -1355 -686
rect -1301 -310 -1267 -294
rect -1301 -702 -1267 -686
rect -1361 -770 -1345 -736
rect -1311 -770 -1295 -736
rect -1537 -838 -1469 -776
rect -1187 -838 -1153 -776
rect -1537 -872 -1407 -838
rect -1249 -872 -1153 -838
rect -1537 -934 -1469 -872
rect -1537 -1490 -1503 -934
rect -1187 -934 -1153 -872
rect -1389 -1024 -1355 -1008
rect -1389 -1416 -1355 -1400
rect -1301 -1024 -1267 -1008
rect -1301 -1416 -1267 -1400
rect -1361 -1484 -1345 -1450
rect -1311 -1484 -1295 -1450
rect -1537 -1552 -1469 -1490
rect -1187 -1552 -1153 -1490
rect -1537 -1586 -1407 -1552
rect -1249 -1586 -1153 -1552
<< viali >>
rect -1738 3084 -1704 3460
rect -1650 3084 -1616 3460
rect -1536 3078 -1502 3466
rect -1694 3000 -1660 3034
rect -1738 2370 -1704 2746
rect -1650 2370 -1616 2746
rect -1536 2364 -1502 2752
rect -1694 2286 -1660 2320
rect -1070 3078 -1036 3466
rect -956 3084 -922 3460
rect -868 3084 -834 3460
rect -912 3000 -878 3034
rect -1070 2364 -1036 2752
rect -956 2370 -922 2746
rect -868 2370 -834 2746
rect -912 2286 -878 2320
rect -2849 1981 -2815 2015
rect -2753 1981 -2719 2015
rect -2657 1981 -2623 2015
rect -2561 1981 -2527 2015
rect -2465 1981 -2431 2015
rect -2369 1981 -2335 2015
rect -2273 1981 -2239 2015
rect -2177 1981 -2143 2015
rect -2081 1981 -2047 2015
rect -1985 1981 -1951 2015
rect -1889 1981 -1855 2015
rect -1793 1981 -1759 2015
rect -1697 1981 -1663 2015
rect -1601 1981 -1567 2015
rect -1505 1981 -1471 2015
rect -1409 1981 -1375 2015
rect -1313 1981 -1279 2015
rect -1217 1981 -1183 2015
rect -1121 1981 -1087 2015
rect -1025 1981 -991 2015
rect -929 1981 -895 2015
rect -833 1981 -799 2015
rect -737 1981 -703 2015
rect -641 1981 -607 2015
rect -545 1981 -511 2015
rect -449 1981 -415 2015
rect -353 1981 -319 2015
rect -257 1981 -223 2015
rect -161 1981 -127 2015
rect -65 1981 -31 2015
rect 31 1981 65 2015
rect 127 1981 161 2015
rect 223 1981 257 2015
rect 319 1981 353 2015
rect 415 1981 449 2015
rect 511 1981 545 2015
rect 607 1981 641 2015
rect 703 1981 737 2015
rect 799 1981 833 2015
rect 895 1981 929 2015
rect 991 1981 1025 2015
rect 1087 1981 1121 2015
rect 1183 1981 1217 2015
rect 1279 1981 1313 2015
rect 1375 1981 1409 2015
rect 1471 1981 1505 2015
rect 1567 1981 1601 2015
rect 1663 1981 1697 2015
rect 1759 1981 1793 2015
rect 1855 1981 1889 2015
rect 1951 1981 1985 2015
rect 2047 1981 2081 2015
rect 2143 1981 2177 2015
rect 2239 1981 2273 2015
rect 2335 1981 2369 2015
rect 2431 1981 2465 2015
rect 2527 1981 2561 2015
rect 2623 1981 2657 2015
rect 2719 1981 2753 2015
rect 2815 1981 2849 2015
rect 2911 1981 2945 2015
rect 3007 1981 3041 2015
rect 3103 1981 3137 2015
rect 3199 1981 3233 2015
rect 3295 1981 3329 2015
rect 3391 1981 3425 2015
rect 3487 1981 3521 2015
rect 3583 1981 3617 2015
rect 3679 1981 3713 2015
rect 3775 1981 3809 2015
rect 3871 1981 3905 2015
rect 3967 1981 4001 2015
rect 4063 1981 4097 2015
rect 4159 1981 4193 2015
rect 4255 1981 4289 2015
rect 4351 1981 4385 2015
rect 4447 1981 4481 2015
rect 4543 1981 4577 2015
rect 4639 1981 4673 2015
rect 4735 1981 4769 2015
rect 4831 1981 4865 2015
rect -2839 1608 -2835 1642
rect -2835 1608 -2805 1642
rect -2767 1608 -2733 1642
rect -2498 1483 -2101 1733
rect -1967 1483 -1570 1733
rect -1223 1592 -1189 1626
rect -1233 1452 -1199 1458
rect -1233 1424 -1200 1452
rect -1200 1424 -1199 1452
rect 127 1876 161 1904
rect 127 1870 161 1876
rect 31 1454 65 1460
rect 31 1426 65 1454
rect -2849 1315 -2815 1349
rect -2753 1315 -2719 1349
rect -2657 1315 -2623 1349
rect -2561 1315 -2527 1349
rect -2465 1315 -2431 1349
rect -2369 1315 -2335 1349
rect -2273 1315 -2239 1349
rect -2177 1315 -2143 1349
rect -2081 1315 -2047 1349
rect -1985 1315 -1951 1349
rect -1889 1315 -1855 1349
rect -1793 1315 -1759 1349
rect -1697 1315 -1663 1349
rect -1601 1315 -1567 1349
rect -1505 1315 -1471 1349
rect -1409 1315 -1375 1349
rect -1313 1315 -1279 1349
rect -1217 1315 -1183 1349
rect -1121 1315 -1087 1349
rect -1025 1315 -991 1349
rect -929 1315 -895 1349
rect -833 1315 -799 1349
rect -737 1315 -703 1349
rect -641 1315 -607 1349
rect -545 1315 -511 1349
rect -449 1315 -415 1349
rect -353 1315 -319 1349
rect -257 1315 -223 1349
rect -161 1315 -127 1349
rect -65 1315 -31 1349
rect 31 1315 65 1349
rect 127 1315 161 1349
rect 223 1315 257 1349
rect 319 1315 353 1349
rect 415 1315 449 1349
rect 511 1315 545 1349
rect 607 1315 641 1349
rect 703 1315 737 1349
rect 799 1315 833 1349
rect 895 1315 929 1349
rect 991 1315 1025 1349
rect 1087 1315 1121 1349
rect 1183 1315 1217 1349
rect 1279 1315 1313 1349
rect 1375 1315 1409 1349
rect 1471 1315 1505 1349
rect 1567 1315 1601 1349
rect 1663 1315 1697 1349
rect 1759 1315 1793 1349
rect 1855 1315 1889 1349
rect 1951 1315 1985 1349
rect 2047 1315 2081 1349
rect 2143 1315 2177 1349
rect 2239 1315 2273 1349
rect 2335 1315 2369 1349
rect 2431 1315 2465 1349
rect 2527 1315 2561 1349
rect 2623 1315 2657 1349
rect 2719 1315 2753 1349
rect 2815 1315 2849 1349
rect 2911 1315 2945 1349
rect 3007 1315 3041 1349
rect 3103 1315 3137 1349
rect 3199 1315 3233 1349
rect 3295 1315 3329 1349
rect 3391 1315 3425 1349
rect 3487 1315 3521 1349
rect 3583 1315 3617 1349
rect 3679 1315 3713 1349
rect 3775 1315 3809 1349
rect 3871 1315 3905 1349
rect 3967 1315 4001 1349
rect 4063 1315 4097 1349
rect 4159 1315 4193 1349
rect 4255 1315 4289 1349
rect 4351 1315 4385 1349
rect 4447 1315 4481 1349
rect 4543 1315 4577 1349
rect 4639 1315 4673 1349
rect 4735 1315 4769 1349
rect 4831 1315 4865 1349
rect -2839 1022 -2835 1056
rect -2835 1022 -2805 1056
rect -2767 1022 -2733 1056
rect -2498 931 -2101 1181
rect -1967 931 -1570 1181
rect -1233 1212 -1200 1240
rect -1200 1212 -1199 1240
rect -1233 1206 -1199 1212
rect -1223 1038 -1189 1072
rect -1036 1046 -1002 1049
rect -1036 1015 -1035 1046
rect -1035 1015 -1002 1046
rect -759 1038 -725 1072
rect 31 1210 65 1238
rect 31 1204 65 1210
rect -645 1072 -611 1074
rect -645 1040 -611 1072
rect -252 1056 -218 1061
rect -252 1027 -251 1056
rect -251 1027 -218 1056
rect -360 869 -326 887
rect -360 853 -343 869
rect -343 853 -326 869
rect -158 786 -124 815
rect -158 781 -127 786
rect -127 781 -124 786
rect 509 1024 543 1025
rect 509 991 539 1024
rect 539 991 543 1024
rect 917 1012 921 1046
rect 921 1012 951 1046
rect 127 788 161 794
rect 127 760 161 788
rect 1375 1056 1409 1090
rect 2239 1056 2273 1090
rect 2047 982 2081 1016
rect 2623 982 2657 1016
rect 2996 981 2997 1014
rect 2997 981 3030 1014
rect 2996 980 3030 981
rect 4282 1012 4286 1046
rect 4286 1012 4316 1046
rect 4354 1012 4388 1046
rect 4669 1012 4673 1046
rect 4673 1012 4703 1046
rect 4741 1012 4775 1046
rect 3680 918 3711 943
rect 3711 918 3714 943
rect 3680 909 3714 918
rect 3680 869 3714 871
rect 3680 837 3711 869
rect 3711 837 3714 869
rect -2849 649 -2815 683
rect -2753 649 -2719 683
rect -2657 649 -2623 683
rect -2561 649 -2527 683
rect -2465 649 -2431 683
rect -2369 649 -2335 683
rect -2273 649 -2239 683
rect -2177 649 -2143 683
rect -2081 649 -2047 683
rect -1985 649 -1951 683
rect -1889 649 -1855 683
rect -1793 649 -1759 683
rect -1697 649 -1663 683
rect -1601 649 -1567 683
rect -1505 649 -1471 683
rect -1409 649 -1375 683
rect -1313 649 -1279 683
rect -1217 649 -1183 683
rect -1121 649 -1087 683
rect -1025 649 -991 683
rect -929 649 -895 683
rect -833 649 -799 683
rect -737 649 -703 683
rect -641 649 -607 683
rect -545 649 -511 683
rect -449 649 -415 683
rect -353 649 -319 683
rect -257 649 -223 683
rect -161 649 -127 683
rect -65 649 -31 683
rect 31 649 65 683
rect 127 649 161 683
rect 223 649 257 683
rect 319 649 353 683
rect 415 649 449 683
rect 511 649 545 683
rect 607 649 641 683
rect 703 649 737 683
rect 799 649 833 683
rect 895 649 929 683
rect 991 649 1025 683
rect 1087 649 1121 683
rect 1183 649 1217 683
rect 1279 649 1313 683
rect 1375 649 1409 683
rect 1471 649 1505 683
rect 1567 649 1601 683
rect 1663 649 1697 683
rect 1759 649 1793 683
rect 1855 649 1889 683
rect 1951 649 1985 683
rect 2047 649 2081 683
rect 2143 649 2177 683
rect 2239 649 2273 683
rect 2335 649 2369 683
rect 2431 649 2465 683
rect 2527 649 2561 683
rect 2623 649 2657 683
rect 2719 649 2753 683
rect 2815 649 2849 683
rect 2911 649 2945 683
rect 3007 649 3041 683
rect 3103 649 3137 683
rect 3199 649 3233 683
rect 3295 649 3329 683
rect 3391 649 3425 683
rect 3487 649 3521 683
rect 3583 649 3617 683
rect 3679 649 3713 683
rect 3775 649 3809 683
rect 3871 649 3905 683
rect 3967 649 4001 683
rect 4063 649 4097 683
rect 4159 649 4193 683
rect 4255 649 4289 683
rect 4351 649 4385 683
rect 4447 649 4481 683
rect 4543 649 4577 683
rect 4639 649 4673 683
rect 4735 649 4769 683
rect 4831 649 4865 683
rect -1687 276 -1683 310
rect -1683 276 -1653 310
rect -1615 276 -1581 310
rect -1346 151 -949 401
rect -815 151 -418 401
rect 127 544 161 572
rect 127 538 161 544
rect -71 260 -37 294
rect 505 308 539 342
rect -81 120 -47 126
rect -81 92 -48 120
rect -48 92 -47 120
rect 31 122 65 128
rect 31 94 65 122
rect 921 286 955 320
rect 1375 242 1409 276
rect 2047 316 2081 350
rect 2239 242 2273 276
rect 2623 316 2657 350
rect 2998 351 3032 353
rect 2998 319 3031 351
rect 3031 319 3032 351
rect 3274 463 3283 490
rect 3283 463 3308 490
rect 3274 456 3308 463
rect 3274 414 3308 418
rect 3274 384 3283 414
rect 3283 384 3308 414
rect 3683 463 3711 486
rect 3711 463 3717 486
rect 3683 452 3717 463
rect 3683 380 3711 414
rect 3711 380 3717 414
rect 4262 340 4296 341
rect 4262 307 4295 340
rect 4295 307 4296 340
rect 4387 319 4421 334
rect 4387 300 4395 319
rect 4395 300 4421 319
rect -1697 -17 -1663 17
rect -1601 -17 -1567 17
rect -1505 -17 -1471 17
rect -1409 -17 -1375 17
rect -1313 -17 -1279 17
rect -1217 -17 -1183 17
rect -1121 -17 -1087 17
rect -1025 -17 -991 17
rect -929 -17 -895 17
rect -833 -17 -799 17
rect -737 -17 -703 17
rect -641 -17 -607 17
rect -545 -17 -511 17
rect -449 -17 -415 17
rect -353 -17 -319 17
rect -257 -17 -223 17
rect -161 -17 -127 17
rect -65 -17 -31 17
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
rect 3199 -17 3233 17
rect 3295 -17 3329 17
rect 3391 -17 3425 17
rect 3487 -17 3521 17
rect 3583 -17 3617 17
rect 3679 -17 3713 17
rect 3775 -17 3809 17
rect 3871 -17 3905 17
rect 3967 -17 4001 17
rect 4063 -17 4097 17
rect 4159 -17 4193 17
rect 4255 -17 4289 17
rect 4351 -17 4385 17
rect 4447 -17 4481 17
rect 4543 -17 4577 17
rect 4639 -17 4673 17
rect 4735 -17 4769 17
rect 4831 -17 4865 17
rect -1503 -692 -1469 -304
rect -1389 -686 -1355 -310
rect -1301 -686 -1267 -310
rect -1345 -770 -1311 -736
rect -1503 -1406 -1469 -1018
rect -1389 -1400 -1355 -1024
rect -1301 -1400 -1267 -1024
rect -1345 -1484 -1311 -1450
<< metal1 >>
rect -1859 3472 -1739 3475
rect -833 3472 -713 3475
rect -1859 3465 -1698 3472
rect -1859 3095 -1849 3465
rect -1749 3460 -1698 3465
rect -1749 3095 -1738 3460
rect -1859 3085 -1738 3095
rect -1744 3084 -1738 3085
rect -1704 3084 -1698 3460
rect -1744 3072 -1698 3084
rect -1656 3466 -1468 3472
rect -1656 3460 -1536 3466
rect -1656 3084 -1650 3460
rect -1616 3452 -1536 3460
rect -1566 3092 -1536 3452
rect -1616 3084 -1536 3092
rect -1656 3078 -1536 3084
rect -1502 3078 -1468 3466
rect -1656 3072 -1468 3078
rect -1104 3466 -916 3472
rect -1104 3078 -1070 3466
rect -1036 3460 -916 3466
rect -1036 3452 -956 3460
rect -1036 3092 -1006 3452
rect -1036 3084 -956 3092
rect -922 3084 -916 3460
rect -1036 3078 -916 3084
rect -1104 3072 -916 3078
rect -874 3465 -713 3472
rect -874 3460 -823 3465
rect -874 3084 -868 3460
rect -834 3095 -823 3460
rect -723 3095 -713 3465
rect -834 3085 -713 3095
rect -834 3084 -828 3085
rect -874 3072 -828 3084
rect -1710 3034 -1564 3040
rect -1710 3000 -1694 3034
rect -1660 3026 -1564 3034
rect -1660 3000 -1630 3026
rect -1710 2984 -1630 3000
rect -1644 2974 -1630 2984
rect -1578 2974 -1564 3026
rect -1644 2960 -1564 2974
rect -1008 3034 -862 3040
rect -1008 3026 -912 3034
rect -1008 2974 -994 3026
rect -942 3000 -912 3026
rect -878 3000 -862 3034
rect -942 2984 -862 3000
rect -942 2974 -928 2984
rect -1008 2960 -928 2974
rect -1744 2751 -1698 2758
rect -1859 2746 -1698 2751
rect -1859 2741 -1738 2746
rect -1859 2371 -1849 2741
rect -1749 2371 -1738 2741
rect -1859 2370 -1738 2371
rect -1704 2370 -1698 2746
rect -1859 2361 -1698 2370
rect -1744 2358 -1698 2361
rect -1656 2752 -1468 2758
rect -1656 2746 -1536 2752
rect -1656 2370 -1650 2746
rect -1616 2734 -1536 2746
rect -1616 2370 -1536 2384
rect -1656 2364 -1536 2370
rect -1502 2364 -1468 2752
rect -1656 2358 -1468 2364
rect -1104 2752 -916 2758
rect -1104 2364 -1070 2752
rect -1036 2746 -916 2752
rect -1036 2734 -956 2746
rect -1036 2370 -956 2384
rect -922 2370 -916 2746
rect -1036 2364 -916 2370
rect -1104 2358 -916 2364
rect -874 2751 -828 2758
rect -874 2746 -713 2751
rect -874 2370 -868 2746
rect -834 2741 -713 2746
rect -834 2371 -823 2741
rect -723 2371 -713 2741
rect -834 2370 -713 2371
rect -874 2361 -713 2370
rect -874 2358 -828 2361
rect -1710 2320 -1564 2326
rect -1710 2286 -1694 2320
rect -1660 2312 -1564 2320
rect -1660 2286 -1630 2312
rect -1710 2270 -1630 2286
rect -1644 2260 -1630 2270
rect -1578 2260 -1564 2312
rect -1644 2246 -1564 2260
rect -1008 2320 -862 2326
rect -1008 2312 -912 2320
rect -1008 2260 -994 2312
rect -942 2286 -912 2312
rect -878 2286 -862 2320
rect -942 2270 -862 2286
rect -942 2260 -928 2270
rect -1008 2246 -928 2260
rect -2880 2040 4896 2047
rect -2880 2015 240 2040
rect 660 2015 1440 2040
rect 1860 2015 2640 2040
rect 3060 2015 3840 2040
rect 4260 2015 4896 2040
rect -2880 1981 -2849 2015
rect -2815 1981 -2753 2015
rect -2719 1981 -2657 2015
rect -2623 1981 -2561 2015
rect -2527 1981 -2465 2015
rect -2431 1981 -2369 2015
rect -2335 1981 -2273 2015
rect -2239 1981 -2177 2015
rect -2143 1981 -2081 2015
rect -2047 1981 -1985 2015
rect -1951 1981 -1889 2015
rect -1855 1981 -1793 2015
rect -1759 1981 -1697 2015
rect -1663 1981 -1601 2015
rect -1567 1981 -1505 2015
rect -1471 1981 -1409 2015
rect -1375 1981 -1313 2015
rect -1279 1981 -1217 2015
rect -1183 1981 -1121 2015
rect -1087 1981 -1025 2015
rect -991 1981 -929 2015
rect -895 1981 -833 2015
rect -799 1981 -737 2015
rect -703 1981 -641 2015
rect -607 1981 -545 2015
rect -511 1981 -449 2015
rect -415 1981 -353 2015
rect -319 1981 -257 2015
rect -223 1981 -161 2015
rect -127 1981 -65 2015
rect -31 1981 31 2015
rect 65 1981 127 2015
rect 161 1981 223 2015
rect 660 1981 703 2015
rect 737 1981 799 2015
rect 833 1981 895 2015
rect 929 1981 991 2015
rect 1025 1981 1087 2015
rect 1121 1981 1183 2015
rect 1217 1981 1279 2015
rect 1313 1981 1375 2015
rect 1409 1981 1440 2015
rect 1889 1981 1951 2015
rect 1985 1981 2047 2015
rect 2081 1981 2143 2015
rect 2177 1981 2239 2015
rect 2273 1981 2335 2015
rect 2369 1981 2431 2015
rect 2465 1981 2527 2015
rect 2561 1981 2623 2015
rect 3060 1981 3103 2015
rect 3137 1981 3199 2015
rect 3233 1981 3295 2015
rect 3329 1981 3391 2015
rect 3425 1981 3487 2015
rect 3521 1981 3583 2015
rect 3617 1981 3679 2015
rect 3713 1981 3775 2015
rect 3809 1981 3840 2015
rect 4289 1981 4351 2015
rect 4385 1981 4447 2015
rect 4481 1981 4543 2015
rect 4577 1981 4639 2015
rect 4673 1981 4735 2015
rect 4769 1981 4831 2015
rect 4865 1981 4896 2015
rect -2880 1960 240 1981
rect 660 1960 1440 1981
rect 1860 1960 2640 1981
rect 3060 1960 3840 1981
rect 4260 1960 4896 1981
rect -2880 1949 4896 1960
rect 112 1904 176 1913
rect 112 1870 127 1904
rect 161 1870 176 1904
rect 112 1861 176 1870
rect -2677 1790 -1173 1856
rect -2677 1673 -2611 1790
rect -2781 1651 -2611 1673
rect -2854 1599 -2848 1651
rect -2796 1599 -2776 1651
rect -2724 1607 -2611 1651
rect -2510 1733 -2089 1739
rect -2724 1599 -2718 1607
rect -2510 1483 -2498 1733
rect -2101 1483 -2089 1733
rect -2510 1477 -2089 1483
rect -1979 1733 -1558 1739
rect -1979 1483 -1967 1733
rect -1570 1483 -1558 1733
rect -1239 1626 -1173 1790
rect -1239 1592 -1223 1626
rect -1189 1592 -1173 1626
rect -1239 1576 -1173 1592
rect -1979 1477 -1558 1483
rect -1242 1467 -1190 1478
rect 16 1460 80 1469
rect 16 1426 31 1460
rect 65 1426 80 1460
rect 16 1417 80 1426
rect -1242 1409 -1190 1415
rect -2880 1380 4896 1381
rect -2880 1349 -460 1380
rect -40 1360 4896 1380
rect -40 1349 840 1360
rect 1260 1349 2040 1360
rect 2460 1349 3240 1360
rect 3660 1349 4440 1360
rect 4860 1349 4896 1360
rect -2880 1315 -2849 1349
rect -2815 1315 -2753 1349
rect -2719 1315 -2657 1349
rect -2623 1315 -2561 1349
rect -2527 1315 -2465 1349
rect -2431 1315 -2369 1349
rect -2335 1315 -2273 1349
rect -2239 1315 -2177 1349
rect -2143 1315 -2081 1349
rect -2047 1315 -1985 1349
rect -1951 1315 -1889 1349
rect -1855 1315 -1793 1349
rect -1759 1315 -1697 1349
rect -1663 1315 -1601 1349
rect -1567 1315 -1505 1349
rect -1471 1315 -1409 1349
rect -1375 1315 -1313 1349
rect -1279 1315 -1217 1349
rect -1183 1315 -1121 1349
rect -1087 1315 -1025 1349
rect -991 1315 -929 1349
rect -895 1315 -833 1349
rect -799 1315 -737 1349
rect -703 1315 -641 1349
rect -607 1315 -545 1349
rect -511 1315 -460 1349
rect -31 1315 31 1349
rect 65 1315 127 1349
rect 161 1315 223 1349
rect 257 1315 319 1349
rect 353 1315 415 1349
rect 449 1315 511 1349
rect 545 1315 607 1349
rect 641 1315 703 1349
rect 737 1315 799 1349
rect 833 1315 840 1349
rect 1260 1315 1279 1349
rect 1313 1315 1375 1349
rect 1409 1315 1471 1349
rect 1505 1315 1567 1349
rect 1601 1315 1663 1349
rect 1697 1315 1759 1349
rect 1793 1315 1855 1349
rect 1889 1315 1951 1349
rect 1985 1315 2040 1349
rect 2465 1315 2527 1349
rect 2561 1315 2623 1349
rect 2657 1315 2719 1349
rect 2753 1315 2815 1349
rect 2849 1315 2911 1349
rect 2945 1315 3007 1349
rect 3041 1315 3103 1349
rect 3137 1315 3199 1349
rect 3233 1315 3240 1349
rect 3660 1315 3679 1349
rect 3713 1315 3775 1349
rect 3809 1315 3871 1349
rect 3905 1315 3967 1349
rect 4001 1315 4063 1349
rect 4097 1315 4159 1349
rect 4193 1315 4255 1349
rect 4289 1315 4351 1349
rect 4385 1315 4440 1349
rect 4865 1315 4896 1349
rect -2880 1300 -460 1315
rect -40 1300 840 1315
rect 1260 1300 2040 1315
rect 2460 1300 3240 1315
rect 3660 1300 4440 1315
rect 4860 1300 4896 1315
rect -2880 1283 4896 1300
rect -1242 1249 -1190 1255
rect -2510 1181 -2089 1187
rect -2854 1013 -2848 1065
rect -2796 1013 -2776 1065
rect -2724 1057 -2718 1065
rect -2724 1013 -2611 1057
rect -2781 991 -2611 1013
rect -2677 874 -2611 991
rect -2510 931 -2498 1181
rect -2101 931 -2089 1181
rect -2510 925 -2089 931
rect -1979 1181 -1558 1187
rect -1242 1186 -1190 1197
rect 16 1238 80 1247
rect 16 1204 31 1238
rect 65 1204 80 1238
rect 16 1195 80 1204
rect -1979 931 -1967 1181
rect -1570 931 -1558 1181
rect 1363 1090 1421 1096
rect -1979 925 -1558 931
rect -1239 1072 -1173 1088
rect -1239 1038 -1223 1072
rect -1189 1038 -1173 1072
rect -1239 874 -1173 1038
rect -1051 1006 -1045 1058
rect -993 1006 -987 1058
rect -774 1029 -768 1081
rect -716 1029 -710 1081
rect -660 1031 -654 1083
rect -602 1031 -596 1083
rect -267 1018 -261 1070
rect -209 1018 -203 1070
rect 1363 1056 1375 1090
rect 1409 1087 1421 1090
rect 2227 1090 2285 1096
rect 2227 1087 2239 1090
rect 1409 1059 2239 1087
rect 1409 1056 1421 1059
rect 497 1025 555 1034
rect 497 991 509 1025
rect 543 991 555 1025
rect 902 1003 908 1055
rect 960 1003 966 1055
rect 1363 1050 1421 1056
rect 2227 1056 2239 1059
rect 2273 1056 2285 1090
rect 2227 1050 2285 1056
rect 2035 1016 2093 1022
rect 497 982 555 991
rect 2035 982 2047 1016
rect 2081 1013 2093 1016
rect 2611 1016 2669 1022
rect 2611 1013 2623 1016
rect 2081 985 2623 1013
rect 2081 982 2093 985
rect -2677 808 -1173 874
rect -375 844 -369 896
rect -317 844 -311 896
rect -167 824 -115 830
rect -167 766 -115 772
rect 112 794 176 803
rect 112 760 127 794
rect 161 760 176 794
rect 112 751 176 760
rect 501 715 547 982
rect 2035 976 2093 982
rect 2611 982 2623 985
rect 2657 982 2669 1016
rect 2611 976 2669 982
rect 2632 715 2660 976
rect 2981 971 2987 1023
rect 3039 971 3045 1023
rect 4267 1003 4273 1055
rect 4325 1003 4345 1055
rect 4397 1003 4403 1055
rect 4654 1003 4660 1055
rect 4712 1003 4732 1055
rect 4784 1003 4790 1055
rect 3671 952 3723 958
rect 3671 880 3723 900
rect 3671 822 3723 828
rect -2880 700 4896 715
rect -2880 683 240 700
rect 660 683 1440 700
rect 1860 683 2640 700
rect 3060 683 3840 700
rect 4260 683 4896 700
rect -2880 649 -2849 683
rect -2815 649 -2753 683
rect -2719 649 -2657 683
rect -2623 649 -2561 683
rect -2527 649 -2465 683
rect -2431 649 -2369 683
rect -2335 649 -2273 683
rect -2239 649 -2177 683
rect -2143 649 -2081 683
rect -2047 649 -1985 683
rect -1951 649 -1889 683
rect -1855 649 -1793 683
rect -1759 649 -1697 683
rect -1663 649 -1601 683
rect -1567 649 -1505 683
rect -1471 649 -1409 683
rect -1375 649 -1313 683
rect -1279 649 -1217 683
rect -1183 649 -1121 683
rect -1087 649 -1025 683
rect -991 649 -929 683
rect -895 649 -833 683
rect -799 649 -737 683
rect -703 649 -641 683
rect -607 649 -545 683
rect -511 649 -449 683
rect -415 649 -353 683
rect -319 649 -257 683
rect -223 649 -161 683
rect -127 649 -65 683
rect -31 649 31 683
rect 65 649 127 683
rect 161 649 223 683
rect 660 649 703 683
rect 737 649 799 683
rect 833 649 895 683
rect 929 649 991 683
rect 1025 649 1087 683
rect 1121 649 1183 683
rect 1217 649 1279 683
rect 1313 649 1375 683
rect 1409 649 1440 683
rect 1889 649 1951 683
rect 1985 649 2047 683
rect 2081 649 2143 683
rect 2177 649 2239 683
rect 2273 649 2335 683
rect 2369 649 2431 683
rect 2465 649 2527 683
rect 2561 649 2623 683
rect 3060 649 3103 683
rect 3137 649 3199 683
rect 3233 649 3295 683
rect 3329 649 3391 683
rect 3425 649 3487 683
rect 3521 649 3583 683
rect 3617 649 3679 683
rect 3713 649 3775 683
rect 3809 649 3840 683
rect 4289 649 4351 683
rect 4385 649 4447 683
rect 4481 649 4543 683
rect 4577 649 4639 683
rect 4673 649 4735 683
rect 4769 649 4831 683
rect 4865 649 4896 683
rect -2880 640 240 649
rect 660 640 1440 649
rect 1860 640 2640 649
rect 3060 640 3840 649
rect 4260 640 4896 649
rect -2880 617 4896 640
rect 112 572 176 581
rect 112 538 127 572
rect 161 538 176 572
rect 112 529 176 538
rect -1525 458 -21 524
rect -1525 341 -1459 458
rect -1629 319 -1459 341
rect -1702 267 -1696 319
rect -1644 267 -1624 319
rect -1572 275 -1459 319
rect -1358 401 -937 407
rect -1572 267 -1566 275
rect -1358 151 -1346 401
rect -949 151 -937 401
rect -1358 145 -937 151
rect -827 401 -406 407
rect -827 151 -815 401
rect -418 151 -406 401
rect -87 294 -21 458
rect 2632 356 2660 617
rect 3265 499 3317 505
rect 3265 427 3317 447
rect 3265 369 3317 375
rect 3674 495 3726 501
rect 3674 423 3726 443
rect 3674 365 3726 371
rect 490 299 496 351
rect 548 299 554 351
rect 2035 350 2093 356
rect -87 260 -71 294
rect -37 260 -21 294
rect 906 277 912 329
rect 964 277 970 329
rect 2035 316 2047 350
rect 2081 347 2093 350
rect 2611 350 2669 356
rect 2611 347 2623 350
rect 2081 319 2623 347
rect 2081 316 2093 319
rect 2035 310 2093 316
rect 2611 316 2623 319
rect 2657 316 2669 350
rect 2611 310 2669 316
rect 2983 310 2989 362
rect 3041 310 3047 362
rect 4245 350 4311 356
rect 4245 298 4253 350
rect 4305 298 4311 350
rect 4245 290 4311 298
rect 4372 291 4378 343
rect 4430 291 4450 343
rect -87 244 -21 260
rect 1363 276 1421 282
rect 1363 242 1375 276
rect 1409 273 1421 276
rect 2227 276 2285 282
rect 2227 273 2239 276
rect 1409 245 2239 273
rect 1409 242 1421 245
rect 1363 236 1421 242
rect 2227 242 2239 245
rect 2273 242 2285 276
rect 2227 236 2285 242
rect -827 145 -406 151
rect -90 135 -38 146
rect 16 128 80 137
rect 16 94 31 128
rect 65 94 80 128
rect 16 85 80 94
rect -90 77 -38 83
rect -1728 20 4896 49
rect -1728 17 840 20
rect 1260 17 2040 20
rect 2460 17 3240 20
rect 3660 17 4440 20
rect 4860 17 4896 20
rect -1728 -17 -1697 17
rect -1663 -17 -1601 17
rect -1567 -17 -1505 17
rect -1471 -17 -1409 17
rect -1375 -17 -1313 17
rect -1279 -17 -1217 17
rect -1183 -17 -1121 17
rect -1087 -17 -1025 17
rect -991 -17 -929 17
rect -895 -17 -833 17
rect -799 -17 -737 17
rect -703 -17 -641 17
rect -607 -17 -545 17
rect -511 -17 -449 17
rect -415 -17 -353 17
rect -319 -17 -257 17
rect -223 -17 -161 17
rect -127 -17 -65 17
rect -31 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 840 17
rect 1260 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2040 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3240 17
rect 3660 -17 3679 17
rect 3713 -17 3775 17
rect 3809 -17 3871 17
rect 3905 -17 3967 17
rect 4001 -17 4063 17
rect 4097 -17 4159 17
rect 4193 -17 4255 17
rect 4289 -17 4351 17
rect 4385 -17 4440 17
rect 4865 -17 4896 17
rect -1728 -40 840 -17
rect 1260 -40 2040 -17
rect 2460 -40 3240 -17
rect 3660 -40 4440 -17
rect 4860 -40 4896 -17
rect -1728 -49 4896 -40
rect -1266 -298 -1146 -295
rect -1537 -304 -1349 -298
rect -1537 -692 -1503 -304
rect -1469 -310 -1349 -304
rect -1469 -318 -1389 -310
rect -1469 -678 -1439 -318
rect -1469 -686 -1389 -678
rect -1355 -686 -1349 -310
rect -1469 -692 -1349 -686
rect -1537 -698 -1349 -692
rect -1307 -305 -1146 -298
rect -1307 -310 -1256 -305
rect -1307 -686 -1301 -310
rect -1267 -675 -1256 -310
rect -1156 -675 -1146 -305
rect -1267 -685 -1146 -675
rect -1267 -686 -1261 -685
rect -1307 -698 -1261 -686
rect -1441 -736 -1295 -730
rect -1441 -744 -1345 -736
rect -1441 -796 -1427 -744
rect -1375 -770 -1345 -744
rect -1311 -770 -1295 -736
rect -1375 -786 -1295 -770
rect -1375 -796 -1361 -786
rect -1441 -810 -1361 -796
rect -1537 -1018 -1349 -1012
rect -1537 -1406 -1503 -1018
rect -1469 -1024 -1349 -1018
rect -1469 -1036 -1389 -1024
rect -1469 -1400 -1389 -1386
rect -1355 -1400 -1349 -1024
rect -1469 -1406 -1349 -1400
rect -1537 -1412 -1349 -1406
rect -1307 -1019 -1261 -1012
rect -1307 -1024 -1146 -1019
rect -1307 -1400 -1301 -1024
rect -1267 -1029 -1146 -1024
rect -1267 -1399 -1256 -1029
rect -1156 -1399 -1146 -1029
rect -1267 -1400 -1146 -1399
rect -1307 -1409 -1146 -1400
rect -1307 -1412 -1261 -1409
rect -1441 -1450 -1295 -1444
rect -1441 -1458 -1345 -1450
rect -1441 -1510 -1427 -1458
rect -1375 -1484 -1345 -1458
rect -1311 -1484 -1295 -1450
rect -1375 -1500 -1295 -1484
rect -1375 -1510 -1361 -1500
rect -1441 -1524 -1361 -1510
<< via1 >>
rect -1849 3095 -1749 3465
rect -1636 3092 -1616 3452
rect -1616 3092 -1566 3452
rect -1006 3092 -956 3452
rect -956 3092 -936 3452
rect -823 3095 -723 3465
rect -1630 2974 -1578 3026
rect -994 2974 -942 3026
rect -1849 2371 -1749 2741
rect -1636 2384 -1616 2734
rect -1616 2384 -1536 2734
rect -1536 2384 -1526 2734
rect -1046 2384 -1036 2734
rect -1036 2384 -956 2734
rect -956 2384 -936 2734
rect -823 2371 -723 2741
rect -1630 2260 -1578 2312
rect -994 2260 -942 2312
rect 240 2015 660 2040
rect 1440 2015 1860 2040
rect 2640 2015 3060 2040
rect 3840 2015 4260 2040
rect 240 1981 257 2015
rect 257 1981 319 2015
rect 319 1981 353 2015
rect 353 1981 415 2015
rect 415 1981 449 2015
rect 449 1981 511 2015
rect 511 1981 545 2015
rect 545 1981 607 2015
rect 607 1981 641 2015
rect 641 1981 660 2015
rect 1440 1981 1471 2015
rect 1471 1981 1505 2015
rect 1505 1981 1567 2015
rect 1567 1981 1601 2015
rect 1601 1981 1663 2015
rect 1663 1981 1697 2015
rect 1697 1981 1759 2015
rect 1759 1981 1793 2015
rect 1793 1981 1855 2015
rect 1855 1981 1860 2015
rect 2640 1981 2657 2015
rect 2657 1981 2719 2015
rect 2719 1981 2753 2015
rect 2753 1981 2815 2015
rect 2815 1981 2849 2015
rect 2849 1981 2911 2015
rect 2911 1981 2945 2015
rect 2945 1981 3007 2015
rect 3007 1981 3041 2015
rect 3041 1981 3060 2015
rect 3840 1981 3871 2015
rect 3871 1981 3905 2015
rect 3905 1981 3967 2015
rect 3967 1981 4001 2015
rect 4001 1981 4063 2015
rect 4063 1981 4097 2015
rect 4097 1981 4159 2015
rect 4159 1981 4193 2015
rect 4193 1981 4255 2015
rect 4255 1981 4260 2015
rect 240 1960 660 1981
rect 1440 1960 1860 1981
rect 2640 1960 3060 1981
rect 3840 1960 4260 1981
rect -2848 1642 -2796 1651
rect -2848 1608 -2839 1642
rect -2839 1608 -2805 1642
rect -2805 1608 -2796 1642
rect -2848 1599 -2796 1608
rect -2776 1642 -2724 1651
rect -2776 1608 -2767 1642
rect -2767 1608 -2733 1642
rect -2733 1608 -2724 1642
rect -2776 1599 -2724 1608
rect -1957 1488 -1577 1728
rect -1242 1458 -1190 1467
rect -1242 1424 -1233 1458
rect -1233 1424 -1199 1458
rect -1199 1424 -1190 1458
rect -1242 1415 -1190 1424
rect -460 1349 -40 1380
rect 840 1349 1260 1360
rect 2040 1349 2460 1360
rect 3240 1349 3660 1360
rect 4440 1349 4860 1360
rect -460 1315 -449 1349
rect -449 1315 -415 1349
rect -415 1315 -353 1349
rect -353 1315 -319 1349
rect -319 1315 -257 1349
rect -257 1315 -223 1349
rect -223 1315 -161 1349
rect -161 1315 -127 1349
rect -127 1315 -65 1349
rect -65 1315 -40 1349
rect 840 1315 895 1349
rect 895 1315 929 1349
rect 929 1315 991 1349
rect 991 1315 1025 1349
rect 1025 1315 1087 1349
rect 1087 1315 1121 1349
rect 1121 1315 1183 1349
rect 1183 1315 1217 1349
rect 1217 1315 1260 1349
rect 2040 1315 2047 1349
rect 2047 1315 2081 1349
rect 2081 1315 2143 1349
rect 2143 1315 2177 1349
rect 2177 1315 2239 1349
rect 2239 1315 2273 1349
rect 2273 1315 2335 1349
rect 2335 1315 2369 1349
rect 2369 1315 2431 1349
rect 2431 1315 2460 1349
rect 3240 1315 3295 1349
rect 3295 1315 3329 1349
rect 3329 1315 3391 1349
rect 3391 1315 3425 1349
rect 3425 1315 3487 1349
rect 3487 1315 3521 1349
rect 3521 1315 3583 1349
rect 3583 1315 3617 1349
rect 3617 1315 3660 1349
rect 4440 1315 4447 1349
rect 4447 1315 4481 1349
rect 4481 1315 4543 1349
rect 4543 1315 4577 1349
rect 4577 1315 4639 1349
rect 4639 1315 4673 1349
rect 4673 1315 4735 1349
rect 4735 1315 4769 1349
rect 4769 1315 4831 1349
rect 4831 1315 4860 1349
rect -460 1300 -40 1315
rect 840 1300 1260 1315
rect 2040 1300 2460 1315
rect 3240 1300 3660 1315
rect 4440 1300 4860 1315
rect -1242 1240 -1190 1249
rect -1242 1206 -1233 1240
rect -1233 1206 -1199 1240
rect -1199 1206 -1190 1240
rect -1242 1197 -1190 1206
rect -2848 1056 -2796 1065
rect -2848 1022 -2839 1056
rect -2839 1022 -2805 1056
rect -2805 1022 -2796 1056
rect -2848 1013 -2796 1022
rect -2776 1056 -2724 1065
rect -2776 1022 -2767 1056
rect -2767 1022 -2733 1056
rect -2733 1022 -2724 1056
rect -2776 1013 -2724 1022
rect -1957 936 -1577 1176
rect -1045 1049 -993 1058
rect -1045 1015 -1036 1049
rect -1036 1015 -1002 1049
rect -1002 1015 -993 1049
rect -1045 1006 -993 1015
rect -768 1072 -716 1081
rect -768 1038 -759 1072
rect -759 1038 -725 1072
rect -725 1038 -716 1072
rect -768 1029 -716 1038
rect -654 1074 -602 1083
rect -654 1040 -645 1074
rect -645 1040 -611 1074
rect -611 1040 -602 1074
rect -654 1031 -602 1040
rect -261 1061 -209 1070
rect -261 1027 -252 1061
rect -252 1027 -218 1061
rect -218 1027 -209 1061
rect -261 1018 -209 1027
rect 908 1046 960 1055
rect 908 1012 917 1046
rect 917 1012 951 1046
rect 951 1012 960 1046
rect 908 1003 960 1012
rect -369 887 -317 896
rect -369 853 -360 887
rect -360 853 -326 887
rect -326 853 -317 887
rect -369 844 -317 853
rect -167 815 -115 824
rect -167 781 -158 815
rect -158 781 -124 815
rect -124 781 -115 815
rect -167 772 -115 781
rect 2987 1014 3039 1023
rect 2987 980 2996 1014
rect 2996 980 3030 1014
rect 3030 980 3039 1014
rect 2987 971 3039 980
rect 4273 1046 4325 1055
rect 4273 1012 4282 1046
rect 4282 1012 4316 1046
rect 4316 1012 4325 1046
rect 4273 1003 4325 1012
rect 4345 1046 4397 1055
rect 4345 1012 4354 1046
rect 4354 1012 4388 1046
rect 4388 1012 4397 1046
rect 4345 1003 4397 1012
rect 4660 1046 4712 1055
rect 4660 1012 4669 1046
rect 4669 1012 4703 1046
rect 4703 1012 4712 1046
rect 4660 1003 4712 1012
rect 4732 1046 4784 1055
rect 4732 1012 4741 1046
rect 4741 1012 4775 1046
rect 4775 1012 4784 1046
rect 4732 1003 4784 1012
rect 3671 943 3723 952
rect 3671 909 3680 943
rect 3680 909 3714 943
rect 3714 909 3723 943
rect 3671 900 3723 909
rect 3671 871 3723 880
rect 3671 837 3680 871
rect 3680 837 3714 871
rect 3714 837 3723 871
rect 3671 828 3723 837
rect 240 683 660 700
rect 1440 683 1860 700
rect 2640 683 3060 700
rect 3840 683 4260 700
rect 240 649 257 683
rect 257 649 319 683
rect 319 649 353 683
rect 353 649 415 683
rect 415 649 449 683
rect 449 649 511 683
rect 511 649 545 683
rect 545 649 607 683
rect 607 649 641 683
rect 641 649 660 683
rect 1440 649 1471 683
rect 1471 649 1505 683
rect 1505 649 1567 683
rect 1567 649 1601 683
rect 1601 649 1663 683
rect 1663 649 1697 683
rect 1697 649 1759 683
rect 1759 649 1793 683
rect 1793 649 1855 683
rect 1855 649 1860 683
rect 2640 649 2657 683
rect 2657 649 2719 683
rect 2719 649 2753 683
rect 2753 649 2815 683
rect 2815 649 2849 683
rect 2849 649 2911 683
rect 2911 649 2945 683
rect 2945 649 3007 683
rect 3007 649 3041 683
rect 3041 649 3060 683
rect 3840 649 3871 683
rect 3871 649 3905 683
rect 3905 649 3967 683
rect 3967 649 4001 683
rect 4001 649 4063 683
rect 4063 649 4097 683
rect 4097 649 4159 683
rect 4159 649 4193 683
rect 4193 649 4255 683
rect 4255 649 4260 683
rect 240 640 660 649
rect 1440 640 1860 649
rect 2640 640 3060 649
rect 3840 640 4260 649
rect -1696 310 -1644 319
rect -1696 276 -1687 310
rect -1687 276 -1653 310
rect -1653 276 -1644 310
rect -1696 267 -1644 276
rect -1624 310 -1572 319
rect -1624 276 -1615 310
rect -1615 276 -1581 310
rect -1581 276 -1572 310
rect -1624 267 -1572 276
rect -805 156 -425 396
rect 3265 490 3317 499
rect 3265 456 3274 490
rect 3274 456 3308 490
rect 3308 456 3317 490
rect 3265 447 3317 456
rect 3265 418 3317 427
rect 3265 384 3274 418
rect 3274 384 3308 418
rect 3308 384 3317 418
rect 3265 375 3317 384
rect 3674 486 3726 495
rect 3674 452 3683 486
rect 3683 452 3717 486
rect 3717 452 3726 486
rect 3674 443 3726 452
rect 3674 414 3726 423
rect 3674 380 3683 414
rect 3683 380 3717 414
rect 3717 380 3726 414
rect 3674 371 3726 380
rect 496 342 548 351
rect 496 308 505 342
rect 505 308 539 342
rect 539 308 548 342
rect 496 299 548 308
rect 912 320 964 329
rect 912 286 921 320
rect 921 286 955 320
rect 955 286 964 320
rect 912 277 964 286
rect 2989 353 3041 362
rect 2989 319 2998 353
rect 2998 319 3032 353
rect 3032 319 3041 353
rect 2989 310 3041 319
rect 4253 341 4305 350
rect 4253 307 4262 341
rect 4262 307 4296 341
rect 4296 307 4305 341
rect 4253 298 4305 307
rect 4378 334 4430 343
rect 4378 300 4387 334
rect 4387 300 4421 334
rect 4421 300 4430 334
rect 4378 291 4430 300
rect -90 126 -38 135
rect -90 92 -81 126
rect -81 92 -47 126
rect -47 92 -38 126
rect -90 83 -38 92
rect 840 17 1260 20
rect 2040 17 2460 20
rect 3240 17 3660 20
rect 4440 17 4860 20
rect 840 -17 895 17
rect 895 -17 929 17
rect 929 -17 991 17
rect 991 -17 1025 17
rect 1025 -17 1087 17
rect 1087 -17 1121 17
rect 1121 -17 1183 17
rect 1183 -17 1217 17
rect 1217 -17 1260 17
rect 2040 -17 2047 17
rect 2047 -17 2081 17
rect 2081 -17 2143 17
rect 2143 -17 2177 17
rect 2177 -17 2239 17
rect 2239 -17 2273 17
rect 2273 -17 2335 17
rect 2335 -17 2369 17
rect 2369 -17 2431 17
rect 2431 -17 2460 17
rect 3240 -17 3295 17
rect 3295 -17 3329 17
rect 3329 -17 3391 17
rect 3391 -17 3425 17
rect 3425 -17 3487 17
rect 3487 -17 3521 17
rect 3521 -17 3583 17
rect 3583 -17 3617 17
rect 3617 -17 3660 17
rect 4440 -17 4447 17
rect 4447 -17 4481 17
rect 4481 -17 4543 17
rect 4543 -17 4577 17
rect 4577 -17 4639 17
rect 4639 -17 4673 17
rect 4673 -17 4735 17
rect 4735 -17 4769 17
rect 4769 -17 4831 17
rect 4831 -17 4860 17
rect 840 -40 1260 -17
rect 2040 -40 2460 -17
rect 3240 -40 3660 -17
rect 4440 -40 4860 -17
rect -1439 -678 -1389 -318
rect -1389 -678 -1369 -318
rect -1256 -675 -1156 -305
rect -1427 -796 -1375 -744
rect -1479 -1386 -1469 -1036
rect -1469 -1386 -1389 -1036
rect -1389 -1386 -1369 -1036
rect -1256 -1399 -1156 -1029
rect -1427 -1510 -1375 -1458
<< metal2 >>
rect -1859 3465 -1739 3475
rect -1859 3095 -1849 3465
rect -1749 3095 -1739 3465
rect -833 3465 -713 3475
rect -1859 3085 -1739 3095
rect -1646 3452 -1556 3462
rect -1646 3092 -1636 3452
rect -1566 3092 -1556 3452
rect -1646 3082 -1556 3092
rect -1016 3452 -926 3462
rect -1016 3092 -1006 3452
rect -936 3092 -926 3452
rect -1016 3082 -926 3092
rect -833 3095 -823 3465
rect -723 3095 -713 3465
rect -833 3085 -713 3095
rect -2280 3026 -928 3040
rect -2280 2974 -1630 3026
rect -1578 2974 -994 3026
rect -942 2974 -928 3026
rect -2280 2960 -928 2974
rect -2920 1651 -2820 1660
rect -2920 1599 -2848 1651
rect -2796 1599 -2776 1651
rect -2724 1599 -2718 1651
rect -2920 1580 -2820 1599
rect -2940 1065 -2840 1080
rect -2940 1013 -2848 1065
rect -2796 1013 -2776 1065
rect -2724 1013 -2718 1065
rect -2940 1000 -2840 1013
rect -2280 180 -2200 2960
rect -1859 2741 -1739 2751
rect -1859 2371 -1849 2741
rect -1749 2371 -1739 2741
rect -1646 2734 -1516 2744
rect -1646 2384 -1636 2734
rect -1526 2384 -1516 2734
rect -1646 2374 -1516 2384
rect -1056 2734 -926 2744
rect -1056 2384 -1046 2734
rect -936 2384 -926 2734
rect -1056 2374 -926 2384
rect -833 2741 -713 2751
rect -1859 2361 -1739 2371
rect -833 2371 -823 2741
rect -723 2371 -713 2741
rect -833 2361 -713 2371
rect -2320 160 -2200 180
rect -2320 80 -2300 160
rect -2220 80 -2200 160
rect -2320 60 -2200 80
rect -2280 -1460 -2200 60
rect -2140 2312 -928 2326
rect -2140 2260 -1630 2312
rect -1578 2260 -994 2312
rect -942 2260 -928 2312
rect -2140 2246 -928 2260
rect -2140 0 -2060 2246
rect 220 2040 680 2060
rect 220 1960 240 2040
rect 660 1960 680 2040
rect 220 1940 680 1960
rect 1420 2040 1880 2060
rect 1420 1960 1440 2040
rect 1860 1960 1880 2040
rect 1420 1940 1880 1960
rect 2620 2040 3080 2060
rect 2620 1960 2640 2040
rect 3060 1960 3080 2040
rect 2620 1940 3080 1960
rect 3820 2040 4280 2060
rect 3820 1960 3840 2040
rect 4260 1960 4280 2040
rect 3820 1940 4280 1960
rect -1967 1728 -1567 1738
rect -1967 1720 -1957 1728
rect -1967 1500 -1960 1720
rect -1967 1488 -1957 1500
rect -1577 1488 -1567 1728
rect -1967 1478 -1567 1488
rect -1242 1467 -1190 1478
rect -1190 1439 -1141 1461
rect -1190 1415 -613 1439
rect -1242 1409 -613 1415
rect -1242 1249 -1190 1255
rect -1190 1238 -1141 1249
rect -1190 1208 -726 1238
rect -1190 1197 -1141 1208
rect -1242 1186 -1190 1197
rect -1967 1176 -1567 1186
rect -1967 1160 -1957 1176
rect -1967 940 -1960 1160
rect -1967 936 -1957 940
rect -1577 936 -1567 1176
rect -1967 926 -1567 936
rect -1144 1128 -910 1165
rect -1493 550 -1441 552
rect -1144 550 -1107 1128
rect -1051 1006 -1045 1058
rect -993 1006 -987 1058
rect -1045 970 -993 1006
rect -947 977 -910 1128
rect -756 1081 -726 1208
rect -643 1083 -613 1409
rect -480 1380 -20 1400
rect -480 1300 -460 1380
rect -40 1300 -20 1380
rect -480 1280 -20 1300
rect 820 1360 1280 1380
rect 820 1280 840 1360
rect 1260 1280 1280 1360
rect 820 1260 1280 1280
rect 2020 1360 2480 1380
rect 2020 1280 2040 1360
rect 2460 1280 2480 1360
rect 2020 1260 2480 1280
rect 3220 1360 3680 1380
rect 3220 1280 3240 1360
rect 3660 1280 3680 1360
rect 3220 1260 3680 1280
rect 4420 1360 4880 1380
rect 4420 1280 4440 1360
rect 4860 1280 4880 1360
rect 4420 1260 4880 1280
rect 767 1101 3033 1141
rect -774 1029 -768 1081
rect -716 1029 -710 1081
rect -660 1031 -654 1083
rect -602 1031 -596 1083
rect -267 1018 -261 1070
rect -209 1018 -203 1070
rect -259 977 -222 1018
rect -1038 581 -997 970
rect -947 940 -222 977
rect 767 908 807 1101
rect 902 1041 908 1055
rect -375 896 807 908
rect -375 844 -369 896
rect -317 868 807 896
rect 856 1003 908 1041
rect 960 1003 966 1055
rect 2993 1023 3033 1101
rect 4049 1107 4714 1144
rect -317 844 -310 868
rect 856 830 894 1003
rect 2981 971 2987 1023
rect 3039 971 3045 1023
rect -167 824 894 830
rect -115 792 894 824
rect 3671 952 3723 958
rect 3723 943 3740 952
rect 4049 943 4086 1107
rect 4677 1055 4714 1107
rect 4267 1003 4273 1055
rect 4325 1003 4345 1055
rect 4397 1003 4403 1055
rect 4654 1003 4660 1055
rect 4712 1003 4732 1055
rect 4784 1003 4790 1055
rect 3723 906 4086 943
rect 3723 900 3740 906
rect 3671 880 3723 900
rect 3671 822 3723 828
rect -167 766 -115 772
rect 220 720 680 740
rect 220 640 240 720
rect 660 640 680 720
rect 220 620 680 640
rect 1420 720 1880 740
rect 1420 640 1440 720
rect 1860 640 1880 720
rect 1420 620 1880 640
rect 2620 720 3080 740
rect 2620 640 2640 720
rect 3060 640 3080 720
rect 2620 620 3080 640
rect 3820 720 4280 740
rect 3820 640 3840 720
rect 4260 640 4280 720
rect 3820 620 4280 640
rect -1493 498 -1100 550
rect -1038 540 3370 581
rect -1980 340 -1860 360
rect -1980 260 -1960 340
rect -1880 319 -1640 340
rect -1493 319 -1441 498
rect -1880 267 -1696 319
rect -1644 267 -1624 319
rect -1572 267 -1441 319
rect -820 400 -400 420
rect -820 396 -800 400
rect -1880 260 -1640 267
rect -1980 240 -1860 260
rect -820 156 -805 396
rect -420 160 -400 400
rect 502 351 543 540
rect 3265 499 3370 540
rect 3317 447 3370 499
rect 3265 427 3370 447
rect 3317 416 3370 427
rect 3674 495 3726 501
rect 3674 423 3726 443
rect 4330 423 4363 1003
rect 3317 375 3594 416
rect 3265 369 3317 375
rect 490 299 496 351
rect 548 299 554 351
rect 906 325 912 329
rect -425 156 -400 160
rect -820 140 -400 156
rect 784 277 912 325
rect 964 277 970 329
rect 2983 310 2989 362
rect 3041 310 3047 362
rect -90 135 -38 146
rect 784 131 832 277
rect 2983 274 3047 310
rect 3549 327 3590 375
rect 3726 390 4363 423
rect 3726 371 3759 390
rect 3674 365 3726 371
rect 4205 350 4311 356
rect 4205 327 4253 350
rect 3549 298 4253 327
rect 4305 298 4311 350
rect 4700 343 4733 1003
rect 3549 290 4311 298
rect 4372 291 4378 343
rect 4430 291 4733 343
rect 3549 286 4205 290
rect -38 83 832 131
rect -90 77 -38 83
rect 820 20 1280 40
rect -2140 -20 -2020 0
rect -2140 -100 -2120 -20
rect -2040 -100 -2020 -20
rect 820 -60 840 20
rect 1260 -60 1280 20
rect 820 -80 1280 -60
rect 2020 20 2480 40
rect 2020 -60 2040 20
rect 2460 -60 2480 20
rect 2020 -80 2480 -60
rect 3220 20 3680 40
rect 3220 -60 3240 20
rect 3660 -60 3680 20
rect 3220 -80 3680 -60
rect 4420 20 4880 40
rect 4420 -60 4440 20
rect 4860 -60 4880 20
rect 4420 -80 4880 -60
rect -2140 -120 -2020 -100
rect -2140 -740 -2060 -120
rect -1266 -305 -1146 -295
rect -1449 -318 -1359 -308
rect -1449 -678 -1439 -318
rect -1369 -678 -1359 -318
rect -1449 -688 -1359 -678
rect -1266 -675 -1256 -305
rect -1156 -675 -1146 -305
rect -1266 -685 -1146 -675
rect -1441 -735 -1361 -730
rect -1446 -740 -1361 -735
rect -2140 -744 -1361 -740
rect -2140 -796 -1427 -744
rect -1375 -796 -1361 -744
rect -2140 -810 -1361 -796
rect -2140 -820 -1440 -810
rect -1489 -1036 -1359 -1026
rect -1489 -1386 -1479 -1036
rect -1369 -1386 -1359 -1036
rect -1489 -1396 -1359 -1386
rect -1266 -1029 -1146 -1019
rect -1266 -1399 -1256 -1029
rect -1156 -1399 -1146 -1029
rect -1266 -1409 -1146 -1399
rect -1441 -1449 -1361 -1444
rect -1446 -1458 -1361 -1449
rect -1446 -1460 -1427 -1458
rect -2280 -1510 -1427 -1460
rect -1375 -1510 -1361 -1458
rect -2280 -1524 -1361 -1510
rect -2280 -1540 -1380 -1524
<< via2 >>
rect -1849 3095 -1749 3465
rect -1626 3092 -1566 3452
rect -1006 3092 -946 3452
rect -823 3095 -723 3465
rect -1849 2371 -1749 2741
rect -1626 2384 -1526 2734
rect -1046 2384 -946 2734
rect -823 2371 -723 2741
rect -2300 80 -2220 160
rect 240 1960 660 2040
rect 1440 1960 1860 2040
rect 2640 1960 3060 2040
rect 3840 1960 4260 2040
rect -1960 1500 -1957 1720
rect -1957 1500 -1580 1720
rect -1960 940 -1957 1160
rect -1957 940 -1580 1160
rect -460 1300 -40 1380
rect 840 1300 1260 1360
rect 840 1280 1260 1300
rect 2040 1300 2460 1360
rect 2040 1280 2460 1300
rect 3240 1300 3660 1360
rect 3240 1280 3660 1300
rect 4440 1300 4860 1360
rect 4440 1280 4860 1300
rect 240 700 660 720
rect 240 640 660 700
rect 1440 700 1860 720
rect 1440 640 1860 700
rect 2640 700 3060 720
rect 2640 640 3060 700
rect 3840 700 4260 720
rect 3840 640 4260 700
rect -1960 260 -1880 340
rect -800 396 -420 400
rect -800 160 -425 396
rect -425 160 -420 396
rect -2120 -100 -2040 -20
rect 840 -40 1260 20
rect 840 -60 1260 -40
rect 2040 -40 2460 20
rect 2040 -60 2460 -40
rect 3240 -40 3660 20
rect 3240 -60 3660 -40
rect 4440 -40 4860 20
rect 4440 -60 4860 -40
rect -1439 -678 -1379 -318
rect -1256 -675 -1156 -305
rect -1479 -1386 -1379 -1036
rect -1256 -1399 -1156 -1029
<< metal3 >>
rect -3729 3465 -1699 3475
rect -3729 3435 -1849 3465
rect -1749 3435 -1699 3465
rect -3729 3115 -1979 3435
rect -1739 3115 -1699 3435
rect -3729 3095 -1849 3115
rect -1749 3095 -1699 3115
rect -3729 3081 -1699 3095
rect -1636 3452 -936 3472
rect -1636 3092 -1626 3452
rect -1566 3332 -1006 3452
rect -1566 3232 -1556 3332
rect -1420 3232 -1260 3332
rect -1016 3232 -1006 3332
rect -1566 3092 -1006 3232
rect -946 3092 -936 3452
rect -1636 3082 -1556 3092
rect -5299 2741 -1699 2761
rect -1420 2754 -1260 3092
rect -1016 3082 -936 3092
rect -873 3465 1157 3475
rect -873 3435 -823 3465
rect -723 3435 1157 3465
rect -873 3115 -833 3435
rect -593 3115 1157 3435
rect -873 3095 -823 3115
rect -723 3095 1157 3115
rect -873 3081 1157 3095
rect -5299 2721 -1849 2741
rect -1749 2721 -1699 2741
rect -5299 2401 -1979 2721
rect -1739 2401 -1699 2721
rect -5299 2371 -1849 2401
rect -1749 2371 -1699 2401
rect -1636 2734 -936 2754
rect -1636 2384 -1626 2734
rect -1526 2614 -1046 2734
rect -1526 2514 -1516 2614
rect -1420 2514 -1260 2614
rect -1056 2514 -1046 2614
rect -1526 2384 -1046 2514
rect -946 2384 -936 2734
rect -1636 2374 -936 2384
rect -873 2741 2727 2761
rect -873 2721 -823 2741
rect -723 2721 2727 2741
rect -873 2401 -833 2721
rect -593 2401 2727 2721
rect -5299 2367 -1699 2371
rect -1859 2361 -1739 2367
rect -1980 1720 -1560 1740
rect -1980 1500 -1960 1720
rect -1580 1500 -1560 1720
rect -1980 1480 -1560 1500
rect -1420 1420 -1260 2374
rect -873 2371 -823 2401
rect -723 2371 2727 2401
rect -873 2367 2727 2371
rect -833 2361 -713 2367
rect 220 2040 4280 2060
rect 220 1960 240 2040
rect 660 1960 1440 2040
rect 1860 1960 2640 2040
rect 3060 1960 3840 2040
rect 4260 1960 4280 2040
rect 220 1940 4280 1960
rect -1420 1380 40 1420
rect -1420 1300 -460 1380
rect -40 1300 40 1380
rect -1420 1260 40 1300
rect -1980 1160 -1560 1180
rect -1980 940 -1960 1160
rect -1580 940 -1560 1160
rect -1980 920 -1560 940
rect -1420 820 -1260 1260
rect -1780 660 -1260 820
rect 220 740 340 1940
rect 560 740 680 1940
rect 220 720 680 740
rect -2480 340 -1860 360
rect -2480 260 -1960 340
rect -1880 260 -1860 340
rect -2480 240 -1860 260
rect -2480 160 -2200 180
rect -2480 80 -2300 160
rect -2220 80 -2200 160
rect -2480 60 -2200 80
rect -1780 40 -1620 660
rect 220 640 240 720
rect 660 640 680 720
rect 220 620 680 640
rect 820 1360 1280 1380
rect 820 1280 840 1360
rect 1260 1280 1280 1360
rect 820 1260 1280 1280
rect -820 400 -400 420
rect -820 160 -800 400
rect -420 160 -400 400
rect -820 140 -400 160
rect 820 40 940 1260
rect 1160 40 1280 1260
rect 1420 740 1540 1940
rect 1760 740 1880 1940
rect 1420 720 1880 740
rect 1420 640 1440 720
rect 1860 640 1880 720
rect 1420 620 1880 640
rect 2020 1360 2480 1380
rect 2020 1280 2040 1360
rect 2460 1280 2480 1360
rect 2020 1260 2480 1280
rect 2020 40 2140 1260
rect 2360 40 2480 1260
rect 2620 740 2740 1940
rect 2960 740 3080 1940
rect 2620 720 3080 740
rect 2620 640 2640 720
rect 3060 640 3080 720
rect 2620 620 3080 640
rect 3220 1360 3680 1380
rect 3220 1280 3240 1360
rect 3660 1280 3680 1360
rect 3220 1260 3680 1280
rect 3220 40 3340 1260
rect 3560 40 3680 1260
rect 3820 740 3940 1940
rect 4160 740 4280 1940
rect 3820 720 4280 740
rect 3820 640 3840 720
rect 4260 640 4280 720
rect 3820 620 4280 640
rect 4420 1360 4880 1380
rect 4420 1280 4440 1360
rect 4860 1280 4880 1360
rect 4420 1260 4880 1280
rect 4420 40 4540 1260
rect 4760 40 4880 1260
rect -1780 20 4880 40
rect -2480 -20 -2020 0
rect -2480 -100 -2120 -20
rect -2040 -100 -2020 -20
rect -2480 -120 -2020 -100
rect -1780 -60 840 20
rect 1260 -60 2040 20
rect 2460 -60 3240 20
rect 3660 -60 4440 20
rect 4860 -60 4880 20
rect -1780 -80 4880 -60
rect -1780 -298 -1620 -80
rect -1780 -318 -1369 -298
rect -1780 -438 -1439 -318
rect -1780 -538 -1620 -438
rect -1449 -538 -1439 -438
rect -1780 -678 -1439 -538
rect -1379 -678 -1369 -318
rect -1780 -1016 -1620 -678
rect -1449 -688 -1369 -678
rect -1306 -305 724 -295
rect -1306 -335 -1256 -305
rect -1156 -335 724 -305
rect -1306 -655 -1266 -335
rect -1026 -655 724 -335
rect -1306 -675 -1256 -655
rect -1156 -675 724 -655
rect -1306 -689 724 -675
rect -1780 -1036 -1369 -1016
rect -1780 -1156 -1479 -1036
rect -1780 -1256 -1620 -1156
rect -1489 -1256 -1479 -1156
rect -1780 -1386 -1479 -1256
rect -1379 -1386 -1369 -1036
rect -1780 -1396 -1369 -1386
rect -1306 -1029 2294 -1009
rect -1306 -1049 -1256 -1029
rect -1156 -1049 2294 -1029
rect -1306 -1369 -1266 -1049
rect -1026 -1369 2294 -1049
rect -1780 -1580 -1620 -1396
rect -1306 -1399 -1256 -1369
rect -1156 -1399 2294 -1369
rect -1306 -1403 2294 -1399
rect -1266 -1409 -1146 -1403
<< via3 >>
rect -1979 3115 -1849 3435
rect -1849 3115 -1749 3435
rect -1749 3115 -1739 3435
rect -833 3115 -823 3435
rect -823 3115 -723 3435
rect -723 3115 -593 3435
rect -1979 2401 -1849 2721
rect -1849 2401 -1749 2721
rect -1749 2401 -1739 2721
rect -833 2401 -823 2721
rect -823 2401 -723 2721
rect -723 2401 -593 2721
rect -1960 1500 -1580 1720
rect -1960 940 -1580 1160
rect -800 160 -420 400
rect -1266 -655 -1256 -335
rect -1256 -655 -1156 -335
rect -1156 -655 -1026 -335
rect -1266 -1369 -1256 -1049
rect -1256 -1369 -1156 -1049
rect -1156 -1369 -1026 -1049
<< mimcap >>
rect -3689 3415 -2119 3435
rect -3689 3135 -3669 3415
rect -2139 3135 -2119 3415
rect -3689 3115 -2119 3135
rect -453 3415 1117 3435
rect -453 3135 -433 3415
rect 1097 3135 1117 3415
rect -453 3115 1117 3135
rect -5259 2701 -2119 2721
rect -5259 2421 -5239 2701
rect -2139 2421 -2119 2701
rect -5259 2401 -2119 2421
rect -453 2701 2687 2721
rect -453 2421 -433 2701
rect 2667 2421 2687 2701
rect -453 2401 2687 2421
rect -886 -355 684 -335
rect -886 -635 -866 -355
rect 664 -635 684 -355
rect -886 -655 684 -635
rect -886 -1069 2254 -1049
rect -886 -1349 -866 -1069
rect 2234 -1349 2254 -1069
rect -886 -1369 2254 -1349
<< mimcapcontact >>
rect -3669 3135 -2139 3415
rect -433 3135 1097 3415
rect -5239 2421 -2139 2701
rect -433 2421 2667 2701
rect -866 -635 664 -355
rect -866 -1349 2234 -1069
<< metal4 >>
rect -3729 3465 -2079 3475
rect -3739 3415 -2079 3465
rect -3739 3135 -3669 3415
rect -2139 3135 -2079 3415
rect -3739 3085 -2079 3135
rect -3729 3081 -2079 3085
rect -2019 3435 -1699 3475
rect -2019 3115 -1979 3435
rect -1739 3115 -1699 3435
rect -2019 3081 -1699 3115
rect -873 3435 -553 3475
rect -873 3115 -833 3435
rect -593 3115 -553 3435
rect -873 3081 -553 3115
rect -493 3465 1157 3475
rect -493 3415 1167 3465
rect -493 3135 -433 3415
rect 1097 3135 1167 3415
rect -493 3085 1167 3135
rect -493 3081 1157 3085
rect -2400 2761 -2200 3081
rect -360 2761 -160 3081
rect -5299 2751 -2079 2761
rect -5309 2701 -2079 2751
rect -5309 2421 -5239 2701
rect -2139 2421 -2079 2701
rect -5309 2371 -2079 2421
rect -5299 2367 -2079 2371
rect -2019 2721 -1699 2761
rect -2019 2401 -1979 2721
rect -1739 2401 -1699 2721
rect -2019 2367 -1699 2401
rect -873 2721 -553 2761
rect -873 2401 -833 2721
rect -593 2401 -553 2721
rect -873 2367 -553 2401
rect -493 2751 2727 2761
rect -493 2701 2737 2751
rect -493 2421 -433 2701
rect 2667 2421 2737 2701
rect -493 2371 2737 2421
rect -493 2367 2727 2371
rect -2400 1200 -2200 2367
rect -360 1760 -160 2367
rect -2000 1720 -160 1760
rect -2000 1500 -1960 1720
rect -1580 1560 -160 1720
rect -1580 1500 -1500 1560
rect -2000 1460 -1500 1500
rect -2400 1160 -1500 1200
rect -2400 1000 -1960 1160
rect -2000 940 -1960 1000
rect -1580 940 -1500 1160
rect -2000 900 -1500 940
rect -820 400 -400 420
rect -820 160 -800 400
rect -420 160 -400 400
rect -820 140 -400 160
rect -680 -295 -480 140
rect -1306 -335 -986 -295
rect -1306 -655 -1266 -335
rect -1026 -655 -986 -335
rect -1306 -689 -986 -655
rect -926 -305 724 -295
rect -926 -355 734 -305
rect -926 -635 -866 -355
rect 664 -635 734 -355
rect -926 -685 734 -635
rect -926 -689 724 -685
rect -680 -1009 -480 -689
rect -1306 -1049 -986 -1009
rect -1306 -1369 -1266 -1049
rect -1026 -1369 -986 -1049
rect -1306 -1403 -986 -1369
rect -926 -1019 2294 -1009
rect -926 -1069 2304 -1019
rect -926 -1349 -866 -1069
rect 2234 -1349 2304 -1069
rect -926 -1399 2304 -1349
rect -926 -1403 2294 -1399
<< via4 >>
rect -1979 3115 -1739 3435
rect -833 3115 -593 3435
rect -1979 2401 -1739 2721
rect -833 2401 -593 2721
rect -1266 -655 -1026 -335
rect -1266 -1369 -1026 -1049
<< mimcap2 >>
rect -3689 3415 -2119 3435
rect -3689 3135 -3669 3415
rect -2139 3135 -2119 3415
rect -3689 3115 -2119 3135
rect -453 3415 1117 3435
rect -453 3135 -433 3415
rect 1097 3135 1117 3415
rect -453 3115 1117 3135
rect -5259 2701 -2119 2721
rect -5259 2421 -5239 2701
rect -2139 2421 -2119 2701
rect -5259 2401 -2119 2421
rect -453 2701 2687 2721
rect -453 2421 -433 2701
rect 2667 2421 2687 2701
rect -453 2401 2687 2421
rect -886 -355 684 -335
rect -886 -635 -866 -355
rect 664 -635 684 -355
rect -886 -655 684 -635
rect -886 -1069 2254 -1049
rect -886 -1349 -866 -1069
rect 2234 -1349 2254 -1069
rect -886 -1369 2254 -1349
<< mimcap2contact >>
rect -3669 3135 -2139 3415
rect -433 3135 1097 3415
rect -5239 2421 -2139 2701
rect -433 2421 2667 2701
rect -866 -635 664 -355
rect -866 -1349 2234 -1069
<< metal5 >>
rect -3729 3435 -1699 3475
rect -3729 3415 -1979 3435
rect -3729 3135 -3669 3415
rect -2139 3135 -1979 3415
rect -3729 3115 -1979 3135
rect -1739 3115 -1699 3435
rect -3729 3081 -1699 3115
rect -873 3435 1157 3475
rect -873 3115 -833 3435
rect -593 3415 1157 3435
rect -593 3135 -433 3415
rect 1097 3135 1157 3415
rect -593 3115 1157 3135
rect -873 3081 1157 3115
rect -5299 2721 -1699 2761
rect -5299 2701 -1979 2721
rect -5299 2421 -5239 2701
rect -2139 2421 -1979 2701
rect -5299 2401 -1979 2421
rect -1739 2401 -1699 2721
rect -5299 2367 -1699 2401
rect -873 2721 2727 2761
rect -873 2401 -833 2721
rect -593 2701 2727 2721
rect -593 2421 -433 2701
rect 2667 2421 2727 2701
rect -593 2401 2727 2421
rect -873 2367 2727 2401
rect -1306 -335 724 -295
rect -1306 -655 -1266 -335
rect -1026 -355 724 -335
rect -1026 -635 -866 -355
rect 664 -635 724 -355
rect -1026 -655 724 -635
rect -1306 -689 724 -655
rect -1306 -1049 2294 -1009
rect -1306 -1369 -1266 -1049
rect -1026 -1069 2294 -1049
rect -1026 -1349 -866 -1069
rect 2234 -1349 2294 -1069
rect -1026 -1369 2294 -1349
rect -1306 -1403 2294 -1369
<< res1p41 >>
rect -2086 1465 -1982 1751
rect -2086 913 -1982 1199
rect -934 133 -830 419
<< labels >>
rlabel metal2 3720 371 3759 423 1 UPDN
rlabel metal3 -2480 240 -2420 360 1 CLKIN
rlabel metal2 -2940 1000 -2840 1080 1 A0
rlabel metal2 -2920 1580 -2820 1660 1 A1
rlabel locali 4900 1000 4940 1080 1 GP
rlabel metal2 2983 274 3047 362 1 RSTB
rlabel metal3 720 2037 788 2060 1 VHI
rlabel metal3 -439 1396 -371 1419 1 VLO
rlabel metal3 -2480 60 -2420 180 1 C100
rlabel metal3 -2480 -120 -2420 0 1 C50
rlabel metal2 2 870 32 906 1 MUX_OUT
rlabel metal2 180 792 210 828 1 ENCLK
rlabel locali 4934 265 4974 345 1 GN
rlabel metal2 174 92 209 121 1 UDCLK
<< end >>