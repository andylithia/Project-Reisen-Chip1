magic
tech sky130A
magscale 1 2
timestamp 1672019510
<< metal3 >>
rect 46000 46560 286000 46600
rect 46000 46240 47000 46560
rect 55000 46240 57000 46560
rect 65000 46240 67000 46560
rect 75000 46240 77000 46560
rect 85000 46240 87000 46560
rect 95000 46240 97000 46560
rect 105000 46240 107000 46560
rect 115000 46240 117000 46560
rect 125000 46240 127000 46560
rect 135000 46240 137000 46560
rect 145000 46240 147000 46560
rect 155000 46240 157000 46560
rect 165000 46240 167000 46560
rect 175000 46240 177000 46560
rect 185000 46240 187000 46560
rect 195000 46240 197000 46560
rect 205000 46240 207000 46560
rect 215000 46240 217000 46560
rect 225000 46240 227000 46560
rect 235000 46240 237000 46560
rect 245000 46240 247000 46560
rect 255000 46240 257000 46560
rect 265000 46240 267000 46560
rect 275000 46240 277000 46560
rect 285000 46240 286000 46560
rect 46000 46000 286000 46240
rect 46000 27000 51000 46000
rect 56000 27000 61000 46000
rect 66000 27000 71000 46000
rect 76000 27000 81000 46000
rect 86000 27000 91000 46000
rect 96000 27000 101000 46000
rect 106000 27000 111000 46000
rect 116000 27000 121000 46000
rect 126000 27000 131000 46000
rect 136000 27000 141000 46000
rect 146000 27000 151000 46000
rect 156000 27000 161000 46000
rect 166000 27000 171000 46000
rect 176000 27000 181000 46000
rect 186000 27000 191000 46000
rect 196000 27000 201000 46000
rect 206000 27000 211000 46000
rect 216000 27000 221000 46000
rect 226000 27000 231000 46000
rect 236000 27000 241000 46000
rect 246000 27000 251000 46000
rect 256000 27000 261000 46000
rect 266000 27000 271000 46000
rect 276000 27000 281000 46000
rect 46000 26000 52000 27000
rect 50000 25900 52000 26000
rect 55000 26000 62000 27000
rect 55000 25900 57000 26000
rect 50000 25000 57000 25900
rect 60000 25900 62000 26000
rect 65000 26000 72000 27000
rect 65000 25900 67000 26000
rect 60000 25000 67000 25900
rect 70000 25900 72000 26000
rect 75000 26000 82000 27000
rect 75000 25900 77000 26000
rect 70000 25000 77000 25900
rect 80000 25900 82000 26000
rect 85000 26000 92000 27000
rect 85000 25900 87000 26000
rect 80000 25000 87000 25900
rect 90000 25900 92000 26000
rect 95000 26000 102000 27000
rect 95000 25900 97000 26000
rect 90000 25000 97000 25900
rect 100000 25900 102000 26000
rect 105000 26000 112000 27000
rect 105000 25900 107000 26000
rect 100000 25000 107000 25900
rect 110000 25900 112000 26000
rect 115000 26000 122000 27000
rect 115000 25900 117000 26000
rect 110000 25000 117000 25900
rect 120000 25900 122000 26000
rect 125000 26000 132000 27000
rect 125000 25900 127000 26000
rect 120000 25000 127000 25900
rect 130000 25900 132000 26000
rect 135000 26000 142000 27000
rect 135000 25900 137000 26000
rect 130000 25000 137000 25900
rect 140000 25900 142000 26000
rect 145000 26000 152000 27000
rect 145000 25900 147000 26000
rect 140000 25000 147000 25900
rect 150000 25900 152000 26000
rect 155000 26000 162000 27000
rect 155000 25900 157000 26000
rect 150000 25000 157000 25900
rect 160000 25900 162000 26000
rect 165000 26000 172000 27000
rect 165000 25900 167000 26000
rect 160000 25000 167000 25900
rect 170000 25900 172000 26000
rect 175000 26000 182000 27000
rect 175000 25900 177000 26000
rect 170000 25000 177000 25900
rect 180000 25900 182000 26000
rect 185000 26000 192000 27000
rect 185000 25900 187000 26000
rect 180000 25000 187000 25900
rect 190000 25900 192000 26000
rect 195000 26000 202000 27000
rect 195000 25900 197000 26000
rect 190000 25000 197000 25900
rect 200000 25900 202000 26000
rect 205000 26000 212000 27000
rect 205000 25900 207000 26000
rect 200000 25000 207000 25900
rect 210000 25900 212000 26000
rect 215000 26000 222000 27000
rect 215000 25900 217000 26000
rect 210000 25000 217000 25900
rect 220000 25900 222000 26000
rect 225000 26000 232000 27000
rect 225000 25900 227000 26000
rect 220000 25000 227000 25900
rect 230000 25900 232000 26000
rect 235000 26000 242000 27000
rect 235000 25900 237000 26000
rect 230000 25000 237000 25900
rect 240000 25900 242000 26000
rect 245000 26000 252000 27000
rect 245000 25900 247000 26000
rect 240000 25000 247000 25900
rect 250000 25900 252000 26000
rect 255000 26000 262000 27000
rect 255000 25900 257000 26000
rect 250000 25000 257000 25900
rect 260000 25900 262000 26000
rect 265000 26000 272000 27000
rect 265000 25900 267000 26000
rect 260000 25000 267000 25900
rect 270000 25900 272000 26000
rect 275000 26000 282000 27000
rect 275000 25900 277000 26000
rect 270000 25000 277000 25900
rect 280000 25900 282000 26000
rect 285000 25900 287000 27000
rect 280000 25000 287000 25900
rect 51000 5900 56000 25000
rect 61000 5900 66000 25000
rect 71000 5900 76000 25000
rect 81000 5900 86000 25000
rect 91000 5900 96000 25000
rect 101000 5900 106000 25000
rect 111000 5900 116000 25000
rect 121000 5900 126000 25000
rect 131000 5900 136000 25000
rect 141000 5900 146000 25000
rect 151000 5900 156000 25000
rect 161000 5900 166000 25000
rect 171000 5900 176000 25000
rect 181000 5900 186000 25000
rect 191000 5900 196000 25000
rect 201000 5900 206000 25000
rect 211000 5900 216000 25000
rect 221000 5900 226000 25000
rect 231000 5900 236000 25000
rect 241000 5900 246000 25000
rect 251000 5900 256000 25000
rect 261000 5900 266000 25000
rect 271000 5900 276000 25000
rect 281000 5900 286000 25000
rect 46000 5660 286000 5900
rect 46000 5340 47000 5660
rect 55960 5340 57000 5660
rect 65960 5340 67000 5660
rect 75960 5340 77000 5660
rect 85960 5340 87000 5660
rect 95960 5340 97000 5660
rect 105960 5340 107000 5660
rect 115960 5340 117000 5660
rect 125960 5340 127000 5660
rect 135960 5340 137000 5660
rect 145960 5340 147000 5660
rect 155960 5340 157000 5660
rect 165960 5340 167000 5660
rect 175960 5340 177000 5660
rect 185960 5340 187000 5660
rect 195960 5340 197000 5660
rect 205960 5340 207000 5660
rect 215960 5340 217000 5660
rect 225960 5340 227000 5660
rect 235960 5340 237000 5660
rect 245960 5340 247000 5660
rect 255960 5340 257000 5660
rect 265960 5340 267000 5660
rect 275960 5340 277000 5660
rect 285960 5340 286000 5660
rect 46000 5300 286000 5340
<< via3 >>
rect 47000 46240 55000 46560
rect 57000 46240 65000 46560
rect 67000 46240 75000 46560
rect 77000 46240 85000 46560
rect 87000 46240 95000 46560
rect 97000 46240 105000 46560
rect 107000 46240 115000 46560
rect 117000 46240 125000 46560
rect 127000 46240 135000 46560
rect 137000 46240 145000 46560
rect 147000 46240 155000 46560
rect 157000 46240 165000 46560
rect 167000 46240 175000 46560
rect 177000 46240 185000 46560
rect 187000 46240 195000 46560
rect 197000 46240 205000 46560
rect 207000 46240 215000 46560
rect 217000 46240 225000 46560
rect 227000 46240 235000 46560
rect 237000 46240 245000 46560
rect 247000 46240 255000 46560
rect 257000 46240 265000 46560
rect 267000 46240 275000 46560
rect 277000 46240 285000 46560
rect 47000 5340 55960 5660
rect 57000 5340 65960 5660
rect 67000 5340 75960 5660
rect 77000 5340 85960 5660
rect 87000 5340 95960 5660
rect 97000 5340 105960 5660
rect 107000 5340 115960 5660
rect 117000 5340 125960 5660
rect 127000 5340 135960 5660
rect 137000 5340 145960 5660
rect 147000 5340 155960 5660
rect 157000 5340 165960 5660
rect 167000 5340 175960 5660
rect 177000 5340 185960 5660
rect 187000 5340 195960 5660
rect 197000 5340 205960 5660
rect 207000 5340 215960 5660
rect 217000 5340 225960 5660
rect 227000 5340 235960 5660
rect 237000 5340 245960 5660
rect 247000 5340 255960 5660
rect 257000 5340 265960 5660
rect 267000 5340 275960 5660
rect 277000 5340 285960 5660
<< mimcap >>
rect 46040 45940 50960 45960
rect 46040 26060 46060 45940
rect 50940 26060 50960 45940
rect 46040 26040 50960 26060
rect 56040 45940 60960 45960
rect 56040 26060 56060 45940
rect 60940 26060 60960 45940
rect 56040 26040 60960 26060
rect 66040 45940 70960 45960
rect 66040 26060 66060 45940
rect 70940 26060 70960 45940
rect 66040 26040 70960 26060
rect 76040 45940 80960 45960
rect 76040 26060 76060 45940
rect 80940 26060 80960 45940
rect 76040 26040 80960 26060
rect 86040 45940 90960 45960
rect 86040 26060 86060 45940
rect 90940 26060 90960 45940
rect 86040 26040 90960 26060
rect 96040 45940 100960 45960
rect 96040 26060 96060 45940
rect 100940 26060 100960 45940
rect 96040 26040 100960 26060
rect 106040 45940 110960 45960
rect 106040 26060 106060 45940
rect 110940 26060 110960 45940
rect 106040 26040 110960 26060
rect 116040 45940 120960 45960
rect 116040 26060 116060 45940
rect 120940 26060 120960 45940
rect 116040 26040 120960 26060
rect 126040 45940 130960 45960
rect 126040 26060 126060 45940
rect 130940 26060 130960 45940
rect 126040 26040 130960 26060
rect 136040 45940 140960 45960
rect 136040 26060 136060 45940
rect 140940 26060 140960 45940
rect 136040 26040 140960 26060
rect 146040 45940 150960 45960
rect 146040 26060 146060 45940
rect 150940 26060 150960 45940
rect 146040 26040 150960 26060
rect 156040 45940 160960 45960
rect 156040 26060 156060 45940
rect 160940 26060 160960 45940
rect 156040 26040 160960 26060
rect 166040 45940 170960 45960
rect 166040 26060 166060 45940
rect 170940 26060 170960 45940
rect 166040 26040 170960 26060
rect 176040 45940 180960 45960
rect 176040 26060 176060 45940
rect 180940 26060 180960 45940
rect 176040 26040 180960 26060
rect 186040 45940 190960 45960
rect 186040 26060 186060 45940
rect 190940 26060 190960 45940
rect 186040 26040 190960 26060
rect 196040 45940 200960 45960
rect 196040 26060 196060 45940
rect 200940 26060 200960 45940
rect 196040 26040 200960 26060
rect 206040 45940 210960 45960
rect 206040 26060 206060 45940
rect 210940 26060 210960 45940
rect 206040 26040 210960 26060
rect 216040 45940 220960 45960
rect 216040 26060 216060 45940
rect 220940 26060 220960 45940
rect 216040 26040 220960 26060
rect 226040 45940 230960 45960
rect 226040 26060 226060 45940
rect 230940 26060 230960 45940
rect 226040 26040 230960 26060
rect 236040 45940 240960 45960
rect 236040 26060 236060 45940
rect 240940 26060 240960 45940
rect 236040 26040 240960 26060
rect 246040 45940 250960 45960
rect 246040 26060 246060 45940
rect 250940 26060 250960 45940
rect 246040 26040 250960 26060
rect 256040 45940 260960 45960
rect 256040 26060 256060 45940
rect 260940 26060 260960 45940
rect 256040 26040 260960 26060
rect 266040 45940 270960 45960
rect 266040 26060 266060 45940
rect 270940 26060 270960 45940
rect 266040 26040 270960 26060
rect 276040 45940 280960 45960
rect 276040 26060 276060 45940
rect 280940 26060 280960 45940
rect 276040 26040 280960 26060
rect 51040 25840 55960 25860
rect 51040 5960 51060 25840
rect 55940 5960 55960 25840
rect 51040 5940 55960 5960
rect 61040 25840 65960 25860
rect 61040 5960 61060 25840
rect 65940 5960 65960 25840
rect 61040 5940 65960 5960
rect 71040 25840 75960 25860
rect 71040 5960 71060 25840
rect 75940 5960 75960 25840
rect 71040 5940 75960 5960
rect 81040 25840 85960 25860
rect 81040 5960 81060 25840
rect 85940 5960 85960 25840
rect 81040 5940 85960 5960
rect 91040 25840 95960 25860
rect 91040 5960 91060 25840
rect 95940 5960 95960 25840
rect 91040 5940 95960 5960
rect 101040 25840 105960 25860
rect 101040 5960 101060 25840
rect 105940 5960 105960 25840
rect 101040 5940 105960 5960
rect 111040 25840 115960 25860
rect 111040 5960 111060 25840
rect 115940 5960 115960 25840
rect 111040 5940 115960 5960
rect 121040 25840 125960 25860
rect 121040 5960 121060 25840
rect 125940 5960 125960 25840
rect 121040 5940 125960 5960
rect 131040 25840 135960 25860
rect 131040 5960 131060 25840
rect 135940 5960 135960 25840
rect 131040 5940 135960 5960
rect 141040 25840 145960 25860
rect 141040 5960 141060 25840
rect 145940 5960 145960 25840
rect 141040 5940 145960 5960
rect 151040 25840 155960 25860
rect 151040 5960 151060 25840
rect 155940 5960 155960 25840
rect 151040 5940 155960 5960
rect 161040 25840 165960 25860
rect 161040 5960 161060 25840
rect 165940 5960 165960 25840
rect 161040 5940 165960 5960
rect 171040 25840 175960 25860
rect 171040 5960 171060 25840
rect 175940 5960 175960 25840
rect 171040 5940 175960 5960
rect 181040 25840 185960 25860
rect 181040 5960 181060 25840
rect 185940 5960 185960 25840
rect 181040 5940 185960 5960
rect 191040 25840 195960 25860
rect 191040 5960 191060 25840
rect 195940 5960 195960 25840
rect 191040 5940 195960 5960
rect 201040 25840 205960 25860
rect 201040 5960 201060 25840
rect 205940 5960 205960 25840
rect 201040 5940 205960 5960
rect 211040 25840 215960 25860
rect 211040 5960 211060 25840
rect 215940 5960 215960 25840
rect 211040 5940 215960 5960
rect 221040 25840 225960 25860
rect 221040 5960 221060 25840
rect 225940 5960 225960 25840
rect 221040 5940 225960 5960
rect 231040 25840 235960 25860
rect 231040 5960 231060 25840
rect 235940 5960 235960 25840
rect 231040 5940 235960 5960
rect 241040 25840 245960 25860
rect 241040 5960 241060 25840
rect 245940 5960 245960 25840
rect 241040 5940 245960 5960
rect 251040 25840 255960 25860
rect 251040 5960 251060 25840
rect 255940 5960 255960 25840
rect 251040 5940 255960 5960
rect 261040 25840 265960 25860
rect 261040 5960 261060 25840
rect 265940 5960 265960 25840
rect 261040 5940 265960 5960
rect 271040 25840 275960 25860
rect 271040 5960 271060 25840
rect 275940 5960 275960 25840
rect 271040 5940 275960 5960
rect 281040 25840 285960 25860
rect 281040 5960 281060 25840
rect 285940 5960 285960 25840
rect 281040 5940 285960 5960
<< mimcapcontact >>
rect 46060 26060 50940 45940
rect 56060 26060 60940 45940
rect 66060 26060 70940 45940
rect 76060 26060 80940 45940
rect 86060 26060 90940 45940
rect 96060 26060 100940 45940
rect 106060 26060 110940 45940
rect 116060 26060 120940 45940
rect 126060 26060 130940 45940
rect 136060 26060 140940 45940
rect 146060 26060 150940 45940
rect 156060 26060 160940 45940
rect 166060 26060 170940 45940
rect 176060 26060 180940 45940
rect 186060 26060 190940 45940
rect 196060 26060 200940 45940
rect 206060 26060 210940 45940
rect 216060 26060 220940 45940
rect 226060 26060 230940 45940
rect 236060 26060 240940 45940
rect 246060 26060 250940 45940
rect 256060 26060 260940 45940
rect 266060 26060 270940 45940
rect 276060 26060 280940 45940
rect 51060 5960 55940 25840
rect 61060 5960 65940 25840
rect 71060 5960 75940 25840
rect 81060 5960 85940 25840
rect 91060 5960 95940 25840
rect 101060 5960 105940 25840
rect 111060 5960 115940 25840
rect 121060 5960 125940 25840
rect 131060 5960 135940 25840
rect 141060 5960 145940 25840
rect 151060 5960 155940 25840
rect 161060 5960 165940 25840
rect 171060 5960 175940 25840
rect 181060 5960 185940 25840
rect 191060 5960 195940 25840
rect 201060 5960 205940 25840
rect 211060 5960 215940 25840
rect 221060 5960 225940 25840
rect 231060 5960 235940 25840
rect 241060 5960 245940 25840
rect 251060 5960 255940 25840
rect 261060 5960 265940 25840
rect 271060 5960 275940 25840
rect 281060 5960 285940 25840
<< metal4 >>
rect 46000 46560 286000 46600
rect 46000 46240 47000 46560
rect 55000 46240 57000 46560
rect 65000 46240 67000 46560
rect 75000 46240 77000 46560
rect 85000 46240 87000 46560
rect 95000 46240 97000 46560
rect 105000 46240 107000 46560
rect 115000 46240 117000 46560
rect 125000 46240 127000 46560
rect 135000 46240 137000 46560
rect 145000 46240 147000 46560
rect 155000 46240 157000 46560
rect 165000 46240 167000 46560
rect 175000 46240 177000 46560
rect 185000 46240 187000 46560
rect 195000 46240 197000 46560
rect 205000 46240 207000 46560
rect 215000 46240 217000 46560
rect 225000 46240 227000 46560
rect 235000 46240 237000 46560
rect 245000 46240 247000 46560
rect 255000 46240 257000 46560
rect 265000 46240 267000 46560
rect 275000 46240 277000 46560
rect 285000 46240 286000 46560
rect 46000 46200 286000 46240
rect 46000 45940 51000 46000
rect 46000 26060 46060 45940
rect 50940 27000 51000 45940
rect 56000 45940 61000 46000
rect 56000 27000 56060 45940
rect 50940 26060 52000 27000
rect 46000 26000 52000 26060
rect 50000 25900 52000 26000
rect 55000 26060 56060 27000
rect 60940 27000 61000 45940
rect 66000 45940 71000 46000
rect 66000 27000 66060 45940
rect 60940 26060 62000 27000
rect 55000 26000 62000 26060
rect 55000 25900 57000 26000
rect 50000 25840 57000 25900
rect 50000 25000 51060 25840
rect 51000 5960 51060 25000
rect 55940 25000 57000 25840
rect 60000 25900 62000 26000
rect 65000 26060 66060 27000
rect 70940 27000 71000 45940
rect 76000 45940 81000 46000
rect 76000 27000 76060 45940
rect 70940 26060 72000 27000
rect 65000 26000 72000 26060
rect 65000 25900 67000 26000
rect 60000 25840 67000 25900
rect 60000 25000 61060 25840
rect 55940 5960 56000 25000
rect 51000 5900 56000 5960
rect 61000 5960 61060 25000
rect 65940 25000 67000 25840
rect 70000 25900 72000 26000
rect 75000 26060 76060 27000
rect 80940 27000 81000 45940
rect 86000 45940 91000 46000
rect 86000 27000 86060 45940
rect 80940 26060 82000 27000
rect 75000 26000 82000 26060
rect 75000 25900 77000 26000
rect 70000 25840 77000 25900
rect 70000 25000 71060 25840
rect 65940 5960 66000 25000
rect 61000 5900 66000 5960
rect 71000 5960 71060 25000
rect 75940 25000 77000 25840
rect 80000 25900 82000 26000
rect 85000 26060 86060 27000
rect 90940 27000 91000 45940
rect 96000 45940 101000 46000
rect 96000 27000 96060 45940
rect 90940 26060 92000 27000
rect 85000 26000 92000 26060
rect 85000 25900 87000 26000
rect 80000 25840 87000 25900
rect 80000 25000 81060 25840
rect 75940 5960 76000 25000
rect 71000 5900 76000 5960
rect 81000 5960 81060 25000
rect 85940 25000 87000 25840
rect 90000 25900 92000 26000
rect 95000 26060 96060 27000
rect 100940 27000 101000 45940
rect 106000 45940 111000 46000
rect 106000 27000 106060 45940
rect 100940 26060 102000 27000
rect 95000 26000 102000 26060
rect 95000 25900 97000 26000
rect 90000 25840 97000 25900
rect 90000 25000 91060 25840
rect 85940 5960 86000 25000
rect 81000 5900 86000 5960
rect 91000 5960 91060 25000
rect 95940 25000 97000 25840
rect 100000 25900 102000 26000
rect 105000 26060 106060 27000
rect 110940 27000 111000 45940
rect 116000 45940 121000 46000
rect 116000 27000 116060 45940
rect 110940 26060 112000 27000
rect 105000 26000 112000 26060
rect 105000 25900 107000 26000
rect 100000 25840 107000 25900
rect 100000 25000 101060 25840
rect 95940 5960 96000 25000
rect 91000 5900 96000 5960
rect 101000 5960 101060 25000
rect 105940 25000 107000 25840
rect 110000 25900 112000 26000
rect 115000 26060 116060 27000
rect 120940 27000 121000 45940
rect 126000 45940 131000 46000
rect 126000 27000 126060 45940
rect 120940 26060 122000 27000
rect 115000 26000 122000 26060
rect 115000 25900 117000 26000
rect 110000 25840 117000 25900
rect 110000 25000 111060 25840
rect 105940 5960 106000 25000
rect 101000 5900 106000 5960
rect 111000 5960 111060 25000
rect 115940 25000 117000 25840
rect 120000 25900 122000 26000
rect 125000 26060 126060 27000
rect 130940 27000 131000 45940
rect 136000 45940 141000 46000
rect 136000 27000 136060 45940
rect 130940 26060 132000 27000
rect 125000 26000 132000 26060
rect 125000 25900 127000 26000
rect 120000 25840 127000 25900
rect 120000 25000 121060 25840
rect 115940 5960 116000 25000
rect 111000 5900 116000 5960
rect 121000 5960 121060 25000
rect 125940 25000 127000 25840
rect 130000 25900 132000 26000
rect 135000 26060 136060 27000
rect 140940 27000 141000 45940
rect 146000 45940 151000 46000
rect 146000 27000 146060 45940
rect 140940 26060 142000 27000
rect 135000 26000 142000 26060
rect 135000 25900 137000 26000
rect 130000 25840 137000 25900
rect 130000 25000 131060 25840
rect 125940 5960 126000 25000
rect 121000 5900 126000 5960
rect 131000 5960 131060 25000
rect 135940 25000 137000 25840
rect 140000 25900 142000 26000
rect 145000 26060 146060 27000
rect 150940 27000 151000 45940
rect 156000 45940 161000 46000
rect 156000 27000 156060 45940
rect 150940 26060 152000 27000
rect 145000 26000 152000 26060
rect 145000 25900 147000 26000
rect 140000 25840 147000 25900
rect 140000 25000 141060 25840
rect 135940 5960 136000 25000
rect 131000 5900 136000 5960
rect 141000 5960 141060 25000
rect 145940 25000 147000 25840
rect 150000 25900 152000 26000
rect 155000 26060 156060 27000
rect 160940 27000 161000 45940
rect 166000 45940 171000 46000
rect 166000 27000 166060 45940
rect 160940 26060 162000 27000
rect 155000 26000 162000 26060
rect 155000 25900 157000 26000
rect 150000 25840 157000 25900
rect 150000 25000 151060 25840
rect 145940 5960 146000 25000
rect 141000 5900 146000 5960
rect 151000 5960 151060 25000
rect 155940 25000 157000 25840
rect 160000 25900 162000 26000
rect 165000 26060 166060 27000
rect 170940 27000 171000 45940
rect 176000 45940 181000 46000
rect 176000 27000 176060 45940
rect 170940 26060 172000 27000
rect 165000 26000 172000 26060
rect 165000 25900 167000 26000
rect 160000 25840 167000 25900
rect 160000 25000 161060 25840
rect 155940 5960 156000 25000
rect 151000 5900 156000 5960
rect 161000 5960 161060 25000
rect 165940 25000 167000 25840
rect 170000 25900 172000 26000
rect 175000 26060 176060 27000
rect 180940 27000 181000 45940
rect 186000 45940 191000 46000
rect 186000 27000 186060 45940
rect 180940 26060 182000 27000
rect 175000 26000 182000 26060
rect 175000 25900 177000 26000
rect 170000 25840 177000 25900
rect 170000 25000 171060 25840
rect 165940 5960 166000 25000
rect 161000 5900 166000 5960
rect 171000 5960 171060 25000
rect 175940 25000 177000 25840
rect 180000 25900 182000 26000
rect 185000 26060 186060 27000
rect 190940 27000 191000 45940
rect 196000 45940 201000 46000
rect 196000 27000 196060 45940
rect 190940 26060 192000 27000
rect 185000 26000 192000 26060
rect 185000 25900 187000 26000
rect 180000 25840 187000 25900
rect 180000 25000 181060 25840
rect 175940 5960 176000 25000
rect 171000 5900 176000 5960
rect 181000 5960 181060 25000
rect 185940 25000 187000 25840
rect 190000 25900 192000 26000
rect 195000 26060 196060 27000
rect 200940 27000 201000 45940
rect 206000 45940 211000 46000
rect 206000 27000 206060 45940
rect 200940 26060 202000 27000
rect 195000 26000 202000 26060
rect 195000 25900 197000 26000
rect 190000 25840 197000 25900
rect 190000 25000 191060 25840
rect 185940 5960 186000 25000
rect 181000 5900 186000 5960
rect 191000 5960 191060 25000
rect 195940 25000 197000 25840
rect 200000 25900 202000 26000
rect 205000 26060 206060 27000
rect 210940 27000 211000 45940
rect 216000 45940 221000 46000
rect 216000 27000 216060 45940
rect 210940 26060 212000 27000
rect 205000 26000 212000 26060
rect 205000 25900 207000 26000
rect 200000 25840 207000 25900
rect 200000 25000 201060 25840
rect 195940 5960 196000 25000
rect 191000 5900 196000 5960
rect 201000 5960 201060 25000
rect 205940 25000 207000 25840
rect 210000 25900 212000 26000
rect 215000 26060 216060 27000
rect 220940 27000 221000 45940
rect 226000 45940 231000 46000
rect 226000 27000 226060 45940
rect 220940 26060 222000 27000
rect 215000 26000 222000 26060
rect 215000 25900 217000 26000
rect 210000 25840 217000 25900
rect 210000 25000 211060 25840
rect 205940 5960 206000 25000
rect 201000 5900 206000 5960
rect 211000 5960 211060 25000
rect 215940 25000 217000 25840
rect 220000 25900 222000 26000
rect 225000 26060 226060 27000
rect 230940 27000 231000 45940
rect 236000 45940 241000 46000
rect 236000 27000 236060 45940
rect 230940 26060 232000 27000
rect 225000 26000 232000 26060
rect 225000 25900 227000 26000
rect 220000 25840 227000 25900
rect 220000 25000 221060 25840
rect 215940 5960 216000 25000
rect 211000 5900 216000 5960
rect 221000 5960 221060 25000
rect 225940 25000 227000 25840
rect 230000 25900 232000 26000
rect 235000 26060 236060 27000
rect 240940 27000 241000 45940
rect 246000 45940 251000 46000
rect 246000 27000 246060 45940
rect 240940 26060 242000 27000
rect 235000 26000 242000 26060
rect 235000 25900 237000 26000
rect 230000 25840 237000 25900
rect 230000 25000 231060 25840
rect 225940 5960 226000 25000
rect 221000 5900 226000 5960
rect 231000 5960 231060 25000
rect 235940 25000 237000 25840
rect 240000 25900 242000 26000
rect 245000 26060 246060 27000
rect 250940 27000 251000 45940
rect 256000 45940 261000 46000
rect 256000 27000 256060 45940
rect 250940 26060 252000 27000
rect 245000 26000 252000 26060
rect 245000 25900 247000 26000
rect 240000 25840 247000 25900
rect 240000 25000 241060 25840
rect 235940 5960 236000 25000
rect 231000 5900 236000 5960
rect 241000 5960 241060 25000
rect 245940 25000 247000 25840
rect 250000 25900 252000 26000
rect 255000 26060 256060 27000
rect 260940 27000 261000 45940
rect 266000 45940 271000 46000
rect 266000 27000 266060 45940
rect 260940 26060 262000 27000
rect 255000 26000 262000 26060
rect 255000 25900 257000 26000
rect 250000 25840 257000 25900
rect 250000 25000 251060 25840
rect 245940 5960 246000 25000
rect 241000 5900 246000 5960
rect 251000 5960 251060 25000
rect 255940 25000 257000 25840
rect 260000 25900 262000 26000
rect 265000 26060 266060 27000
rect 270940 27000 271000 45940
rect 276000 45940 281000 46000
rect 276000 27000 276060 45940
rect 270940 26060 272000 27000
rect 265000 26000 272000 26060
rect 265000 25900 267000 26000
rect 260000 25840 267000 25900
rect 260000 25000 261060 25840
rect 255940 5960 256000 25000
rect 251000 5900 256000 5960
rect 261000 5960 261060 25000
rect 265940 25000 267000 25840
rect 270000 25900 272000 26000
rect 275000 26060 276060 27000
rect 280940 27000 281000 45940
rect 280940 26060 282000 27000
rect 275000 26000 282000 26060
rect 275000 25900 277000 26000
rect 270000 25840 277000 25900
rect 270000 25000 271060 25840
rect 265940 5960 266000 25000
rect 261000 5900 266000 5960
rect 271000 5960 271060 25000
rect 275940 25000 277000 25840
rect 280000 25900 282000 26000
rect 285000 25900 287000 27000
rect 280000 25840 287000 25900
rect 280000 25000 281060 25840
rect 275940 5960 276000 25000
rect 271000 5900 276000 5960
rect 281000 5960 281060 25000
rect 285940 25000 287000 25840
rect 285940 5960 286000 25000
rect 281000 5900 286000 5960
rect 46000 5660 286000 5700
rect 46000 5340 47000 5660
rect 55960 5340 57000 5660
rect 65960 5340 67000 5660
rect 75960 5340 77000 5660
rect 85960 5340 87000 5660
rect 95960 5340 97000 5660
rect 105960 5340 107000 5660
rect 115960 5340 117000 5660
rect 125960 5340 127000 5660
rect 135960 5340 137000 5660
rect 145960 5340 147000 5660
rect 155960 5340 157000 5660
rect 165960 5340 167000 5660
rect 175960 5340 177000 5660
rect 185960 5340 187000 5660
rect 195960 5340 197000 5660
rect 205960 5340 207000 5660
rect 215960 5340 217000 5660
rect 225960 5340 227000 5660
rect 235960 5340 237000 5660
rect 245960 5340 247000 5660
rect 255960 5340 257000 5660
rect 265960 5340 267000 5660
rect 275960 5340 277000 5660
rect 285960 5340 286000 5660
rect 46000 5300 286000 5340
<< via4 >>
rect 47000 46240 55000 46560
rect 57000 46240 65000 46560
rect 67000 46240 75000 46560
rect 77000 46240 85000 46560
rect 87000 46240 95000 46560
rect 97000 46240 105000 46560
rect 107000 46240 115000 46560
rect 117000 46240 125000 46560
rect 127000 46240 135000 46560
rect 137000 46240 145000 46560
rect 147000 46240 155000 46560
rect 157000 46240 165000 46560
rect 167000 46240 175000 46560
rect 177000 46240 185000 46560
rect 187000 46240 195000 46560
rect 197000 46240 205000 46560
rect 207000 46240 215000 46560
rect 217000 46240 225000 46560
rect 227000 46240 235000 46560
rect 237000 46240 245000 46560
rect 247000 46240 255000 46560
rect 257000 46240 265000 46560
rect 267000 46240 275000 46560
rect 277000 46240 285000 46560
rect 47000 5340 55000 5660
rect 57000 5340 65000 5660
rect 67000 5340 75000 5660
rect 77000 5340 85000 5660
rect 87000 5340 95000 5660
rect 97000 5340 105000 5660
rect 107000 5340 115000 5660
rect 117000 5340 125000 5660
rect 127000 5340 135000 5660
rect 137000 5340 145000 5660
rect 147000 5340 155000 5660
rect 157000 5340 165000 5660
rect 167000 5340 175000 5660
rect 177000 5340 185000 5660
rect 187000 5340 195000 5660
rect 197000 5340 205000 5660
rect 207000 5340 215000 5660
rect 217000 5340 225000 5660
rect 227000 5340 235000 5660
rect 237000 5340 245000 5660
rect 247000 5340 255000 5660
rect 257000 5340 265000 5660
rect 267000 5340 275000 5660
rect 277000 5340 285000 5660
<< mimcap2 >>
rect 46040 45940 50960 45960
rect 46040 26060 46060 45940
rect 50940 26060 50960 45940
rect 46040 26040 50960 26060
rect 56040 45940 60960 45960
rect 56040 26060 56060 45940
rect 60940 26060 60960 45940
rect 56040 26040 60960 26060
rect 66040 45940 70960 45960
rect 66040 26060 66060 45940
rect 70940 26060 70960 45940
rect 66040 26040 70960 26060
rect 76040 45940 80960 45960
rect 76040 26060 76060 45940
rect 80940 26060 80960 45940
rect 76040 26040 80960 26060
rect 86040 45940 90960 45960
rect 86040 26060 86060 45940
rect 90940 26060 90960 45940
rect 86040 26040 90960 26060
rect 96040 45940 100960 45960
rect 96040 26060 96060 45940
rect 100940 26060 100960 45940
rect 96040 26040 100960 26060
rect 106040 45940 110960 45960
rect 106040 26060 106060 45940
rect 110940 26060 110960 45940
rect 106040 26040 110960 26060
rect 116040 45940 120960 45960
rect 116040 26060 116060 45940
rect 120940 26060 120960 45940
rect 116040 26040 120960 26060
rect 126040 45940 130960 45960
rect 126040 26060 126060 45940
rect 130940 26060 130960 45940
rect 126040 26040 130960 26060
rect 136040 45940 140960 45960
rect 136040 26060 136060 45940
rect 140940 26060 140960 45940
rect 136040 26040 140960 26060
rect 146040 45940 150960 45960
rect 146040 26060 146060 45940
rect 150940 26060 150960 45940
rect 146040 26040 150960 26060
rect 156040 45940 160960 45960
rect 156040 26060 156060 45940
rect 160940 26060 160960 45940
rect 156040 26040 160960 26060
rect 166040 45940 170960 45960
rect 166040 26060 166060 45940
rect 170940 26060 170960 45940
rect 166040 26040 170960 26060
rect 176040 45940 180960 45960
rect 176040 26060 176060 45940
rect 180940 26060 180960 45940
rect 176040 26040 180960 26060
rect 186040 45940 190960 45960
rect 186040 26060 186060 45940
rect 190940 26060 190960 45940
rect 186040 26040 190960 26060
rect 196040 45940 200960 45960
rect 196040 26060 196060 45940
rect 200940 26060 200960 45940
rect 196040 26040 200960 26060
rect 206040 45940 210960 45960
rect 206040 26060 206060 45940
rect 210940 26060 210960 45940
rect 206040 26040 210960 26060
rect 216040 45940 220960 45960
rect 216040 26060 216060 45940
rect 220940 26060 220960 45940
rect 216040 26040 220960 26060
rect 226040 45940 230960 45960
rect 226040 26060 226060 45940
rect 230940 26060 230960 45940
rect 226040 26040 230960 26060
rect 236040 45940 240960 45960
rect 236040 26060 236060 45940
rect 240940 26060 240960 45940
rect 236040 26040 240960 26060
rect 246040 45940 250960 45960
rect 246040 26060 246060 45940
rect 250940 26060 250960 45940
rect 246040 26040 250960 26060
rect 256040 45940 260960 45960
rect 256040 26060 256060 45940
rect 260940 26060 260960 45940
rect 256040 26040 260960 26060
rect 266040 45940 270960 45960
rect 266040 26060 266060 45940
rect 270940 26060 270960 45940
rect 266040 26040 270960 26060
rect 276040 45940 280960 45960
rect 276040 26060 276060 45940
rect 280940 26060 280960 45940
rect 276040 26040 280960 26060
rect 51040 25840 55960 25860
rect 51040 5960 51060 25840
rect 55940 5960 55960 25840
rect 51040 5940 55960 5960
rect 61040 25840 65960 25860
rect 61040 5960 61060 25840
rect 65940 5960 65960 25840
rect 61040 5940 65960 5960
rect 71040 25840 75960 25860
rect 71040 5960 71060 25840
rect 75940 5960 75960 25840
rect 71040 5940 75960 5960
rect 81040 25840 85960 25860
rect 81040 5960 81060 25840
rect 85940 5960 85960 25840
rect 81040 5940 85960 5960
rect 91040 25840 95960 25860
rect 91040 5960 91060 25840
rect 95940 5960 95960 25840
rect 91040 5940 95960 5960
rect 101040 25840 105960 25860
rect 101040 5960 101060 25840
rect 105940 5960 105960 25840
rect 101040 5940 105960 5960
rect 111040 25840 115960 25860
rect 111040 5960 111060 25840
rect 115940 5960 115960 25840
rect 111040 5940 115960 5960
rect 121040 25840 125960 25860
rect 121040 5960 121060 25840
rect 125940 5960 125960 25840
rect 121040 5940 125960 5960
rect 131040 25840 135960 25860
rect 131040 5960 131060 25840
rect 135940 5960 135960 25840
rect 131040 5940 135960 5960
rect 141040 25840 145960 25860
rect 141040 5960 141060 25840
rect 145940 5960 145960 25840
rect 141040 5940 145960 5960
rect 151040 25840 155960 25860
rect 151040 5960 151060 25840
rect 155940 5960 155960 25840
rect 151040 5940 155960 5960
rect 161040 25840 165960 25860
rect 161040 5960 161060 25840
rect 165940 5960 165960 25840
rect 161040 5940 165960 5960
rect 171040 25840 175960 25860
rect 171040 5960 171060 25840
rect 175940 5960 175960 25840
rect 171040 5940 175960 5960
rect 181040 25840 185960 25860
rect 181040 5960 181060 25840
rect 185940 5960 185960 25840
rect 181040 5940 185960 5960
rect 191040 25840 195960 25860
rect 191040 5960 191060 25840
rect 195940 5960 195960 25840
rect 191040 5940 195960 5960
rect 201040 25840 205960 25860
rect 201040 5960 201060 25840
rect 205940 5960 205960 25840
rect 201040 5940 205960 5960
rect 211040 25840 215960 25860
rect 211040 5960 211060 25840
rect 215940 5960 215960 25840
rect 211040 5940 215960 5960
rect 221040 25840 225960 25860
rect 221040 5960 221060 25840
rect 225940 5960 225960 25840
rect 221040 5940 225960 5960
rect 231040 25840 235960 25860
rect 231040 5960 231060 25840
rect 235940 5960 235960 25840
rect 231040 5940 235960 5960
rect 241040 25840 245960 25860
rect 241040 5960 241060 25840
rect 245940 5960 245960 25840
rect 241040 5940 245960 5960
rect 251040 25840 255960 25860
rect 251040 5960 251060 25840
rect 255940 5960 255960 25840
rect 251040 5940 255960 5960
rect 261040 25840 265960 25860
rect 261040 5960 261060 25840
rect 265940 5960 265960 25840
rect 261040 5940 265960 5960
rect 271040 25840 275960 25860
rect 271040 5960 271060 25840
rect 275940 5960 275960 25840
rect 271040 5940 275960 5960
rect 281040 25840 285960 25860
rect 281040 5960 281060 25840
rect 285940 5960 285960 25840
rect 281040 5940 285960 5960
<< mimcap2contact >>
rect 46060 26060 50940 45940
rect 56060 26060 60940 45940
rect 66060 26060 70940 45940
rect 76060 26060 80940 45940
rect 86060 26060 90940 45940
rect 96060 26060 100940 45940
rect 106060 26060 110940 45940
rect 116060 26060 120940 45940
rect 126060 26060 130940 45940
rect 136060 26060 140940 45940
rect 146060 26060 150940 45940
rect 156060 26060 160940 45940
rect 166060 26060 170940 45940
rect 176060 26060 180940 45940
rect 186060 26060 190940 45940
rect 196060 26060 200940 45940
rect 206060 26060 210940 45940
rect 216060 26060 220940 45940
rect 226060 26060 230940 45940
rect 236060 26060 240940 45940
rect 246060 26060 250940 45940
rect 256060 26060 260940 45940
rect 266060 26060 270940 45940
rect 276060 26060 280940 45940
rect 51060 5960 55940 25840
rect 61060 5960 65940 25840
rect 71060 5960 75940 25840
rect 81060 5960 85940 25840
rect 91060 5960 95940 25840
rect 101060 5960 105940 25840
rect 111060 5960 115940 25840
rect 121060 5960 125940 25840
rect 131060 5960 135940 25840
rect 141060 5960 145940 25840
rect 151060 5960 155940 25840
rect 161060 5960 165940 25840
rect 171060 5960 175940 25840
rect 181060 5960 185940 25840
rect 191060 5960 195940 25840
rect 201060 5960 205940 25840
rect 211060 5960 215940 25840
rect 221060 5960 225940 25840
rect 231060 5960 235940 25840
rect 241060 5960 245940 25840
rect 251060 5960 255940 25840
rect 261060 5960 265940 25840
rect 271060 5960 275940 25840
rect 281060 5960 285940 25840
<< metal5 >>
rect 46000 46560 286000 46600
rect 46000 46240 47000 46560
rect 55000 46240 57000 46560
rect 65000 46240 67000 46560
rect 75000 46240 77000 46560
rect 85000 46240 87000 46560
rect 95000 46240 97000 46560
rect 105000 46240 107000 46560
rect 115000 46240 117000 46560
rect 125000 46240 127000 46560
rect 135000 46240 137000 46560
rect 145000 46240 147000 46560
rect 155000 46240 157000 46560
rect 165000 46240 167000 46560
rect 175000 46240 177000 46560
rect 185000 46240 187000 46560
rect 195000 46240 197000 46560
rect 205000 46240 207000 46560
rect 215000 46240 217000 46560
rect 225000 46240 227000 46560
rect 235000 46240 237000 46560
rect 245000 46240 247000 46560
rect 255000 46240 257000 46560
rect 265000 46240 267000 46560
rect 275000 46240 277000 46560
rect 285000 46240 286000 46560
rect 46000 46000 286000 46240
rect 46000 45940 51000 46000
rect 46000 26060 46060 45940
rect 50940 27000 51000 45940
rect 56000 45940 61000 46000
rect 56000 27000 56060 45940
rect 50940 26060 52000 27000
rect 46000 26000 52000 26060
rect 50000 25900 52000 26000
rect 55000 26060 56060 27000
rect 60940 27000 61000 45940
rect 66000 45940 71000 46000
rect 66000 27000 66060 45940
rect 60940 26060 62000 27000
rect 55000 26000 62000 26060
rect 55000 25900 57000 26000
rect 50000 25840 57000 25900
rect 50000 25000 51060 25840
rect 51000 5960 51060 25000
rect 55940 25000 57000 25840
rect 60000 25900 62000 26000
rect 65000 26060 66060 27000
rect 70940 27000 71000 45940
rect 76000 45940 81000 46000
rect 76000 27000 76060 45940
rect 70940 26060 72000 27000
rect 65000 26000 72000 26060
rect 65000 25900 67000 26000
rect 60000 25840 67000 25900
rect 60000 25000 61060 25840
rect 55940 5960 56000 25000
rect 51000 5900 56000 5960
rect 61000 5960 61060 25000
rect 65940 25000 67000 25840
rect 70000 25900 72000 26000
rect 75000 26060 76060 27000
rect 80940 27000 81000 45940
rect 86000 45940 91000 46000
rect 86000 27000 86060 45940
rect 80940 26060 82000 27000
rect 75000 26000 82000 26060
rect 75000 25900 77000 26000
rect 70000 25840 77000 25900
rect 70000 25000 71060 25840
rect 65940 5960 66000 25000
rect 61000 5900 66000 5960
rect 71000 5960 71060 25000
rect 75940 25000 77000 25840
rect 80000 25900 82000 26000
rect 85000 26060 86060 27000
rect 90940 27000 91000 45940
rect 96000 45940 101000 46000
rect 96000 27000 96060 45940
rect 90940 26060 92000 27000
rect 85000 26000 92000 26060
rect 85000 25900 87000 26000
rect 80000 25840 87000 25900
rect 80000 25000 81060 25840
rect 75940 5960 76000 25000
rect 71000 5900 76000 5960
rect 81000 5960 81060 25000
rect 85940 25000 87000 25840
rect 90000 25900 92000 26000
rect 95000 26060 96060 27000
rect 100940 27000 101000 45940
rect 106000 45940 111000 46000
rect 106000 27000 106060 45940
rect 100940 26060 102000 27000
rect 95000 26000 102000 26060
rect 95000 25900 97000 26000
rect 90000 25840 97000 25900
rect 90000 25000 91060 25840
rect 85940 5960 86000 25000
rect 81000 5900 86000 5960
rect 91000 5960 91060 25000
rect 95940 25000 97000 25840
rect 100000 25900 102000 26000
rect 105000 26060 106060 27000
rect 110940 27000 111000 45940
rect 116000 45940 121000 46000
rect 116000 27000 116060 45940
rect 110940 26060 112000 27000
rect 105000 26000 112000 26060
rect 105000 25900 107000 26000
rect 100000 25840 107000 25900
rect 100000 25000 101060 25840
rect 95940 5960 96000 25000
rect 91000 5900 96000 5960
rect 101000 5960 101060 25000
rect 105940 25000 107000 25840
rect 110000 25900 112000 26000
rect 115000 26060 116060 27000
rect 120940 27000 121000 45940
rect 126000 45940 131000 46000
rect 126000 27000 126060 45940
rect 120940 26060 122000 27000
rect 115000 26000 122000 26060
rect 115000 25900 117000 26000
rect 110000 25840 117000 25900
rect 110000 25000 111060 25840
rect 105940 5960 106000 25000
rect 101000 5900 106000 5960
rect 111000 5960 111060 25000
rect 115940 25000 117000 25840
rect 120000 25900 122000 26000
rect 125000 26060 126060 27000
rect 130940 27000 131000 45940
rect 136000 45940 141000 46000
rect 136000 27000 136060 45940
rect 130940 26060 132000 27000
rect 125000 26000 132000 26060
rect 125000 25900 127000 26000
rect 120000 25840 127000 25900
rect 120000 25000 121060 25840
rect 115940 5960 116000 25000
rect 111000 5900 116000 5960
rect 121000 5960 121060 25000
rect 125940 25000 127000 25840
rect 130000 25900 132000 26000
rect 135000 26060 136060 27000
rect 140940 27000 141000 45940
rect 146000 45940 151000 46000
rect 146000 27000 146060 45940
rect 140940 26060 142000 27000
rect 135000 26000 142000 26060
rect 135000 25900 137000 26000
rect 130000 25840 137000 25900
rect 130000 25000 131060 25840
rect 125940 5960 126000 25000
rect 121000 5900 126000 5960
rect 131000 5960 131060 25000
rect 135940 25000 137000 25840
rect 140000 25900 142000 26000
rect 145000 26060 146060 27000
rect 150940 27000 151000 45940
rect 156000 45940 161000 46000
rect 156000 27000 156060 45940
rect 150940 26060 152000 27000
rect 145000 26000 152000 26060
rect 145000 25900 147000 26000
rect 140000 25840 147000 25900
rect 140000 25000 141060 25840
rect 135940 5960 136000 25000
rect 131000 5900 136000 5960
rect 141000 5960 141060 25000
rect 145940 25000 147000 25840
rect 150000 25900 152000 26000
rect 155000 26060 156060 27000
rect 160940 27000 161000 45940
rect 166000 45940 171000 46000
rect 166000 27000 166060 45940
rect 160940 26060 162000 27000
rect 155000 26000 162000 26060
rect 155000 25900 157000 26000
rect 150000 25840 157000 25900
rect 150000 25000 151060 25840
rect 145940 5960 146000 25000
rect 141000 5900 146000 5960
rect 151000 5960 151060 25000
rect 155940 25000 157000 25840
rect 160000 25900 162000 26000
rect 165000 26060 166060 27000
rect 170940 27000 171000 45940
rect 176000 45940 181000 46000
rect 176000 27000 176060 45940
rect 170940 26060 172000 27000
rect 165000 26000 172000 26060
rect 165000 25900 167000 26000
rect 160000 25840 167000 25900
rect 160000 25000 161060 25840
rect 155940 5960 156000 25000
rect 151000 5900 156000 5960
rect 161000 5960 161060 25000
rect 165940 25000 167000 25840
rect 170000 25900 172000 26000
rect 175000 26060 176060 27000
rect 180940 27000 181000 45940
rect 186000 45940 191000 46000
rect 186000 27000 186060 45940
rect 180940 26060 182000 27000
rect 175000 26000 182000 26060
rect 175000 25900 177000 26000
rect 170000 25840 177000 25900
rect 170000 25000 171060 25840
rect 165940 5960 166000 25000
rect 161000 5900 166000 5960
rect 171000 5960 171060 25000
rect 175940 25000 177000 25840
rect 180000 25900 182000 26000
rect 185000 26060 186060 27000
rect 190940 27000 191000 45940
rect 196000 45940 201000 46000
rect 196000 27000 196060 45940
rect 190940 26060 192000 27000
rect 185000 26000 192000 26060
rect 185000 25900 187000 26000
rect 180000 25840 187000 25900
rect 180000 25000 181060 25840
rect 175940 5960 176000 25000
rect 171000 5900 176000 5960
rect 181000 5960 181060 25000
rect 185940 25000 187000 25840
rect 190000 25900 192000 26000
rect 195000 26060 196060 27000
rect 200940 27000 201000 45940
rect 206000 45940 211000 46000
rect 206000 27000 206060 45940
rect 200940 26060 202000 27000
rect 195000 26000 202000 26060
rect 195000 25900 197000 26000
rect 190000 25840 197000 25900
rect 190000 25000 191060 25840
rect 185940 5960 186000 25000
rect 181000 5900 186000 5960
rect 191000 5960 191060 25000
rect 195940 25000 197000 25840
rect 200000 25900 202000 26000
rect 205000 26060 206060 27000
rect 210940 27000 211000 45940
rect 216000 45940 221000 46000
rect 216000 27000 216060 45940
rect 210940 26060 212000 27000
rect 205000 26000 212000 26060
rect 205000 25900 207000 26000
rect 200000 25840 207000 25900
rect 200000 25000 201060 25840
rect 195940 5960 196000 25000
rect 191000 5900 196000 5960
rect 201000 5960 201060 25000
rect 205940 25000 207000 25840
rect 210000 25900 212000 26000
rect 215000 26060 216060 27000
rect 220940 27000 221000 45940
rect 226000 45940 231000 46000
rect 226000 27000 226060 45940
rect 220940 26060 222000 27000
rect 215000 26000 222000 26060
rect 215000 25900 217000 26000
rect 210000 25840 217000 25900
rect 210000 25000 211060 25840
rect 205940 5960 206000 25000
rect 201000 5900 206000 5960
rect 211000 5960 211060 25000
rect 215940 25000 217000 25840
rect 220000 25900 222000 26000
rect 225000 26060 226060 27000
rect 230940 27000 231000 45940
rect 236000 45940 241000 46000
rect 236000 27000 236060 45940
rect 230940 26060 232000 27000
rect 225000 26000 232000 26060
rect 225000 25900 227000 26000
rect 220000 25840 227000 25900
rect 220000 25000 221060 25840
rect 215940 5960 216000 25000
rect 211000 5900 216000 5960
rect 221000 5960 221060 25000
rect 225940 25000 227000 25840
rect 230000 25900 232000 26000
rect 235000 26060 236060 27000
rect 240940 27000 241000 45940
rect 246000 45940 251000 46000
rect 246000 27000 246060 45940
rect 240940 26060 242000 27000
rect 235000 26000 242000 26060
rect 235000 25900 237000 26000
rect 230000 25840 237000 25900
rect 230000 25000 231060 25840
rect 225940 5960 226000 25000
rect 221000 5900 226000 5960
rect 231000 5960 231060 25000
rect 235940 25000 237000 25840
rect 240000 25900 242000 26000
rect 245000 26060 246060 27000
rect 250940 27000 251000 45940
rect 256000 45940 261000 46000
rect 256000 27000 256060 45940
rect 250940 26060 252000 27000
rect 245000 26000 252000 26060
rect 245000 25900 247000 26000
rect 240000 25840 247000 25900
rect 240000 25000 241060 25840
rect 235940 5960 236000 25000
rect 231000 5900 236000 5960
rect 241000 5960 241060 25000
rect 245940 25000 247000 25840
rect 250000 25900 252000 26000
rect 255000 26060 256060 27000
rect 260940 27000 261000 45940
rect 266000 45940 271000 46000
rect 266000 27000 266060 45940
rect 260940 26060 262000 27000
rect 255000 26000 262000 26060
rect 255000 25900 257000 26000
rect 250000 25840 257000 25900
rect 250000 25000 251060 25840
rect 245940 5960 246000 25000
rect 241000 5900 246000 5960
rect 251000 5960 251060 25000
rect 255940 25000 257000 25840
rect 260000 25900 262000 26000
rect 265000 26060 266060 27000
rect 270940 27000 271000 45940
rect 276000 45940 281000 46000
rect 276000 27000 276060 45940
rect 270940 26060 272000 27000
rect 265000 26000 272000 26060
rect 265000 25900 267000 26000
rect 260000 25840 267000 25900
rect 260000 25000 261060 25840
rect 255940 5960 256000 25000
rect 251000 5900 256000 5960
rect 261000 5960 261060 25000
rect 265940 25000 267000 25840
rect 270000 25900 272000 26000
rect 275000 26060 276060 27000
rect 280940 27000 281000 45940
rect 280940 26060 282000 27000
rect 275000 26000 282000 26060
rect 275000 25900 277000 26000
rect 270000 25840 277000 25900
rect 270000 25000 271060 25840
rect 265940 5960 266000 25000
rect 261000 5900 266000 5960
rect 271000 5960 271060 25000
rect 275940 25000 277000 25840
rect 280000 25900 282000 26000
rect 285000 25900 287000 27000
rect 280000 25840 287000 25900
rect 280000 25000 281060 25840
rect 275940 5960 276000 25000
rect 271000 5900 276000 5960
rect 281000 5960 281060 25000
rect 285940 25000 287000 25840
rect 285940 5960 286000 25000
rect 281000 5900 286000 5960
rect 46000 5660 286000 5900
rect 46000 5340 47000 5660
rect 55000 5340 57000 5660
rect 65000 5340 67000 5660
rect 75000 5340 77000 5660
rect 85000 5340 87000 5660
rect 95000 5340 97000 5660
rect 105000 5340 107000 5660
rect 115000 5340 117000 5660
rect 125000 5340 127000 5660
rect 135000 5340 137000 5660
rect 145000 5340 147000 5660
rect 155000 5340 157000 5660
rect 165000 5340 167000 5660
rect 175000 5340 177000 5660
rect 185000 5340 187000 5660
rect 195000 5340 197000 5660
rect 205000 5340 207000 5660
rect 215000 5340 217000 5660
rect 225000 5340 227000 5660
rect 235000 5340 237000 5660
rect 245000 5340 247000 5660
rect 255000 5340 257000 5660
rect 265000 5340 267000 5660
rect 275000 5340 277000 5660
rect 285000 5340 286000 5660
rect 46000 5300 286000 5340
use sky130_fd_pr__res_xhigh_po_0p35_FE9J4G  sky130_fd_pr__res_xhigh_po_0p35_FE9J4G_0
timestamp 1672019510
transform 0 1 56598 -1 0 48201
box -201 -10598 201 10598
<< end >>
