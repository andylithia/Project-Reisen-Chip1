** sch_path: /home/andylithia/openmpw/Project-Reisen-Chip1/xschem/CML_latch_1mA_transient_tb.sch
**.subckt CML_latch_1mA_transient_tb
V1 VDD GND 1.8
XM6 net1 vref GND GND sky130_fd_pr__nfet_01v8 L=1.2 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
I0 VDD vref 0.05m
XM3 vref vbias net1 GND sky130_fd_pr__nfet_01v8 L=1.2 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 net2 net2 GND GND sky130_fd_pr__nfet_01v8 L=1.2 W=0.7 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM7 vbias net3 net2 GND sky130_fd_pr__nfet_01v8 L=1.2 W=0.7 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM9 net3 net3 vbias GND sky130_fd_pr__nfet_01v8 L=1.2 W=0.7 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
R4 VDD net3 1k m=1
V8 cki GND PULSE(0 1.8 0 0.01n 0.01n 0.1n 0.2n)
x4 cki gnd gnd vdd vdd net4 sky130_fd_sc_hs__clkinv_8
x3 cki gnd gnd vdd vdd net5 sky130_fd_sc_hs__clkinv_4
x5 net5 gnd gnd vdd vdd ckbuf_p sky130_fd_sc_hs__clkinv_16
x6 net4 gnd gnd vdd vdd net6 sky130_fd_sc_hs__clkinv_8
x7 net6 gnd gnd vdd vdd ckbuf_n sky130_fd_sc_hs__clkinv_16
V4 vin GND PULSE(1.35 1.25 0 10n 0 1 2)
x1 VDD vop_i von_i vip vin ckbuf_p ckbuf_n vbias vref GND CML_latch_1mA
V2 vip GND PULSE(1.25 1.35 0 10n 0 1 2)
x2 VDD vop1_i von1_i vop_i von_i ckbuf_n ckbuf_p vbias vref GND CML_latch_1mA
x8 VDD vop2_i von2_i vop1_i von1_i ckbuf_p ckbuf_n vbias vref GND CML_latch_1mA
x9 VDD vop3_i von3_i vop2_i von2_i ckbuf_n ckbuf_p vbias vref GND CML_latch_1mA
**** begin user architecture code
.lib /home/andylithia/openmpw/pdk_1/sky130B/libs.tech/ngspice/sky130.lib.spice tt
.include /home/andylithia/openmpw/pdk_1/sky130B/libs.ref/sky130_fd_sc_hs/spice/sky130_fd_sc_hs.spice


.tran 100ps 10ns
.control
run
display
plot vop_i von_i
plot vop_i vop1_i vop2_i vop3_i ckbuf_p
plot ckbuf_p ckbuf_n
.endc


**** end user architecture code
**.ends

* expanding   symbol:  CML_latch_1mA.sym # of pins=10
** sym_path: /home/andylithia/openmpw/Project-Reisen-Chip1/xschem/CML_latch_1mA.sym
** sch_path: /home/andylithia/openmpw/Project-Reisen-Chip1/xschem/CML_latch_1mA.sch
.subckt CML_latch_1mA  vhi cml_q cml_qn vip vin ckin_amp ckin_hold vref_cas vref vlo
*.opin cml_q
*.opin cml_qn
*.iopin vhi
*.ipin ckin_amp
*.ipin ckin_hold
*.ipin vref_cas
*.ipin vref
*.iopin vlo
*.ipin vip
*.ipin vin
XM5 net1 vref vlo vlo sky130_fd_pr__nfet_01v8 L=1.2 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=20 m=20
XM2 vcenter vref_cas net1 vlo sky130_fd_pr__nfet_01v8 L=1.2 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=20 m=20
XM1 vmid_amp ckin_amp vcenter vlo sky130_fd_pr__nfet_01v8 L=0.15 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM8 vmid_hold ckin_hold vcenter vlo sky130_fd_pr__nfet_01v8 L=0.15 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM10 cml_qn vip vmid_amp vlo sky130_fd_pr__nfet_01v8 L=0.15 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM11 cml_q vin vmid_amp vlo sky130_fd_pr__nfet_01v8 L=0.15 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM12 cml_q cml_qn vmid_hold vlo sky130_fd_pr__nfet_01v8 L=0.15 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM13 cml_qn cml_q vmid_hold vlo sky130_fd_pr__nfet_01v8 L=0.15 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
R1 vhi cml_qn 1k m=1
R2 vhi cml_q 1k m=1
.ends

.GLOBAL GND
.GLOBAL VDD
.end
