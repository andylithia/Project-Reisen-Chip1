* NGSPICE file created from test_123.ext - technology: sky130A

X0 VSUBS G2 A VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X1 A G1 VSUBS VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
C0 G1 G2 0.01fF
C1 A G2 0.01fF
C2 G1 A 0.02fF
C3 A VSUBS 3.23fF $ **FLOATING
C4 G1 VSUBS 0.26fF $ **FLOATING
C5 G2 VSUBS 0.27fF $ **FLOATING
