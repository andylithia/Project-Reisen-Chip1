magic
tech sky130A
magscale 1 2
timestamp 1671381513
<< pwell >>
rect -307 -898 307 898
<< psubdiff >>
rect -271 828 -175 862
rect 175 828 271 862
rect -271 766 -237 828
rect 237 766 271 828
rect -271 -828 -237 -766
rect 237 -828 271 -766
rect -271 -862 -175 -828
rect 175 -862 271 -828
<< psubdiffcont >>
rect -175 828 175 862
rect -271 -766 -237 766
rect 237 -766 271 766
rect -175 -862 175 -828
<< xpolycontact >>
rect -141 300 141 732
rect -141 -732 141 -300
<< ppolyres >>
rect -141 -300 141 300
<< locali >>
rect -271 828 -175 862
rect 175 828 271 862
rect -271 766 -237 828
rect 237 766 271 828
rect -271 -828 -237 -766
rect 237 -828 271 -766
rect -271 -862 -175 -828
rect 175 -862 271 -828
<< viali >>
rect -125 317 125 714
rect -125 -714 125 -317
<< metal1 >>
rect -131 714 131 726
rect -131 317 -125 714
rect 125 317 131 714
rect -131 305 131 317
rect -131 -317 131 -305
rect -131 -714 -125 -317
rect 125 -714 131 -317
rect -131 -726 131 -714
<< res1p41 >>
rect -143 -302 143 302
<< properties >>
string FIXED_BBOX -254 -845 254 845
string gencell sky130_fd_pr__res_high_po_1p41
string library sky130
string parameters w 1.410 l 3 m 1 nx 1 wmin 1.410 lmin 0.50 rho 319.8 val 956.765 dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 1.410 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
