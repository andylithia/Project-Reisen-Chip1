magic
tech sky130A
magscale 1 2
timestamp 1672473348
<< obsli1 >>
rect 1104 2159 14812 27761
<< obsm1 >>
rect 750 2128 15166 27792
<< metal2 >>
rect 1766 29200 1822 30000
rect 2042 29200 2098 30000
rect 2318 29200 2374 30000
rect 2594 29200 2650 30000
rect 2870 29200 2926 30000
rect 3146 29200 3202 30000
rect 3422 29200 3478 30000
rect 3698 29200 3754 30000
rect 3974 29200 4030 30000
rect 4250 29200 4306 30000
rect 4526 29200 4582 30000
rect 4802 29200 4858 30000
rect 5078 29200 5134 30000
rect 5354 29200 5410 30000
rect 5630 29200 5686 30000
rect 5906 29200 5962 30000
rect 6182 29200 6238 30000
rect 6458 29200 6514 30000
rect 6734 29200 6790 30000
rect 7010 29200 7066 30000
rect 7286 29200 7342 30000
rect 7562 29200 7618 30000
rect 7838 29200 7894 30000
rect 8114 29200 8170 30000
rect 8390 29200 8446 30000
rect 8666 29200 8722 30000
rect 8942 29200 8998 30000
rect 9218 29200 9274 30000
rect 9494 29200 9550 30000
rect 9770 29200 9826 30000
rect 10046 29200 10102 30000
rect 10322 29200 10378 30000
rect 10598 29200 10654 30000
rect 10874 29200 10930 30000
rect 11150 29200 11206 30000
rect 11426 29200 11482 30000
rect 11702 29200 11758 30000
rect 11978 29200 12034 30000
rect 12254 29200 12310 30000
rect 12530 29200 12586 30000
rect 12806 29200 12862 30000
rect 13082 29200 13138 30000
rect 13358 29200 13414 30000
rect 13634 29200 13690 30000
rect 13910 29200 13966 30000
rect 14186 29200 14242 30000
rect 754 0 810 800
rect 1858 0 1914 800
rect 2962 0 3018 800
rect 4066 0 4122 800
rect 5170 0 5226 800
rect 6274 0 6330 800
rect 7378 0 7434 800
rect 8482 0 8538 800
rect 9586 0 9642 800
rect 10690 0 10746 800
rect 11794 0 11850 800
rect 12898 0 12954 800
rect 14002 0 14058 800
rect 15106 0 15162 800
<< obsm2 >>
rect 756 29144 1710 29322
rect 1878 29144 1986 29322
rect 2154 29144 2262 29322
rect 2430 29144 2538 29322
rect 2706 29144 2814 29322
rect 2982 29144 3090 29322
rect 3258 29144 3366 29322
rect 3534 29144 3642 29322
rect 3810 29144 3918 29322
rect 4086 29144 4194 29322
rect 4362 29144 4470 29322
rect 4638 29144 4746 29322
rect 4914 29144 5022 29322
rect 5190 29144 5298 29322
rect 5466 29144 5574 29322
rect 5742 29144 5850 29322
rect 6018 29144 6126 29322
rect 6294 29144 6402 29322
rect 6570 29144 6678 29322
rect 6846 29144 6954 29322
rect 7122 29144 7230 29322
rect 7398 29144 7506 29322
rect 7674 29144 7782 29322
rect 7950 29144 8058 29322
rect 8226 29144 8334 29322
rect 8502 29144 8610 29322
rect 8778 29144 8886 29322
rect 9054 29144 9162 29322
rect 9330 29144 9438 29322
rect 9606 29144 9714 29322
rect 9882 29144 9990 29322
rect 10158 29144 10266 29322
rect 10434 29144 10542 29322
rect 10710 29144 10818 29322
rect 10986 29144 11094 29322
rect 11262 29144 11370 29322
rect 11538 29144 11646 29322
rect 11814 29144 11922 29322
rect 12090 29144 12198 29322
rect 12366 29144 12474 29322
rect 12642 29144 12750 29322
rect 12918 29144 13026 29322
rect 13194 29144 13302 29322
rect 13470 29144 13578 29322
rect 13746 29144 13854 29322
rect 14022 29144 14130 29322
rect 14298 29144 15160 29322
rect 756 856 15160 29144
rect 866 800 1802 856
rect 1970 800 2906 856
rect 3074 800 4010 856
rect 4178 800 5114 856
rect 5282 800 6218 856
rect 6386 800 7322 856
rect 7490 800 8426 856
rect 8594 800 9530 856
rect 9698 800 10634 856
rect 10802 800 11738 856
rect 11906 800 12842 856
rect 13010 800 13946 856
rect 14114 800 15050 856
<< obsm3 >>
rect 2659 2143 14969 27777
<< metal4 >>
rect 2657 2128 2977 27792
rect 4370 2128 4690 27792
rect 6084 2128 6404 27792
rect 7797 2128 8117 27792
rect 9511 2128 9831 27792
rect 11224 2128 11544 27792
rect 12938 2128 13258 27792
rect 14651 2128 14971 27792
<< obsm4 >>
rect 7419 2483 7485 11117
<< labels >>
rlabel metal2 s 2962 0 3018 800 6 clk
port 1 nsew signal input
rlabel metal2 s 14002 0 14058 800 6 dac_in[0]
port 2 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 dac_in[1]
port 3 nsew signal input
rlabel metal2 s 11794 0 11850 800 6 dac_in[2]
port 4 nsew signal input
rlabel metal2 s 10690 0 10746 800 6 dac_in[3]
port 5 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 dac_in[4]
port 6 nsew signal input
rlabel metal2 s 8482 0 8538 800 6 dac_in[5]
port 7 nsew signal input
rlabel metal2 s 7378 0 7434 800 6 dac_in[6]
port 8 nsew signal input
rlabel metal2 s 6274 0 6330 800 6 dac_in[7]
port 9 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 dac_in[8]
port 10 nsew signal input
rlabel metal2 s 4066 0 4122 800 6 dac_in[9]
port 11 nsew signal input
rlabel metal2 s 15106 0 15162 800 6 dummy
port 12 nsew signal input
rlabel metal2 s 14186 29200 14242 30000 6 llsb
port 13 nsew signal output
rlabel metal2 s 13910 29200 13966 30000 6 llsb_n
port 14 nsew signal output
rlabel metal2 s 13634 29200 13690 30000 6 lsb[0]
port 15 nsew signal output
rlabel metal2 s 13082 29200 13138 30000 6 lsb[1]
port 16 nsew signal output
rlabel metal2 s 12530 29200 12586 30000 6 lsb[2]
port 17 nsew signal output
rlabel metal2 s 11978 29200 12034 30000 6 lsb[3]
port 18 nsew signal output
rlabel metal2 s 11426 29200 11482 30000 6 lsb[4]
port 19 nsew signal output
rlabel metal2 s 10874 29200 10930 30000 6 lsb[5]
port 20 nsew signal output
rlabel metal2 s 13358 29200 13414 30000 6 lsb_n[0]
port 21 nsew signal output
rlabel metal2 s 12806 29200 12862 30000 6 lsb_n[1]
port 22 nsew signal output
rlabel metal2 s 12254 29200 12310 30000 6 lsb_n[2]
port 23 nsew signal output
rlabel metal2 s 11702 29200 11758 30000 6 lsb_n[3]
port 24 nsew signal output
rlabel metal2 s 11150 29200 11206 30000 6 lsb_n[4]
port 25 nsew signal output
rlabel metal2 s 10598 29200 10654 30000 6 lsb_n[5]
port 26 nsew signal output
rlabel metal2 s 10322 29200 10378 30000 6 msb[0]
port 27 nsew signal output
rlabel metal2 s 4802 29200 4858 30000 6 msb[10]
port 28 nsew signal output
rlabel metal2 s 4250 29200 4306 30000 6 msb[11]
port 29 nsew signal output
rlabel metal2 s 3698 29200 3754 30000 6 msb[12]
port 30 nsew signal output
rlabel metal2 s 3146 29200 3202 30000 6 msb[13]
port 31 nsew signal output
rlabel metal2 s 2594 29200 2650 30000 6 msb[14]
port 32 nsew signal output
rlabel metal2 s 2042 29200 2098 30000 6 msb[15]
port 33 nsew signal output
rlabel metal2 s 9770 29200 9826 30000 6 msb[1]
port 34 nsew signal output
rlabel metal2 s 9218 29200 9274 30000 6 msb[2]
port 35 nsew signal output
rlabel metal2 s 8666 29200 8722 30000 6 msb[3]
port 36 nsew signal output
rlabel metal2 s 8114 29200 8170 30000 6 msb[4]
port 37 nsew signal output
rlabel metal2 s 7562 29200 7618 30000 6 msb[5]
port 38 nsew signal output
rlabel metal2 s 7010 29200 7066 30000 6 msb[6]
port 39 nsew signal output
rlabel metal2 s 6458 29200 6514 30000 6 msb[7]
port 40 nsew signal output
rlabel metal2 s 5906 29200 5962 30000 6 msb[8]
port 41 nsew signal output
rlabel metal2 s 5354 29200 5410 30000 6 msb[9]
port 42 nsew signal output
rlabel metal2 s 10046 29200 10102 30000 6 msb_n[0]
port 43 nsew signal output
rlabel metal2 s 4526 29200 4582 30000 6 msb_n[10]
port 44 nsew signal output
rlabel metal2 s 3974 29200 4030 30000 6 msb_n[11]
port 45 nsew signal output
rlabel metal2 s 3422 29200 3478 30000 6 msb_n[12]
port 46 nsew signal output
rlabel metal2 s 2870 29200 2926 30000 6 msb_n[13]
port 47 nsew signal output
rlabel metal2 s 2318 29200 2374 30000 6 msb_n[14]
port 48 nsew signal output
rlabel metal2 s 1766 29200 1822 30000 6 msb_n[15]
port 49 nsew signal output
rlabel metal2 s 9494 29200 9550 30000 6 msb_n[1]
port 50 nsew signal output
rlabel metal2 s 8942 29200 8998 30000 6 msb_n[2]
port 51 nsew signal output
rlabel metal2 s 8390 29200 8446 30000 6 msb_n[3]
port 52 nsew signal output
rlabel metal2 s 7838 29200 7894 30000 6 msb_n[4]
port 53 nsew signal output
rlabel metal2 s 7286 29200 7342 30000 6 msb_n[5]
port 54 nsew signal output
rlabel metal2 s 6734 29200 6790 30000 6 msb_n[6]
port 55 nsew signal output
rlabel metal2 s 6182 29200 6238 30000 6 msb_n[7]
port 56 nsew signal output
rlabel metal2 s 5630 29200 5686 30000 6 msb_n[8]
port 57 nsew signal output
rlabel metal2 s 5078 29200 5134 30000 6 msb_n[9]
port 58 nsew signal output
rlabel metal2 s 1858 0 1914 800 6 rst_n
port 59 nsew signal input
rlabel metal2 s 754 0 810 800 6 test_mode
port 60 nsew signal input
rlabel metal4 s 2657 2128 2977 27792 6 vccd1
port 61 nsew power bidirectional
rlabel metal4 s 6084 2128 6404 27792 6 vccd1
port 61 nsew power bidirectional
rlabel metal4 s 9511 2128 9831 27792 6 vccd1
port 61 nsew power bidirectional
rlabel metal4 s 12938 2128 13258 27792 6 vccd1
port 61 nsew power bidirectional
rlabel metal4 s 4370 2128 4690 27792 6 vssd1
port 62 nsew ground bidirectional
rlabel metal4 s 7797 2128 8117 27792 6 vssd1
port 62 nsew ground bidirectional
rlabel metal4 s 11224 2128 11544 27792 6 vssd1
port 62 nsew ground bidirectional
rlabel metal4 s 14651 2128 14971 27792 6 vssd1
port 62 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 16000 30000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 820498
string GDS_FILE /home/andylithia/openmpw/Project-Reisen-Chip1_digital/openlane/dac_con/runs/22_12_31_02_55/results/signoff/dac_con.magic.gds
string GDS_START 157264
<< end >>

