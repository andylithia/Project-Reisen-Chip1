magic
tech sky130A
magscale 1 2
timestamp 1671823962
<< nwell >>
rect 96 284 1708 656
<< pwell >>
rect 139 -10 225 207
rect 231 1 421 228
rect 423 1 613 228
rect 619 1 1093 200
rect 1095 1 1573 200
rect 230 -48 1574 1
rect 1579 -10 1665 207
<< scpmos >>
rect 699 344 729 544
rect 789 344 819 544
rect 890 320 920 544
rect 980 320 1010 544
rect 1181 320 1211 544
rect 1271 320 1301 544
rect 1363 320 1393 544
rect 1453 320 1483 544
<< nmoslvt >>
rect 702 26 732 174
rect 780 26 810 174
rect 882 26 912 174
rect 968 26 998 174
rect 1178 26 1208 174
rect 1274 26 1304 174
rect 1360 26 1390 174
rect 1456 26 1486 174
<< ndiff >>
rect 645 162 702 174
rect 645 128 657 162
rect 691 128 702 162
rect 645 72 702 128
rect 645 38 657 72
rect 691 38 702 72
rect 645 26 702 38
rect 732 26 780 174
rect 810 83 882 174
rect 810 49 821 83
rect 855 49 882 83
rect 810 26 882 49
rect 912 83 968 174
rect 912 49 923 83
rect 957 49 968 83
rect 912 26 968 49
rect 998 72 1067 174
rect 998 38 1015 72
rect 1049 38 1067 72
rect 998 26 1067 38
rect 1121 162 1178 174
rect 1121 128 1133 162
rect 1167 128 1178 162
rect 1121 72 1178 128
rect 1121 38 1133 72
rect 1167 38 1178 72
rect 1121 26 1178 38
rect 1208 88 1274 174
rect 1208 54 1219 88
rect 1253 54 1274 88
rect 1208 26 1274 54
rect 1304 162 1360 174
rect 1304 128 1315 162
rect 1349 128 1360 162
rect 1304 72 1360 128
rect 1304 38 1315 72
rect 1349 38 1360 72
rect 1304 26 1360 38
rect 1390 141 1456 174
rect 1390 107 1401 141
rect 1435 107 1456 141
rect 1390 26 1456 107
rect 1486 88 1547 174
rect 1486 54 1501 88
rect 1535 54 1547 88
rect 1486 26 1547 54
<< pdiff >>
rect 641 532 699 544
rect 641 498 652 532
rect 686 498 699 532
rect 641 462 699 498
rect 641 428 652 462
rect 686 428 699 462
rect 641 392 699 428
rect 641 358 652 392
rect 686 358 699 392
rect 641 344 699 358
rect 729 532 789 544
rect 729 498 742 532
rect 776 498 789 532
rect 729 462 789 498
rect 729 428 742 462
rect 776 428 789 462
rect 729 392 789 428
rect 729 358 742 392
rect 776 358 789 392
rect 729 344 789 358
rect 819 532 890 544
rect 819 498 842 532
rect 876 498 890 532
rect 819 460 890 498
rect 819 426 842 460
rect 876 426 890 460
rect 819 344 890 426
rect 837 320 890 344
rect 920 532 980 544
rect 920 498 933 532
rect 967 498 980 532
rect 920 449 980 498
rect 920 415 933 449
rect 967 415 980 449
rect 920 366 980 415
rect 920 332 933 366
rect 967 332 980 366
rect 920 320 980 332
rect 1010 532 1067 544
rect 1010 498 1023 532
rect 1057 498 1067 532
rect 1010 414 1067 498
rect 1010 380 1023 414
rect 1057 380 1067 414
rect 1010 320 1067 380
rect 1122 532 1181 544
rect 1122 498 1134 532
rect 1168 498 1181 532
rect 1122 449 1181 498
rect 1122 415 1134 449
rect 1168 415 1181 449
rect 1122 366 1181 415
rect 1122 332 1134 366
rect 1168 332 1181 366
rect 1122 320 1181 332
rect 1211 532 1271 544
rect 1211 498 1224 532
rect 1258 498 1271 532
rect 1211 462 1271 498
rect 1211 428 1224 462
rect 1258 428 1271 462
rect 1211 392 1271 428
rect 1211 358 1224 392
rect 1258 358 1271 392
rect 1211 320 1271 358
rect 1301 532 1363 544
rect 1301 498 1314 532
rect 1348 498 1363 532
rect 1301 460 1363 498
rect 1301 426 1314 460
rect 1348 426 1363 460
rect 1301 320 1363 426
rect 1393 532 1453 544
rect 1393 498 1406 532
rect 1440 498 1453 532
rect 1393 462 1453 498
rect 1393 428 1406 462
rect 1440 428 1453 462
rect 1393 392 1453 428
rect 1393 358 1406 392
rect 1440 358 1453 392
rect 1393 320 1453 358
rect 1483 532 1542 544
rect 1483 498 1496 532
rect 1530 498 1542 532
rect 1483 460 1542 498
rect 1483 426 1496 460
rect 1530 426 1542 460
rect 1483 320 1542 426
<< ndiffc >>
rect 657 128 691 162
rect 657 38 691 72
rect 821 49 855 83
rect 923 49 957 83
rect 1015 38 1049 72
rect 1133 128 1167 162
rect 1133 38 1167 72
rect 1219 54 1253 88
rect 1315 128 1349 162
rect 1315 38 1349 72
rect 1401 107 1435 141
rect 1501 54 1535 88
<< pdiffc >>
rect 652 498 686 532
rect 652 428 686 462
rect 652 358 686 392
rect 742 498 776 532
rect 742 428 776 462
rect 742 358 776 392
rect 842 498 876 532
rect 842 426 876 460
rect 933 498 967 532
rect 933 415 967 449
rect 933 332 967 366
rect 1023 498 1057 532
rect 1023 380 1057 414
rect 1134 498 1168 532
rect 1134 415 1168 449
rect 1134 332 1168 366
rect 1224 498 1258 532
rect 1224 428 1258 462
rect 1224 358 1258 392
rect 1314 498 1348 532
rect 1314 426 1348 460
rect 1406 498 1440 532
rect 1406 428 1440 462
rect 1406 358 1440 392
rect 1496 498 1530 532
rect 1496 426 1530 460
<< psubdiff >>
rect 165 157 199 181
rect 165 74 199 123
rect 165 16 199 40
rect 1605 157 1639 181
rect 1605 74 1639 123
rect 1605 16 1639 40
<< nsubdiff >>
rect 165 530 199 554
rect 165 444 199 496
rect 165 386 199 410
rect 1605 530 1639 554
rect 1605 444 1639 496
rect 1605 386 1639 410
<< psubdiffcont >>
rect 165 123 199 157
rect 165 40 199 74
rect 1605 123 1639 157
rect 1605 40 1639 74
<< nsubdiffcont >>
rect 165 496 199 530
rect 165 410 199 444
rect 1605 496 1639 530
rect 1605 410 1639 444
<< poly >>
rect 699 544 729 570
rect 789 544 819 570
rect 890 544 920 570
rect 980 544 1010 570
rect 1181 544 1211 570
rect 1271 544 1301 570
rect 1363 544 1393 570
rect 1453 544 1483 570
rect 699 329 729 344
rect 789 329 819 344
rect 696 278 732 329
rect 786 278 822 329
rect 890 305 920 320
rect 980 305 1010 320
rect 1181 305 1211 320
rect 1271 305 1301 320
rect 1363 305 1393 320
rect 1453 305 1483 320
rect 635 262 732 278
rect 635 228 651 262
rect 685 228 732 262
rect 635 212 732 228
rect 774 262 840 278
rect 887 262 923 305
rect 977 262 1013 305
rect 774 228 790 262
rect 824 228 840 262
rect 774 212 840 228
rect 882 246 1013 262
rect 882 212 898 246
rect 932 212 1013 246
rect 702 174 732 212
rect 780 174 810 212
rect 882 196 1013 212
rect 1178 288 1214 305
rect 1268 288 1304 305
rect 1178 272 1304 288
rect 1178 238 1231 272
rect 1265 238 1304 272
rect 1178 222 1304 238
rect 882 174 912 196
rect 968 174 998 196
rect 1178 174 1208 222
rect 1274 174 1304 222
rect 1360 288 1396 305
rect 1450 288 1486 305
rect 1360 272 1486 288
rect 1360 238 1407 272
rect 1441 238 1486 272
rect 1360 222 1486 238
rect 1360 174 1390 222
rect 1456 174 1486 222
rect 702 0 732 26
rect 780 0 810 26
rect 882 0 912 26
rect 968 0 998 26
rect 1178 0 1208 26
rect 1274 0 1304 26
rect 1360 0 1390 26
rect 1456 0 1486 26
<< polycont >>
rect 651 228 685 262
rect 790 228 824 262
rect 898 212 932 246
rect 1231 238 1265 272
rect 1407 238 1441 272
<< ndiode >>
rect 257 194 395 202
rect 257 160 269 194
rect 303 160 349 194
rect 383 160 395 194
rect 257 126 395 160
rect 257 92 269 126
rect 303 92 349 126
rect 383 92 395 126
rect 257 58 395 92
rect 257 24 269 58
rect 303 24 349 58
rect 383 24 395 58
rect 257 16 395 24
rect 449 194 587 202
rect 449 160 461 194
rect 495 160 541 194
rect 575 160 587 194
rect 449 126 587 160
rect 449 92 461 126
rect 495 92 541 126
rect 575 92 587 126
rect 449 58 587 92
rect 449 24 461 58
rect 495 24 541 58
rect 575 24 587 58
rect 449 16 587 24
<< ndiodec >>
rect 269 160 303 194
rect 349 160 383 194
rect 269 92 303 126
rect 349 92 383 126
rect 269 24 303 58
rect 349 24 383 58
rect 461 160 495 194
rect 541 160 575 194
rect 461 92 495 126
rect 541 92 575 126
rect 461 24 495 58
rect 541 24 575 58
<< locali >>
rect 134 601 165 635
rect 199 601 261 635
rect 295 601 357 635
rect 391 601 453 635
rect 487 601 549 635
rect 583 601 645 635
rect 679 601 741 635
rect 775 601 837 635
rect 871 601 933 635
rect 967 601 1029 635
rect 1063 601 1125 635
rect 1159 601 1221 635
rect 1255 601 1317 635
rect 1351 601 1413 635
rect 1447 601 1509 635
rect 1543 601 1605 635
rect 1639 601 1670 635
rect 152 530 212 601
rect 152 496 165 530
rect 199 496 212 530
rect 152 444 212 496
rect 152 410 165 444
rect 199 410 212 444
rect 152 393 212 410
rect 249 300 403 565
rect 441 310 595 565
rect 636 532 702 601
rect 636 498 652 532
rect 686 498 702 532
rect 636 462 702 498
rect 636 428 652 462
rect 686 428 702 462
rect 636 392 702 428
rect 636 358 652 392
rect 686 358 702 392
rect 636 342 702 358
rect 742 532 792 548
rect 776 498 792 532
rect 742 462 792 498
rect 776 428 792 462
rect 742 392 792 428
rect 826 532 892 601
rect 826 498 842 532
rect 876 498 892 532
rect 826 460 892 498
rect 826 426 842 460
rect 876 426 892 460
rect 826 410 892 426
rect 933 532 983 548
rect 967 498 983 532
rect 933 449 983 498
rect 967 415 983 449
rect 776 376 792 392
rect 776 358 899 376
rect 742 342 899 358
rect 249 220 270 300
rect 380 220 403 300
rect 249 194 403 220
rect 440 300 595 310
rect 440 220 460 300
rect 570 220 595 300
rect 440 210 595 220
rect 635 262 701 308
rect 635 261 651 262
rect 635 227 644 261
rect 685 228 701 262
rect 678 227 701 228
rect 635 212 701 227
rect 735 262 831 308
rect 735 261 790 262
rect 735 227 788 261
rect 824 228 831 262
rect 822 227 831 228
rect 735 212 831 227
rect 865 262 899 342
rect 933 366 983 415
rect 967 332 983 366
rect 1023 532 1073 601
rect 1057 498 1073 532
rect 1023 414 1073 498
rect 1057 380 1073 414
rect 1023 364 1073 380
rect 1118 532 1168 601
rect 1118 498 1134 532
rect 1118 449 1168 498
rect 1118 415 1134 449
rect 1118 366 1168 415
rect 933 330 983 332
rect 1118 332 1134 366
rect 1208 532 1258 548
rect 1208 498 1224 532
rect 1208 462 1258 498
rect 1208 428 1224 462
rect 1208 392 1258 428
rect 1298 532 1364 601
rect 1298 498 1314 532
rect 1348 498 1364 532
rect 1298 460 1364 498
rect 1298 426 1314 460
rect 1348 426 1364 460
rect 1298 410 1364 426
rect 1406 532 1440 548
rect 1406 462 1440 498
rect 1208 358 1224 392
rect 1406 392 1440 428
rect 1480 532 1546 601
rect 1480 498 1496 532
rect 1530 498 1546 532
rect 1480 460 1546 498
rect 1480 426 1496 460
rect 1530 426 1546 460
rect 1480 410 1546 426
rect 1592 530 1652 601
rect 1592 496 1605 530
rect 1639 496 1652 530
rect 1592 444 1652 496
rect 1592 410 1605 444
rect 1639 410 1652 444
rect 1592 393 1652 410
rect 1258 358 1406 376
rect 1440 358 1549 376
rect 1208 342 1549 358
rect 933 296 1016 330
rect 1118 316 1168 332
rect 982 277 1016 296
rect 865 246 948 262
rect 865 212 898 246
rect 932 212 948 246
rect 152 157 212 173
rect 152 123 165 157
rect 199 123 212 157
rect 152 74 212 123
rect 152 40 165 74
rect 199 40 212 74
rect 152 -31 212 40
rect 249 160 269 194
rect 303 160 349 194
rect 383 160 403 194
rect 249 126 403 160
rect 249 92 269 126
rect 303 92 349 126
rect 383 92 403 126
rect 249 58 403 92
rect 249 24 269 58
rect 303 24 349 58
rect 383 24 403 58
rect 249 5 403 24
rect 441 194 595 210
rect 441 160 461 194
rect 495 160 541 194
rect 575 160 595 194
rect 865 196 948 212
rect 982 261 1034 277
rect 982 227 991 261
rect 1025 227 1034 261
rect 982 212 1034 227
rect 1215 272 1357 308
rect 1215 271 1231 272
rect 1215 237 1224 271
rect 1265 238 1357 272
rect 1258 237 1357 238
rect 1215 222 1357 237
rect 1391 272 1457 308
rect 1391 271 1407 272
rect 1391 237 1400 271
rect 1441 238 1457 272
rect 1434 237 1457 238
rect 1391 222 1457 237
rect 1503 287 1549 342
rect 1503 271 1555 287
rect 1503 237 1512 271
rect 1546 237 1555 271
rect 1503 222 1555 237
rect 865 178 899 196
rect 441 126 595 160
rect 441 92 461 126
rect 495 92 541 126
rect 575 92 595 126
rect 441 58 595 92
rect 441 24 461 58
rect 495 24 541 58
rect 575 24 595 58
rect 441 5 595 24
rect 641 162 899 178
rect 641 128 657 162
rect 691 144 899 162
rect 982 156 1016 212
rect 1503 188 1549 222
rect 691 128 707 144
rect 641 72 707 128
rect 939 122 1016 156
rect 1117 162 1349 188
rect 1117 128 1133 162
rect 1167 154 1315 162
rect 939 110 973 122
rect 641 38 657 72
rect 691 38 707 72
rect 641 22 707 38
rect 805 83 871 110
rect 805 49 821 83
rect 855 49 871 83
rect 805 -31 871 49
rect 907 83 973 110
rect 907 49 923 83
rect 957 49 973 83
rect 907 22 973 49
rect 1009 72 1071 88
rect 1009 38 1015 72
rect 1049 38 1071 72
rect 1009 -31 1071 38
rect 1117 72 1167 128
rect 1117 38 1133 72
rect 1117 22 1167 38
rect 1203 88 1269 120
rect 1203 54 1219 88
rect 1253 54 1269 88
rect 1203 -31 1269 54
rect 1315 72 1349 128
rect 1385 154 1549 188
rect 1592 157 1652 173
rect 1385 141 1451 154
rect 1385 107 1401 141
rect 1435 107 1451 141
rect 1592 123 1605 157
rect 1639 123 1652 157
rect 1385 71 1451 107
rect 1485 88 1551 120
rect 1315 37 1349 38
rect 1485 54 1501 88
rect 1535 54 1551 88
rect 1485 37 1551 54
rect 1315 3 1551 37
rect 1592 74 1652 123
rect 1592 40 1605 74
rect 1639 40 1652 74
rect 1592 -31 1652 40
rect 134 -65 165 -31
rect 199 -65 261 -31
rect 295 -65 357 -31
rect 391 -65 453 -31
rect 487 -65 549 -31
rect 583 -65 645 -31
rect 679 -65 741 -31
rect 775 -65 837 -31
rect 871 -65 933 -31
rect 967 -65 1029 -31
rect 1063 -65 1125 -31
rect 1159 -65 1221 -31
rect 1255 -65 1317 -31
rect 1351 -65 1413 -31
rect 1447 -65 1509 -31
rect 1543 -65 1605 -31
rect 1639 -65 1670 -31
<< viali >>
rect 165 601 199 635
rect 261 601 295 635
rect 357 601 391 635
rect 453 601 487 635
rect 549 601 583 635
rect 645 601 679 635
rect 741 601 775 635
rect 837 601 871 635
rect 933 601 967 635
rect 1029 601 1063 635
rect 1125 601 1159 635
rect 1221 601 1255 635
rect 1317 601 1351 635
rect 1413 601 1447 635
rect 1509 601 1543 635
rect 1605 601 1639 635
rect 270 220 380 300
rect 460 220 570 300
rect 644 228 651 261
rect 651 228 678 261
rect 644 227 678 228
rect 788 228 790 261
rect 790 228 822 261
rect 788 227 822 228
rect 991 227 1025 261
rect 1224 238 1231 271
rect 1231 238 1258 271
rect 1224 237 1258 238
rect 1400 238 1407 271
rect 1407 238 1434 271
rect 1400 237 1434 238
rect 1512 237 1546 271
rect 165 -65 199 -31
rect 261 -65 295 -31
rect 357 -65 391 -31
rect 453 -65 487 -31
rect 549 -65 583 -31
rect 645 -65 679 -31
rect 741 -65 775 -31
rect 837 -65 871 -31
rect 933 -65 967 -31
rect 1029 -65 1063 -31
rect 1125 -65 1159 -31
rect 1221 -65 1255 -31
rect 1317 -65 1351 -31
rect 1413 -65 1447 -31
rect 1509 -65 1543 -31
rect 1605 -65 1639 -31
<< metal1 >>
rect 134 650 1670 667
rect 134 635 240 650
rect 780 635 1670 650
rect 134 601 165 635
rect 199 601 240 635
rect 780 601 837 635
rect 871 601 933 635
rect 967 601 1029 635
rect 1063 601 1125 635
rect 1159 601 1221 635
rect 1255 601 1317 635
rect 1351 601 1413 635
rect 1447 601 1509 635
rect 1543 601 1605 635
rect 1639 601 1670 635
rect 134 580 240 601
rect 780 580 1670 601
rect 134 569 1670 580
rect 250 300 400 310
rect 250 220 260 300
rect 390 220 400 300
rect 250 210 400 220
rect 440 300 590 310
rect 440 220 450 300
rect 580 270 590 300
rect 1215 280 1267 287
rect 635 270 687 277
rect 580 220 635 270
rect 440 210 590 220
rect 635 212 687 218
rect 779 270 831 277
rect 779 212 831 218
rect 982 270 1034 277
rect 1215 222 1267 228
rect 1391 280 1443 287
rect 1391 222 1443 228
rect 1503 280 1555 287
rect 1503 222 1555 228
rect 982 212 1034 218
rect 134 -10 1670 1
rect 134 -31 1020 -10
rect 1560 -31 1670 -10
rect 134 -65 165 -31
rect 199 -65 261 -31
rect 295 -65 357 -31
rect 391 -65 453 -31
rect 487 -65 549 -31
rect 583 -65 645 -31
rect 679 -65 741 -31
rect 775 -65 837 -31
rect 871 -65 933 -31
rect 967 -65 1020 -31
rect 1560 -65 1605 -31
rect 1639 -65 1670 -31
rect 134 -80 1020 -65
rect 1560 -80 1670 -65
rect 134 -97 1670 -80
<< via1 >>
rect 240 635 780 650
rect 240 601 261 635
rect 261 601 295 635
rect 295 601 357 635
rect 357 601 391 635
rect 391 601 453 635
rect 453 601 487 635
rect 487 601 549 635
rect 549 601 583 635
rect 583 601 645 635
rect 645 601 679 635
rect 679 601 741 635
rect 741 601 775 635
rect 775 601 780 635
rect 240 580 780 601
rect 260 220 270 300
rect 270 220 380 300
rect 380 220 390 300
rect 450 220 460 300
rect 460 220 570 300
rect 570 220 580 300
rect 635 261 687 270
rect 635 227 644 261
rect 644 227 678 261
rect 678 227 687 261
rect 635 218 687 227
rect 779 261 831 270
rect 779 227 788 261
rect 788 227 822 261
rect 822 227 831 261
rect 779 218 831 227
rect 982 261 1034 270
rect 982 227 991 261
rect 991 227 1025 261
rect 1025 227 1034 261
rect 982 218 1034 227
rect 1215 271 1267 280
rect 1215 237 1224 271
rect 1224 237 1258 271
rect 1258 237 1267 271
rect 1215 228 1267 237
rect 1391 271 1443 280
rect 1391 237 1400 271
rect 1400 237 1434 271
rect 1434 237 1443 271
rect 1391 228 1443 237
rect 1503 271 1555 280
rect 1503 237 1512 271
rect 1512 237 1546 271
rect 1546 237 1555 271
rect 1503 228 1555 237
rect 1020 -31 1560 -10
rect 1020 -65 1029 -31
rect 1029 -65 1063 -31
rect 1063 -65 1125 -31
rect 1125 -65 1159 -31
rect 1159 -65 1221 -31
rect 1221 -65 1255 -31
rect 1255 -65 1317 -31
rect 1317 -65 1351 -31
rect 1351 -65 1413 -31
rect 1413 -65 1447 -31
rect 1447 -65 1509 -31
rect 1509 -65 1543 -31
rect 1543 -65 1560 -31
rect 1020 -80 1560 -65
<< metal2 >>
rect 230 650 790 660
rect 230 580 240 650
rect 780 580 790 650
rect 230 570 790 580
rect 650 363 1255 393
rect 250 300 400 310
rect 250 220 260 300
rect 390 220 400 300
rect 250 210 400 220
rect 440 300 590 310
rect 440 220 450 300
rect 580 220 590 300
rect 650 277 680 363
rect 790 305 1135 335
rect 790 277 820 305
rect 440 210 590 220
rect 635 270 687 277
rect 635 212 687 218
rect 779 270 831 277
rect 779 212 831 218
rect 982 270 1034 277
rect 982 212 1034 218
rect 325 182 355 210
rect 790 182 820 212
rect 325 152 820 182
rect 1105 194 1135 305
rect 1225 287 1255 363
rect 1215 280 1267 287
rect 1215 222 1267 228
rect 1391 280 1443 287
rect 1391 222 1443 228
rect 1503 280 1555 287
rect 1503 222 1555 228
rect 1405 194 1435 222
rect 1105 164 1435 194
rect 1010 -10 1570 0
rect 1010 -80 1020 -10
rect 1560 -80 1570 -10
rect 1010 -90 1570 -80
<< via2 >>
rect 240 580 780 650
rect 260 220 370 300
rect 470 220 580 300
rect 1020 -80 1560 -10
<< metal3 >>
rect 230 650 790 660
rect 230 580 240 650
rect 780 580 790 650
rect 230 570 790 580
rect 250 300 380 310
rect 250 220 260 300
rect 370 220 380 300
rect 250 210 380 220
rect 460 300 590 310
rect 460 220 470 300
rect 580 220 590 300
rect 460 210 590 220
rect 1010 -10 1570 0
rect 1010 -80 1020 -10
rect 1560 -80 1570 -10
rect 1010 -90 1570 -80
<< labels >>
rlabel locali 250 210 400 310 1 S1
rlabel locali 440 210 590 310 1 S2
rlabel metal2 982 212 1034 277 1 YAND
rlabel metal2 1503 222 1555 287 1 YNAND
rlabel metal3 230 570 790 660 1 VHI
rlabel metal3 1010 -90 1570 0 1 VLO
<< end >>
