magic
tech sky130A
magscale 1 2
timestamp 1671898674
<< nwell >>
rect -2999 -3134 2527 -696
<< pwell >>
rect -3000 -5634 -1486 -3214
rect -1363 -4310 891 -3390
rect -4360 -6214 -3440 -5748
rect -4360 -6218 -3602 -6214
rect -3556 -6218 -3440 -6214
rect -4360 -6534 -3440 -6218
rect -4360 -6640 -3528 -6534
rect -3519 -6640 -3440 -6534
rect -4360 -6882 -3440 -6640
rect -1319 -6750 847 -4330
rect 1013 -4342 3231 -3214
rect 1013 -5634 2527 -4342
<< nmos >>
rect -2804 -5424 -2744 -3424
rect -2686 -5424 -2626 -3424
rect -2568 -5424 -2508 -3424
rect -2450 -5424 -2390 -3424
rect -2332 -5424 -2272 -3424
rect -2214 -5424 -2154 -3424
rect -2096 -5424 -2036 -3424
rect -1978 -5424 -1918 -3424
rect -1860 -5424 -1800 -3424
rect -1742 -5424 -1682 -3424
rect -4150 -5978 -3650 -5948
rect -4150 -6074 -3650 -6044
rect -4150 -6170 -3650 -6140
rect -4150 -6266 -3650 -6236
rect -1123 -6540 -723 -4540
rect -665 -6540 -265 -4540
rect -207 -6540 193 -4540
rect 251 -6540 651 -4540
rect 1209 -5424 1269 -3424
rect 1327 -5424 1387 -3424
rect 1445 -5424 1505 -3424
rect 1563 -5424 1623 -3424
rect 1681 -5424 1741 -3424
rect 1799 -5424 1859 -3424
rect 1917 -5424 1977 -3424
rect 2035 -5424 2095 -3424
rect 2153 -5424 2213 -3424
rect 2271 -5424 2331 -3424
<< pmos >>
rect -2803 -2915 -2743 -915
rect -2685 -2915 -2625 -915
rect -2567 -2915 -2507 -915
rect -2449 -2915 -2389 -915
rect -2331 -2915 -2271 -915
rect -2213 -2915 -2153 -915
rect -2095 -2915 -2035 -915
rect -1977 -2915 -1917 -915
rect -1859 -2915 -1799 -915
rect -1741 -2915 -1681 -915
rect -1623 -2915 -1563 -915
rect -1505 -2915 -1445 -915
rect -1387 -2915 -1327 -915
rect -1269 -2915 -1209 -915
rect -1151 -2915 -1091 -915
rect -1033 -2915 -973 -915
rect -915 -2915 -855 -915
rect -797 -2915 -737 -915
rect -679 -2915 -619 -915
rect -561 -2915 -501 -915
rect -443 -2915 -383 -915
rect -325 -2915 -265 -915
rect -207 -2915 -147 -915
rect -89 -2915 -29 -915
rect 29 -2915 89 -915
rect 147 -2915 207 -915
rect 265 -2915 325 -915
rect 383 -2915 443 -915
rect 501 -2915 561 -915
rect 619 -2915 679 -915
rect 737 -2915 797 -915
rect 855 -2915 915 -915
rect 973 -2915 1033 -915
rect 1091 -2915 1151 -915
rect 1209 -2915 1269 -915
rect 1327 -2915 1387 -915
rect 1445 -2915 1505 -915
rect 1563 -2915 1623 -915
rect 1681 -2915 1741 -915
rect 1799 -2915 1859 -915
rect 1917 -2915 1977 -915
rect 2035 -2915 2095 -915
rect 2153 -2915 2213 -915
rect 2271 -2915 2331 -915
<< nmoslvt >>
rect -1163 -4100 -1133 -3600
rect -1067 -4100 -1037 -3600
rect -971 -4100 -941 -3600
rect -875 -4100 -845 -3600
rect -779 -4100 -749 -3600
rect -683 -4100 -653 -3600
rect -587 -4100 -557 -3600
rect -491 -4100 -461 -3600
rect -395 -4100 -365 -3600
rect -299 -4100 -269 -3600
rect -203 -4100 -173 -3600
rect -107 -4100 -77 -3600
rect -11 -4100 19 -3600
rect 85 -4100 115 -3600
rect 181 -4100 211 -3600
rect 277 -4100 307 -3600
rect 373 -4100 403 -3600
rect 469 -4100 499 -3600
rect 565 -4100 595 -3600
rect 661 -4100 691 -3600
<< ndiff >>
rect -2862 -3436 -2804 -3424
rect -2862 -5412 -2850 -3436
rect -2816 -5412 -2804 -3436
rect -2862 -5424 -2804 -5412
rect -2744 -3436 -2686 -3424
rect -2744 -5412 -2732 -3436
rect -2698 -5412 -2686 -3436
rect -2744 -5424 -2686 -5412
rect -2626 -3436 -2568 -3424
rect -2626 -5412 -2614 -3436
rect -2580 -5412 -2568 -3436
rect -2626 -5424 -2568 -5412
rect -2508 -3436 -2450 -3424
rect -2508 -5412 -2496 -3436
rect -2462 -5412 -2450 -3436
rect -2508 -5424 -2450 -5412
rect -2390 -3436 -2332 -3424
rect -2390 -5412 -2378 -3436
rect -2344 -5412 -2332 -3436
rect -2390 -5424 -2332 -5412
rect -2272 -3436 -2214 -3424
rect -2272 -5412 -2260 -3436
rect -2226 -5412 -2214 -3436
rect -2272 -5424 -2214 -5412
rect -2154 -3436 -2096 -3424
rect -2154 -5412 -2142 -3436
rect -2108 -5412 -2096 -3436
rect -2154 -5424 -2096 -5412
rect -2036 -3436 -1978 -3424
rect -2036 -5412 -2024 -3436
rect -1990 -5412 -1978 -3436
rect -2036 -5424 -1978 -5412
rect -1918 -3436 -1860 -3424
rect -1918 -5412 -1906 -3436
rect -1872 -5412 -1860 -3436
rect -1918 -5424 -1860 -5412
rect -1800 -3436 -1742 -3424
rect -1800 -5412 -1788 -3436
rect -1754 -5412 -1742 -3436
rect -1800 -5424 -1742 -5412
rect -1682 -3436 -1624 -3424
rect -1682 -5412 -1670 -3436
rect -1636 -5412 -1624 -3436
rect -1682 -5424 -1624 -5412
rect -1225 -3612 -1163 -3600
rect -1225 -4088 -1213 -3612
rect -1179 -4088 -1163 -3612
rect -1225 -4100 -1163 -4088
rect -1133 -3612 -1067 -3600
rect -1133 -4088 -1117 -3612
rect -1083 -4088 -1067 -3612
rect -1133 -4100 -1067 -4088
rect -1037 -3612 -971 -3600
rect -1037 -4088 -1021 -3612
rect -987 -4088 -971 -3612
rect -1037 -4100 -971 -4088
rect -941 -3612 -875 -3600
rect -941 -4088 -925 -3612
rect -891 -4088 -875 -3612
rect -941 -4100 -875 -4088
rect -845 -3612 -779 -3600
rect -845 -4088 -829 -3612
rect -795 -4088 -779 -3612
rect -845 -4100 -779 -4088
rect -749 -3612 -683 -3600
rect -749 -4088 -733 -3612
rect -699 -4088 -683 -3612
rect -749 -4100 -683 -4088
rect -653 -3612 -587 -3600
rect -653 -4088 -637 -3612
rect -603 -4088 -587 -3612
rect -653 -4100 -587 -4088
rect -557 -3612 -491 -3600
rect -557 -4088 -541 -3612
rect -507 -4088 -491 -3612
rect -557 -4100 -491 -4088
rect -461 -3612 -395 -3600
rect -461 -4088 -445 -3612
rect -411 -4088 -395 -3612
rect -461 -4100 -395 -4088
rect -365 -3612 -299 -3600
rect -365 -4088 -349 -3612
rect -315 -4088 -299 -3612
rect -365 -4100 -299 -4088
rect -269 -3612 -203 -3600
rect -269 -4088 -253 -3612
rect -219 -4088 -203 -3612
rect -269 -4100 -203 -4088
rect -173 -3612 -107 -3600
rect -173 -4088 -157 -3612
rect -123 -4088 -107 -3612
rect -173 -4100 -107 -4088
rect -77 -3612 -11 -3600
rect -77 -4088 -61 -3612
rect -27 -4088 -11 -3612
rect -77 -4100 -11 -4088
rect 19 -3612 85 -3600
rect 19 -4088 35 -3612
rect 69 -4088 85 -3612
rect 19 -4100 85 -4088
rect 115 -3612 181 -3600
rect 115 -4088 131 -3612
rect 165 -4088 181 -3612
rect 115 -4100 181 -4088
rect 211 -3612 277 -3600
rect 211 -4088 227 -3612
rect 261 -4088 277 -3612
rect 211 -4100 277 -4088
rect 307 -3612 373 -3600
rect 307 -4088 323 -3612
rect 357 -4088 373 -3612
rect 307 -4100 373 -4088
rect 403 -3612 469 -3600
rect 403 -4088 419 -3612
rect 453 -4088 469 -3612
rect 403 -4100 469 -4088
rect 499 -3612 565 -3600
rect 499 -4088 515 -3612
rect 549 -4088 565 -3612
rect 499 -4100 565 -4088
rect 595 -3612 661 -3600
rect 595 -4088 611 -3612
rect 645 -4088 661 -3612
rect 595 -4100 661 -4088
rect 691 -3612 753 -3600
rect 691 -4088 707 -3612
rect 741 -4088 753 -3612
rect 691 -4100 753 -4088
rect -4150 -5898 -3650 -5886
rect -4150 -5932 -4138 -5898
rect -3662 -5932 -3650 -5898
rect -4150 -5948 -3650 -5932
rect -4150 -5994 -3650 -5978
rect -4150 -6028 -4138 -5994
rect -3662 -6028 -3650 -5994
rect -4150 -6044 -3650 -6028
rect -4150 -6090 -3650 -6074
rect -4150 -6124 -4138 -6090
rect -3662 -6124 -3650 -6090
rect -4150 -6140 -3650 -6124
rect -4150 -6186 -3650 -6170
rect -4150 -6220 -4138 -6186
rect -3662 -6220 -3650 -6186
rect -4150 -6236 -3650 -6220
rect -4150 -6282 -3650 -6266
rect -4150 -6316 -4138 -6282
rect -3662 -6316 -3650 -6282
rect -4150 -6328 -3650 -6316
rect -1181 -4552 -1123 -4540
rect -1181 -6528 -1169 -4552
rect -1135 -6528 -1123 -4552
rect -1181 -6540 -1123 -6528
rect -723 -4552 -665 -4540
rect -723 -6528 -711 -4552
rect -677 -6528 -665 -4552
rect -723 -6540 -665 -6528
rect -265 -4552 -207 -4540
rect -265 -6528 -253 -4552
rect -219 -6528 -207 -4552
rect -265 -6540 -207 -6528
rect 193 -4552 251 -4540
rect 193 -6528 205 -4552
rect 239 -6528 251 -4552
rect 193 -6540 251 -6528
rect 651 -4552 709 -4540
rect 651 -6528 663 -4552
rect 697 -6528 709 -4552
rect 651 -6540 709 -6528
rect 1151 -3436 1209 -3424
rect 1151 -5412 1163 -3436
rect 1197 -5412 1209 -3436
rect 1151 -5424 1209 -5412
rect 1269 -3436 1327 -3424
rect 1269 -5412 1281 -3436
rect 1315 -5412 1327 -3436
rect 1269 -5424 1327 -5412
rect 1387 -3436 1445 -3424
rect 1387 -5412 1399 -3436
rect 1433 -5412 1445 -3436
rect 1387 -5424 1445 -5412
rect 1505 -3436 1563 -3424
rect 1505 -5412 1517 -3436
rect 1551 -5412 1563 -3436
rect 1505 -5424 1563 -5412
rect 1623 -3436 1681 -3424
rect 1623 -5412 1635 -3436
rect 1669 -5412 1681 -3436
rect 1623 -5424 1681 -5412
rect 1741 -3436 1799 -3424
rect 1741 -5412 1753 -3436
rect 1787 -5412 1799 -3436
rect 1741 -5424 1799 -5412
rect 1859 -3436 1917 -3424
rect 1859 -5412 1871 -3436
rect 1905 -5412 1917 -3436
rect 1859 -5424 1917 -5412
rect 1977 -3436 2035 -3424
rect 1977 -5412 1989 -3436
rect 2023 -5412 2035 -3436
rect 1977 -5424 2035 -5412
rect 2095 -3436 2153 -3424
rect 2095 -5412 2107 -3436
rect 2141 -5412 2153 -3436
rect 2095 -5424 2153 -5412
rect 2213 -3436 2271 -3424
rect 2213 -5412 2225 -3436
rect 2259 -5412 2271 -3436
rect 2213 -5424 2271 -5412
rect 2331 -3436 2389 -3424
rect 2331 -5412 2343 -3436
rect 2377 -5412 2389 -3436
rect 2331 -5424 2389 -5412
<< pdiff >>
rect -2861 -927 -2803 -915
rect -2861 -2903 -2849 -927
rect -2815 -2903 -2803 -927
rect -2861 -2915 -2803 -2903
rect -2743 -927 -2685 -915
rect -2743 -2903 -2731 -927
rect -2697 -2903 -2685 -927
rect -2743 -2915 -2685 -2903
rect -2625 -927 -2567 -915
rect -2625 -2903 -2613 -927
rect -2579 -2903 -2567 -927
rect -2625 -2915 -2567 -2903
rect -2507 -927 -2449 -915
rect -2507 -2903 -2495 -927
rect -2461 -2903 -2449 -927
rect -2507 -2915 -2449 -2903
rect -2389 -927 -2331 -915
rect -2389 -2903 -2377 -927
rect -2343 -2903 -2331 -927
rect -2389 -2915 -2331 -2903
rect -2271 -927 -2213 -915
rect -2271 -2903 -2259 -927
rect -2225 -2903 -2213 -927
rect -2271 -2915 -2213 -2903
rect -2153 -927 -2095 -915
rect -2153 -2903 -2141 -927
rect -2107 -2903 -2095 -927
rect -2153 -2915 -2095 -2903
rect -2035 -927 -1977 -915
rect -2035 -2903 -2023 -927
rect -1989 -2903 -1977 -927
rect -2035 -2915 -1977 -2903
rect -1917 -927 -1859 -915
rect -1917 -2903 -1905 -927
rect -1871 -2903 -1859 -927
rect -1917 -2915 -1859 -2903
rect -1799 -927 -1741 -915
rect -1799 -2903 -1787 -927
rect -1753 -2903 -1741 -927
rect -1799 -2915 -1741 -2903
rect -1681 -927 -1623 -915
rect -1681 -2903 -1669 -927
rect -1635 -2903 -1623 -927
rect -1681 -2915 -1623 -2903
rect -1563 -927 -1505 -915
rect -1563 -2903 -1551 -927
rect -1517 -2903 -1505 -927
rect -1563 -2915 -1505 -2903
rect -1445 -927 -1387 -915
rect -1445 -2903 -1433 -927
rect -1399 -2903 -1387 -927
rect -1445 -2915 -1387 -2903
rect -1327 -927 -1269 -915
rect -1327 -2903 -1315 -927
rect -1281 -2903 -1269 -927
rect -1327 -2915 -1269 -2903
rect -1209 -927 -1151 -915
rect -1209 -2903 -1197 -927
rect -1163 -2903 -1151 -927
rect -1209 -2915 -1151 -2903
rect -1091 -927 -1033 -915
rect -1091 -2903 -1079 -927
rect -1045 -2903 -1033 -927
rect -1091 -2915 -1033 -2903
rect -973 -927 -915 -915
rect -973 -2903 -961 -927
rect -927 -2903 -915 -927
rect -973 -2915 -915 -2903
rect -855 -927 -797 -915
rect -855 -2903 -843 -927
rect -809 -2903 -797 -927
rect -855 -2915 -797 -2903
rect -737 -927 -679 -915
rect -737 -2903 -725 -927
rect -691 -2903 -679 -927
rect -737 -2915 -679 -2903
rect -619 -927 -561 -915
rect -619 -2903 -607 -927
rect -573 -2903 -561 -927
rect -619 -2915 -561 -2903
rect -501 -927 -443 -915
rect -501 -2903 -489 -927
rect -455 -2903 -443 -927
rect -501 -2915 -443 -2903
rect -383 -927 -325 -915
rect -383 -2903 -371 -927
rect -337 -2903 -325 -927
rect -383 -2915 -325 -2903
rect -265 -927 -207 -915
rect -265 -2903 -253 -927
rect -219 -2903 -207 -927
rect -265 -2915 -207 -2903
rect -147 -927 -89 -915
rect -147 -2903 -135 -927
rect -101 -2903 -89 -927
rect -147 -2915 -89 -2903
rect -29 -927 29 -915
rect -29 -2903 -17 -927
rect 17 -2903 29 -927
rect -29 -2915 29 -2903
rect 89 -927 147 -915
rect 89 -2903 101 -927
rect 135 -2903 147 -927
rect 89 -2915 147 -2903
rect 207 -927 265 -915
rect 207 -2903 219 -927
rect 253 -2903 265 -927
rect 207 -2915 265 -2903
rect 325 -927 383 -915
rect 325 -2903 337 -927
rect 371 -2903 383 -927
rect 325 -2915 383 -2903
rect 443 -927 501 -915
rect 443 -2903 455 -927
rect 489 -2903 501 -927
rect 443 -2915 501 -2903
rect 561 -927 619 -915
rect 561 -2903 573 -927
rect 607 -2903 619 -927
rect 561 -2915 619 -2903
rect 679 -927 737 -915
rect 679 -2903 691 -927
rect 725 -2903 737 -927
rect 679 -2915 737 -2903
rect 797 -927 855 -915
rect 797 -2903 809 -927
rect 843 -2903 855 -927
rect 797 -2915 855 -2903
rect 915 -927 973 -915
rect 915 -2903 927 -927
rect 961 -2903 973 -927
rect 915 -2915 973 -2903
rect 1033 -927 1091 -915
rect 1033 -2903 1045 -927
rect 1079 -2903 1091 -927
rect 1033 -2915 1091 -2903
rect 1151 -927 1209 -915
rect 1151 -2903 1163 -927
rect 1197 -2903 1209 -927
rect 1151 -2915 1209 -2903
rect 1269 -927 1327 -915
rect 1269 -2903 1281 -927
rect 1315 -2903 1327 -927
rect 1269 -2915 1327 -2903
rect 1387 -927 1445 -915
rect 1387 -2903 1399 -927
rect 1433 -2903 1445 -927
rect 1387 -2915 1445 -2903
rect 1505 -927 1563 -915
rect 1505 -2903 1517 -927
rect 1551 -2903 1563 -927
rect 1505 -2915 1563 -2903
rect 1623 -927 1681 -915
rect 1623 -2903 1635 -927
rect 1669 -2903 1681 -927
rect 1623 -2915 1681 -2903
rect 1741 -927 1799 -915
rect 1741 -2903 1753 -927
rect 1787 -2903 1799 -927
rect 1741 -2915 1799 -2903
rect 1859 -927 1917 -915
rect 1859 -2903 1871 -927
rect 1905 -2903 1917 -927
rect 1859 -2915 1917 -2903
rect 1977 -927 2035 -915
rect 1977 -2903 1989 -927
rect 2023 -2903 2035 -927
rect 1977 -2915 2035 -2903
rect 2095 -927 2153 -915
rect 2095 -2903 2107 -927
rect 2141 -2903 2153 -927
rect 2095 -2915 2153 -2903
rect 2213 -927 2271 -915
rect 2213 -2903 2225 -927
rect 2259 -2903 2271 -927
rect 2213 -2915 2271 -2903
rect 2331 -927 2389 -915
rect 2331 -2903 2343 -927
rect 2377 -2903 2389 -927
rect 2331 -2915 2389 -2903
<< ndiffc >>
rect -2850 -5412 -2816 -3436
rect -2732 -5412 -2698 -3436
rect -2614 -5412 -2580 -3436
rect -2496 -5412 -2462 -3436
rect -2378 -5412 -2344 -3436
rect -2260 -5412 -2226 -3436
rect -2142 -5412 -2108 -3436
rect -2024 -5412 -1990 -3436
rect -1906 -5412 -1872 -3436
rect -1788 -5412 -1754 -3436
rect -1670 -5412 -1636 -3436
rect -1213 -4088 -1179 -3612
rect -1117 -4088 -1083 -3612
rect -1021 -4088 -987 -3612
rect -925 -4088 -891 -3612
rect -829 -4088 -795 -3612
rect -733 -4088 -699 -3612
rect -637 -4088 -603 -3612
rect -541 -4088 -507 -3612
rect -445 -4088 -411 -3612
rect -349 -4088 -315 -3612
rect -253 -4088 -219 -3612
rect -157 -4088 -123 -3612
rect -61 -4088 -27 -3612
rect 35 -4088 69 -3612
rect 131 -4088 165 -3612
rect 227 -4088 261 -3612
rect 323 -4088 357 -3612
rect 419 -4088 453 -3612
rect 515 -4088 549 -3612
rect 611 -4088 645 -3612
rect 707 -4088 741 -3612
rect -4138 -5932 -3662 -5898
rect -4138 -6028 -3662 -5994
rect -4138 -6124 -3662 -6090
rect -4138 -6220 -3662 -6186
rect -4138 -6316 -3662 -6282
rect -1169 -6528 -1135 -4552
rect -711 -6528 -677 -4552
rect -253 -6528 -219 -4552
rect 205 -6528 239 -4552
rect 663 -6528 697 -4552
rect 1163 -5412 1197 -3436
rect 1281 -5412 1315 -3436
rect 1399 -5412 1433 -3436
rect 1517 -5412 1551 -3436
rect 1635 -5412 1669 -3436
rect 1753 -5412 1787 -3436
rect 1871 -5412 1905 -3436
rect 1989 -5412 2023 -3436
rect 2107 -5412 2141 -3436
rect 2225 -5412 2259 -3436
rect 2343 -5412 2377 -3436
<< pdiffc >>
rect -2849 -2903 -2815 -927
rect -2731 -2903 -2697 -927
rect -2613 -2903 -2579 -927
rect -2495 -2903 -2461 -927
rect -2377 -2903 -2343 -927
rect -2259 -2903 -2225 -927
rect -2141 -2903 -2107 -927
rect -2023 -2903 -1989 -927
rect -1905 -2903 -1871 -927
rect -1787 -2903 -1753 -927
rect -1669 -2903 -1635 -927
rect -1551 -2903 -1517 -927
rect -1433 -2903 -1399 -927
rect -1315 -2903 -1281 -927
rect -1197 -2903 -1163 -927
rect -1079 -2903 -1045 -927
rect -961 -2903 -927 -927
rect -843 -2903 -809 -927
rect -725 -2903 -691 -927
rect -607 -2903 -573 -927
rect -489 -2903 -455 -927
rect -371 -2903 -337 -927
rect -253 -2903 -219 -927
rect -135 -2903 -101 -927
rect -17 -2903 17 -927
rect 101 -2903 135 -927
rect 219 -2903 253 -927
rect 337 -2903 371 -927
rect 455 -2903 489 -927
rect 573 -2903 607 -927
rect 691 -2903 725 -927
rect 809 -2903 843 -927
rect 927 -2903 961 -927
rect 1045 -2903 1079 -927
rect 1163 -2903 1197 -927
rect 1281 -2903 1315 -927
rect 1399 -2903 1433 -927
rect 1517 -2903 1551 -927
rect 1635 -2903 1669 -927
rect 1753 -2903 1787 -927
rect 1871 -2903 1905 -927
rect 1989 -2903 2023 -927
rect 2107 -2903 2141 -927
rect 2225 -2903 2259 -927
rect 2343 -2903 2377 -927
<< psubdiff >>
rect -2964 -3284 -2868 -3250
rect -1618 -3284 -1522 -3250
rect -2964 -3346 -2930 -3284
rect -1556 -3346 -1522 -3284
rect -2964 -5564 -2930 -5502
rect 1049 -3284 1145 -3250
rect 2395 -3284 2491 -3250
rect 1049 -3346 1083 -3284
rect -1327 -3460 -1231 -3426
rect 759 -3460 855 -3426
rect -1327 -3522 -1293 -3460
rect 821 -3522 855 -3460
rect -1327 -4240 -1293 -4178
rect 821 -4240 855 -4178
rect -1327 -4274 -1231 -4240
rect 759 -4274 855 -4240
rect -1556 -5564 -1522 -5502
rect -2964 -5598 -2868 -5564
rect -1618 -5598 -1522 -5564
rect -1283 -4400 -1187 -4366
rect 715 -4400 811 -4366
rect -1283 -4462 -1249 -4400
rect -4324 -5818 -4228 -5784
rect -3572 -5818 -3476 -5784
rect -4324 -5880 -4290 -5818
rect -3510 -5880 -3476 -5818
rect -4324 -6812 -4290 -6730
rect 777 -4462 811 -4400
rect -1283 -6680 -1249 -6618
rect 2457 -3346 2491 -3284
rect 1049 -5564 1083 -5502
rect 2563 -3284 2659 -3250
rect 3099 -3284 3195 -3250
rect 2563 -3346 2597 -3284
rect 3161 -3346 3195 -3284
rect 2563 -4272 2597 -4210
rect 3161 -4272 3195 -4210
rect 2563 -4306 2659 -4272
rect 3099 -4306 3195 -4272
rect 2457 -5564 2491 -5502
rect 1049 -5598 1145 -5564
rect 2395 -5598 2491 -5564
rect 777 -6680 811 -6618
rect -1283 -6714 -1187 -6680
rect 715 -6714 811 -6680
rect -3510 -6812 -3476 -6730
rect -4324 -6846 -4228 -6812
rect -3572 -6846 -3476 -6812
<< nsubdiff >>
rect -2963 -766 -2867 -732
rect 2395 -766 2491 -732
rect -2963 -828 -2929 -766
rect 2457 -828 2491 -766
rect -2963 -3064 -2929 -3002
rect 2457 -3064 2491 -3002
rect -2963 -3098 -2867 -3064
rect 2395 -3098 2491 -3064
<< psubdiffcont >>
rect -2868 -3284 -1618 -3250
rect -2964 -5502 -2930 -3346
rect -1556 -5502 -1522 -3346
rect 1145 -3284 2395 -3250
rect -1231 -3460 759 -3426
rect -1327 -4178 -1293 -3522
rect 821 -4178 855 -3522
rect -1231 -4274 759 -4240
rect -2868 -5598 -1618 -5564
rect -1187 -4400 715 -4366
rect -4228 -5818 -3572 -5784
rect -4324 -6730 -4290 -5880
rect -3510 -6730 -3476 -5880
rect -1283 -6618 -1249 -4462
rect 777 -6618 811 -4462
rect 1049 -5502 1083 -3346
rect 2457 -5502 2491 -3346
rect 2659 -3284 3099 -3250
rect 2563 -4210 2597 -3346
rect 3161 -4210 3195 -3346
rect 2659 -4306 3099 -4272
rect 1145 -5598 2395 -5564
rect -1187 -6714 715 -6680
rect -4228 -6846 -3572 -6812
<< nsubdiffcont >>
rect -2867 -766 2395 -732
rect -2963 -3002 -2929 -828
rect 2457 -3002 2491 -828
rect -2867 -3098 2395 -3064
<< poly >>
rect -2806 -834 -2740 -818
rect -2806 -868 -2790 -834
rect -2756 -868 -2740 -834
rect -2806 -884 -2740 -868
rect -2688 -834 -2622 -818
rect -2688 -868 -2672 -834
rect -2638 -868 -2622 -834
rect -2688 -884 -2622 -868
rect -2570 -834 -2504 -818
rect -2570 -868 -2554 -834
rect -2520 -868 -2504 -834
rect -2570 -884 -2504 -868
rect -2452 -834 -2386 -818
rect -2452 -868 -2436 -834
rect -2402 -868 -2386 -834
rect -2452 -884 -2386 -868
rect -2334 -834 -2268 -818
rect -2334 -868 -2318 -834
rect -2284 -868 -2268 -834
rect -2334 -884 -2268 -868
rect -2216 -834 -2150 -818
rect -2216 -868 -2200 -834
rect -2166 -868 -2150 -834
rect -2216 -884 -2150 -868
rect -2098 -834 -2032 -818
rect -2098 -868 -2082 -834
rect -2048 -868 -2032 -834
rect -2098 -884 -2032 -868
rect -1980 -834 -1914 -818
rect -1980 -868 -1964 -834
rect -1930 -868 -1914 -834
rect -1980 -884 -1914 -868
rect -1862 -834 -1796 -818
rect -1862 -868 -1846 -834
rect -1812 -868 -1796 -834
rect -1862 -884 -1796 -868
rect -1744 -834 -1678 -818
rect -1744 -868 -1728 -834
rect -1694 -868 -1678 -834
rect -1744 -884 -1678 -868
rect -1626 -834 -1560 -818
rect -1626 -868 -1610 -834
rect -1576 -868 -1560 -834
rect -1626 -884 -1560 -868
rect -1508 -834 -1442 -818
rect -1508 -868 -1492 -834
rect -1458 -868 -1442 -834
rect -1508 -884 -1442 -868
rect -1390 -834 -1324 -818
rect -1390 -868 -1374 -834
rect -1340 -868 -1324 -834
rect -1390 -884 -1324 -868
rect -1272 -834 -1206 -818
rect -1272 -868 -1256 -834
rect -1222 -868 -1206 -834
rect -1272 -884 -1206 -868
rect -1154 -834 -1088 -818
rect -1154 -868 -1138 -834
rect -1104 -868 -1088 -834
rect -1154 -884 -1088 -868
rect -1036 -834 -970 -818
rect -1036 -868 -1020 -834
rect -986 -868 -970 -834
rect -1036 -884 -970 -868
rect -918 -834 -852 -818
rect -918 -868 -902 -834
rect -868 -868 -852 -834
rect -918 -884 -852 -868
rect -800 -834 -734 -818
rect -800 -868 -784 -834
rect -750 -868 -734 -834
rect -800 -884 -734 -868
rect -682 -834 -616 -818
rect -682 -868 -666 -834
rect -632 -868 -616 -834
rect -682 -884 -616 -868
rect -564 -834 -498 -818
rect -564 -868 -548 -834
rect -514 -868 -498 -834
rect -564 -884 -498 -868
rect -446 -884 -380 -818
rect -328 -884 -262 -818
rect -210 -884 -144 -818
rect -92 -884 -26 -818
rect 26 -834 92 -818
rect 26 -868 42 -834
rect 76 -868 92 -834
rect 26 -884 92 -868
rect 144 -834 210 -818
rect 144 -868 160 -834
rect 194 -868 210 -834
rect 144 -884 210 -868
rect 262 -834 328 -818
rect 262 -868 278 -834
rect 312 -868 328 -834
rect 262 -884 328 -868
rect 380 -834 446 -818
rect 380 -868 396 -834
rect 430 -868 446 -834
rect 380 -884 446 -868
rect 498 -834 564 -818
rect 498 -868 514 -834
rect 548 -868 564 -834
rect 498 -884 564 -868
rect 616 -834 682 -818
rect 616 -868 632 -834
rect 666 -868 682 -834
rect 616 -884 682 -868
rect 734 -834 800 -818
rect 734 -868 750 -834
rect 784 -868 800 -834
rect 734 -884 800 -868
rect 852 -834 918 -818
rect 852 -868 868 -834
rect 902 -868 918 -834
rect 852 -884 918 -868
rect 970 -834 1036 -818
rect 970 -868 986 -834
rect 1020 -868 1036 -834
rect 970 -884 1036 -868
rect 1088 -834 1154 -818
rect 1088 -868 1104 -834
rect 1138 -868 1154 -834
rect 1088 -884 1154 -868
rect 1206 -834 1272 -818
rect 1206 -868 1222 -834
rect 1256 -868 1272 -834
rect 1206 -884 1272 -868
rect 1324 -834 1390 -818
rect 1324 -868 1340 -834
rect 1374 -868 1390 -834
rect 1324 -884 1390 -868
rect 1442 -834 1508 -818
rect 1442 -868 1458 -834
rect 1492 -868 1508 -834
rect 1442 -884 1508 -868
rect 1560 -834 1626 -818
rect 1560 -868 1576 -834
rect 1610 -868 1626 -834
rect 1560 -884 1626 -868
rect 1678 -834 1744 -818
rect 1678 -868 1694 -834
rect 1728 -868 1744 -834
rect 1678 -884 1744 -868
rect 1796 -834 1862 -818
rect 1796 -868 1812 -834
rect 1846 -868 1862 -834
rect 1796 -884 1862 -868
rect 1914 -834 1980 -818
rect 1914 -868 1930 -834
rect 1964 -868 1980 -834
rect 1914 -884 1980 -868
rect 2032 -834 2098 -818
rect 2032 -868 2048 -834
rect 2082 -868 2098 -834
rect 2032 -884 2098 -868
rect 2150 -834 2216 -818
rect 2150 -868 2166 -834
rect 2200 -868 2216 -834
rect 2150 -884 2216 -868
rect 2268 -834 2334 -818
rect 2268 -868 2284 -834
rect 2318 -868 2334 -834
rect 2268 -884 2334 -868
rect -2803 -915 -2743 -884
rect -2685 -915 -2625 -884
rect -2567 -915 -2507 -884
rect -2449 -915 -2389 -884
rect -2331 -915 -2271 -884
rect -2213 -915 -2153 -884
rect -2095 -915 -2035 -884
rect -1977 -915 -1917 -884
rect -1859 -915 -1799 -884
rect -1741 -915 -1681 -884
rect -1623 -915 -1563 -884
rect -1505 -915 -1445 -884
rect -1387 -915 -1327 -884
rect -1269 -915 -1209 -884
rect -1151 -915 -1091 -884
rect -1033 -915 -973 -884
rect -915 -915 -855 -884
rect -797 -915 -737 -884
rect -679 -915 -619 -884
rect -561 -915 -501 -884
rect -443 -915 -383 -884
rect -325 -915 -265 -884
rect -207 -915 -147 -884
rect -89 -915 -29 -884
rect 29 -915 89 -884
rect 147 -915 207 -884
rect 265 -915 325 -884
rect 383 -915 443 -884
rect 501 -915 561 -884
rect 619 -915 679 -884
rect 737 -915 797 -884
rect 855 -915 915 -884
rect 973 -915 1033 -884
rect 1091 -915 1151 -884
rect 1209 -915 1269 -884
rect 1327 -915 1387 -884
rect 1445 -915 1505 -884
rect 1563 -915 1623 -884
rect 1681 -915 1741 -884
rect 1799 -915 1859 -884
rect 1917 -915 1977 -884
rect 2035 -915 2095 -884
rect 2153 -915 2213 -884
rect 2271 -915 2331 -884
rect -2803 -2946 -2743 -2915
rect -2685 -2946 -2625 -2915
rect -2567 -2946 -2507 -2915
rect -2449 -2946 -2389 -2915
rect -2331 -2946 -2271 -2915
rect -2213 -2946 -2153 -2915
rect -2095 -2946 -2035 -2915
rect -1977 -2946 -1917 -2915
rect -1859 -2946 -1799 -2915
rect -1741 -2946 -1681 -2915
rect -1623 -2946 -1563 -2915
rect -1505 -2946 -1445 -2915
rect -1387 -2946 -1327 -2915
rect -1269 -2946 -1209 -2915
rect -1151 -2946 -1091 -2915
rect -1033 -2946 -973 -2915
rect -915 -2946 -855 -2915
rect -797 -2946 -737 -2915
rect -679 -2946 -619 -2915
rect -561 -2946 -501 -2915
rect -443 -2946 -383 -2915
rect -325 -2946 -265 -2915
rect -207 -2946 -147 -2915
rect -89 -2946 -29 -2915
rect 29 -2946 89 -2915
rect 147 -2946 207 -2915
rect 265 -2946 325 -2915
rect 383 -2946 443 -2915
rect 501 -2946 561 -2915
rect 619 -2946 679 -2915
rect 737 -2946 797 -2915
rect 855 -2946 915 -2915
rect 973 -2946 1033 -2915
rect 1091 -2946 1151 -2915
rect 1209 -2946 1269 -2915
rect 1327 -2946 1387 -2915
rect 1445 -2946 1505 -2915
rect 1563 -2946 1623 -2915
rect 1681 -2946 1741 -2915
rect 1799 -2946 1859 -2915
rect 1917 -2946 1977 -2915
rect 2035 -2946 2095 -2915
rect 2153 -2946 2213 -2915
rect 2271 -2946 2331 -2915
rect -2806 -2962 -2740 -2946
rect -2806 -2996 -2790 -2962
rect -2756 -2996 -2740 -2962
rect -2806 -3012 -2740 -2996
rect -2688 -2962 -2622 -2946
rect -2688 -2996 -2672 -2962
rect -2638 -2996 -2622 -2962
rect -2688 -3012 -2622 -2996
rect -2570 -2962 -2504 -2946
rect -2570 -2996 -2554 -2962
rect -2520 -2996 -2504 -2962
rect -2570 -3012 -2504 -2996
rect -2452 -2962 -2386 -2946
rect -2452 -2996 -2436 -2962
rect -2402 -2996 -2386 -2962
rect -2452 -3012 -2386 -2996
rect -2334 -2962 -2268 -2946
rect -2334 -2996 -2318 -2962
rect -2284 -2996 -2268 -2962
rect -2334 -3012 -2268 -2996
rect -2216 -2962 -2150 -2946
rect -2216 -2996 -2200 -2962
rect -2166 -2996 -2150 -2962
rect -2216 -3012 -2150 -2996
rect -2098 -2962 -2032 -2946
rect -2098 -2996 -2082 -2962
rect -2048 -2996 -2032 -2962
rect -2098 -3012 -2032 -2996
rect -1980 -2962 -1914 -2946
rect -1980 -2996 -1964 -2962
rect -1930 -2996 -1914 -2962
rect -1980 -3012 -1914 -2996
rect -1862 -2962 -1796 -2946
rect -1862 -2996 -1846 -2962
rect -1812 -2996 -1796 -2962
rect -1862 -3012 -1796 -2996
rect -1744 -2962 -1678 -2946
rect -1744 -2996 -1728 -2962
rect -1694 -2996 -1678 -2962
rect -1744 -3012 -1678 -2996
rect -1626 -2962 -1560 -2946
rect -1626 -2996 -1610 -2962
rect -1576 -2996 -1560 -2962
rect -1626 -3012 -1560 -2996
rect -1508 -2962 -1442 -2946
rect -1508 -2996 -1492 -2962
rect -1458 -2996 -1442 -2962
rect -1508 -3012 -1442 -2996
rect -1390 -2962 -1324 -2946
rect -1390 -2996 -1374 -2962
rect -1340 -2996 -1324 -2962
rect -1390 -3012 -1324 -2996
rect -1272 -2962 -1206 -2946
rect -1272 -2996 -1256 -2962
rect -1222 -2996 -1206 -2962
rect -1272 -3012 -1206 -2996
rect -1154 -2962 -1088 -2946
rect -1154 -2996 -1138 -2962
rect -1104 -2996 -1088 -2962
rect -1154 -3012 -1088 -2996
rect -1036 -2962 -970 -2946
rect -1036 -2996 -1020 -2962
rect -986 -2996 -970 -2962
rect -1036 -3012 -970 -2996
rect -918 -2962 -852 -2946
rect -918 -2996 -902 -2962
rect -868 -2996 -852 -2962
rect -918 -3012 -852 -2996
rect -800 -2962 -734 -2946
rect -800 -2996 -784 -2962
rect -750 -2996 -734 -2962
rect -800 -3012 -734 -2996
rect -682 -2962 -616 -2946
rect -682 -2996 -666 -2962
rect -632 -2996 -616 -2962
rect -682 -3012 -616 -2996
rect -564 -2962 -498 -2946
rect -564 -2996 -548 -2962
rect -514 -2996 -498 -2962
rect -564 -3012 -498 -2996
rect -446 -2962 -380 -2946
rect -446 -2996 -430 -2962
rect -396 -2996 -380 -2962
rect -446 -3012 -380 -2996
rect -328 -2962 -262 -2946
rect -328 -2996 -312 -2962
rect -278 -2996 -262 -2962
rect -328 -3012 -262 -2996
rect -210 -2962 -144 -2946
rect -210 -2996 -194 -2962
rect -160 -2996 -144 -2962
rect -210 -3012 -144 -2996
rect -92 -2962 -26 -2946
rect -92 -2996 -76 -2962
rect -42 -2996 -26 -2962
rect -92 -3012 -26 -2996
rect 26 -2962 92 -2946
rect 26 -2996 42 -2962
rect 76 -2996 92 -2962
rect 26 -3012 92 -2996
rect 144 -2962 210 -2946
rect 144 -2996 160 -2962
rect 194 -2996 210 -2962
rect 144 -3012 210 -2996
rect 262 -2962 328 -2946
rect 262 -2996 278 -2962
rect 312 -2996 328 -2962
rect 262 -3012 328 -2996
rect 380 -2962 446 -2946
rect 380 -2996 396 -2962
rect 430 -2996 446 -2962
rect 380 -3012 446 -2996
rect 498 -2962 564 -2946
rect 498 -2996 514 -2962
rect 548 -2996 564 -2962
rect 498 -3012 564 -2996
rect 616 -2962 682 -2946
rect 616 -2996 632 -2962
rect 666 -2996 682 -2962
rect 616 -3012 682 -2996
rect 734 -2962 800 -2946
rect 734 -2996 750 -2962
rect 784 -2996 800 -2962
rect 734 -3012 800 -2996
rect 852 -2962 918 -2946
rect 852 -2996 868 -2962
rect 902 -2996 918 -2962
rect 852 -3012 918 -2996
rect 970 -2962 1036 -2946
rect 970 -2996 986 -2962
rect 1020 -2996 1036 -2962
rect 970 -3012 1036 -2996
rect 1088 -2962 1154 -2946
rect 1088 -2996 1104 -2962
rect 1138 -2996 1154 -2962
rect 1088 -3012 1154 -2996
rect 1206 -2962 1272 -2946
rect 1206 -2996 1222 -2962
rect 1256 -2996 1272 -2962
rect 1206 -3012 1272 -2996
rect 1324 -2962 1390 -2946
rect 1324 -2996 1340 -2962
rect 1374 -2996 1390 -2962
rect 1324 -3012 1390 -2996
rect 1442 -2962 1508 -2946
rect 1442 -2996 1458 -2962
rect 1492 -2996 1508 -2962
rect 1442 -3012 1508 -2996
rect 1560 -2962 1626 -2946
rect 1560 -2996 1576 -2962
rect 1610 -2996 1626 -2962
rect 1560 -3012 1626 -2996
rect 1678 -2962 1744 -2946
rect 1678 -2996 1694 -2962
rect 1728 -2996 1744 -2962
rect 1678 -3012 1744 -2996
rect 1796 -2962 1862 -2946
rect 1796 -2996 1812 -2962
rect 1846 -2996 1862 -2962
rect 1796 -3012 1862 -2996
rect 1914 -2962 1980 -2946
rect 1914 -2996 1930 -2962
rect 1964 -2996 1980 -2962
rect 1914 -3012 1980 -2996
rect 2032 -2962 2098 -2946
rect 2032 -2996 2048 -2962
rect 2082 -2996 2098 -2962
rect 2032 -3012 2098 -2996
rect 2150 -2962 2216 -2946
rect 2150 -2996 2166 -2962
rect 2200 -2996 2216 -2962
rect 2150 -3012 2216 -2996
rect 2268 -2962 2334 -2946
rect 2268 -2996 2284 -2962
rect 2318 -2996 2334 -2962
rect 2268 -3012 2334 -2996
rect -2807 -3352 -2741 -3336
rect -2807 -3386 -2791 -3352
rect -2757 -3386 -2741 -3352
rect -2807 -3402 -2741 -3386
rect -2689 -3352 -2623 -3336
rect -2689 -3386 -2673 -3352
rect -2639 -3386 -2623 -3352
rect -2689 -3402 -2623 -3386
rect -2571 -3352 -2505 -3336
rect -2571 -3386 -2555 -3352
rect -2521 -3386 -2505 -3352
rect -2571 -3402 -2505 -3386
rect -2453 -3352 -2387 -3336
rect -2453 -3386 -2437 -3352
rect -2403 -3386 -2387 -3352
rect -2453 -3402 -2387 -3386
rect -2335 -3352 -2269 -3336
rect -2335 -3386 -2319 -3352
rect -2285 -3386 -2269 -3352
rect -2335 -3402 -2269 -3386
rect -2217 -3352 -2151 -3336
rect -2217 -3386 -2201 -3352
rect -2167 -3386 -2151 -3352
rect -2217 -3402 -2151 -3386
rect -2099 -3352 -2033 -3336
rect -2099 -3386 -2083 -3352
rect -2049 -3386 -2033 -3352
rect -2099 -3402 -2033 -3386
rect -1981 -3352 -1915 -3336
rect -1981 -3386 -1965 -3352
rect -1931 -3386 -1915 -3352
rect -1981 -3402 -1915 -3386
rect -1863 -3352 -1797 -3336
rect -1863 -3386 -1847 -3352
rect -1813 -3386 -1797 -3352
rect -1863 -3402 -1797 -3386
rect -1745 -3352 -1679 -3336
rect -1745 -3386 -1729 -3352
rect -1695 -3386 -1679 -3352
rect -1745 -3402 -1679 -3386
rect -2804 -3424 -2744 -3402
rect -2686 -3424 -2626 -3402
rect -2568 -3424 -2508 -3402
rect -2450 -3424 -2390 -3402
rect -2332 -3424 -2272 -3402
rect -2214 -3424 -2154 -3402
rect -2096 -3424 -2036 -3402
rect -1978 -3424 -1918 -3402
rect -1860 -3424 -1800 -3402
rect -1742 -3424 -1682 -3402
rect -2804 -5446 -2744 -5424
rect -2686 -5446 -2626 -5424
rect -2568 -5446 -2508 -5424
rect -2450 -5446 -2390 -5424
rect -2332 -5446 -2272 -5424
rect -2214 -5446 -2154 -5424
rect -2096 -5446 -2036 -5424
rect -1978 -5446 -1918 -5424
rect -1860 -5446 -1800 -5424
rect -1742 -5446 -1682 -5424
rect -2807 -5462 -2741 -5446
rect -2807 -5496 -2791 -5462
rect -2757 -5496 -2741 -5462
rect -2807 -5512 -2741 -5496
rect -2689 -5462 -2623 -5446
rect -2689 -5496 -2673 -5462
rect -2639 -5496 -2623 -5462
rect -2689 -5512 -2623 -5496
rect -2571 -5462 -2505 -5446
rect -2571 -5496 -2555 -5462
rect -2521 -5496 -2505 -5462
rect -2571 -5512 -2505 -5496
rect -2453 -5462 -2387 -5446
rect -2453 -5496 -2437 -5462
rect -2403 -5496 -2387 -5462
rect -2453 -5512 -2387 -5496
rect -2335 -5462 -2269 -5446
rect -2335 -5496 -2319 -5462
rect -2285 -5496 -2269 -5462
rect -2335 -5512 -2269 -5496
rect -2217 -5462 -2151 -5446
rect -2217 -5496 -2201 -5462
rect -2167 -5496 -2151 -5462
rect -2217 -5512 -2151 -5496
rect -2099 -5462 -2033 -5446
rect -2099 -5496 -2083 -5462
rect -2049 -5496 -2033 -5462
rect -2099 -5512 -2033 -5496
rect -1981 -5462 -1915 -5446
rect -1981 -5496 -1965 -5462
rect -1931 -5496 -1915 -5462
rect -1981 -5512 -1915 -5496
rect -1863 -5462 -1797 -5446
rect -1863 -5496 -1847 -5462
rect -1813 -5496 -1797 -5462
rect -1863 -5512 -1797 -5496
rect -1745 -5462 -1679 -5446
rect -1745 -5496 -1729 -5462
rect -1695 -5496 -1679 -5462
rect -1745 -5512 -1679 -5496
rect -1163 -3524 -1037 -3496
rect -1163 -3558 -1117 -3524
rect -1083 -3558 -1037 -3524
rect -1163 -3574 -1037 -3558
rect 565 -3524 691 -3496
rect 565 -3558 611 -3524
rect 645 -3558 691 -3524
rect 565 -3574 691 -3558
rect -1163 -3600 -1133 -3574
rect -1067 -3600 -1037 -3574
rect -971 -3600 -941 -3574
rect -875 -3600 -845 -3574
rect -779 -3600 -749 -3574
rect -683 -3600 -653 -3574
rect -587 -3600 -557 -3574
rect -491 -3600 -461 -3574
rect -395 -3600 -365 -3574
rect -299 -3600 -269 -3574
rect -203 -3600 -173 -3574
rect -107 -3600 -77 -3574
rect -11 -3600 19 -3574
rect 85 -3600 115 -3574
rect 181 -3600 211 -3574
rect 277 -3600 307 -3574
rect 373 -3600 403 -3574
rect 469 -3600 499 -3574
rect 565 -3600 595 -3574
rect 661 -3600 691 -3574
rect -1163 -4126 -1133 -4100
rect -1067 -4126 -1037 -4100
rect -971 -4122 -941 -4100
rect -875 -4122 -845 -4100
rect -971 -4150 -845 -4122
rect -971 -4184 -925 -4150
rect -891 -4184 -845 -4150
rect -971 -4200 -845 -4184
rect -779 -4122 -749 -4100
rect -683 -4122 -653 -4100
rect -779 -4150 -653 -4122
rect -779 -4184 -733 -4150
rect -699 -4184 -653 -4150
rect -779 -4200 -653 -4184
rect -587 -4122 -557 -4100
rect -491 -4122 -461 -4100
rect -587 -4150 -461 -4122
rect -587 -4184 -541 -4150
rect -507 -4184 -461 -4150
rect -587 -4200 -461 -4184
rect -395 -4122 -365 -4100
rect -299 -4122 -269 -4100
rect -395 -4150 -269 -4122
rect -395 -4184 -349 -4150
rect -315 -4184 -269 -4150
rect -395 -4200 -269 -4184
rect -203 -4122 -173 -4100
rect -107 -4122 -77 -4100
rect -203 -4150 -77 -4122
rect -203 -4184 -157 -4150
rect -123 -4184 -77 -4150
rect -203 -4200 -77 -4184
rect -11 -4122 19 -4100
rect 85 -4122 115 -4100
rect -11 -4150 115 -4122
rect -11 -4184 35 -4150
rect 69 -4184 115 -4150
rect -11 -4200 115 -4184
rect 181 -4122 211 -4100
rect 277 -4122 307 -4100
rect 181 -4150 307 -4122
rect 181 -4184 227 -4150
rect 261 -4184 307 -4150
rect 181 -4200 307 -4184
rect 373 -4122 403 -4100
rect 469 -4122 499 -4100
rect 373 -4150 499 -4122
rect 565 -4126 595 -4100
rect 661 -4126 691 -4100
rect 373 -4184 419 -4150
rect 453 -4184 499 -4150
rect 373 -4200 499 -4184
rect -4238 -5964 -4150 -5948
rect -4238 -5998 -4222 -5964
rect -4188 -5978 -4150 -5964
rect -3650 -5978 -3624 -5948
rect -4188 -5998 -4172 -5978
rect -4238 -6044 -4172 -5998
rect -4238 -6074 -4150 -6044
rect -3650 -6074 -3624 -6044
rect -4238 -6156 -4150 -6140
rect -4238 -6190 -4222 -6156
rect -4188 -6170 -4150 -6156
rect -3650 -6170 -3624 -6140
rect -4188 -6190 -4172 -6170
rect -4238 -6236 -4172 -6190
rect -4238 -6266 -4150 -6236
rect -3650 -6266 -3624 -6236
rect -1123 -4468 -723 -4452
rect -1123 -4502 -1107 -4468
rect -739 -4502 -723 -4468
rect -1123 -4540 -723 -4502
rect -665 -4468 -265 -4452
rect -665 -4502 -649 -4468
rect -281 -4502 -265 -4468
rect -665 -4540 -265 -4502
rect -207 -4468 193 -4452
rect -207 -4502 -191 -4468
rect 177 -4502 193 -4468
rect -207 -4540 193 -4502
rect 251 -4468 651 -4452
rect 251 -4502 267 -4468
rect 635 -4502 651 -4468
rect 251 -4540 651 -4502
rect -1123 -6578 -723 -6540
rect -1123 -6612 -1107 -6578
rect -739 -6612 -723 -6578
rect -1123 -6628 -723 -6612
rect -665 -6578 -265 -6540
rect -665 -6612 -649 -6578
rect -281 -6612 -265 -6578
rect -665 -6628 -265 -6612
rect -207 -6578 193 -6540
rect -207 -6612 -191 -6578
rect 177 -6612 193 -6578
rect -207 -6628 193 -6612
rect 251 -6578 651 -6540
rect 251 -6612 267 -6578
rect 635 -6612 651 -6578
rect 251 -6628 651 -6612
rect 1206 -3352 1272 -3336
rect 1206 -3386 1222 -3352
rect 1256 -3386 1272 -3352
rect 1206 -3402 1272 -3386
rect 1324 -3352 1390 -3336
rect 1324 -3386 1340 -3352
rect 1374 -3386 1390 -3352
rect 1324 -3402 1390 -3386
rect 1442 -3352 1508 -3336
rect 1442 -3386 1458 -3352
rect 1492 -3386 1508 -3352
rect 1442 -3402 1508 -3386
rect 1560 -3352 1626 -3336
rect 1560 -3386 1576 -3352
rect 1610 -3386 1626 -3352
rect 1560 -3402 1626 -3386
rect 1678 -3352 1744 -3336
rect 1678 -3386 1694 -3352
rect 1728 -3386 1744 -3352
rect 1678 -3402 1744 -3386
rect 1796 -3352 1862 -3336
rect 1796 -3386 1812 -3352
rect 1846 -3386 1862 -3352
rect 1796 -3402 1862 -3386
rect 1914 -3352 1980 -3336
rect 1914 -3386 1930 -3352
rect 1964 -3386 1980 -3352
rect 1914 -3402 1980 -3386
rect 2032 -3352 2098 -3336
rect 2032 -3386 2048 -3352
rect 2082 -3386 2098 -3352
rect 2032 -3402 2098 -3386
rect 2150 -3352 2216 -3336
rect 2150 -3386 2166 -3352
rect 2200 -3386 2216 -3352
rect 2150 -3402 2216 -3386
rect 2268 -3352 2334 -3336
rect 2268 -3386 2284 -3352
rect 2318 -3386 2334 -3352
rect 2268 -3402 2334 -3386
rect 1209 -3424 1269 -3402
rect 1327 -3424 1387 -3402
rect 1445 -3424 1505 -3402
rect 1563 -3424 1623 -3402
rect 1681 -3424 1741 -3402
rect 1799 -3424 1859 -3402
rect 1917 -3424 1977 -3402
rect 2035 -3424 2095 -3402
rect 2153 -3424 2213 -3402
rect 2271 -3424 2331 -3402
rect 1209 -5446 1269 -5424
rect 1327 -5446 1387 -5424
rect 1445 -5446 1505 -5424
rect 1563 -5446 1623 -5424
rect 1681 -5446 1741 -5424
rect 1799 -5446 1859 -5424
rect 1917 -5446 1977 -5424
rect 2035 -5446 2095 -5424
rect 2153 -5446 2213 -5424
rect 2271 -5446 2331 -5424
rect 1206 -5462 1272 -5446
rect 1206 -5496 1222 -5462
rect 1256 -5496 1272 -5462
rect 1206 -5512 1272 -5496
rect 1324 -5462 1390 -5446
rect 1324 -5496 1340 -5462
rect 1374 -5496 1390 -5462
rect 1324 -5512 1390 -5496
rect 1442 -5462 1508 -5446
rect 1442 -5496 1458 -5462
rect 1492 -5496 1508 -5462
rect 1442 -5512 1508 -5496
rect 1560 -5462 1626 -5446
rect 1560 -5496 1576 -5462
rect 1610 -5496 1626 -5462
rect 1560 -5512 1626 -5496
rect 1678 -5462 1744 -5446
rect 1678 -5496 1694 -5462
rect 1728 -5496 1744 -5462
rect 1678 -5512 1744 -5496
rect 1796 -5462 1862 -5446
rect 1796 -5496 1812 -5462
rect 1846 -5496 1862 -5462
rect 1796 -5512 1862 -5496
rect 1914 -5462 1980 -5446
rect 1914 -5496 1930 -5462
rect 1964 -5496 1980 -5462
rect 1914 -5512 1980 -5496
rect 2032 -5462 2098 -5446
rect 2032 -5496 2048 -5462
rect 2082 -5496 2098 -5462
rect 2032 -5512 2098 -5496
rect 2150 -5462 2216 -5446
rect 2150 -5496 2166 -5462
rect 2200 -5496 2216 -5462
rect 2150 -5512 2216 -5496
rect 2268 -5462 2334 -5446
rect 2268 -5496 2284 -5462
rect 2318 -5496 2334 -5462
rect 2268 -5512 2334 -5496
<< polycont >>
rect -2790 -868 -2756 -834
rect -2672 -868 -2638 -834
rect -2554 -868 -2520 -834
rect -2436 -868 -2402 -834
rect -2318 -868 -2284 -834
rect -2200 -868 -2166 -834
rect -2082 -868 -2048 -834
rect -1964 -868 -1930 -834
rect -1846 -868 -1812 -834
rect -1728 -868 -1694 -834
rect -1610 -868 -1576 -834
rect -1492 -868 -1458 -834
rect -1374 -868 -1340 -834
rect -1256 -868 -1222 -834
rect -1138 -868 -1104 -834
rect -1020 -868 -986 -834
rect -902 -868 -868 -834
rect -784 -868 -750 -834
rect -666 -868 -632 -834
rect -548 -868 -514 -834
rect 42 -868 76 -834
rect 160 -868 194 -834
rect 278 -868 312 -834
rect 396 -868 430 -834
rect 514 -868 548 -834
rect 632 -868 666 -834
rect 750 -868 784 -834
rect 868 -868 902 -834
rect 986 -868 1020 -834
rect 1104 -868 1138 -834
rect 1222 -868 1256 -834
rect 1340 -868 1374 -834
rect 1458 -868 1492 -834
rect 1576 -868 1610 -834
rect 1694 -868 1728 -834
rect 1812 -868 1846 -834
rect 1930 -868 1964 -834
rect 2048 -868 2082 -834
rect 2166 -868 2200 -834
rect 2284 -868 2318 -834
rect -2790 -2996 -2756 -2962
rect -2672 -2996 -2638 -2962
rect -2554 -2996 -2520 -2962
rect -2436 -2996 -2402 -2962
rect -2318 -2996 -2284 -2962
rect -2200 -2996 -2166 -2962
rect -2082 -2996 -2048 -2962
rect -1964 -2996 -1930 -2962
rect -1846 -2996 -1812 -2962
rect -1728 -2996 -1694 -2962
rect -1610 -2996 -1576 -2962
rect -1492 -2996 -1458 -2962
rect -1374 -2996 -1340 -2962
rect -1256 -2996 -1222 -2962
rect -1138 -2996 -1104 -2962
rect -1020 -2996 -986 -2962
rect -902 -2996 -868 -2962
rect -784 -2996 -750 -2962
rect -666 -2996 -632 -2962
rect -548 -2996 -514 -2962
rect -430 -2996 -396 -2962
rect -312 -2996 -278 -2962
rect -194 -2996 -160 -2962
rect -76 -2996 -42 -2962
rect 42 -2996 76 -2962
rect 160 -2996 194 -2962
rect 278 -2996 312 -2962
rect 396 -2996 430 -2962
rect 514 -2996 548 -2962
rect 632 -2996 666 -2962
rect 750 -2996 784 -2962
rect 868 -2996 902 -2962
rect 986 -2996 1020 -2962
rect 1104 -2996 1138 -2962
rect 1222 -2996 1256 -2962
rect 1340 -2996 1374 -2962
rect 1458 -2996 1492 -2962
rect 1576 -2996 1610 -2962
rect 1694 -2996 1728 -2962
rect 1812 -2996 1846 -2962
rect 1930 -2996 1964 -2962
rect 2048 -2996 2082 -2962
rect 2166 -2996 2200 -2962
rect 2284 -2996 2318 -2962
rect -2791 -3386 -2757 -3352
rect -2673 -3386 -2639 -3352
rect -2555 -3386 -2521 -3352
rect -2437 -3386 -2403 -3352
rect -2319 -3386 -2285 -3352
rect -2201 -3386 -2167 -3352
rect -2083 -3386 -2049 -3352
rect -1965 -3386 -1931 -3352
rect -1847 -3386 -1813 -3352
rect -1729 -3386 -1695 -3352
rect -2791 -5496 -2757 -5462
rect -2673 -5496 -2639 -5462
rect -2555 -5496 -2521 -5462
rect -2437 -5496 -2403 -5462
rect -2319 -5496 -2285 -5462
rect -2201 -5496 -2167 -5462
rect -2083 -5496 -2049 -5462
rect -1965 -5496 -1931 -5462
rect -1847 -5496 -1813 -5462
rect -1729 -5496 -1695 -5462
rect -1117 -3558 -1083 -3524
rect 611 -3558 645 -3524
rect -925 -4184 -891 -4150
rect -733 -4184 -699 -4150
rect -541 -4184 -507 -4150
rect -349 -4184 -315 -4150
rect -157 -4184 -123 -4150
rect 35 -4184 69 -4150
rect 227 -4184 261 -4150
rect 419 -4184 453 -4150
rect -4222 -5998 -4188 -5964
rect -4222 -6190 -4188 -6156
rect -1107 -4502 -739 -4468
rect -649 -4502 -281 -4468
rect -191 -4502 177 -4468
rect 267 -4502 635 -4468
rect -1107 -6612 -739 -6578
rect -649 -6612 -281 -6578
rect -191 -6612 177 -6578
rect 267 -6612 635 -6578
rect 1222 -3386 1256 -3352
rect 1340 -3386 1374 -3352
rect 1458 -3386 1492 -3352
rect 1576 -3386 1610 -3352
rect 1694 -3386 1728 -3352
rect 1812 -3386 1846 -3352
rect 1930 -3386 1964 -3352
rect 2048 -3386 2082 -3352
rect 2166 -3386 2200 -3352
rect 2284 -3386 2318 -3352
rect 1222 -5496 1256 -5462
rect 1340 -5496 1374 -5462
rect 1458 -5496 1492 -5462
rect 1576 -5496 1610 -5462
rect 1694 -5496 1728 -5462
rect 1812 -5496 1846 -5462
rect 1930 -5496 1964 -5462
rect 2048 -5496 2082 -5462
rect 2166 -5496 2200 -5462
rect 2284 -5496 2318 -5462
<< xpolycontact >>
rect -4194 -6504 -3762 -6434
rect -4194 -6670 -3762 -6600
rect 2693 -3812 2831 -3380
rect 2927 -3812 3065 -3380
<< ppolyres >>
rect 2693 -4038 2831 -3812
rect 2927 -4038 3065 -3812
rect 2693 -4176 3065 -4038
<< xpolyres >>
rect -3762 -6504 -3626 -6434
rect -3696 -6600 -3626 -6504
rect -3762 -6670 -3626 -6600
<< locali >>
rect -2963 -766 -2867 -732
rect 2395 -766 2491 -732
rect -2963 -828 -2929 -766
rect 2457 -828 2491 -766
rect -2806 -868 -2790 -834
rect -2756 -868 -2740 -834
rect -2688 -868 -2672 -834
rect -2638 -868 -2622 -834
rect -2570 -868 -2554 -834
rect -2520 -868 -2504 -834
rect -2452 -868 -2436 -834
rect -2402 -868 -2386 -834
rect -2334 -868 -2318 -834
rect -2284 -868 -2268 -834
rect -2216 -868 -2200 -834
rect -2166 -868 -2150 -834
rect -2098 -868 -2082 -834
rect -2048 -868 -2032 -834
rect -1980 -868 -1964 -834
rect -1930 -868 -1914 -834
rect -1862 -868 -1846 -834
rect -1812 -868 -1796 -834
rect -1744 -868 -1728 -834
rect -1694 -868 -1678 -834
rect -1626 -868 -1610 -834
rect -1576 -868 -1560 -834
rect -1508 -868 -1492 -834
rect -1458 -868 -1442 -834
rect -1390 -868 -1374 -834
rect -1340 -868 -1324 -834
rect -1272 -868 -1256 -834
rect -1222 -868 -1206 -834
rect -1154 -868 -1138 -834
rect -1104 -868 -1088 -834
rect -1036 -868 -1020 -834
rect -986 -868 -970 -834
rect -918 -868 -902 -834
rect -868 -868 -852 -834
rect -800 -868 -784 -834
rect -750 -868 -734 -834
rect -682 -868 -666 -834
rect -632 -868 -616 -834
rect -564 -868 -548 -834
rect -514 -868 -498 -834
rect 26 -868 42 -834
rect 76 -868 92 -834
rect 144 -868 160 -834
rect 194 -868 210 -834
rect 262 -868 278 -834
rect 312 -868 328 -834
rect 380 -868 396 -834
rect 430 -868 446 -834
rect 498 -868 514 -834
rect 548 -868 564 -834
rect 616 -868 632 -834
rect 666 -868 682 -834
rect 734 -868 750 -834
rect 784 -868 800 -834
rect 852 -868 868 -834
rect 902 -868 918 -834
rect 970 -868 986 -834
rect 1020 -868 1036 -834
rect 1088 -868 1104 -834
rect 1138 -868 1154 -834
rect 1206 -868 1222 -834
rect 1256 -868 1272 -834
rect 1324 -868 1340 -834
rect 1374 -868 1390 -834
rect 1442 -868 1458 -834
rect 1492 -868 1508 -834
rect 1560 -868 1576 -834
rect 1610 -868 1626 -834
rect 1678 -868 1694 -834
rect 1728 -868 1744 -834
rect 1796 -868 1812 -834
rect 1846 -868 1862 -834
rect 1914 -868 1930 -834
rect 1964 -868 1980 -834
rect 2032 -868 2048 -834
rect 2082 -868 2098 -834
rect 2150 -868 2166 -834
rect 2200 -868 2216 -834
rect 2268 -868 2284 -834
rect 2318 -868 2334 -834
rect -2849 -927 -2815 -911
rect -2849 -2919 -2815 -2903
rect -2731 -927 -2697 -911
rect -2731 -2919 -2697 -2903
rect -2613 -927 -2579 -911
rect -2613 -2919 -2579 -2903
rect -2495 -927 -2461 -911
rect -2495 -2919 -2461 -2903
rect -2377 -927 -2343 -911
rect -2377 -2919 -2343 -2903
rect -2259 -927 -2225 -911
rect -2259 -2919 -2225 -2903
rect -2141 -927 -2107 -911
rect -2141 -2919 -2107 -2903
rect -2023 -927 -1989 -911
rect -2023 -2919 -1989 -2903
rect -1905 -927 -1871 -911
rect -1905 -2919 -1871 -2903
rect -1787 -927 -1753 -911
rect -1787 -2919 -1753 -2903
rect -1669 -927 -1635 -911
rect -1669 -2919 -1635 -2903
rect -1551 -927 -1517 -911
rect -1551 -2919 -1517 -2903
rect -1433 -927 -1399 -911
rect -1433 -2919 -1399 -2903
rect -1315 -927 -1281 -911
rect -1315 -2919 -1281 -2903
rect -1197 -927 -1163 -911
rect -1197 -2919 -1163 -2903
rect -1079 -927 -1045 -911
rect -1079 -2919 -1045 -2903
rect -961 -927 -927 -911
rect -961 -2919 -927 -2903
rect -843 -927 -809 -911
rect -843 -2919 -809 -2903
rect -725 -927 -691 -911
rect -725 -2919 -691 -2903
rect -607 -927 -573 -911
rect -607 -2919 -573 -2903
rect -489 -927 -455 -911
rect -489 -2919 -455 -2903
rect -371 -927 -337 -911
rect -371 -2919 -337 -2903
rect -253 -927 -219 -911
rect -253 -2919 -219 -2903
rect -135 -927 -101 -911
rect -135 -2919 -101 -2903
rect -17 -927 17 -911
rect -17 -2919 17 -2903
rect 101 -927 135 -911
rect 101 -2919 135 -2903
rect 219 -927 253 -911
rect 219 -2919 253 -2903
rect 337 -927 371 -911
rect 337 -2919 371 -2903
rect 455 -927 489 -911
rect 455 -2919 489 -2903
rect 573 -927 607 -911
rect 573 -2919 607 -2903
rect 691 -927 725 -911
rect 691 -2919 725 -2903
rect 809 -927 843 -911
rect 809 -2919 843 -2903
rect 927 -927 961 -911
rect 927 -2919 961 -2903
rect 1045 -927 1079 -911
rect 1045 -2919 1079 -2903
rect 1163 -927 1197 -911
rect 1163 -2919 1197 -2903
rect 1281 -927 1315 -911
rect 1281 -2919 1315 -2903
rect 1399 -927 1433 -911
rect 1399 -2919 1433 -2903
rect 1517 -927 1551 -911
rect 1517 -2919 1551 -2903
rect 1635 -927 1669 -911
rect 1635 -2919 1669 -2903
rect 1753 -927 1787 -911
rect 1753 -2919 1787 -2903
rect 1871 -927 1905 -911
rect 1871 -2919 1905 -2903
rect 1989 -927 2023 -911
rect 1989 -2919 2023 -2903
rect 2107 -927 2141 -911
rect 2107 -2919 2141 -2903
rect 2225 -927 2259 -911
rect 2225 -2919 2259 -2903
rect 2343 -927 2377 -911
rect 2343 -2919 2377 -2903
rect -2806 -2996 -2790 -2962
rect -2756 -2996 -2740 -2962
rect -2688 -2996 -2672 -2962
rect -2638 -2996 -2622 -2962
rect -2570 -2996 -2554 -2962
rect -2520 -2996 -2504 -2962
rect -2452 -2996 -2436 -2962
rect -2402 -2996 -2386 -2962
rect -2334 -2996 -2318 -2962
rect -2284 -2996 -2268 -2962
rect -2216 -2996 -2200 -2962
rect -2166 -2996 -2150 -2962
rect -2098 -2996 -2082 -2962
rect -2048 -2996 -2032 -2962
rect -1980 -2996 -1964 -2962
rect -1930 -2996 -1914 -2962
rect -1862 -2996 -1846 -2962
rect -1812 -2996 -1796 -2962
rect -1744 -2996 -1728 -2962
rect -1694 -2996 -1678 -2962
rect -1626 -2996 -1610 -2962
rect -1576 -2996 -1560 -2962
rect -1508 -2996 -1492 -2962
rect -1458 -2996 -1442 -2962
rect -1390 -2996 -1374 -2962
rect -1340 -2996 -1324 -2962
rect -1272 -2996 -1256 -2962
rect -1222 -2996 -1206 -2962
rect -1154 -2996 -1138 -2962
rect -1104 -2996 -1088 -2962
rect -1036 -2996 -1020 -2962
rect -986 -2996 -970 -2962
rect -918 -2996 -902 -2962
rect -868 -2996 -852 -2962
rect -800 -2996 -784 -2962
rect -750 -2996 -734 -2962
rect -682 -2996 -666 -2962
rect -632 -2996 -616 -2962
rect -564 -2996 -548 -2962
rect -514 -2996 -498 -2962
rect -446 -2996 -430 -2962
rect -396 -2996 -380 -2962
rect -328 -2996 -312 -2962
rect -278 -2996 -262 -2962
rect -210 -2996 -194 -2962
rect -160 -2996 -144 -2962
rect -92 -2996 -76 -2962
rect -42 -2996 -26 -2962
rect 26 -2996 42 -2962
rect 76 -2996 92 -2962
rect 144 -2996 160 -2962
rect 194 -2996 210 -2962
rect 262 -2996 278 -2962
rect 312 -2996 328 -2962
rect 380 -2996 396 -2962
rect 430 -2996 446 -2962
rect 498 -2996 514 -2962
rect 548 -2996 564 -2962
rect 616 -2996 632 -2962
rect 666 -2996 682 -2962
rect 734 -2996 750 -2962
rect 784 -2996 800 -2962
rect 852 -2996 868 -2962
rect 902 -2996 918 -2962
rect 970 -2996 986 -2962
rect 1020 -2996 1036 -2962
rect 1088 -2996 1104 -2962
rect 1138 -2996 1154 -2962
rect 1206 -2996 1222 -2962
rect 1256 -2996 1272 -2962
rect 1324 -2996 1340 -2962
rect 1374 -2996 1390 -2962
rect 1442 -2996 1458 -2962
rect 1492 -2996 1508 -2962
rect 1560 -2996 1576 -2962
rect 1610 -2996 1626 -2962
rect 1678 -2996 1694 -2962
rect 1728 -2996 1744 -2962
rect 1796 -2996 1812 -2962
rect 1846 -2996 1862 -2962
rect 1914 -2996 1930 -2962
rect 1964 -2996 1980 -2962
rect 2032 -2996 2048 -2962
rect 2082 -2996 2098 -2962
rect 2150 -2996 2166 -2962
rect 2200 -2996 2216 -2962
rect 2268 -2996 2284 -2962
rect 2318 -2996 2334 -2962
rect -2963 -3064 -2929 -3002
rect 2457 -3064 2491 -3002
rect -2963 -3098 -2867 -3064
rect 2395 -3098 2491 -3064
rect -2964 -3284 -2868 -3250
rect -1618 -3284 -1522 -3250
rect -2964 -3346 -2930 -3284
rect -1556 -3346 -1522 -3284
rect -2807 -3386 -2791 -3352
rect -2757 -3386 -2741 -3352
rect -2689 -3386 -2673 -3352
rect -2639 -3386 -2623 -3352
rect -2571 -3386 -2555 -3352
rect -2521 -3386 -2505 -3352
rect -2453 -3386 -2437 -3352
rect -2403 -3386 -2387 -3352
rect -2335 -3386 -2319 -3352
rect -2285 -3386 -2269 -3352
rect -2217 -3386 -2201 -3352
rect -2167 -3386 -2151 -3352
rect -2099 -3386 -2083 -3352
rect -2049 -3386 -2033 -3352
rect -1981 -3386 -1965 -3352
rect -1931 -3386 -1915 -3352
rect -1863 -3386 -1847 -3352
rect -1813 -3386 -1797 -3352
rect -1745 -3386 -1729 -3352
rect -1695 -3386 -1679 -3352
rect -2850 -3436 -2816 -3420
rect -2850 -5428 -2816 -5412
rect -2732 -3436 -2698 -3420
rect -2732 -5428 -2698 -5412
rect -2614 -3436 -2580 -3420
rect -2614 -5428 -2580 -5412
rect -2496 -3436 -2462 -3420
rect -2496 -5428 -2462 -5412
rect -2378 -3436 -2344 -3420
rect -2378 -5428 -2344 -5412
rect -2260 -3436 -2226 -3420
rect -2260 -5428 -2226 -5412
rect -2142 -3436 -2108 -3420
rect -2142 -5428 -2108 -5412
rect -2024 -3436 -1990 -3420
rect -2024 -5428 -1990 -5412
rect -1906 -3436 -1872 -3420
rect -1906 -5428 -1872 -5412
rect -1788 -3436 -1754 -3420
rect -1788 -5428 -1754 -5412
rect -1670 -3436 -1636 -3420
rect -1670 -5428 -1636 -5412
rect 1049 -3284 1145 -3250
rect 2395 -3284 2491 -3250
rect 1049 -3346 1083 -3284
rect 2457 -3346 2491 -3284
rect 1206 -3386 1222 -3352
rect 1256 -3386 1272 -3352
rect 1324 -3386 1340 -3352
rect 1374 -3386 1390 -3352
rect 1442 -3386 1458 -3352
rect 1492 -3386 1508 -3352
rect 1560 -3386 1576 -3352
rect 1610 -3386 1626 -3352
rect 1678 -3386 1694 -3352
rect 1728 -3386 1744 -3352
rect 1796 -3386 1812 -3352
rect 1846 -3386 1862 -3352
rect 1914 -3386 1930 -3352
rect 1964 -3386 1980 -3352
rect 2032 -3386 2048 -3352
rect 2082 -3386 2098 -3352
rect 2150 -3386 2166 -3352
rect 2200 -3386 2216 -3352
rect 2268 -3386 2284 -3352
rect 2318 -3386 2334 -3352
rect -1327 -3460 -1231 -3426
rect 759 -3460 855 -3426
rect -1327 -3522 -1293 -3460
rect 821 -3522 855 -3460
rect -1133 -3558 -1117 -3524
rect -1083 -3558 -1067 -3524
rect 595 -3558 611 -3524
rect 645 -3558 661 -3524
rect -1213 -3612 -1179 -3596
rect -1213 -4104 -1179 -4088
rect -1117 -3612 -1083 -3596
rect -1117 -4104 -1083 -4088
rect -1021 -3612 -987 -3596
rect -1021 -4104 -987 -4088
rect -925 -3612 -891 -3596
rect -925 -4104 -891 -4088
rect -829 -3612 -795 -3596
rect -829 -4104 -795 -4088
rect -733 -3612 -699 -3596
rect -733 -4104 -699 -4088
rect -637 -3612 -603 -3596
rect -637 -4104 -603 -4088
rect -541 -3612 -507 -3596
rect -541 -4104 -507 -4088
rect -445 -3612 -411 -3596
rect -445 -4104 -411 -4088
rect -349 -3612 -315 -3596
rect -349 -4104 -315 -4088
rect -253 -3612 -219 -3596
rect -253 -4104 -219 -4088
rect -157 -3612 -123 -3596
rect -157 -4104 -123 -4088
rect -61 -3612 -27 -3596
rect -61 -4104 -27 -4088
rect 35 -3612 69 -3596
rect 35 -4104 69 -4088
rect 131 -3612 165 -3596
rect 131 -4104 165 -4088
rect 227 -3612 261 -3596
rect 227 -4104 261 -4088
rect 323 -3612 357 -3596
rect 323 -4104 357 -4088
rect 419 -3612 453 -3596
rect 419 -4104 453 -4088
rect 515 -3612 549 -3596
rect 515 -4104 549 -4088
rect 611 -3612 645 -3596
rect 611 -4104 645 -4088
rect 707 -3612 741 -3596
rect 707 -4104 741 -4088
rect -1327 -4240 -1293 -4178
rect -941 -4184 -925 -4150
rect -891 -4184 -875 -4150
rect -749 -4184 -733 -4150
rect -699 -4184 -683 -4150
rect -557 -4184 -541 -4150
rect -507 -4184 -491 -4150
rect -365 -4184 -349 -4150
rect -315 -4184 -299 -4150
rect -173 -4184 -157 -4150
rect -123 -4184 -107 -4150
rect 19 -4184 35 -4150
rect 69 -4184 85 -4150
rect 211 -4184 227 -4150
rect 261 -4184 277 -4150
rect 403 -4184 419 -4150
rect 453 -4184 469 -4150
rect 821 -4240 855 -4178
rect -1327 -4274 -1231 -4240
rect 759 -4274 855 -4240
rect -2807 -5496 -2791 -5462
rect -2757 -5496 -2741 -5462
rect -2689 -5496 -2673 -5462
rect -2639 -5496 -2623 -5462
rect -2571 -5496 -2555 -5462
rect -2521 -5496 -2505 -5462
rect -2453 -5496 -2437 -5462
rect -2403 -5496 -2387 -5462
rect -2335 -5496 -2319 -5462
rect -2285 -5496 -2269 -5462
rect -2217 -5496 -2201 -5462
rect -2167 -5496 -2151 -5462
rect -2099 -5496 -2083 -5462
rect -2049 -5496 -2033 -5462
rect -1981 -5496 -1965 -5462
rect -1931 -5496 -1915 -5462
rect -1863 -5496 -1847 -5462
rect -1813 -5496 -1797 -5462
rect -1745 -5496 -1729 -5462
rect -1695 -5496 -1679 -5462
rect -2964 -5564 -2930 -5502
rect -1556 -5564 -1522 -5502
rect -2964 -5598 -2868 -5564
rect -1618 -5598 -1522 -5564
rect -1283 -4400 -1187 -4366
rect 715 -4400 811 -4366
rect -1283 -4462 -1249 -4400
rect 777 -4462 811 -4400
rect -1123 -4502 -1107 -4468
rect -739 -4502 -723 -4468
rect -665 -4502 -649 -4468
rect -281 -4502 -265 -4468
rect -207 -4502 -191 -4468
rect 177 -4502 193 -4468
rect 251 -4502 267 -4468
rect 635 -4502 651 -4468
rect -4358 -5784 -3442 -5750
rect -4358 -5818 -4228 -5784
rect -3572 -5818 -3442 -5784
rect -4358 -5880 -4290 -5818
rect -4358 -6730 -4324 -5880
rect -3510 -5880 -3442 -5818
rect -4154 -5932 -4138 -5898
rect -3662 -5932 -3646 -5898
rect -4222 -5964 -4188 -5948
rect -4222 -6014 -4188 -5998
rect -4154 -6028 -4138 -5994
rect -3662 -6028 -3646 -5994
rect -4154 -6124 -4138 -6090
rect -3662 -6124 -3646 -6090
rect -4222 -6156 -4188 -6140
rect -4222 -6206 -4188 -6190
rect -4154 -6220 -4138 -6186
rect -3662 -6220 -3510 -6186
rect -4233 -6316 -4138 -6282
rect -3662 -6316 -3646 -6282
rect -4233 -6434 -4182 -6316
rect -4233 -6504 -4194 -6434
rect -4233 -6608 -4194 -6600
rect -4233 -6661 -4210 -6608
rect -4233 -6670 -4194 -6661
rect -4358 -6812 -4290 -6730
rect -3476 -5920 -3442 -5880
rect -3476 -5940 -3320 -5920
rect -3476 -6730 -3400 -5940
rect -3510 -6812 -3400 -6730
rect -4358 -6846 -4228 -6812
rect -3572 -6846 -3400 -6812
rect -4358 -6860 -3400 -6846
rect -3340 -6860 -3320 -5940
rect -1169 -4552 -1135 -4536
rect -1169 -6544 -1135 -6528
rect -711 -4552 -677 -4536
rect -711 -6544 -677 -6528
rect -253 -4552 -219 -4536
rect -253 -6544 -219 -6528
rect 205 -4552 239 -4536
rect 205 -6544 239 -6528
rect 663 -4552 697 -4536
rect 663 -6544 697 -6528
rect 1163 -3436 1197 -3420
rect 1163 -5428 1197 -5412
rect 1281 -3436 1315 -3420
rect 1281 -5428 1315 -5412
rect 1399 -3436 1433 -3420
rect 1399 -5428 1433 -5412
rect 1517 -3436 1551 -3420
rect 1517 -5428 1551 -5412
rect 1635 -3436 1669 -3420
rect 1635 -5428 1669 -5412
rect 1753 -3436 1787 -3420
rect 1753 -5428 1787 -5412
rect 1871 -3436 1905 -3420
rect 1871 -5428 1905 -5412
rect 1989 -3436 2023 -3420
rect 1989 -5428 2023 -5412
rect 2107 -3436 2141 -3420
rect 2107 -5428 2141 -5412
rect 2225 -3436 2259 -3420
rect 2225 -5428 2259 -5412
rect 2343 -3436 2377 -3420
rect 2343 -5428 2377 -5412
rect 2563 -3284 2659 -3250
rect 3099 -3284 3195 -3250
rect 2563 -3346 2597 -3284
rect 3161 -3346 3195 -3284
rect 2563 -4272 2597 -4210
rect 3161 -4272 3195 -4210
rect 2563 -4306 2659 -4272
rect 3099 -4306 3195 -4272
rect 1206 -5496 1222 -5462
rect 1256 -5496 1272 -5462
rect 1324 -5496 1340 -5462
rect 1374 -5496 1390 -5462
rect 1442 -5496 1458 -5462
rect 1492 -5496 1508 -5462
rect 1560 -5496 1576 -5462
rect 1610 -5496 1626 -5462
rect 1678 -5496 1694 -5462
rect 1728 -5496 1744 -5462
rect 1796 -5496 1812 -5462
rect 1846 -5496 1862 -5462
rect 1914 -5496 1930 -5462
rect 1964 -5496 1980 -5462
rect 2032 -5496 2048 -5462
rect 2082 -5496 2098 -5462
rect 2150 -5496 2166 -5462
rect 2200 -5496 2216 -5462
rect 2268 -5496 2284 -5462
rect 2318 -5496 2334 -5462
rect 1049 -5564 1083 -5502
rect 2457 -5564 2491 -5502
rect 1049 -5598 1145 -5564
rect 2395 -5598 2491 -5564
rect -1123 -6612 -1107 -6578
rect -739 -6612 -723 -6578
rect -665 -6612 -649 -6578
rect -281 -6612 -265 -6578
rect -207 -6612 -191 -6578
rect 177 -6612 193 -6578
rect 251 -6612 267 -6578
rect 635 -6612 651 -6578
rect -1283 -6680 -1249 -6618
rect 777 -6680 811 -6618
rect -1283 -6714 -1187 -6680
rect 715 -6714 811 -6680
rect -4358 -6880 -3320 -6860
<< viali >>
rect -2790 -868 -2756 -834
rect -2672 -868 -2638 -834
rect -2554 -868 -2520 -834
rect -2436 -868 -2402 -834
rect -2318 -868 -2284 -834
rect -2200 -868 -2166 -834
rect -2082 -868 -2048 -834
rect -1964 -868 -1930 -834
rect -1846 -868 -1812 -834
rect -1728 -868 -1694 -834
rect -1610 -868 -1576 -834
rect -1492 -868 -1458 -834
rect -1374 -868 -1340 -834
rect -1256 -868 -1222 -834
rect -1138 -868 -1104 -834
rect -1020 -868 -986 -834
rect -902 -868 -868 -834
rect -784 -868 -750 -834
rect -666 -868 -632 -834
rect -548 -868 -514 -834
rect 42 -868 76 -834
rect 160 -868 194 -834
rect 278 -868 312 -834
rect 396 -868 430 -834
rect 514 -868 548 -834
rect 632 -868 666 -834
rect 750 -868 784 -834
rect 868 -868 902 -834
rect 986 -868 1020 -834
rect 1104 -868 1138 -834
rect 1222 -868 1256 -834
rect 1340 -868 1374 -834
rect 1458 -868 1492 -834
rect 1576 -868 1610 -834
rect 1694 -868 1728 -834
rect 1812 -868 1846 -834
rect 1930 -868 1964 -834
rect 2048 -868 2082 -834
rect 2166 -868 2200 -834
rect 2284 -868 2318 -834
rect -2963 -1315 -2929 -915
rect -2963 -2915 -2929 -2515
rect -2849 -2903 -2815 -927
rect -2731 -2903 -2697 -927
rect -2613 -2903 -2579 -927
rect -2495 -2903 -2461 -927
rect -2377 -2903 -2343 -927
rect -2259 -2903 -2225 -927
rect -2141 -2903 -2107 -927
rect -2023 -2903 -1989 -927
rect -1905 -2903 -1871 -927
rect -1787 -2903 -1753 -927
rect -1669 -2903 -1635 -927
rect -1551 -2903 -1517 -927
rect -1433 -2903 -1399 -927
rect -1315 -2903 -1281 -927
rect -1197 -2903 -1163 -927
rect -1079 -2903 -1045 -927
rect -961 -2903 -927 -927
rect -843 -2903 -809 -927
rect -725 -2903 -691 -927
rect -607 -2903 -573 -927
rect -489 -2903 -455 -927
rect -371 -2903 -337 -927
rect -253 -2903 -219 -927
rect -135 -2903 -101 -927
rect -17 -2903 17 -927
rect 101 -2903 135 -927
rect 219 -2903 253 -927
rect 337 -2903 371 -927
rect 455 -2903 489 -927
rect 573 -2903 607 -927
rect 691 -2903 725 -927
rect 809 -2903 843 -927
rect 927 -2903 961 -927
rect 1045 -2903 1079 -927
rect 1163 -2903 1197 -927
rect 1281 -2903 1315 -927
rect 1399 -2903 1433 -927
rect 1517 -2903 1551 -927
rect 1635 -2903 1669 -927
rect 1753 -2903 1787 -927
rect 1871 -2903 1905 -927
rect 1989 -2903 2023 -927
rect 2107 -2903 2141 -927
rect 2225 -2903 2259 -927
rect 2343 -2903 2377 -927
rect 2457 -1315 2491 -915
rect 2457 -2915 2491 -2515
rect -2790 -2996 -2756 -2962
rect -2672 -2996 -2638 -2962
rect -2554 -2996 -2520 -2962
rect -2436 -2996 -2402 -2962
rect -2318 -2996 -2284 -2962
rect -2200 -2996 -2166 -2962
rect -2082 -2996 -2048 -2962
rect -1964 -2996 -1930 -2962
rect -1846 -2996 -1812 -2962
rect -1728 -2996 -1694 -2962
rect -1610 -2996 -1576 -2962
rect -1492 -2996 -1458 -2962
rect -1374 -2996 -1340 -2962
rect -1256 -2996 -1222 -2962
rect -1138 -2996 -1104 -2962
rect -1020 -2996 -986 -2962
rect -902 -2996 -868 -2962
rect -784 -2996 -750 -2962
rect -666 -2996 -632 -2962
rect -548 -2996 -514 -2962
rect -430 -2996 -396 -2962
rect -312 -2996 -278 -2962
rect -194 -2996 -160 -2962
rect -76 -2996 -42 -2962
rect 42 -2996 76 -2962
rect 160 -2996 194 -2962
rect 278 -2996 312 -2962
rect 396 -2996 430 -2962
rect 514 -2996 548 -2962
rect 632 -2996 666 -2962
rect 750 -2996 784 -2962
rect 868 -2996 902 -2962
rect 986 -2996 1020 -2962
rect 1104 -2996 1138 -2962
rect 1222 -2996 1256 -2962
rect 1340 -2996 1374 -2962
rect 1458 -2996 1492 -2962
rect 1576 -2996 1610 -2962
rect 1694 -2996 1728 -2962
rect 1812 -2996 1846 -2962
rect 1930 -2996 1964 -2962
rect 2048 -2996 2082 -2962
rect 2166 -2996 2200 -2962
rect 2284 -2996 2318 -2962
rect -2791 -3386 -2757 -3352
rect -2673 -3386 -2639 -3352
rect -2555 -3386 -2521 -3352
rect -2437 -3386 -2403 -3352
rect -2319 -3386 -2285 -3352
rect -2201 -3386 -2167 -3352
rect -2083 -3386 -2049 -3352
rect -1965 -3386 -1931 -3352
rect -1847 -3386 -1813 -3352
rect -1729 -3386 -1695 -3352
rect -2964 -3824 -2930 -3424
rect -2964 -5424 -2930 -5024
rect -2850 -5412 -2816 -3436
rect -2732 -5412 -2698 -3436
rect -2614 -5412 -2580 -3436
rect -2496 -5412 -2462 -3436
rect -2378 -5412 -2344 -3436
rect -2260 -5412 -2226 -3436
rect -2142 -5412 -2108 -3436
rect -2024 -5412 -1990 -3436
rect -1906 -5412 -1872 -3436
rect -1788 -5412 -1754 -3436
rect -1670 -5412 -1636 -3436
rect -1556 -3824 -1522 -3424
rect 1222 -3386 1256 -3352
rect 1340 -3386 1374 -3352
rect 1458 -3386 1492 -3352
rect 1576 -3386 1610 -3352
rect 1694 -3386 1728 -3352
rect 1812 -3386 1846 -3352
rect 1930 -3386 1964 -3352
rect 2048 -3386 2082 -3352
rect 2166 -3386 2200 -3352
rect 2284 -3386 2318 -3352
rect -1117 -3558 -1083 -3524
rect 611 -3558 645 -3524
rect -1327 -4100 -1293 -3600
rect -1213 -4088 -1179 -3612
rect -1117 -4088 -1083 -3612
rect -1021 -4088 -987 -3612
rect -925 -4088 -891 -3612
rect -829 -4088 -795 -3612
rect -733 -4088 -699 -3612
rect -637 -4088 -603 -3612
rect -541 -4088 -507 -3612
rect -445 -4088 -411 -3612
rect -349 -4088 -315 -3612
rect -253 -4088 -219 -3612
rect -157 -4088 -123 -3612
rect -61 -4088 -27 -3612
rect 35 -4088 69 -3612
rect 131 -4088 165 -3612
rect 227 -4088 261 -3612
rect 323 -4088 357 -3612
rect 419 -4088 453 -3612
rect 515 -4088 549 -3612
rect 611 -4088 645 -3612
rect 707 -4088 741 -3612
rect 821 -4100 855 -3600
rect -925 -4184 -891 -4150
rect -733 -4184 -699 -4150
rect -541 -4184 -507 -4150
rect -349 -4184 -315 -4150
rect -157 -4184 -123 -4150
rect 35 -4184 69 -4150
rect 227 -4184 261 -4150
rect 419 -4184 453 -4150
rect 1049 -3824 1083 -3424
rect -1556 -5424 -1522 -5024
rect -2791 -5496 -2757 -5462
rect -2673 -5496 -2639 -5462
rect -2555 -5496 -2521 -5462
rect -2437 -5496 -2403 -5462
rect -2319 -5496 -2285 -5462
rect -2201 -5496 -2167 -5462
rect -2083 -5496 -2049 -5462
rect -1965 -5496 -1931 -5462
rect -1847 -5496 -1813 -5462
rect -1729 -5496 -1695 -5462
rect -1107 -4502 -739 -4468
rect -649 -4502 -281 -4468
rect -191 -4502 177 -4468
rect 267 -4502 635 -4468
rect -1283 -4940 -1249 -4540
rect -4138 -5932 -3662 -5898
rect -4222 -5998 -4188 -5964
rect -4138 -6028 -3662 -5994
rect -4138 -6124 -3662 -6090
rect -4222 -6190 -4188 -6156
rect -4138 -6220 -3662 -6186
rect -4138 -6316 -3662 -6282
rect -4210 -6661 -4194 -6608
rect -4194 -6661 -3778 -6608
rect -3400 -6860 -3340 -5940
rect -1283 -6540 -1249 -6140
rect -1169 -6528 -1135 -4552
rect -711 -6528 -677 -4552
rect -253 -6528 -219 -4552
rect 205 -6528 239 -4552
rect 663 -6528 697 -4552
rect 777 -4940 811 -4540
rect 1049 -5424 1083 -5024
rect 1163 -5412 1197 -3436
rect 1281 -5412 1315 -3436
rect 1399 -5412 1433 -3436
rect 1517 -5412 1551 -3436
rect 1635 -5412 1669 -3436
rect 1753 -5412 1787 -3436
rect 1871 -5412 1905 -3436
rect 1989 -5412 2023 -3436
rect 2107 -5412 2141 -3436
rect 2225 -5412 2259 -3436
rect 2343 -5412 2377 -3436
rect 2457 -3824 2491 -3424
rect 2720 -3780 2800 -3420
rect 2960 -3780 3040 -3420
rect 2457 -5424 2491 -5024
rect 1222 -5496 1256 -5462
rect 1340 -5496 1374 -5462
rect 1458 -5496 1492 -5462
rect 1576 -5496 1610 -5462
rect 1694 -5496 1728 -5462
rect 1812 -5496 1846 -5462
rect 1930 -5496 1964 -5462
rect 2048 -5496 2082 -5462
rect 2166 -5496 2200 -5462
rect 2284 -5496 2318 -5462
rect 777 -6540 811 -6140
rect -1107 -6612 -739 -6578
rect -649 -6612 -281 -6578
rect -191 -6612 177 -6578
rect 267 -6612 635 -6578
<< metal1 >>
rect -2858 -834 -2626 -828
rect -2858 -868 -2790 -834
rect -2756 -868 -2672 -834
rect -2638 -868 -2626 -834
rect -2858 -874 -2626 -868
rect -2566 -834 -502 -828
rect -2566 -868 -2554 -834
rect -2520 -868 -2436 -834
rect -2402 -868 -2318 -834
rect -2284 -868 -2200 -834
rect -2166 -868 -2082 -834
rect -2048 -868 -1964 -834
rect -1930 -868 -1846 -834
rect -1812 -868 -1728 -834
rect -1694 -868 -1610 -834
rect -1576 -868 -1492 -834
rect -1458 -868 -1374 -834
rect -1340 -868 -1256 -834
rect -1222 -868 -1138 -834
rect -1104 -868 -1020 -834
rect -986 -868 -902 -834
rect -868 -868 -784 -834
rect -750 -868 -666 -834
rect -632 -868 -548 -834
rect -514 -868 -502 -834
rect -2566 -874 -502 -868
rect 30 -834 2094 -828
rect 30 -868 42 -834
rect 76 -868 160 -834
rect 194 -868 278 -834
rect 312 -868 396 -834
rect 430 -868 514 -834
rect 548 -868 632 -834
rect 666 -868 750 -834
rect 784 -868 868 -834
rect 902 -868 986 -834
rect 1020 -868 1104 -834
rect 1138 -868 1222 -834
rect 1256 -868 1340 -834
rect 1374 -868 1458 -834
rect 1492 -868 1576 -834
rect 1610 -868 1694 -834
rect 1728 -868 1812 -834
rect 1846 -868 1930 -834
rect 1964 -868 2048 -834
rect 2082 -868 2094 -834
rect 30 -874 2094 -868
rect 2154 -834 2386 -828
rect 2154 -868 2166 -834
rect 2200 -868 2284 -834
rect 2318 -868 2386 -834
rect 2154 -874 2386 -868
rect -2969 -915 -2923 -903
rect -2858 -915 -2806 -874
rect -2969 -1315 -2963 -915
rect -2929 -927 -2806 -915
rect -2929 -1315 -2858 -927
rect -2969 -1327 -2923 -1315
rect -2969 -2515 -2923 -2503
rect -2969 -2915 -2963 -2515
rect -2929 -2903 -2858 -2515
rect -2929 -2915 -2806 -2903
rect -2969 -2927 -2923 -2915
rect -2858 -2956 -2806 -2915
rect -2740 -927 -2688 -874
rect -2740 -2956 -2688 -2903
rect -2622 -927 -2570 -915
rect -2622 -2915 -2570 -2903
rect -2504 -927 -2452 -915
rect -2504 -2915 -2452 -2903
rect -2386 -927 -2334 -915
rect -2386 -2915 -2334 -2903
rect -2268 -927 -2216 -915
rect -2268 -2915 -2216 -2903
rect -2150 -927 -2098 -915
rect -2150 -2915 -2098 -2903
rect -2032 -927 -1980 -915
rect -2032 -2915 -1980 -2903
rect -1914 -927 -1862 -915
rect -1914 -2915 -1862 -2903
rect -1796 -927 -1744 -915
rect -1796 -2915 -1744 -2903
rect -1678 -927 -1626 -915
rect -1678 -2915 -1626 -2903
rect -1560 -927 -1508 -915
rect -1560 -2915 -1508 -2903
rect -1442 -927 -1390 -915
rect -1442 -2915 -1390 -2903
rect -1324 -927 -1272 -915
rect -1324 -2915 -1272 -2903
rect -1206 -927 -1154 -915
rect -1206 -2915 -1154 -2903
rect -1088 -927 -1036 -915
rect -1088 -2915 -1036 -2903
rect -970 -927 -918 -915
rect -970 -2915 -918 -2903
rect -852 -927 -800 -915
rect -852 -2915 -800 -2903
rect -734 -927 -682 -915
rect -734 -2915 -682 -2903
rect -616 -927 -564 -874
rect -616 -2956 -564 -2903
rect -498 -927 -446 -915
rect -498 -2915 -446 -2903
rect -380 -927 -328 -915
rect -380 -2950 -328 -2903
rect -262 -927 -210 -915
rect -262 -2915 -210 -2903
rect -144 -927 -92 -915
rect -380 -2956 -262 -2950
rect -144 -2956 -92 -2903
rect -26 -927 26 -915
rect -26 -2915 26 -2903
rect 92 -927 144 -874
rect 92 -2956 144 -2903
rect 210 -927 262 -915
rect 210 -2915 262 -2903
rect 328 -927 380 -915
rect 328 -2915 380 -2903
rect 446 -927 498 -915
rect 446 -2915 498 -2903
rect 564 -927 616 -915
rect 564 -2915 616 -2903
rect 682 -927 734 -915
rect 682 -2915 734 -2903
rect 800 -927 852 -915
rect 800 -2915 852 -2903
rect 918 -927 970 -915
rect 918 -2915 970 -2903
rect 1036 -927 1088 -915
rect 1036 -2915 1088 -2903
rect 1154 -927 1206 -915
rect 1154 -2915 1206 -2903
rect 1272 -927 1324 -915
rect 1272 -2915 1324 -2903
rect 1390 -927 1442 -915
rect 1390 -2915 1442 -2903
rect 1508 -927 1560 -915
rect 1508 -2915 1560 -2903
rect 1626 -927 1678 -915
rect 1626 -2915 1678 -2903
rect 1744 -927 1796 -915
rect 1744 -2915 1796 -2903
rect 1862 -927 1914 -915
rect 1862 -2915 1914 -2903
rect 1980 -927 2032 -915
rect 1980 -2915 2032 -2903
rect 2098 -927 2150 -915
rect 2098 -2915 2150 -2903
rect 2216 -927 2268 -874
rect 2216 -2956 2268 -2903
rect 2334 -915 2386 -874
rect 2451 -915 2497 -903
rect 2334 -927 2457 -915
rect 2386 -1315 2457 -927
rect 2491 -1315 2497 -915
rect 2451 -1327 2497 -1315
rect 2451 -2515 2497 -2503
rect 2386 -2903 2457 -2515
rect 2334 -2915 2457 -2903
rect 2491 -2915 2497 -2515
rect 2334 -2956 2386 -2915
rect 2451 -2927 2497 -2915
rect -2858 -2962 -2626 -2956
rect -2858 -2996 -2790 -2962
rect -2756 -2996 -2672 -2962
rect -2638 -2996 -2626 -2962
rect -2858 -3002 -2626 -2996
rect -2566 -2962 -262 -2956
rect -2566 -2996 -2554 -2962
rect -2520 -2996 -2436 -2962
rect -2402 -2996 -2318 -2962
rect -2284 -2996 -2200 -2962
rect -2166 -2996 -2082 -2962
rect -2048 -2996 -1964 -2962
rect -1930 -2996 -1846 -2962
rect -1812 -2996 -1728 -2962
rect -1694 -2996 -1610 -2962
rect -1576 -2996 -1492 -2962
rect -1458 -2996 -1374 -2962
rect -1340 -2996 -1256 -2962
rect -1222 -2996 -1138 -2962
rect -1104 -2996 -1020 -2962
rect -986 -2996 -902 -2962
rect -868 -2996 -784 -2962
rect -750 -2996 -666 -2962
rect -632 -2996 -548 -2962
rect -514 -2996 -430 -2962
rect -396 -2996 -312 -2962
rect -278 -2996 -262 -2962
rect -2566 -3002 -262 -2996
rect -328 -3019 -262 -3002
rect -206 -2962 2094 -2956
rect -206 -2996 -194 -2962
rect -160 -2996 -76 -2962
rect -42 -2996 42 -2962
rect 76 -2996 160 -2962
rect 194 -2996 278 -2962
rect 312 -2996 396 -2962
rect 430 -2996 514 -2962
rect 548 -2996 632 -2962
rect 666 -2996 750 -2962
rect 784 -2996 868 -2962
rect 902 -2996 986 -2962
rect 1020 -2996 1104 -2962
rect 1138 -2996 1222 -2962
rect 1256 -2996 1340 -2962
rect 1374 -2996 1458 -2962
rect 1492 -2996 1576 -2962
rect 1610 -2996 1694 -2962
rect 1728 -2996 1812 -2962
rect 1846 -2996 1930 -2962
rect 1964 -2996 2048 -2962
rect 2082 -2996 2094 -2962
rect -206 -3002 2094 -2996
rect 2154 -2962 2386 -2956
rect 2154 -2996 2166 -2962
rect 2200 -2996 2284 -2962
rect 2318 -2996 2386 -2962
rect 2154 -3002 2386 -2996
rect -206 -3013 -147 -3002
rect -2505 -3242 -2453 -3236
rect -2505 -3346 -2453 -3294
rect -2269 -3242 -2217 -3236
rect -2269 -3346 -2217 -3294
rect -2033 -3242 -1981 -3236
rect -2033 -3346 -1981 -3294
rect 1508 -3242 1560 -3236
rect 1508 -3346 1560 -3294
rect 1744 -3242 1796 -3236
rect 1744 -3346 1796 -3294
rect 1980 -3242 2032 -3236
rect 1980 -3346 2032 -3294
rect -2859 -3352 -2745 -3346
rect -2859 -3386 -2791 -3352
rect -2757 -3386 -2745 -3352
rect -2859 -3392 -2745 -3386
rect -2685 -3352 -1801 -3346
rect -2685 -3386 -2673 -3352
rect -2639 -3386 -2555 -3352
rect -2521 -3386 -2437 -3352
rect -2403 -3386 -2319 -3352
rect -2285 -3386 -2201 -3352
rect -2167 -3386 -2083 -3352
rect -2049 -3386 -1965 -3352
rect -1931 -3386 -1847 -3352
rect -1813 -3386 -1801 -3352
rect -2685 -3392 -1801 -3386
rect -1741 -3352 -1627 -3346
rect -1741 -3386 -1729 -3352
rect -1695 -3386 -1627 -3352
rect -1741 -3392 -1627 -3386
rect -2970 -3424 -2924 -3412
rect -2859 -3424 -2807 -3392
rect -1679 -3424 -1627 -3392
rect 1154 -3352 1268 -3346
rect 1154 -3386 1222 -3352
rect 1256 -3386 1268 -3352
rect 1154 -3392 1268 -3386
rect 1328 -3352 2212 -3346
rect 1328 -3386 1340 -3352
rect 1374 -3386 1458 -3352
rect 1492 -3386 1576 -3352
rect 1610 -3386 1694 -3352
rect 1728 -3386 1812 -3352
rect 1846 -3386 1930 -3352
rect 1964 -3386 2048 -3352
rect 2082 -3386 2166 -3352
rect 2200 -3386 2212 -3352
rect 1328 -3392 2212 -3386
rect 2272 -3352 2386 -3346
rect 2272 -3386 2284 -3352
rect 2318 -3386 2386 -3352
rect 2272 -3392 2386 -3386
rect -1536 -3412 -1436 -3400
rect -1562 -3424 -1436 -3412
rect -2970 -3824 -2964 -3424
rect -2930 -3436 -2807 -3424
rect -2930 -3824 -2859 -3436
rect -2970 -3836 -2924 -3824
rect -2970 -5024 -2924 -5012
rect -2970 -5424 -2964 -5024
rect -2930 -5412 -2859 -5024
rect -2930 -5424 -2807 -5412
rect -2741 -3436 -2689 -3424
rect -2741 -5424 -2689 -5412
rect -2623 -3436 -2571 -3424
rect -2623 -5424 -2571 -5412
rect -2505 -3436 -2453 -3424
rect -2505 -5424 -2453 -5412
rect -2387 -3436 -2335 -3424
rect -2387 -5424 -2335 -5412
rect -2269 -3436 -2217 -3424
rect -2269 -5424 -2217 -5412
rect -2151 -3436 -2099 -3424
rect -2151 -5424 -2099 -5412
rect -2033 -3436 -1981 -3424
rect -2033 -5424 -1981 -5412
rect -1915 -3436 -1863 -3424
rect -1915 -5424 -1863 -5412
rect -1797 -3436 -1745 -3424
rect -1797 -5424 -1745 -5412
rect -1679 -3436 -1556 -3424
rect -1627 -3824 -1556 -3436
rect -1522 -3500 -1436 -3424
rect 964 -3412 1064 -3400
rect 964 -3424 1089 -3412
rect 1154 -3424 1206 -3392
rect 2334 -3424 2386 -3392
rect 2451 -3424 2497 -3412
rect 964 -3500 1049 -3424
rect -1522 -3600 -1276 -3500
rect -1219 -3524 -1067 -3518
rect -1219 -3558 -1117 -3524
rect -1083 -3558 -1067 -3524
rect -1219 -3564 -1067 -3558
rect 595 -3524 747 -3518
rect 595 -3558 611 -3524
rect 645 -3558 747 -3524
rect 595 -3564 747 -3558
rect -1219 -3600 -1173 -3564
rect -1123 -3600 -1077 -3564
rect 605 -3600 651 -3564
rect 701 -3600 747 -3564
rect 804 -3600 1049 -3500
rect -1522 -3824 -1327 -3600
rect -1562 -3836 -1327 -3824
rect -1536 -4000 -1327 -3836
rect -1436 -4100 -1327 -4000
rect -1293 -4100 -1223 -3600
rect -1169 -4100 -1163 -3600
rect -1133 -4100 -1127 -3600
rect -1073 -4100 -1067 -3600
rect -1037 -4100 -1031 -3600
rect -977 -4100 -971 -3600
rect -941 -4100 -935 -3600
rect -881 -4100 -875 -3600
rect -845 -4100 -839 -3600
rect -785 -4100 -779 -3600
rect -749 -4100 -743 -3600
rect -689 -4100 -683 -3600
rect -653 -4100 -647 -3600
rect -593 -4100 -587 -3600
rect -557 -4100 -551 -3600
rect -497 -4100 -491 -3600
rect -461 -4100 -455 -3600
rect -401 -4100 -395 -3600
rect -365 -4100 -359 -3600
rect -305 -4100 -299 -3600
rect -269 -4100 -263 -3600
rect -209 -4100 -203 -3600
rect -173 -4100 -167 -3600
rect -113 -4100 -107 -3600
rect -77 -4100 -71 -3600
rect -17 -4100 -11 -3600
rect 19 -4100 25 -3600
rect 79 -4100 85 -3600
rect 115 -4100 121 -3600
rect 175 -4100 181 -3600
rect 211 -4100 217 -3600
rect 271 -4100 277 -3600
rect 307 -4100 313 -3600
rect 367 -4100 373 -3600
rect 403 -4100 409 -3600
rect 463 -4100 469 -3600
rect 499 -4100 505 -3600
rect 559 -4100 565 -3600
rect 595 -4100 601 -3600
rect 655 -4100 661 -3600
rect 691 -4100 697 -3600
rect 751 -4100 821 -3600
rect 855 -3824 1049 -3600
rect 1083 -3436 1206 -3424
rect 1083 -3824 1154 -3436
rect 855 -3836 1089 -3824
rect 855 -4000 1064 -3836
rect 855 -4100 964 -4000
rect -1436 -4400 -1276 -4100
rect -947 -4200 -941 -4144
rect -875 -4200 -869 -4144
rect -755 -4200 -749 -4144
rect -683 -4200 -677 -4144
rect -563 -4200 -557 -4144
rect -491 -4200 -485 -4144
rect -371 -4200 -365 -4144
rect -299 -4200 -293 -4144
rect -179 -4200 -173 -4144
rect -107 -4200 -101 -4144
rect 13 -4200 19 -4144
rect 85 -4200 91 -4144
rect 205 -4200 211 -4144
rect 277 -4200 283 -4144
rect 397 -4200 403 -4144
rect 469 -4200 475 -4144
rect -1436 -4540 -1236 -4400
rect -1200 -4440 -1120 -4430
rect -1200 -4500 -1190 -4440
rect -1130 -4462 -1120 -4440
rect -1130 -4468 647 -4462
rect -1130 -4500 -1107 -4468
rect -1200 -4502 -1107 -4500
rect -739 -4502 -649 -4468
rect -281 -4502 -191 -4468
rect 177 -4502 267 -4468
rect 635 -4502 647 -4468
rect -1200 -4508 647 -4502
rect -1200 -4510 -1120 -4508
rect 804 -4528 964 -4100
rect 771 -4540 964 -4528
rect -1436 -4900 -1283 -4540
rect -1536 -4940 -1283 -4900
rect -1249 -4552 -1126 -4540
rect -1249 -4940 -1178 -4552
rect -1536 -5000 -1236 -4940
rect -1536 -5012 -1276 -5000
rect -1562 -5024 -1276 -5012
rect -1627 -5412 -1556 -5024
rect -1679 -5424 -1556 -5412
rect -1522 -5424 -1276 -5024
rect -2970 -5436 -2924 -5424
rect -2859 -5456 -2807 -5424
rect -1679 -5456 -1627 -5424
rect -1562 -5436 -1276 -5424
rect -2859 -5462 -2745 -5456
rect -2859 -5496 -2791 -5462
rect -2757 -5496 -2745 -5462
rect -2859 -5502 -2745 -5496
rect -2685 -5462 -1801 -5456
rect -2685 -5496 -2673 -5462
rect -2639 -5496 -2555 -5462
rect -2521 -5496 -2437 -5462
rect -2403 -5496 -2319 -5462
rect -2285 -5496 -2201 -5462
rect -2167 -5496 -2083 -5462
rect -2049 -5496 -1965 -5462
rect -1931 -5496 -1847 -5462
rect -1813 -5496 -1801 -5462
rect -2685 -5502 -1801 -5496
rect -1741 -5462 -1627 -5456
rect -1741 -5496 -1729 -5462
rect -1695 -5496 -1627 -5462
rect -1741 -5502 -1627 -5496
rect -1536 -5500 -1276 -5436
rect -1436 -5560 -1276 -5500
rect -4150 -5898 -3542 -5892
rect -4150 -5932 -4138 -5898
rect -3662 -5932 -3542 -5898
rect -4150 -5938 -3542 -5932
rect -4228 -5964 -4182 -5948
rect -4228 -5994 -4222 -5964
rect -4363 -5998 -4222 -5994
rect -4188 -5998 -4182 -5964
rect -4363 -6028 -4182 -5998
rect -4151 -5994 -4134 -5985
rect -3665 -5994 -3650 -5985
rect -4151 -6028 -4138 -5994
rect -3662 -6028 -3650 -5994
rect -4363 -6884 -4329 -6028
rect -4151 -6037 -4134 -6028
rect -3665 -6037 -3650 -6028
rect -3582 -6084 -3542 -5938
rect -4150 -6090 -3542 -6084
rect -4150 -6124 -4138 -6090
rect -3662 -6124 -3542 -6090
rect -4150 -6130 -3542 -6124
rect -4228 -6156 -4182 -6140
rect -4228 -6186 -4222 -6156
rect -4369 -7084 -4329 -6884
rect -4301 -6190 -4222 -6186
rect -4188 -6190 -4182 -6156
rect -4301 -6220 -4182 -6190
rect -4150 -6186 -3650 -6180
rect -4150 -6220 -4138 -6186
rect -3662 -6220 -3650 -6186
rect -4301 -6884 -4267 -6220
rect -4150 -6226 -3650 -6220
rect -3582 -6276 -3542 -6130
rect -4150 -6282 -3542 -6276
rect -4150 -6316 -4138 -6282
rect -3662 -6316 -3542 -6282
rect -4150 -6322 -3542 -6316
rect -3420 -5940 -3180 -5920
rect -4233 -6670 -4210 -6600
rect -3781 -6608 -3762 -6600
rect -3778 -6661 -3762 -6608
rect -3781 -6670 -3762 -6661
rect -3420 -6860 -3400 -5940
rect -3200 -6860 -3180 -5940
rect -1436 -6780 -1416 -5560
rect -1356 -6128 -1276 -5560
rect -1356 -6140 -1243 -6128
rect -1356 -6540 -1283 -6140
rect -1249 -6528 -1178 -6140
rect -1249 -6540 -1126 -6528
rect -720 -4552 -668 -4540
rect -720 -6540 -668 -6528
rect -262 -4552 -210 -4540
rect -262 -6540 -210 -6528
rect 196 -4552 248 -4540
rect 196 -6540 248 -6528
rect 654 -4552 777 -4540
rect 706 -4940 777 -4552
rect 811 -4900 964 -4540
rect 811 -4940 1064 -4900
rect 771 -4952 1064 -4940
rect 804 -5012 1064 -4952
rect 804 -5024 1089 -5012
rect 804 -5424 1049 -5024
rect 1083 -5412 1154 -5024
rect 1083 -5424 1206 -5412
rect 1272 -3436 1324 -3424
rect 1272 -5424 1324 -5412
rect 1390 -3436 1442 -3424
rect 1390 -5424 1442 -5412
rect 1508 -3436 1560 -3424
rect 1508 -5424 1560 -5412
rect 1626 -3436 1678 -3424
rect 1626 -5424 1678 -5412
rect 1744 -3436 1796 -3424
rect 1744 -5424 1796 -5412
rect 1862 -3436 1914 -3424
rect 1862 -5424 1914 -5412
rect 1980 -3436 2032 -3424
rect 1980 -5424 2032 -5412
rect 2098 -3436 2150 -3424
rect 2098 -5424 2150 -5412
rect 2216 -3436 2268 -3424
rect 2216 -5424 2268 -5412
rect 2334 -3436 2457 -3424
rect 2386 -3824 2457 -3436
rect 2491 -3824 2497 -3424
rect 2700 -3420 2820 -3400
rect 2700 -3780 2720 -3420
rect 2800 -3780 2820 -3420
rect 2700 -3800 2820 -3780
rect 2940 -3420 3060 -3400
rect 2940 -3780 2960 -3420
rect 3040 -3780 3060 -3420
rect 2940 -3800 3060 -3780
rect 2451 -3836 2497 -3824
rect 2451 -5024 2497 -5012
rect 2386 -5412 2457 -5024
rect 2334 -5424 2457 -5412
rect 2491 -5424 2497 -5024
rect 804 -5436 1089 -5424
rect 804 -5500 1064 -5436
rect 1154 -5456 1206 -5424
rect 2334 -5456 2386 -5424
rect 2451 -5436 2497 -5424
rect 1154 -5462 1268 -5456
rect 1154 -5496 1222 -5462
rect 1256 -5496 1268 -5462
rect 804 -5560 964 -5500
rect 1154 -5502 1268 -5496
rect 1328 -5462 2212 -5456
rect 1328 -5496 1340 -5462
rect 1374 -5496 1458 -5462
rect 1492 -5496 1576 -5462
rect 1610 -5496 1694 -5462
rect 1728 -5496 1812 -5462
rect 1846 -5496 1930 -5462
rect 1964 -5496 2048 -5462
rect 2082 -5496 2166 -5462
rect 2200 -5496 2212 -5462
rect 1328 -5502 2212 -5496
rect 2272 -5462 2386 -5456
rect 2272 -5496 2284 -5462
rect 2318 -5496 2386 -5462
rect 2272 -5502 2386 -5496
rect 804 -6128 884 -5560
rect 771 -6140 884 -6128
rect 706 -6528 777 -6140
rect 654 -6540 777 -6528
rect 811 -6540 884 -6140
rect -1356 -6552 -1243 -6540
rect 771 -6552 884 -6540
rect -1356 -6780 -1276 -6552
rect -1119 -6578 647 -6572
rect -1119 -6612 -1107 -6578
rect -739 -6612 -649 -6578
rect -281 -6612 -191 -6578
rect 177 -6612 267 -6578
rect 635 -6612 647 -6578
rect -1119 -6618 647 -6612
rect -1436 -6800 -1276 -6780
rect 804 -6780 884 -6552
rect 944 -6780 964 -5560
rect 804 -6800 964 -6780
rect -3420 -6880 -3180 -6860
rect -4301 -7084 -4261 -6884
<< via1 >>
rect -2858 -2903 -2849 -927
rect -2849 -2903 -2815 -927
rect -2815 -2903 -2806 -927
rect -2740 -2903 -2731 -927
rect -2731 -2903 -2697 -927
rect -2697 -2903 -2688 -927
rect -2622 -2903 -2613 -927
rect -2613 -2903 -2579 -927
rect -2579 -2903 -2570 -927
rect -2504 -2903 -2495 -927
rect -2495 -2903 -2461 -927
rect -2461 -2903 -2452 -927
rect -2386 -2903 -2377 -927
rect -2377 -2903 -2343 -927
rect -2343 -2903 -2334 -927
rect -2268 -2903 -2259 -927
rect -2259 -2903 -2225 -927
rect -2225 -2903 -2216 -927
rect -2150 -2903 -2141 -927
rect -2141 -2903 -2107 -927
rect -2107 -2903 -2098 -927
rect -2032 -2903 -2023 -927
rect -2023 -2903 -1989 -927
rect -1989 -2903 -1980 -927
rect -1914 -2903 -1905 -927
rect -1905 -2903 -1871 -927
rect -1871 -2903 -1862 -927
rect -1796 -2903 -1787 -927
rect -1787 -2903 -1753 -927
rect -1753 -2903 -1744 -927
rect -1678 -2903 -1669 -927
rect -1669 -2903 -1635 -927
rect -1635 -2903 -1626 -927
rect -1560 -2903 -1551 -927
rect -1551 -2903 -1517 -927
rect -1517 -2903 -1508 -927
rect -1442 -2903 -1433 -927
rect -1433 -2903 -1399 -927
rect -1399 -2903 -1390 -927
rect -1324 -2903 -1315 -927
rect -1315 -2903 -1281 -927
rect -1281 -2903 -1272 -927
rect -1206 -2903 -1197 -927
rect -1197 -2903 -1163 -927
rect -1163 -2903 -1154 -927
rect -1088 -2903 -1079 -927
rect -1079 -2903 -1045 -927
rect -1045 -2903 -1036 -927
rect -970 -2903 -961 -927
rect -961 -2903 -927 -927
rect -927 -2903 -918 -927
rect -852 -2903 -843 -927
rect -843 -2903 -809 -927
rect -809 -2903 -800 -927
rect -734 -2903 -725 -927
rect -725 -2903 -691 -927
rect -691 -2903 -682 -927
rect -616 -2903 -607 -927
rect -607 -2903 -573 -927
rect -573 -2903 -564 -927
rect -498 -2903 -489 -927
rect -489 -2903 -455 -927
rect -455 -2903 -446 -927
rect -380 -2903 -371 -927
rect -371 -2903 -337 -927
rect -337 -2903 -328 -927
rect -262 -2903 -253 -927
rect -253 -2903 -219 -927
rect -219 -2903 -210 -927
rect -144 -2903 -135 -927
rect -135 -2903 -101 -927
rect -101 -2903 -92 -927
rect -26 -2903 -17 -927
rect -17 -2903 17 -927
rect 17 -2903 26 -927
rect 92 -2903 101 -927
rect 101 -2903 135 -927
rect 135 -2903 144 -927
rect 210 -2903 219 -927
rect 219 -2903 253 -927
rect 253 -2903 262 -927
rect 328 -2903 337 -927
rect 337 -2903 371 -927
rect 371 -2903 380 -927
rect 446 -2903 455 -927
rect 455 -2903 489 -927
rect 489 -2903 498 -927
rect 564 -2903 573 -927
rect 573 -2903 607 -927
rect 607 -2903 616 -927
rect 682 -2903 691 -927
rect 691 -2903 725 -927
rect 725 -2903 734 -927
rect 800 -2903 809 -927
rect 809 -2903 843 -927
rect 843 -2903 852 -927
rect 918 -2903 927 -927
rect 927 -2903 961 -927
rect 961 -2903 970 -927
rect 1036 -2903 1045 -927
rect 1045 -2903 1079 -927
rect 1079 -2903 1088 -927
rect 1154 -2903 1163 -927
rect 1163 -2903 1197 -927
rect 1197 -2903 1206 -927
rect 1272 -2903 1281 -927
rect 1281 -2903 1315 -927
rect 1315 -2903 1324 -927
rect 1390 -2903 1399 -927
rect 1399 -2903 1433 -927
rect 1433 -2903 1442 -927
rect 1508 -2903 1517 -927
rect 1517 -2903 1551 -927
rect 1551 -2903 1560 -927
rect 1626 -2903 1635 -927
rect 1635 -2903 1669 -927
rect 1669 -2903 1678 -927
rect 1744 -2903 1753 -927
rect 1753 -2903 1787 -927
rect 1787 -2903 1796 -927
rect 1862 -2903 1871 -927
rect 1871 -2903 1905 -927
rect 1905 -2903 1914 -927
rect 1980 -2903 1989 -927
rect 1989 -2903 2023 -927
rect 2023 -2903 2032 -927
rect 2098 -2903 2107 -927
rect 2107 -2903 2141 -927
rect 2141 -2903 2150 -927
rect 2216 -2903 2225 -927
rect 2225 -2903 2259 -927
rect 2259 -2903 2268 -927
rect 2334 -2903 2343 -927
rect 2343 -2903 2377 -927
rect 2377 -2903 2386 -927
rect -2505 -3294 -2453 -3242
rect -2269 -3294 -2217 -3242
rect -2033 -3294 -1981 -3242
rect 1508 -3294 1560 -3242
rect 1744 -3294 1796 -3242
rect 1980 -3294 2032 -3242
rect -2859 -5412 -2850 -3436
rect -2850 -5412 -2816 -3436
rect -2816 -5412 -2807 -3436
rect -2741 -5412 -2732 -3436
rect -2732 -5412 -2698 -3436
rect -2698 -5412 -2689 -3436
rect -2623 -5412 -2614 -3436
rect -2614 -5412 -2580 -3436
rect -2580 -5412 -2571 -3436
rect -2505 -5412 -2496 -3436
rect -2496 -5412 -2462 -3436
rect -2462 -5412 -2453 -3436
rect -2387 -5412 -2378 -3436
rect -2378 -5412 -2344 -3436
rect -2344 -5412 -2335 -3436
rect -2269 -5412 -2260 -3436
rect -2260 -5412 -2226 -3436
rect -2226 -5412 -2217 -3436
rect -2151 -5412 -2142 -3436
rect -2142 -5412 -2108 -3436
rect -2108 -5412 -2099 -3436
rect -2033 -5412 -2024 -3436
rect -2024 -5412 -1990 -3436
rect -1990 -5412 -1981 -3436
rect -1915 -5412 -1906 -3436
rect -1906 -5412 -1872 -3436
rect -1872 -5412 -1863 -3436
rect -1797 -5412 -1788 -3436
rect -1788 -5412 -1754 -3436
rect -1754 -5412 -1745 -3436
rect -1679 -5412 -1670 -3436
rect -1670 -5412 -1636 -3436
rect -1636 -5412 -1627 -3436
rect -1223 -3612 -1169 -3600
rect -1223 -4088 -1213 -3612
rect -1213 -4088 -1179 -3612
rect -1179 -4088 -1169 -3612
rect -1223 -4100 -1169 -4088
rect -1127 -3612 -1073 -3600
rect -1127 -4088 -1117 -3612
rect -1117 -4088 -1083 -3612
rect -1083 -4088 -1073 -3612
rect -1127 -4100 -1073 -4088
rect -1031 -3612 -977 -3600
rect -1031 -4088 -1021 -3612
rect -1021 -4088 -987 -3612
rect -987 -4088 -977 -3612
rect -1031 -4100 -977 -4088
rect -935 -3612 -881 -3600
rect -935 -4088 -925 -3612
rect -925 -4088 -891 -3612
rect -891 -4088 -881 -3612
rect -935 -4100 -881 -4088
rect -839 -3612 -785 -3600
rect -839 -4088 -829 -3612
rect -829 -4088 -795 -3612
rect -795 -4088 -785 -3612
rect -839 -4100 -785 -4088
rect -743 -3612 -689 -3600
rect -743 -4088 -733 -3612
rect -733 -4088 -699 -3612
rect -699 -4088 -689 -3612
rect -743 -4100 -689 -4088
rect -647 -3612 -593 -3600
rect -647 -4088 -637 -3612
rect -637 -4088 -603 -3612
rect -603 -4088 -593 -3612
rect -647 -4100 -593 -4088
rect -551 -3612 -497 -3600
rect -551 -4088 -541 -3612
rect -541 -4088 -507 -3612
rect -507 -4088 -497 -3612
rect -551 -4100 -497 -4088
rect -455 -3612 -401 -3600
rect -455 -4088 -445 -3612
rect -445 -4088 -411 -3612
rect -411 -4088 -401 -3612
rect -455 -4100 -401 -4088
rect -359 -3612 -305 -3600
rect -359 -4088 -349 -3612
rect -349 -4088 -315 -3612
rect -315 -4088 -305 -3612
rect -359 -4100 -305 -4088
rect -263 -3612 -209 -3600
rect -263 -4088 -253 -3612
rect -253 -4088 -219 -3612
rect -219 -4088 -209 -3612
rect -263 -4100 -209 -4088
rect -167 -3612 -113 -3600
rect -167 -4088 -157 -3612
rect -157 -4088 -123 -3612
rect -123 -4088 -113 -3612
rect -167 -4100 -113 -4088
rect -71 -3612 -17 -3600
rect -71 -4088 -61 -3612
rect -61 -4088 -27 -3612
rect -27 -4088 -17 -3612
rect -71 -4100 -17 -4088
rect 25 -3612 79 -3600
rect 25 -4088 35 -3612
rect 35 -4088 69 -3612
rect 69 -4088 79 -3612
rect 25 -4100 79 -4088
rect 121 -3612 175 -3600
rect 121 -4088 131 -3612
rect 131 -4088 165 -3612
rect 165 -4088 175 -3612
rect 121 -4100 175 -4088
rect 217 -3612 271 -3600
rect 217 -4088 227 -3612
rect 227 -4088 261 -3612
rect 261 -4088 271 -3612
rect 217 -4100 271 -4088
rect 313 -3612 367 -3600
rect 313 -4088 323 -3612
rect 323 -4088 357 -3612
rect 357 -4088 367 -3612
rect 313 -4100 367 -4088
rect 409 -3612 463 -3600
rect 409 -4088 419 -3612
rect 419 -4088 453 -3612
rect 453 -4088 463 -3612
rect 409 -4100 463 -4088
rect 505 -3612 559 -3600
rect 505 -4088 515 -3612
rect 515 -4088 549 -3612
rect 549 -4088 559 -3612
rect 505 -4100 559 -4088
rect 601 -3612 655 -3600
rect 601 -4088 611 -3612
rect 611 -4088 645 -3612
rect 645 -4088 655 -3612
rect 601 -4100 655 -4088
rect 697 -3612 751 -3600
rect 697 -4088 707 -3612
rect 707 -4088 741 -3612
rect 741 -4088 751 -3612
rect 697 -4100 751 -4088
rect -941 -4150 -875 -4144
rect -941 -4184 -925 -4150
rect -925 -4184 -891 -4150
rect -891 -4184 -875 -4150
rect -941 -4200 -875 -4184
rect -749 -4150 -683 -4144
rect -749 -4184 -733 -4150
rect -733 -4184 -699 -4150
rect -699 -4184 -683 -4150
rect -749 -4200 -683 -4184
rect -557 -4150 -491 -4144
rect -557 -4184 -541 -4150
rect -541 -4184 -507 -4150
rect -507 -4184 -491 -4150
rect -557 -4200 -491 -4184
rect -365 -4150 -299 -4144
rect -365 -4184 -349 -4150
rect -349 -4184 -315 -4150
rect -315 -4184 -299 -4150
rect -365 -4200 -299 -4184
rect -173 -4150 -107 -4144
rect -173 -4184 -157 -4150
rect -157 -4184 -123 -4150
rect -123 -4184 -107 -4150
rect -173 -4200 -107 -4184
rect 19 -4150 85 -4144
rect 19 -4184 35 -4150
rect 35 -4184 69 -4150
rect 69 -4184 85 -4150
rect 19 -4200 85 -4184
rect 211 -4150 277 -4144
rect 211 -4184 227 -4150
rect 227 -4184 261 -4150
rect 261 -4184 277 -4150
rect 211 -4200 277 -4184
rect 403 -4150 469 -4144
rect 403 -4184 419 -4150
rect 419 -4184 453 -4150
rect 453 -4184 469 -4150
rect 403 -4200 469 -4184
rect -1190 -4500 -1130 -4440
rect -4134 -5994 -3665 -5985
rect -4134 -6028 -3665 -5994
rect -4134 -6037 -3665 -6028
rect -4210 -6608 -3781 -6600
rect -4210 -6661 -3781 -6608
rect -4210 -6670 -3781 -6661
rect -3400 -6860 -3340 -5940
rect -3340 -6860 -3200 -5940
rect -1416 -6780 -1356 -5560
rect -1178 -6528 -1169 -4552
rect -1169 -6528 -1135 -4552
rect -1135 -6528 -1126 -4552
rect -720 -6528 -711 -4552
rect -711 -6528 -677 -4552
rect -677 -6528 -668 -4552
rect -262 -6528 -253 -4552
rect -253 -6528 -219 -4552
rect -219 -6528 -210 -4552
rect 196 -6528 205 -4552
rect 205 -6528 239 -4552
rect 239 -6528 248 -4552
rect 654 -6528 663 -4552
rect 663 -6528 697 -4552
rect 697 -6528 706 -4552
rect 1154 -5412 1163 -3436
rect 1163 -5412 1197 -3436
rect 1197 -5412 1206 -3436
rect 1272 -5412 1281 -3436
rect 1281 -5412 1315 -3436
rect 1315 -5412 1324 -3436
rect 1390 -5412 1399 -3436
rect 1399 -5412 1433 -3436
rect 1433 -5412 1442 -3436
rect 1508 -5412 1517 -3436
rect 1517 -5412 1551 -3436
rect 1551 -5412 1560 -3436
rect 1626 -5412 1635 -3436
rect 1635 -5412 1669 -3436
rect 1669 -5412 1678 -3436
rect 1744 -5412 1753 -3436
rect 1753 -5412 1787 -3436
rect 1787 -5412 1796 -3436
rect 1862 -5412 1871 -3436
rect 1871 -5412 1905 -3436
rect 1905 -5412 1914 -3436
rect 1980 -5412 1989 -3436
rect 1989 -5412 2023 -3436
rect 2023 -5412 2032 -3436
rect 2098 -5412 2107 -3436
rect 2107 -5412 2141 -3436
rect 2141 -5412 2150 -3436
rect 2216 -5412 2225 -3436
rect 2225 -5412 2259 -3436
rect 2259 -5412 2268 -3436
rect 2334 -5412 2343 -3436
rect 2343 -5412 2377 -3436
rect 2377 -5412 2386 -3436
rect 2720 -3780 2800 -3420
rect 2960 -3780 3040 -3420
rect 884 -6780 944 -5560
<< metal2 >>
rect -2600 0 2000 100
rect -2600 -400 -2500 0
rect -2836 -500 -2500 -400
rect 1900 -400 2000 0
rect 1900 -500 2364 -400
rect -2836 -600 2364 -500
rect -2836 -664 -2736 -600
rect -2436 -664 -2336 -600
rect -2036 -664 -1936 -600
rect -1636 -664 -1536 -600
rect -1236 -664 -1136 -600
rect -836 -664 -736 -600
rect -436 -664 -336 -600
rect -136 -664 -36 -600
rect 264 -664 364 -600
rect 664 -664 764 -600
rect 1064 -664 1164 -600
rect 1464 -664 1564 -600
rect 1864 -664 1964 -600
rect 2264 -664 2364 -600
rect -2858 -766 2386 -664
rect -2858 -927 -2806 -766
rect -2858 -2915 -2806 -2903
rect -2740 -927 -2688 -766
rect -2740 -2915 -2688 -2903
rect -2622 -927 -2570 -766
rect -2622 -2915 -2570 -2903
rect -2504 -927 -2452 -915
rect -2504 -3064 -2452 -2903
rect -2386 -927 -2334 -766
rect -2386 -2915 -2334 -2903
rect -2268 -927 -2216 -915
rect -2268 -3064 -2216 -2903
rect -2150 -927 -2098 -766
rect -2150 -2915 -2098 -2903
rect -2032 -927 -1980 -915
rect -2032 -3064 -1980 -2903
rect -1914 -927 -1862 -766
rect -1914 -2915 -1862 -2903
rect -1796 -927 -1744 -915
rect -1796 -3064 -1744 -2903
rect -1678 -927 -1626 -766
rect -1678 -2915 -1626 -2903
rect -1560 -927 -1508 -915
rect -1560 -3064 -1508 -2903
rect -1442 -927 -1390 -766
rect -1442 -2915 -1390 -2903
rect -1324 -927 -1272 -915
rect -1324 -3064 -1272 -2903
rect -1206 -927 -1154 -766
rect -1206 -2915 -1154 -2903
rect -1088 -927 -1036 -915
rect -1088 -3064 -1036 -2903
rect -970 -927 -918 -766
rect -970 -2915 -918 -2903
rect -852 -927 -800 -915
rect -852 -3064 -800 -2903
rect -734 -927 -682 -766
rect -734 -2915 -682 -2903
rect -616 -927 -564 -915
rect -2623 -3166 -800 -3064
rect -616 -2956 -564 -2903
rect -498 -927 -446 -766
rect -498 -2915 -446 -2903
rect -380 -927 -328 -915
rect -380 -2956 -328 -2903
rect -262 -927 -210 -766
rect -262 -2916 -210 -2903
rect -144 -927 -92 -915
rect -616 -3002 -328 -2956
rect -144 -2956 -92 -2903
rect -26 -927 26 -766
rect -26 -2915 26 -2903
rect 92 -927 144 -915
rect 92 -2956 144 -2903
rect 210 -927 262 -766
rect 328 -927 380 -915
rect 210 -2915 262 -2903
rect 327 -2903 328 -2835
rect 327 -2915 380 -2903
rect 446 -927 498 -766
rect 564 -927 616 -915
rect 446 -2915 498 -2903
rect 563 -2903 564 -2835
rect 563 -2915 616 -2903
rect 682 -927 734 -766
rect 800 -927 852 -915
rect 682 -2915 734 -2903
rect 799 -2903 800 -2835
rect 799 -2915 852 -2903
rect 918 -927 970 -766
rect 1036 -927 1088 -915
rect 918 -2915 970 -2903
rect 1035 -2903 1036 -2835
rect 1035 -2915 1088 -2903
rect 1154 -927 1206 -766
rect 1272 -927 1324 -915
rect 1154 -2915 1206 -2903
rect 1271 -2903 1272 -2835
rect 1271 -2915 1324 -2903
rect 1390 -927 1442 -766
rect 1508 -927 1560 -915
rect 1390 -2915 1442 -2903
rect 1507 -2903 1508 -2835
rect 1507 -2915 1560 -2903
rect 1626 -927 1678 -766
rect 1744 -927 1796 -915
rect 1626 -2915 1678 -2903
rect 1743 -2903 1744 -2835
rect 1743 -2915 1796 -2903
rect 1862 -927 1914 -766
rect 1980 -927 2032 -915
rect 1862 -2915 1914 -2903
rect 1979 -2903 1980 -2835
rect 1979 -2915 2032 -2903
rect 2098 -927 2150 -766
rect 2216 -927 2268 -766
rect 2098 -2915 2150 -2903
rect 2215 -2903 2216 -2835
rect 2215 -2915 2268 -2903
rect 2334 -927 2386 -766
rect 2334 -2915 2386 -2903
rect -144 -3002 144 -2956
rect -616 -3095 -564 -3002
rect 92 -3095 144 -3002
rect -2623 -3231 -2571 -3166
rect -2387 -3231 -2335 -3166
rect -2151 -3231 -2099 -3166
rect -1915 -3231 -1863 -3166
rect -2623 -3240 -1863 -3231
rect -2623 -3296 -2507 -3240
rect -2451 -3296 -2271 -3240
rect -2215 -3296 -2035 -3240
rect -1979 -3296 -1863 -3240
rect -2623 -3305 -1863 -3296
rect -2859 -3436 -2807 -3424
rect -2859 -5564 -2807 -5412
rect -2741 -3436 -2689 -3424
rect -2741 -5564 -2689 -5412
rect -2623 -3436 -2571 -3305
rect -2623 -5424 -2571 -5412
rect -2505 -3436 -2453 -3424
rect -2505 -5564 -2453 -5412
rect -2387 -3436 -2335 -3305
rect -2387 -5424 -2335 -5412
rect -2269 -3436 -2217 -3424
rect -2269 -5564 -2217 -5412
rect -2151 -3436 -2099 -3305
rect -2151 -5424 -2099 -5412
rect -2033 -3436 -1981 -3424
rect -2033 -5564 -1981 -5412
rect -1915 -3436 -1863 -3305
rect -616 -3390 -512 -3095
rect 40 -3390 144 -3095
rect 327 -3064 379 -2915
rect 563 -3064 615 -2915
rect 799 -3064 851 -2915
rect 1035 -3064 1087 -2915
rect 1271 -3064 1323 -2915
rect 1507 -3064 1559 -2915
rect 1743 -3064 1795 -2915
rect 1979 -3064 2031 -2915
rect 2400 -3000 2540 -2980
rect 327 -3080 2150 -3064
rect 2400 -3080 2420 -3000
rect 327 -3140 2420 -3080
rect 2520 -3140 2540 -3000
rect 327 -3160 2540 -3140
rect 327 -3166 2150 -3160
rect -1915 -5424 -1863 -5412
rect -1797 -3436 -1745 -3424
rect -1797 -5540 -1745 -5412
rect -1679 -3436 -1627 -3424
rect -941 -3530 -299 -3390
rect -941 -3600 -875 -3530
rect -749 -3600 -683 -3530
rect -557 -3600 -491 -3530
rect -365 -3600 -299 -3530
rect -173 -3530 469 -3390
rect -173 -3600 -107 -3530
rect 19 -3600 85 -3530
rect 211 -3600 277 -3530
rect 403 -3600 469 -3530
rect 1154 -3436 1206 -3424
rect -1229 -4100 -1223 -3600
rect -1169 -4100 -1163 -3600
rect -1133 -4100 -1127 -3600
rect -1073 -4100 -1067 -3600
rect -1037 -4100 -1031 -3600
rect -977 -4100 -971 -3600
rect -941 -4100 -935 -3600
rect -881 -4100 -875 -3600
rect -845 -4100 -839 -3600
rect -785 -4100 -779 -3600
rect -749 -4100 -743 -3600
rect -689 -4100 -683 -3600
rect -653 -4100 -647 -3600
rect -593 -4100 -587 -3600
rect -557 -4100 -551 -3600
rect -497 -4100 -491 -3600
rect -461 -4100 -455 -3600
rect -401 -4100 -395 -3600
rect -365 -4100 -359 -3600
rect -305 -4100 -299 -3600
rect -269 -4100 -263 -3600
rect -209 -4100 -203 -3600
rect -173 -4100 -167 -3600
rect -113 -4100 -107 -3600
rect -77 -4100 -71 -3600
rect -17 -4100 -11 -3600
rect 19 -4100 25 -3600
rect 79 -4100 85 -3600
rect 115 -4100 121 -3600
rect 175 -4100 181 -3600
rect 211 -4100 217 -3600
rect 271 -4100 277 -3600
rect 307 -4100 313 -3600
rect 367 -4100 373 -3600
rect 403 -4100 409 -3600
rect 463 -4100 469 -3600
rect 499 -4100 505 -3600
rect 559 -4100 565 -3600
rect 595 -4100 601 -3600
rect 655 -4100 661 -3600
rect 691 -4100 697 -3600
rect 751 -4100 757 -3600
rect -1031 -4260 -977 -4100
rect -941 -4144 -875 -4138
rect -941 -4220 -875 -4206
rect -839 -4260 -785 -4100
rect -749 -4144 -683 -4138
rect -749 -4220 -683 -4206
rect -647 -4260 -593 -4100
rect -557 -4144 -491 -4138
rect -557 -4220 -491 -4206
rect -455 -4260 -401 -4100
rect -365 -4144 -299 -4138
rect -365 -4220 -299 -4206
rect -263 -4260 -209 -4100
rect -173 -4144 -107 -4138
rect -173 -4220 -107 -4206
rect -71 -4260 -17 -4100
rect 19 -4144 85 -4138
rect 19 -4220 85 -4206
rect 121 -4260 175 -4100
rect 211 -4144 277 -4138
rect 211 -4220 277 -4206
rect 313 -4260 367 -4100
rect 403 -4144 469 -4138
rect 403 -4220 469 -4206
rect 505 -4260 559 -4100
rect -1031 -4330 559 -4260
rect -1031 -4416 -977 -4330
rect -839 -4416 -785 -4330
rect -647 -4416 -593 -4330
rect -455 -4416 -401 -4330
rect -263 -4416 -209 -4330
rect -71 -4416 -17 -4330
rect 121 -4416 175 -4330
rect 313 -4416 367 -4330
rect 505 -4416 559 -4330
rect -1400 -4440 -1120 -4430
rect -1400 -4500 -1390 -4440
rect -1230 -4500 -1190 -4440
rect -1130 -4500 -1120 -4440
rect -1400 -4510 -1120 -4500
rect -1031 -4508 559 -4416
rect -1679 -5540 -1627 -5412
rect -1178 -4552 -1126 -4540
rect -1797 -5560 -1336 -5540
rect -1797 -5564 -1416 -5560
rect -2859 -5634 -1416 -5564
rect -3900 -5768 -3650 -5749
rect -3900 -5985 -3880 -5768
rect -3670 -5985 -3650 -5768
rect -2836 -5800 -2736 -5634
rect -2636 -5800 -2536 -5634
rect -2436 -5800 -2336 -5634
rect -2236 -5800 -2136 -5634
rect -2036 -5800 -1936 -5634
rect -1836 -5640 -1416 -5634
rect -1836 -5800 -1736 -5640
rect -1636 -5800 -1536 -5640
rect -1436 -5800 -1416 -5640
rect -4151 -6037 -4134 -5985
rect -3665 -6037 -3650 -5985
rect -3420 -5940 -3180 -5920
rect -4233 -6670 -4210 -6600
rect -3781 -6670 -3762 -6600
rect -4200 -6848 -4000 -6670
rect -4200 -7084 -4120 -6848
rect -3420 -6860 -3400 -5940
rect -3200 -6700 -3180 -5940
rect -2840 -6000 -1416 -5800
rect -2840 -6200 -2340 -6000
rect -1736 -6200 -1536 -6000
rect -2840 -6300 -1536 -6200
rect -1436 -6300 -1416 -6000
rect -2840 -6400 -1416 -6300
rect -2840 -6500 -1536 -6400
rect -2840 -6700 -2340 -6500
rect -1736 -6700 -1536 -6500
rect -1436 -6700 -1416 -6400
rect -3200 -6780 -1416 -6700
rect -1356 -6700 -1336 -5560
rect -1178 -6680 -1126 -6528
rect -720 -4552 -668 -4508
rect -720 -6540 -668 -6528
rect -262 -4552 -210 -4540
rect -262 -6680 -210 -6528
rect 196 -4552 248 -4508
rect 196 -6540 248 -6528
rect 654 -4552 706 -4540
rect 1154 -5540 1206 -5412
rect 1272 -3436 1324 -3424
rect 1272 -5540 1324 -5412
rect 1390 -3436 1442 -3166
rect 1503 -3240 1564 -3231
rect 1503 -3296 1506 -3240
rect 1562 -3296 1564 -3240
rect 1503 -3305 1564 -3296
rect 1390 -5424 1442 -5412
rect 1508 -3436 1560 -3424
rect 654 -6680 706 -6528
rect -1178 -6700 706 -6680
rect 864 -5560 1324 -5540
rect 864 -6700 884 -5560
rect -1356 -6780 884 -6700
rect 944 -5564 1324 -5560
rect 1508 -5564 1560 -5412
rect 1626 -3436 1678 -3166
rect 1739 -3240 1800 -3231
rect 1739 -3296 1742 -3240
rect 1798 -3296 1800 -3240
rect 1739 -3305 1800 -3296
rect 1626 -5424 1678 -5412
rect 1744 -3436 1796 -3424
rect 1744 -5564 1796 -5412
rect 1862 -3436 1914 -3166
rect 1975 -3240 2036 -3231
rect 1975 -3296 1978 -3240
rect 2034 -3296 2036 -3240
rect 1975 -3305 2036 -3296
rect 1862 -5424 1914 -5412
rect 1980 -3436 2032 -3424
rect 1980 -5564 2032 -5412
rect 2098 -3436 2150 -3166
rect 2700 -3420 2820 -3400
rect 2098 -5424 2150 -5412
rect 2216 -3436 2268 -3424
rect 2216 -5564 2268 -5412
rect 2334 -3436 2386 -3424
rect 2700 -3780 2720 -3420
rect 2800 -3780 2820 -3420
rect 2700 -3800 2820 -3780
rect 2940 -3420 3060 -3400
rect 2940 -3780 2960 -3420
rect 3040 -3780 3060 -3420
rect 2940 -3800 3060 -3780
rect 2334 -5564 2386 -5412
rect 944 -5634 2386 -5564
rect 944 -5640 1364 -5634
rect 944 -5900 964 -5640
rect 1064 -5800 1164 -5640
rect 1264 -5800 1364 -5640
rect 1464 -5800 1564 -5634
rect 1664 -5800 1764 -5634
rect 1864 -5800 1964 -5634
rect 2064 -5800 2164 -5634
rect 2264 -5800 2364 -5634
rect 1064 -5900 2364 -5800
rect 944 -6000 2364 -5900
rect 944 -6300 964 -6000
rect 1064 -6300 1264 -6000
rect 944 -6400 1264 -6300
rect 944 -6700 964 -6400
rect 1064 -6700 1264 -6400
rect 944 -6780 1264 -6700
rect -3200 -6860 1264 -6780
rect -3420 -6880 1264 -6860
rect -3320 -7000 1264 -6880
rect 1600 -7000 2000 -6000
rect -3000 -7100 -1200 -7000
rect -3000 -7700 -2900 -7100
rect -1300 -7700 -1200 -7100
rect -3000 -7800 -1200 -7700
rect 600 -7100 2000 -7000
rect 600 -7700 700 -7100
rect 1900 -7700 2000 -7100
rect 600 -7800 2000 -7700
<< via2 >>
rect -2500 -500 1900 0
rect -2507 -3242 -2451 -3240
rect -2507 -3294 -2505 -3242
rect -2505 -3294 -2453 -3242
rect -2453 -3294 -2451 -3242
rect -2507 -3296 -2451 -3294
rect -2271 -3242 -2215 -3240
rect -2271 -3294 -2269 -3242
rect -2269 -3294 -2217 -3242
rect -2217 -3294 -2215 -3242
rect -2271 -3296 -2215 -3294
rect -2035 -3242 -1979 -3240
rect -2035 -3294 -2033 -3242
rect -2033 -3294 -1981 -3242
rect -1981 -3294 -1979 -3242
rect -2035 -3296 -1979 -3294
rect 2420 -3140 2520 -3000
rect -941 -4200 -875 -4150
rect -941 -4206 -875 -4200
rect -749 -4200 -683 -4150
rect -749 -4206 -683 -4200
rect -557 -4200 -491 -4150
rect -557 -4206 -491 -4200
rect -365 -4200 -299 -4150
rect -365 -4206 -299 -4200
rect -173 -4200 -107 -4150
rect -173 -4206 -107 -4200
rect 19 -4200 85 -4150
rect 19 -4206 85 -4200
rect 211 -4200 277 -4150
rect 211 -4206 277 -4200
rect 403 -4200 469 -4150
rect 403 -4206 469 -4200
rect -1390 -4500 -1230 -4440
rect -3880 -5985 -3670 -5768
rect -3880 -5988 -3670 -5985
rect -3400 -6860 -3200 -5940
rect 1506 -3242 1562 -3240
rect 1506 -3294 1508 -3242
rect 1508 -3294 1560 -3242
rect 1560 -3294 1562 -3242
rect 1506 -3296 1562 -3294
rect 1742 -3242 1798 -3240
rect 1742 -3294 1744 -3242
rect 1744 -3294 1796 -3242
rect 1796 -3294 1798 -3242
rect 1742 -3296 1798 -3294
rect 1978 -3242 2034 -3240
rect 1978 -3294 1980 -3242
rect 1980 -3294 2032 -3242
rect 2032 -3294 2034 -3242
rect 1978 -3296 2034 -3294
rect 2720 -3780 2800 -3420
rect 2960 -3780 3040 -3420
rect -2900 -7700 -1300 -7100
rect 700 -7700 1900 -7100
<< metal3 >>
rect -2600 0 2000 100
rect -7600 -7100 -4800 -200
rect -4400 -5600 -3100 -148
rect -2600 -500 -2500 0
rect 1900 -500 2000 0
rect -2600 -600 2000 -500
rect 2400 -3000 2540 -2980
rect 2400 -3140 2420 -3000
rect 2520 -3140 2540 -3000
rect 2700 -3100 4300 700
rect 2400 -3160 2540 -3140
rect 2600 -3231 2820 -3220
rect -2512 -3240 2820 -3231
rect -2512 -3296 -2507 -3240
rect -2451 -3296 -2271 -3240
rect -2215 -3296 -2035 -3240
rect -1979 -3296 1506 -3240
rect 1562 -3296 1742 -3240
rect 1798 -3296 1978 -3240
rect 2034 -3296 2820 -3240
rect -2512 -3305 2820 -3296
rect -1976 -3336 1503 -3305
rect 2600 -3320 2820 -3305
rect 2700 -3420 2820 -3320
rect 2700 -3780 2720 -3420
rect 2800 -3780 2820 -3420
rect 2700 -3800 2820 -3780
rect 2940 -3420 3060 -3400
rect 2940 -3780 2960 -3420
rect 3040 -3620 3060 -3420
rect 3380 -3520 4300 -3100
rect 3380 -3620 3400 -3520
rect 3040 -3740 3400 -3620
rect 3040 -3780 3060 -3740
rect 2940 -3800 3060 -3780
rect 3380 -3840 3400 -3740
rect 4280 -3840 4300 -3520
rect 3380 -3860 4300 -3840
rect -947 -4150 -293 -4138
rect -947 -4206 -941 -4150
rect -875 -4206 -749 -4150
rect -683 -4206 -557 -4150
rect -491 -4206 -365 -4150
rect -299 -4206 -293 -4150
rect -947 -4220 -293 -4206
rect -179 -4150 475 -4138
rect -179 -4206 -173 -4150
rect -107 -4206 19 -4150
rect 85 -4206 211 -4150
rect 277 -4206 403 -4150
rect 469 -4206 475 -4150
rect -179 -4220 475 -4206
rect -1400 -4440 -1220 -4430
rect -1400 -4500 -1390 -4440
rect -1230 -4500 -1220 -4440
rect -4400 -5700 -2800 -5600
rect -1400 -5700 -1220 -4500
rect -4400 -5768 -1220 -5700
rect -4400 -5988 -3880 -5768
rect -3670 -5800 -1220 -5768
rect -3670 -5988 -3500 -5800
rect -4400 -6248 -3500 -5988
rect -4400 -6648 -4300 -6248
rect -3600 -6648 -3500 -6248
rect -4400 -6748 -3500 -6648
rect -3420 -5940 -3100 -5920
rect -3420 -6860 -3400 -5940
rect -3120 -6860 -3100 -5940
rect -3000 -6000 -1220 -5800
rect -3420 -6880 -3100 -6860
rect -7600 -7700 -7500 -7100
rect -4900 -7300 -4800 -7100
rect -3000 -7100 -1200 -7000
rect -4900 -7600 -4600 -7300
rect -4900 -7700 -4800 -7600
rect -7600 -7800 -4800 -7700
rect -3000 -7700 -2900 -7100
rect -1300 -7700 -1200 -7100
rect -3000 -7800 -1200 -7700
rect 600 -7100 2000 -7000
rect 600 -7700 700 -7100
rect 1900 -7700 2000 -7100
rect 600 -7800 2000 -7700
<< via3 >>
rect -2500 -500 1900 0
rect 2420 -3140 2520 -3000
rect 3400 -3840 4280 -3520
rect -4300 -6648 -3600 -6248
rect -3320 -6860 -3200 -5940
rect -3200 -6860 -3120 -5940
rect -7500 -7700 -4900 -7100
rect -2900 -7700 -1300 -7100
rect 700 -7700 1900 -7100
<< mimcap >>
rect 2800 560 4200 600
rect -4300 -288 -3200 -248
rect -7500 -340 -4900 -300
rect -7500 -6460 -7460 -340
rect -4940 -6460 -4900 -340
rect -4300 -5608 -4260 -288
rect -3240 -5608 -3200 -288
rect 2800 -2960 2840 560
rect 4160 -2960 4200 560
rect 2800 -3000 4200 -2960
rect -4300 -5648 -3200 -5608
rect -7500 -6500 -4900 -6460
<< mimcapcontact >>
rect -7460 -6460 -4940 -340
rect -4260 -5608 -3240 -288
rect 2840 -2960 4160 560
<< metal4 >>
rect -7400 100 2000 600
rect -7400 -200 -5000 100
rect -2600 0 2000 100
rect -7600 -340 -4800 -200
rect -7600 -6460 -7460 -340
rect -4940 -6460 -4800 -340
rect -4400 -288 -3100 -148
rect -4400 -5608 -4260 -288
rect -3240 -5608 -3100 -288
rect -2600 -500 -2500 0
rect 1900 -500 2000 0
rect -2600 -600 2000 -500
rect 2700 560 4300 700
rect 2700 -2960 2840 560
rect 4160 -2960 4300 560
rect 2700 -2980 4300 -2960
rect 2400 -3000 4300 -2980
rect 2400 -3140 2420 -3000
rect 2520 -3100 4300 -3000
rect 2520 -3140 2540 -3100
rect 2400 -3160 2540 -3140
rect 3380 -3520 4300 -3500
rect 3380 -3840 3400 -3520
rect 4280 -3840 4300 -3520
rect 3380 -3860 4300 -3840
rect -4400 -5748 -3100 -5608
rect -3340 -5940 -3100 -5748
rect -7600 -6600 -4800 -6460
rect -4400 -6248 -3500 -6148
rect -4400 -6648 -4300 -6248
rect -3600 -6648 -3500 -6248
rect -4400 -6748 -3500 -6648
rect -3340 -6860 -3320 -5940
rect -3120 -6860 -3100 -5940
rect -3340 -6880 -3100 -6860
rect -7600 -7100 -4800 -7000
rect -7600 -7700 -7500 -7100
rect -4900 -7300 -4800 -7100
rect -3000 -7100 2000 -7000
rect -3000 -7300 -2900 -7100
rect -4900 -7700 -2900 -7300
rect -1300 -7700 700 -7100
rect 1900 -7700 2000 -7100
rect -7600 -7800 2000 -7700
<< via4 >>
rect 3420 -3820 4260 -3540
rect -4300 -6648 -3600 -6248
rect -7500 -7700 -4900 -7100
<< mimcap2 >>
rect 2800 560 4200 600
rect -4300 -288 -3200 -248
rect -7500 -340 -4900 -300
rect -7500 -6460 -7460 -340
rect -4940 -6460 -4900 -340
rect -4300 -5608 -4260 -288
rect -3240 -5608 -3200 -288
rect 2800 -2960 2840 560
rect 4160 -2960 4200 560
rect 2800 -3000 4200 -2960
rect -4300 -5648 -3200 -5608
rect -7500 -6500 -4900 -6460
<< mimcap2contact >>
rect -7460 -6460 -4940 -340
rect -4260 -5608 -3240 -288
rect 2840 -2960 4160 560
<< metal5 >>
rect 2700 560 4300 700
rect -7600 -340 -4800 -200
rect -7600 -6460 -7460 -340
rect -4940 -6460 -4800 -340
rect -7600 -7100 -4800 -6460
rect -4400 -288 -3100 -148
rect -4400 -5608 -4260 -288
rect -3240 -5608 -3100 -288
rect 2700 -2960 2840 560
rect 4160 -2960 4300 560
rect 2700 -3100 4300 -2960
rect 3380 -3540 4300 -3100
rect 3380 -3820 3420 -3540
rect 4260 -3820 4300 -3540
rect 3380 -3860 4300 -3820
rect -4400 -5748 -3100 -5608
rect -4400 -6248 -3500 -5748
rect -4400 -6648 -4300 -6248
rect -3600 -6648 -3500 -6248
rect -4400 -6748 -3500 -6648
rect -7600 -7700 -7500 -7100
rect -4900 -7700 -4800 -7100
rect -7600 -7800 -4800 -7700
<< comment >>
rect -236 -5100 -233 -560
<< labels >>
rlabel metal4 -3840 -7800 -3660 -7300 1 VLO
rlabel metal4 -4220 320 -3840 600 1 VHI
rlabel metal3 -660 -4200 -620 -4180 1 VIN
rlabel metal3 120 -4200 160 -4180 1 VIP
rlabel metal1 -4369 -7084 -4329 -7044 1 S
rlabel metal1 -4301 -7084 -4261 -7044 1 SBAR
rlabel metal2 -4200 -7084 -4120 -7004 1 VREF
rlabel metal4 2580 -3100 2680 -2980 1 VOP
<< end >>
