magic
tech sky130A
magscale 1 2
timestamp 1671335613
<< pwell >>
rect 948 781 2082 860
rect 948 772 1734 781
rect 1840 772 2082 781
rect 948 744 2082 772
rect 948 698 1414 744
rect 1418 698 2082 744
rect 948 -60 2082 698
<< nmos >>
rect 1148 150 1178 650
rect 1244 150 1274 650
rect 1340 150 1370 650
rect 1436 150 1466 650
<< ndiff >>
rect 1086 638 1148 650
rect 1086 162 1098 638
rect 1132 162 1148 638
rect 1086 150 1148 162
rect 1178 638 1244 650
rect 1178 162 1194 638
rect 1228 162 1244 638
rect 1178 150 1244 162
rect 1274 638 1340 650
rect 1274 162 1290 638
rect 1324 162 1340 638
rect 1274 150 1340 162
rect 1370 638 1436 650
rect 1370 162 1386 638
rect 1420 162 1436 638
rect 1370 150 1436 162
rect 1466 638 1528 650
rect 1466 162 1482 638
rect 1516 162 1528 638
rect 1466 150 1528 162
<< ndiffc >>
rect 1098 162 1132 638
rect 1194 162 1228 638
rect 1290 162 1324 638
rect 1386 162 1420 638
rect 1482 162 1516 638
<< psubdiff >>
rect 984 790 1080 824
rect 1930 790 2046 824
rect 984 728 1018 790
rect 2012 728 2046 790
rect 984 10 1018 72
rect 2012 10 2046 72
rect 984 -24 1080 10
rect 1930 -24 2046 10
<< psubdiffcont >>
rect 1080 790 1930 824
rect 984 72 1018 728
rect 2012 72 2046 728
rect 1080 -24 1930 10
<< poly >>
rect 1148 650 1178 676
rect 1244 650 1274 676
rect 1340 650 1370 676
rect 1436 650 1466 676
rect 1148 128 1178 150
rect 1244 128 1274 150
rect 1148 112 1274 128
rect 1148 78 1164 112
rect 1198 78 1274 112
rect 1148 62 1274 78
rect 1340 128 1370 150
rect 1436 128 1466 150
rect 1340 112 1466 128
rect 1340 78 1356 112
rect 1390 78 1466 112
rect 1340 62 1466 78
<< polycont >>
rect 1164 78 1198 112
rect 1356 78 1390 112
<< xpolycontact >>
rect 1634 106 1704 538
rect 1800 106 1870 538
<< xpolyres >>
rect 1634 604 1870 674
rect 1634 538 1704 604
rect 1800 538 1870 604
<< locali >>
rect 960 858 1920 980
rect 950 824 2080 858
rect 950 790 1080 824
rect 1930 790 2080 824
rect 950 728 1018 790
rect 950 72 984 728
rect 1098 638 1132 654
rect 1098 146 1132 162
rect 1194 638 1228 654
rect 1194 146 1228 162
rect 1290 638 1324 654
rect 1290 146 1324 162
rect 1386 638 1420 790
rect 2012 728 2080 790
rect 1386 146 1420 162
rect 1482 638 1516 654
rect 1482 118 1516 162
rect 1148 78 1164 112
rect 1198 78 1214 112
rect 1340 78 1356 112
rect 1390 78 1406 112
rect 1482 106 1634 118
rect 950 10 1018 72
rect 1482 67 1704 106
rect 1800 90 1808 106
rect 1861 90 1870 106
rect 1800 67 1870 90
rect 2046 72 2080 728
rect 2012 10 2080 72
rect 950 -24 1080 10
rect 1930 -24 2080 10
rect 950 -58 2080 -24
<< viali >>
rect 1098 162 1132 638
rect 1194 162 1228 638
rect 1290 162 1324 638
rect 1386 162 1420 638
rect 1482 162 1516 638
rect 1164 78 1198 112
rect 1356 78 1390 112
rect 1808 106 1861 522
rect 1808 90 1861 106
<< metal1 >>
rect 960 1100 1920 1120
rect 960 900 980 1100
rect 1900 900 1920 1100
rect 960 880 1920 900
rect 1092 718 1522 758
rect 1092 638 1138 718
rect 1092 162 1098 638
rect 1132 162 1138 638
rect 1092 150 1138 162
rect 1185 638 1237 650
rect 1185 635 1194 638
rect 1228 635 1237 638
rect 1185 162 1194 166
rect 1228 162 1237 166
rect 1185 149 1237 162
rect 1284 638 1330 718
rect 1284 162 1290 638
rect 1324 162 1330 638
rect 1284 150 1330 162
rect 1380 638 1426 650
rect 1380 162 1386 638
rect 1420 162 1426 638
rect 1380 150 1426 162
rect 1476 638 1522 718
rect 1476 162 1482 638
rect 1516 162 1522 638
rect 1476 150 1522 162
rect 1800 522 1870 538
rect 1800 519 1808 522
rect 1861 519 1870 522
rect 954 112 1274 118
rect 954 78 1164 112
rect 1198 78 1274 112
rect 954 72 1274 78
rect 1340 112 1466 118
rect 1340 78 1356 112
rect 1390 78 1466 112
rect 1340 72 1466 78
rect 1374 44 1420 72
rect 1800 67 1870 90
rect 954 -2 1420 44
<< via1 >>
rect 980 900 1900 1100
rect 1185 166 1194 635
rect 1194 166 1228 635
rect 1228 166 1237 635
rect 1800 90 1808 519
rect 1808 90 1861 519
rect 1861 90 1870 519
<< metal2 >>
rect 960 1100 1920 1120
rect 960 900 980 1100
rect 1900 900 1920 1100
rect 960 880 1920 900
rect 949 635 1237 650
rect 949 515 1185 635
rect 2000 580 2200 600
rect 2000 538 2020 580
rect 1185 149 1237 166
rect 1800 519 2020 538
rect 1870 460 2020 519
rect 2000 420 2020 460
rect 2180 420 2200 580
rect 2000 400 2200 420
rect 1800 67 1870 90
<< via2 >>
rect 980 900 1900 1100
rect 2020 420 2180 580
<< metal3 >>
rect 960 1180 1920 1200
rect 960 900 980 1180
rect 1900 900 1920 1180
rect 960 880 1920 900
rect 2200 800 7800 1200
rect 1500 700 7800 800
rect 1900 580 7800 700
rect 1900 420 2020 580
rect 2180 420 7800 580
rect 1900 0 7800 420
rect 1448 -24 7800 0
rect 1400 -100 7800 -24
<< via3 >>
rect 980 1100 1900 1180
rect 980 980 1900 1100
rect 1500 0 1900 700
<< mimcap >>
rect 2300 1060 7700 1100
rect 2300 40 2340 1060
rect 7660 40 7700 1060
rect 2300 0 7700 40
<< mimcapcontact >>
rect 2340 40 7660 1060
<< metal4 >>
rect 960 1180 7800 1200
rect 960 980 980 1180
rect 1900 1060 7800 1180
rect 1900 1000 2340 1060
rect 1900 980 1920 1000
rect 960 960 1920 980
rect 1400 700 2000 800
rect 1400 0 1500 700
rect 1900 0 2000 700
rect 1400 -100 2000 0
rect 2200 40 2340 1000
rect 7660 40 7800 1060
rect 2200 -100 7800 40
<< via4 >>
rect 1500 0 1900 700
<< mimcap2 >>
rect 2300 1060 7700 1100
rect 2300 40 2340 1060
rect 7660 40 7700 1060
rect 2300 0 7700 40
<< mimcap2contact >>
rect 2340 40 7660 1060
<< metal5 >>
rect 2200 1060 7800 1200
rect 2200 800 2340 1060
rect 1400 700 2340 800
rect 1400 0 1500 700
rect 1900 40 2340 700
rect 7660 40 7800 1060
rect 1900 0 7800 40
rect 1400 -100 7800 0
<< labels >>
rlabel metal1 954 72 977 118 1 S
rlabel metal1 954 -2 977 44 1 SBAR
rlabel metal2 949 515 973 650 1 IN
rlabel metal3 2200 800 2300 860 1 OUT
rlabel locali 960 820 1080 840 1 VSUB
<< end >>
