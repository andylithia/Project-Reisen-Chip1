magic
tech sky130B
magscale 1 2
timestamp 1668748373
<< dnwell >>
rect 1600 -600 3600 1400
<< nwell >>
rect 1520 1194 3680 1480
rect 1520 -394 1806 1194
rect 2147 611 3053 853
rect 2147 165 2399 611
rect 2801 165 3053 611
rect 2147 -53 3053 165
rect 3394 -394 3680 1194
rect 1520 -680 3680 -394
<< pwell >>
rect 2399 165 2801 611
<< nmos >>
rect 2585 327 2615 411
<< ndiff >>
rect 2527 399 2585 411
rect 2527 339 2539 399
rect 2573 339 2585 399
rect 2527 327 2585 339
rect 2615 399 2673 411
rect 2615 339 2627 399
rect 2661 339 2673 399
rect 2615 327 2673 339
<< ndiffc >>
rect 2539 339 2573 399
rect 2627 339 2661 399
<< psubdiff >>
rect 2425 551 2521 585
rect 2679 551 2775 585
rect 2425 489 2459 551
rect 2741 489 2775 551
rect 2425 249 2459 311
rect 2741 249 2775 311
rect 2425 215 2521 249
rect 2679 215 2775 249
<< nsubdiff >>
rect 1557 1423 3643 1443
rect 1557 1389 1637 1423
rect 3563 1389 3643 1423
rect 1557 1369 3643 1389
rect 1557 1363 1631 1369
rect 1557 -563 1577 1363
rect 1611 -563 1631 1363
rect 3569 1363 3643 1369
rect 2183 783 2243 817
rect 2957 783 3017 817
rect 2183 757 2217 783
rect 2983 757 3017 783
rect 2183 17 2217 43
rect 2983 17 3017 43
rect 2183 -17 2243 17
rect 2957 -17 3017 17
rect 1557 -569 1631 -563
rect 3569 -563 3589 1363
rect 3623 -563 3643 1363
rect 3569 -569 3643 -563
rect 1557 -589 3643 -569
rect 1557 -623 1637 -589
rect 3563 -623 3643 -589
rect 1557 -643 3643 -623
<< psubdiffcont >>
rect 2521 551 2679 585
rect 2425 311 2459 489
rect 2741 311 2775 489
rect 2521 215 2679 249
<< nsubdiffcont >>
rect 1637 1389 3563 1423
rect 1577 -563 1611 1363
rect 2243 783 2957 817
rect 2183 43 2217 757
rect 2983 43 3017 757
rect 2243 -17 2957 17
rect 3589 -563 3623 1363
rect 1637 -623 3563 -589
<< poly >>
rect 2567 483 2633 499
rect 2567 449 2583 483
rect 2617 449 2633 483
rect 2567 433 2633 449
rect 2585 411 2615 433
rect 2585 301 2615 327
<< polycont >>
rect 2583 449 2617 483
<< locali >>
rect 1577 1389 1637 1423
rect 3563 1389 3623 1423
rect 1577 1363 1611 1389
rect 3589 1363 3623 1389
rect 2183 783 2243 817
rect 2957 783 3017 817
rect 2183 757 2217 783
rect 2983 757 3017 783
rect 2425 551 2521 585
rect 2679 551 2775 585
rect 2425 489 2459 551
rect 2741 489 2775 551
rect 2567 449 2583 483
rect 2617 449 2633 483
rect 2539 399 2573 415
rect 2539 323 2573 339
rect 2627 399 2661 415
rect 2627 323 2661 339
rect 2425 249 2459 311
rect 2741 249 2775 311
rect 2425 215 2521 249
rect 2679 215 2775 249
rect 2183 17 2217 43
rect 2983 17 3017 43
rect 2183 -17 2243 17
rect 2957 -17 3017 17
rect 1577 -589 1611 -563
rect 3589 -589 3623 -563
rect 1577 -623 1637 -589
rect 3563 -623 3623 -589
<< viali >>
rect 2583 449 2617 483
rect 2539 339 2573 399
rect 2627 339 2661 399
<< metal1 >>
rect 2407 569 2459 585
rect 2741 569 2793 585
rect 2559 501 2641 507
rect 2559 449 2573 501
rect 2625 449 2641 501
rect 2559 443 2641 449
rect 2519 399 2579 415
rect 2519 395 2539 399
rect 2573 395 2579 399
rect 2519 343 2527 395
rect 2519 339 2539 343
rect 2573 339 2579 343
rect 2519 323 2579 339
rect 2621 399 2681 415
rect 2621 395 2627 399
rect 2661 395 2681 399
rect 2673 343 2681 395
rect 2621 339 2627 343
rect 2661 339 2681 343
rect 2621 323 2681 339
rect 2407 249 2459 265
rect 2741 249 2793 265
rect 2407 197 2475 249
rect 2725 197 2793 249
<< via1 >>
rect 2407 265 2459 569
rect 2573 483 2625 501
rect 2573 449 2583 483
rect 2583 449 2617 483
rect 2617 449 2625 483
rect 2527 343 2539 395
rect 2539 343 2573 395
rect 2573 343 2579 395
rect 2621 343 2627 395
rect 2627 343 2661 395
rect 2661 343 2673 395
rect 2741 265 2793 569
rect 2475 197 2725 249
<< metal2 >>
rect 2407 569 2459 585
rect 2741 569 2793 585
rect 2559 525 2641 527
rect 2559 469 2571 525
rect 2627 469 2641 525
rect 2559 449 2573 469
rect 2625 449 2641 469
rect 2559 443 2641 449
rect 2519 397 2579 415
rect 2519 341 2523 397
rect 2519 323 2579 341
rect 2621 397 2681 415
rect 2677 341 2681 397
rect 2621 323 2681 341
rect 2407 249 2459 265
rect 2741 249 2793 265
rect 2407 241 2475 249
rect 2725 241 2793 249
rect 2407 185 2417 241
rect 2783 185 2793 241
rect 2407 177 2793 185
<< via2 >>
rect 2571 501 2627 525
rect 2571 469 2573 501
rect 2573 469 2625 501
rect 2625 469 2627 501
rect 2523 395 2579 397
rect 2523 343 2527 395
rect 2527 343 2579 395
rect 2523 341 2579 343
rect 2621 395 2677 397
rect 2621 343 2673 395
rect 2673 343 2677 395
rect 2621 341 2677 343
rect 2417 197 2475 241
rect 2475 197 2725 241
rect 2725 197 2783 241
rect 2417 185 2783 197
<< metal3 >>
rect 2559 525 2641 607
rect 2559 469 2571 525
rect 2627 469 2641 525
rect 2559 463 2641 469
rect 2517 397 2683 403
rect 2517 341 2523 397
rect 2579 341 2621 397
rect 2677 341 2683 397
rect 2517 323 2683 341
rect 2407 241 2793 249
rect 2407 185 2417 241
rect 2783 185 2793 241
rect 2407 177 2793 185
<< comment >>
rect 2425 569 2459 585
rect 2741 569 2775 585
rect 2425 249 2459 265
rect 2741 249 2775 265
rect 2459 215 2475 249
rect 2725 215 2741 249
<< end >>
