magic
tech sky130A
magscale 1 2
timestamp 1671941875
<< nwell >>
rect 5945 10066 10055 12504
rect 2001 2544 10237 2916
rect 2001 1488 10237 1880
rect 11224 1518 14480 3956
rect 1729 1212 10237 1488
rect 1729 1167 2909 1212
rect 10210 -1404 10531 -316
rect 5945 -9104 10055 -6666
<< pwell >>
rect 5709 9618 6751 9986
rect 5006 8250 6751 9618
rect 6873 8890 9127 9810
rect 5709 7566 6751 8250
rect 6917 6450 9083 8870
rect 9250 7566 10292 9986
rect 10642 6986 11562 7452
rect 10642 6982 10758 6986
rect 10804 6982 11562 6986
rect 10642 6666 11562 6982
rect 10642 6560 10721 6666
rect 10730 6560 11562 6666
rect 10642 6318 11562 6560
rect 3319 4432 3741 4562
rect 3319 4379 3499 4432
rect 3553 4379 3741 4432
rect 3319 3718 3741 4379
rect 3319 3665 3499 3718
rect 3553 3665 3741 3718
rect 3319 3028 3741 3665
rect 4101 4432 4523 4562
rect 4101 4379 4289 4432
rect 4343 4379 4523 4432
rect 4101 3718 4523 4379
rect 4101 3665 4289 3718
rect 4343 3665 4523 3718
rect 4101 3028 4523 3665
rect 2044 2250 2130 2467
rect 2136 2261 2326 2488
rect 2402 2261 2612 2460
rect 3771 2261 4045 2460
rect 4071 2261 4688 2407
rect 5212 2261 5394 2467
rect 5415 2261 6032 2407
rect 6087 2261 6704 2407
rect 6759 2261 7376 2407
rect 8103 2261 8720 2407
rect 8775 2261 9392 2407
rect 9447 2261 9809 2407
rect 9820 2261 9906 2467
rect 2044 1957 2130 2174
rect 2135 2163 10103 2261
rect 10108 2250 10194 2467
rect 2136 1936 2326 2163
rect 2402 1964 2612 2163
rect 3771 1964 4045 2163
rect 4056 1964 4916 2163
rect 4923 1964 5205 2163
rect 5212 1957 5394 2163
rect 5405 2020 9046 2163
rect 5405 1994 7472 2020
rect 5405 1983 7377 1994
rect 6061 1977 7377 1983
rect 6061 1940 6425 1977
rect 6846 1951 7377 1977
rect 7745 1964 9046 2020
rect 9048 1964 9238 2163
rect 9240 1964 10102 2163
rect 8142 1922 8330 1964
rect 10108 1957 10194 2174
rect 10656 1518 11224 2786
rect 1770 944 1856 1101
rect 1864 919 2042 1109
rect 2046 944 2132 1101
rect 2138 944 2224 1101
rect 2232 919 2410 1109
rect 2414 944 2500 1101
rect 2506 944 2592 1101
rect 2600 919 2778 1109
rect 2782 944 2868 1101
rect 1888 889 1922 919
rect 2256 889 2290 919
rect 2624 889 2658 919
rect 3196 918 3282 1135
rect 3288 929 3478 1156
rect 3554 929 3764 1128
rect 4923 929 5197 1128
rect 5212 929 5394 1135
rect 6061 1115 6425 1152
rect 6846 1115 7377 1141
rect 8142 1128 8330 1170
rect 6061 1109 7377 1115
rect 5405 1098 7377 1109
rect 5405 1072 7472 1098
rect 7745 1072 9046 1128
rect 5405 929 9046 1072
rect 9048 929 9238 1128
rect 9240 929 10102 1153
rect 3287 880 10103 929
rect 10108 918 10194 1135
rect 3668 662 4090 792
rect 3668 609 3856 662
rect 3910 609 4090 662
rect 3668 -52 4090 609
rect 10308 98 14480 1518
rect 15330 871 38998 1051
rect 15330 817 15460 871
rect 15513 817 16174 871
rect 16227 817 16888 871
rect 16941 817 17602 871
rect 17655 817 18316 871
rect 18369 817 19030 871
rect 19083 817 19744 871
rect 19797 817 20458 871
rect 20511 817 21172 871
rect 21225 817 21886 871
rect 21939 817 22600 871
rect 22653 817 23314 871
rect 23367 817 24028 871
rect 24081 817 24742 871
rect 24795 817 25456 871
rect 25509 817 26170 871
rect 26223 817 26884 871
rect 26937 817 27598 871
rect 27651 817 28312 871
rect 28365 817 29026 871
rect 29079 817 29740 871
rect 29793 817 30454 871
rect 30507 817 31168 871
rect 31221 817 31882 871
rect 31935 817 32596 871
rect 32649 817 33310 871
rect 33363 817 34024 871
rect 34077 817 34738 871
rect 34791 817 35452 871
rect 35505 817 36166 871
rect 36219 817 36880 871
rect 36933 817 37594 871
rect 37647 817 38308 871
rect 38361 817 38998 871
rect 15330 629 38998 817
rect 3668 -105 3856 -52
rect 3910 -105 4090 -52
rect 3668 -742 4090 -105
rect 15330 45 38998 233
rect 15330 -9 15460 45
rect 15513 -9 16174 45
rect 16227 -9 16888 45
rect 16941 -9 17602 45
rect 17655 -9 18316 45
rect 18369 -9 19030 45
rect 19083 -9 19744 45
rect 19797 -9 20458 45
rect 20511 -9 21172 45
rect 21225 -9 21886 45
rect 21939 -9 22600 45
rect 22653 -9 23314 45
rect 23367 -9 24028 45
rect 24081 -9 24742 45
rect 24795 -9 25456 45
rect 25509 -9 26170 45
rect 26223 -9 26884 45
rect 26937 -9 27598 45
rect 27651 -9 28312 45
rect 28365 -9 29026 45
rect 29079 -9 29740 45
rect 29793 -9 30454 45
rect 30507 -9 31168 45
rect 31221 -9 31882 45
rect 31935 -9 32596 45
rect 32649 -9 33310 45
rect 33363 -9 34024 45
rect 34077 -9 34738 45
rect 34791 -9 35452 45
rect 35505 -9 36166 45
rect 36219 -9 36880 45
rect 36933 -9 37594 45
rect 37647 -9 38308 45
rect 38361 -9 38998 45
rect 15330 -189 38998 -9
rect 39197 -353 40493 1211
rect 10597 -443 10754 -357
rect 10589 -475 10779 -451
rect 10589 -509 10809 -475
rect 10589 -629 10779 -509
rect 10597 -719 10754 -633
rect 10589 -935 10771 -770
rect 10589 -956 10809 -935
rect 10775 -969 10809 -956
rect 10597 -1087 10754 -1001
rect 10589 -1119 10779 -1095
rect 10589 -1153 10809 -1119
rect 10589 -1273 10779 -1153
rect 10597 -1363 10754 -1277
rect 5709 -4850 6751 -4166
rect 5006 -6218 6751 -4850
rect 6917 -5470 9083 -3050
rect 10642 -3160 11562 -2918
rect 10642 -3266 10721 -3160
rect 10730 -3266 11562 -3160
rect 10642 -3582 11562 -3266
rect 10642 -3586 10758 -3582
rect 10804 -3586 11562 -3582
rect 10642 -4052 11562 -3586
rect 5709 -6586 6751 -6218
rect 6873 -6410 9127 -5490
rect 9250 -6586 10292 -4166
<< nmos >>
rect 5905 7776 5965 9776
rect 6023 7776 6083 9776
rect 6141 7776 6201 9776
rect 6259 7776 6319 9776
rect 6377 7776 6437 9776
rect 6495 7776 6555 9776
rect 7113 6660 7513 8660
rect 7571 6660 7971 8660
rect 8029 6660 8429 8660
rect 8487 6660 8887 8660
rect 9446 7776 9506 9776
rect 9564 7776 9624 9776
rect 9682 7776 9742 9776
rect 9800 7776 9860 9776
rect 9918 7776 9978 9776
rect 10036 7776 10096 9776
rect 10852 7222 11352 7252
rect 10852 7126 11352 7156
rect 10852 7030 11352 7060
rect 10852 6934 11352 6964
rect 3515 3952 3545 4352
rect 3515 3238 3545 3638
rect 4297 3952 4327 4352
rect 4297 3238 4327 3638
rect 3864 182 3894 582
rect 10504 308 10904 1308
rect 10962 308 11362 1308
rect 11420 308 11820 1308
rect 11878 308 12278 1308
rect 12336 308 12736 1308
rect 12794 308 13194 1308
rect 13252 308 13652 1308
rect 13938 308 13968 1308
rect 14254 308 14284 1308
rect 15540 825 15940 855
rect 16254 825 16654 855
rect 16968 825 17368 855
rect 17682 825 18082 855
rect 18396 825 18796 855
rect 19110 825 19510 855
rect 19824 825 20224 855
rect 20538 825 20938 855
rect 21252 825 21652 855
rect 21966 825 22366 855
rect 22680 825 23080 855
rect 23394 825 23794 855
rect 24108 825 24508 855
rect 24822 825 25222 855
rect 25536 825 25936 855
rect 26250 825 26650 855
rect 26964 825 27364 855
rect 27678 825 28078 855
rect 28392 825 28792 855
rect 29106 825 29506 855
rect 29820 825 30220 855
rect 30534 825 30934 855
rect 31248 825 31648 855
rect 31962 825 32362 855
rect 32676 825 33076 855
rect 33390 825 33790 855
rect 34104 825 34504 855
rect 34818 825 35218 855
rect 35532 825 35932 855
rect 36246 825 36646 855
rect 36960 825 37360 855
rect 37674 825 38074 855
rect 38388 825 38788 855
rect 3864 -532 3894 -132
rect 15540 7 15940 37
rect 16254 7 16654 37
rect 16968 7 17368 37
rect 17682 7 18082 37
rect 18396 7 18796 37
rect 19110 7 19510 37
rect 19824 7 20224 37
rect 20538 7 20938 37
rect 21252 7 21652 37
rect 21966 7 22366 37
rect 22680 7 23080 37
rect 23394 7 23794 37
rect 24108 7 24508 37
rect 24822 7 25222 37
rect 25536 7 25936 37
rect 26250 7 26650 37
rect 26964 7 27364 37
rect 27678 7 28078 37
rect 28392 7 28792 37
rect 29106 7 29506 37
rect 29820 7 30220 37
rect 30534 7 30934 37
rect 31248 7 31648 37
rect 31962 7 32362 37
rect 32676 7 33076 37
rect 33390 7 33790 37
rect 34104 7 34504 37
rect 34818 7 35218 37
rect 35532 7 35932 37
rect 36246 7 36646 37
rect 36960 7 37360 37
rect 37674 7 38074 37
rect 38388 7 38788 37
rect 5905 -6376 5965 -4376
rect 6023 -6376 6083 -4376
rect 6141 -6376 6201 -4376
rect 6259 -6376 6319 -4376
rect 6377 -6376 6437 -4376
rect 6495 -6376 6555 -4376
rect 7113 -5260 7513 -3260
rect 7571 -5260 7971 -3260
rect 8029 -5260 8429 -3260
rect 8487 -5260 8887 -3260
rect 10852 -3564 11352 -3534
rect 10852 -3660 11352 -3630
rect 10852 -3756 11352 -3726
rect 10852 -3852 11352 -3822
rect 9446 -6376 9506 -4376
rect 9564 -6376 9624 -4376
rect 9682 -6376 9742 -4376
rect 9800 -6376 9860 -4376
rect 9918 -6376 9978 -4376
rect 10036 -6376 10096 -4376
<< scnmos >>
rect 10615 -878 10745 -848
<< pmos >>
rect 6141 10285 6201 12285
rect 6259 10285 6319 12285
rect 6377 10285 6437 12285
rect 6495 10285 6555 12285
rect 6613 10285 6673 12285
rect 6731 10285 6791 12285
rect 6849 10285 6909 12285
rect 6967 10285 7027 12285
rect 7085 10285 7145 12285
rect 7203 10285 7263 12285
rect 7321 10285 7381 12285
rect 7439 10285 7499 12285
rect 7557 10285 7617 12285
rect 7675 10285 7735 12285
rect 7793 10285 7853 12285
rect 7911 10285 7971 12285
rect 8029 10285 8089 12285
rect 8147 10285 8207 12285
rect 8265 10285 8325 12285
rect 8383 10285 8443 12285
rect 8501 10285 8561 12285
rect 8619 10285 8679 12285
rect 8737 10285 8797 12285
rect 8855 10285 8915 12285
rect 8973 10285 9033 12285
rect 9091 10285 9151 12285
rect 9209 10285 9269 12285
rect 9327 10285 9387 12285
rect 9445 10285 9505 12285
rect 9563 10285 9623 12285
rect 9681 10285 9741 12285
rect 9799 10285 9859 12285
rect 11420 1737 11820 3737
rect 11878 1737 12278 3737
rect 12336 1737 12736 3737
rect 12794 1737 13194 3737
rect 13252 1737 13652 3737
rect 13938 1737 13968 3737
rect 14254 1737 14284 3737
rect 6141 -8885 6201 -6885
rect 6259 -8885 6319 -6885
rect 6377 -8885 6437 -6885
rect 6495 -8885 6555 -6885
rect 6613 -8885 6673 -6885
rect 6731 -8885 6791 -6885
rect 6849 -8885 6909 -6885
rect 6967 -8885 7027 -6885
rect 7085 -8885 7145 -6885
rect 7203 -8885 7263 -6885
rect 7321 -8885 7381 -6885
rect 7439 -8885 7499 -6885
rect 7557 -8885 7617 -6885
rect 7675 -8885 7735 -6885
rect 7793 -8885 7853 -6885
rect 7911 -8885 7971 -6885
rect 8029 -8885 8089 -6885
rect 8147 -8885 8207 -6885
rect 8265 -8885 8325 -6885
rect 8383 -8885 8443 -6885
rect 8501 -8885 8561 -6885
rect 8619 -8885 8679 -6885
rect 8737 -8885 8797 -6885
rect 8855 -8885 8915 -6885
rect 8973 -8885 9033 -6885
rect 9091 -8885 9151 -6885
rect 9209 -8885 9269 -6885
rect 9327 -8885 9387 -6885
rect 9445 -8885 9505 -6885
rect 9563 -8885 9623 -6885
rect 9681 -8885 9741 -6885
rect 9799 -8885 9859 -6885
<< scpmos >>
rect 2497 2580 2527 2804
rect 3851 2580 3881 2804
rect 3941 2580 3971 2804
rect 4137 2604 4337 2804
rect 4392 2604 4592 2804
rect 5481 2604 5681 2804
rect 5736 2604 5936 2804
rect 6153 2604 6353 2804
rect 6408 2604 6608 2804
rect 6825 2604 7025 2804
rect 7080 2604 7280 2804
rect 8169 2604 8369 2804
rect 8424 2604 8624 2804
rect 8841 2604 9041 2804
rect 9096 2604 9296 2804
rect 9513 2604 9713 2804
rect 2497 1620 2527 1844
rect 3851 1620 3881 1844
rect 3941 1620 3971 1844
rect 4141 1676 4171 1844
rect 4248 1644 4278 1844
rect 4441 1644 4471 1844
rect 4549 1644 4579 1844
rect 4663 1644 4693 1844
rect 4787 1620 4817 1844
rect 5003 1620 5033 1844
rect 5093 1620 5123 1844
rect 5485 1620 5515 1748
rect 5575 1620 5605 1748
rect 5653 1620 5683 1748
rect 5743 1620 5773 1748
rect 5945 1620 5975 1748
rect 6147 1620 6177 1844
rect 6237 1620 6267 1844
rect 6439 1664 6469 1748
rect 6523 1664 6553 1748
rect 6630 1620 6660 1748
rect 6961 1620 6991 1788
rect 7045 1620 7075 1788
rect 7153 1620 7183 1788
rect 7355 1620 7385 1788
rect 7433 1620 7463 1788
rect 7540 1620 7570 1704
rect 7618 1620 7648 1704
rect 7823 1620 7853 1820
rect 7925 1620 7955 1820
rect 8009 1620 8039 1820
rect 8211 1685 8241 1813
rect 8447 1620 8477 1844
rect 8537 1620 8567 1844
rect 8736 1628 8766 1828
rect 8841 1620 8871 1844
rect 8931 1620 8961 1844
rect 9326 1620 9356 1844
rect 9578 1620 9608 1844
rect 9678 1620 9708 1844
rect 9977 1620 10007 1844
rect 3649 1248 3679 1472
rect 5003 1248 5033 1472
rect 5093 1248 5123 1472
rect 5485 1344 5515 1472
rect 5575 1344 5605 1472
rect 5653 1344 5683 1472
rect 5743 1344 5773 1472
rect 5945 1344 5975 1472
rect 6147 1248 6177 1472
rect 6237 1248 6267 1472
rect 6439 1344 6469 1428
rect 6523 1344 6553 1428
rect 6630 1344 6660 1472
rect 6961 1304 6991 1472
rect 7045 1304 7075 1472
rect 7153 1304 7183 1472
rect 7355 1304 7385 1472
rect 7433 1304 7463 1472
rect 7540 1388 7570 1472
rect 7618 1388 7648 1472
rect 7823 1272 7853 1472
rect 7925 1272 7955 1472
rect 8009 1272 8039 1472
rect 8211 1279 8241 1407
rect 8447 1248 8477 1472
rect 8537 1248 8567 1472
rect 8736 1264 8766 1464
rect 8841 1248 8871 1472
rect 8931 1248 8961 1472
rect 9326 1289 9356 1457
rect 9416 1289 9446 1457
rect 9511 1289 9541 1457
rect 9606 1289 9636 1457
rect 9713 1248 9743 1472
rect 9807 1248 9837 1472
rect 9897 1248 9927 1472
rect 9987 1248 10017 1472
<< scpmoshvt >>
rect 10295 -878 10495 -848
<< nmoslvt >>
rect 7073 9100 7103 9600
rect 7169 9100 7199 9600
rect 7265 9100 7295 9600
rect 7361 9100 7391 9600
rect 7457 9100 7487 9600
rect 7553 9100 7583 9600
rect 7649 9100 7679 9600
rect 7745 9100 7775 9600
rect 7841 9100 7871 9600
rect 7937 9100 7967 9600
rect 8033 9100 8063 9600
rect 8129 9100 8159 9600
rect 8225 9100 8255 9600
rect 8321 9100 8351 9600
rect 8417 9100 8447 9600
rect 8513 9100 8543 9600
rect 8609 9100 8639 9600
rect 8705 9100 8735 9600
rect 8801 9100 8831 9600
rect 8897 9100 8927 9600
rect 2499 2286 2529 2434
rect 3854 2286 3884 2434
rect 3932 2286 3962 2434
rect 4150 2297 4350 2381
rect 4406 2297 4606 2381
rect 5494 2297 5694 2381
rect 5750 2297 5950 2381
rect 6166 2297 6366 2381
rect 6422 2297 6622 2381
rect 6838 2297 7038 2381
rect 7094 2297 7294 2381
rect 8182 2297 8382 2381
rect 8438 2297 8638 2381
rect 8854 2297 9054 2381
rect 9110 2297 9310 2381
rect 9526 2297 9726 2381
rect 2499 1990 2529 2138
rect 3854 1990 3884 2138
rect 3932 1990 3962 2138
rect 4139 1990 4169 2100
rect 4251 1990 4281 2138
rect 4329 1990 4359 2138
rect 4468 1990 4498 2138
rect 4660 1990 4690 2138
rect 4803 1990 4833 2138
rect 5006 1990 5036 2138
rect 5092 1990 5122 2138
rect 5488 2009 5518 2093
rect 5566 2009 5596 2093
rect 5732 2009 5762 2093
rect 5810 2009 5840 2093
rect 5946 2009 5976 2093
rect 6144 1966 6174 2114
rect 6312 1966 6342 2114
rect 6554 2003 6584 2087
rect 6626 2003 6656 2087
rect 6717 2003 6747 2087
rect 6964 1977 6994 2087
rect 7050 1977 7080 2087
rect 7171 1977 7201 2087
rect 7271 1977 7301 2087
rect 7366 2020 7396 2130
rect 7616 2046 7646 2130
rect 7694 2046 7724 2130
rect 7821 1990 7851 2138
rect 7925 1990 7955 2138
rect 8011 1990 8041 2138
rect 8224 1948 8254 2032
rect 8430 1990 8460 2138
rect 8516 1990 8546 2138
rect 8728 1990 8758 2118
rect 8848 1990 8878 2138
rect 8934 1990 8964 2138
rect 9323 1990 9353 2138
rect 9409 1990 9439 2138
rect 9495 1990 9525 2138
rect 9581 1990 9611 2138
rect 9675 1990 9705 2138
rect 9767 1990 9797 2138
rect 9867 1990 9897 2138
rect 9980 1990 10010 2138
rect 3651 954 3681 1102
rect 5006 954 5036 1102
rect 5084 954 5114 1102
rect 5488 999 5518 1083
rect 5566 999 5596 1083
rect 5732 999 5762 1083
rect 5810 999 5840 1083
rect 5946 999 5976 1083
rect 6144 978 6174 1126
rect 6312 978 6342 1126
rect 6554 1005 6584 1089
rect 6626 1005 6656 1089
rect 6717 1005 6747 1089
rect 6964 1005 6994 1115
rect 7050 1005 7080 1115
rect 7171 1005 7201 1115
rect 7271 1005 7301 1115
rect 7366 962 7396 1072
rect 7616 962 7646 1046
rect 7694 962 7724 1046
rect 7821 954 7851 1102
rect 7925 954 7955 1102
rect 8011 954 8041 1102
rect 8224 1060 8254 1144
rect 8430 954 8460 1102
rect 8516 954 8546 1102
rect 8728 974 8758 1102
rect 8848 954 8878 1102
rect 8934 954 8964 1102
rect 9323 999 9353 1127
rect 9413 999 9443 1127
rect 9508 999 9538 1127
rect 9599 999 9629 1127
rect 9701 979 9731 1127
rect 9817 979 9847 1127
rect 9903 979 9933 1127
rect 9989 979 10019 1127
rect 7073 -6200 7103 -5700
rect 7169 -6200 7199 -5700
rect 7265 -6200 7295 -5700
rect 7361 -6200 7391 -5700
rect 7457 -6200 7487 -5700
rect 7553 -6200 7583 -5700
rect 7649 -6200 7679 -5700
rect 7745 -6200 7775 -5700
rect 7841 -6200 7871 -5700
rect 7937 -6200 7967 -5700
rect 8033 -6200 8063 -5700
rect 8129 -6200 8159 -5700
rect 8225 -6200 8255 -5700
rect 8321 -6200 8351 -5700
rect 8417 -6200 8447 -5700
rect 8513 -6200 8543 -5700
rect 8609 -6200 8639 -5700
rect 8705 -6200 8735 -5700
rect 8801 -6200 8831 -5700
rect 8897 -6200 8927 -5700
<< ndiff >>
rect 5847 9764 5905 9776
rect 5847 7788 5859 9764
rect 5893 7788 5905 9764
rect 5847 7776 5905 7788
rect 5965 9764 6023 9776
rect 5965 7788 5977 9764
rect 6011 7788 6023 9764
rect 5965 7776 6023 7788
rect 6083 9764 6141 9776
rect 6083 7788 6095 9764
rect 6129 7788 6141 9764
rect 6083 7776 6141 7788
rect 6201 9764 6259 9776
rect 6201 7788 6213 9764
rect 6247 7788 6259 9764
rect 6201 7776 6259 7788
rect 6319 9764 6377 9776
rect 6319 7788 6331 9764
rect 6365 7788 6377 9764
rect 6319 7776 6377 7788
rect 6437 9764 6495 9776
rect 6437 7788 6449 9764
rect 6483 7788 6495 9764
rect 6437 7776 6495 7788
rect 6555 9764 6613 9776
rect 6555 7788 6567 9764
rect 6601 7788 6613 9764
rect 6555 7776 6613 7788
rect 7011 9588 7073 9600
rect 7011 9112 7023 9588
rect 7057 9112 7073 9588
rect 7011 9100 7073 9112
rect 7103 9588 7169 9600
rect 7103 9112 7119 9588
rect 7153 9112 7169 9588
rect 7103 9100 7169 9112
rect 7199 9588 7265 9600
rect 7199 9112 7215 9588
rect 7249 9112 7265 9588
rect 7199 9100 7265 9112
rect 7295 9588 7361 9600
rect 7295 9112 7311 9588
rect 7345 9112 7361 9588
rect 7295 9100 7361 9112
rect 7391 9588 7457 9600
rect 7391 9112 7407 9588
rect 7441 9112 7457 9588
rect 7391 9100 7457 9112
rect 7487 9588 7553 9600
rect 7487 9112 7503 9588
rect 7537 9112 7553 9588
rect 7487 9100 7553 9112
rect 7583 9588 7649 9600
rect 7583 9112 7599 9588
rect 7633 9112 7649 9588
rect 7583 9100 7649 9112
rect 7679 9588 7745 9600
rect 7679 9112 7695 9588
rect 7729 9112 7745 9588
rect 7679 9100 7745 9112
rect 7775 9588 7841 9600
rect 7775 9112 7791 9588
rect 7825 9112 7841 9588
rect 7775 9100 7841 9112
rect 7871 9588 7937 9600
rect 7871 9112 7887 9588
rect 7921 9112 7937 9588
rect 7871 9100 7937 9112
rect 7967 9588 8033 9600
rect 7967 9112 7983 9588
rect 8017 9112 8033 9588
rect 7967 9100 8033 9112
rect 8063 9588 8129 9600
rect 8063 9112 8079 9588
rect 8113 9112 8129 9588
rect 8063 9100 8129 9112
rect 8159 9588 8225 9600
rect 8159 9112 8175 9588
rect 8209 9112 8225 9588
rect 8159 9100 8225 9112
rect 8255 9588 8321 9600
rect 8255 9112 8271 9588
rect 8305 9112 8321 9588
rect 8255 9100 8321 9112
rect 8351 9588 8417 9600
rect 8351 9112 8367 9588
rect 8401 9112 8417 9588
rect 8351 9100 8417 9112
rect 8447 9588 8513 9600
rect 8447 9112 8463 9588
rect 8497 9112 8513 9588
rect 8447 9100 8513 9112
rect 8543 9588 8609 9600
rect 8543 9112 8559 9588
rect 8593 9112 8609 9588
rect 8543 9100 8609 9112
rect 8639 9588 8705 9600
rect 8639 9112 8655 9588
rect 8689 9112 8705 9588
rect 8639 9100 8705 9112
rect 8735 9588 8801 9600
rect 8735 9112 8751 9588
rect 8785 9112 8801 9588
rect 8735 9100 8801 9112
rect 8831 9588 8897 9600
rect 8831 9112 8847 9588
rect 8881 9112 8897 9588
rect 8831 9100 8897 9112
rect 8927 9588 8989 9600
rect 8927 9112 8943 9588
rect 8977 9112 8989 9588
rect 8927 9100 8989 9112
rect 7055 8648 7113 8660
rect 7055 6672 7067 8648
rect 7101 6672 7113 8648
rect 7055 6660 7113 6672
rect 7513 8648 7571 8660
rect 7513 6672 7525 8648
rect 7559 6672 7571 8648
rect 7513 6660 7571 6672
rect 7971 8648 8029 8660
rect 7971 6672 7983 8648
rect 8017 6672 8029 8648
rect 7971 6660 8029 6672
rect 8429 8648 8487 8660
rect 8429 6672 8441 8648
rect 8475 6672 8487 8648
rect 8429 6660 8487 6672
rect 8887 8648 8945 8660
rect 8887 6672 8899 8648
rect 8933 6672 8945 8648
rect 8887 6660 8945 6672
rect 9388 9764 9446 9776
rect 9388 7788 9400 9764
rect 9434 7788 9446 9764
rect 9388 7776 9446 7788
rect 9506 9764 9564 9776
rect 9506 7788 9518 9764
rect 9552 7788 9564 9764
rect 9506 7776 9564 7788
rect 9624 9764 9682 9776
rect 9624 7788 9636 9764
rect 9670 7788 9682 9764
rect 9624 7776 9682 7788
rect 9742 9764 9800 9776
rect 9742 7788 9754 9764
rect 9788 7788 9800 9764
rect 9742 7776 9800 7788
rect 9860 9764 9918 9776
rect 9860 7788 9872 9764
rect 9906 7788 9918 9764
rect 9860 7776 9918 7788
rect 9978 9764 10036 9776
rect 9978 7788 9990 9764
rect 10024 7788 10036 9764
rect 9978 7776 10036 7788
rect 10096 9764 10154 9776
rect 10096 7788 10108 9764
rect 10142 7788 10154 9764
rect 10096 7776 10154 7788
rect 10852 7302 11352 7314
rect 10852 7268 10864 7302
rect 11340 7268 11352 7302
rect 10852 7252 11352 7268
rect 10852 7206 11352 7222
rect 10852 7172 10864 7206
rect 11340 7172 11352 7206
rect 10852 7156 11352 7172
rect 10852 7110 11352 7126
rect 10852 7076 10864 7110
rect 11340 7076 11352 7110
rect 10852 7060 11352 7076
rect 10852 7014 11352 7030
rect 10852 6980 10864 7014
rect 11340 6980 11352 7014
rect 10852 6964 11352 6980
rect 10852 6918 11352 6934
rect 10852 6884 10864 6918
rect 11340 6884 11352 6918
rect 10852 6872 11352 6884
rect 3457 4340 3515 4352
rect 3457 3964 3469 4340
rect 3503 3964 3515 4340
rect 3457 3952 3515 3964
rect 3545 4340 3603 4352
rect 3545 3964 3557 4340
rect 3591 3964 3603 4340
rect 3545 3952 3603 3964
rect 3457 3626 3515 3638
rect 3457 3250 3469 3626
rect 3503 3250 3515 3626
rect 3457 3238 3515 3250
rect 3545 3626 3603 3638
rect 3545 3250 3557 3626
rect 3591 3250 3603 3626
rect 3545 3238 3603 3250
rect 4239 4340 4297 4352
rect 4239 3964 4251 4340
rect 4285 3964 4297 4340
rect 4239 3952 4297 3964
rect 4327 4340 4385 4352
rect 4327 3964 4339 4340
rect 4373 3964 4385 4340
rect 4327 3952 4385 3964
rect 4239 3626 4297 3638
rect 4239 3250 4251 3626
rect 4285 3250 4297 3626
rect 4239 3238 4297 3250
rect 4327 3626 4385 3638
rect 4327 3250 4339 3626
rect 4373 3250 4385 3626
rect 4327 3238 4385 3250
rect 2428 2422 2499 2434
rect 2428 2388 2440 2422
rect 2474 2388 2499 2422
rect 2428 2332 2499 2388
rect 2428 2298 2440 2332
rect 2474 2298 2499 2332
rect 2428 2286 2499 2298
rect 2529 2422 2586 2434
rect 2529 2388 2540 2422
rect 2574 2388 2586 2422
rect 2529 2332 2586 2388
rect 3797 2414 3854 2434
rect 3797 2380 3809 2414
rect 3843 2380 3854 2414
rect 2529 2298 2540 2332
rect 2574 2298 2586 2332
rect 2529 2286 2586 2298
rect 3797 2332 3854 2380
rect 3797 2298 3809 2332
rect 3843 2298 3854 2332
rect 3797 2286 3854 2298
rect 3884 2286 3932 2434
rect 3962 2414 4019 2434
rect 3962 2380 3973 2414
rect 4007 2380 4019 2414
rect 3962 2332 4019 2380
rect 3962 2298 3973 2332
rect 4007 2298 4019 2332
rect 3962 2286 4019 2298
rect 4097 2357 4150 2381
rect 4097 2323 4105 2357
rect 4139 2323 4150 2357
rect 4097 2297 4150 2323
rect 4350 2357 4406 2381
rect 4350 2323 4361 2357
rect 4395 2323 4406 2357
rect 4350 2297 4406 2323
rect 4606 2357 4662 2381
rect 4606 2323 4617 2357
rect 4651 2323 4662 2357
rect 4606 2297 4662 2323
rect 5441 2357 5494 2381
rect 5441 2323 5449 2357
rect 5483 2323 5494 2357
rect 5441 2297 5494 2323
rect 5694 2357 5750 2381
rect 5694 2323 5705 2357
rect 5739 2323 5750 2357
rect 5694 2297 5750 2323
rect 5950 2357 6006 2381
rect 5950 2323 5961 2357
rect 5995 2323 6006 2357
rect 5950 2297 6006 2323
rect 6113 2357 6166 2381
rect 6113 2323 6121 2357
rect 6155 2323 6166 2357
rect 6113 2297 6166 2323
rect 6366 2357 6422 2381
rect 6366 2323 6377 2357
rect 6411 2323 6422 2357
rect 6366 2297 6422 2323
rect 6622 2357 6678 2381
rect 6622 2323 6633 2357
rect 6667 2323 6678 2357
rect 6622 2297 6678 2323
rect 6785 2357 6838 2381
rect 6785 2323 6793 2357
rect 6827 2323 6838 2357
rect 6785 2297 6838 2323
rect 7038 2357 7094 2381
rect 7038 2323 7049 2357
rect 7083 2323 7094 2357
rect 7038 2297 7094 2323
rect 7294 2357 7350 2381
rect 7294 2323 7305 2357
rect 7339 2323 7350 2357
rect 7294 2297 7350 2323
rect 8129 2357 8182 2381
rect 8129 2323 8137 2357
rect 8171 2323 8182 2357
rect 8129 2297 8182 2323
rect 8382 2357 8438 2381
rect 8382 2323 8393 2357
rect 8427 2323 8438 2357
rect 8382 2297 8438 2323
rect 8638 2357 8694 2381
rect 8638 2323 8649 2357
rect 8683 2323 8694 2357
rect 8638 2297 8694 2323
rect 8801 2357 8854 2381
rect 8801 2323 8809 2357
rect 8843 2323 8854 2357
rect 8801 2297 8854 2323
rect 9054 2357 9110 2381
rect 9054 2323 9065 2357
rect 9099 2323 9110 2357
rect 9054 2297 9110 2323
rect 9310 2357 9366 2381
rect 9310 2323 9321 2357
rect 9355 2323 9366 2357
rect 9310 2297 9366 2323
rect 9473 2357 9526 2381
rect 9473 2323 9481 2357
rect 9515 2323 9526 2357
rect 9473 2297 9526 2323
rect 9726 2357 9783 2381
rect 9726 2323 9737 2357
rect 9771 2323 9783 2357
rect 9726 2297 9783 2323
rect 2428 2126 2499 2138
rect 2428 2092 2440 2126
rect 2474 2092 2499 2126
rect 2428 2036 2499 2092
rect 2428 2002 2440 2036
rect 2474 2002 2499 2036
rect 2428 1990 2499 2002
rect 2529 2126 2586 2138
rect 2529 2092 2540 2126
rect 2574 2092 2586 2126
rect 2529 2036 2586 2092
rect 3797 2126 3854 2138
rect 3797 2092 3809 2126
rect 3843 2092 3854 2126
rect 2529 2002 2540 2036
rect 2574 2002 2586 2036
rect 2529 1990 2586 2002
rect 3797 2044 3854 2092
rect 3797 2010 3809 2044
rect 3843 2010 3854 2044
rect 3797 1990 3854 2010
rect 3884 1990 3932 2138
rect 3962 2126 4019 2138
rect 4184 2126 4251 2138
rect 3962 2092 3973 2126
rect 4007 2092 4019 2126
rect 4184 2100 4201 2126
rect 3962 2044 4019 2092
rect 3962 2010 3973 2044
rect 4007 2010 4019 2044
rect 3962 1990 4019 2010
rect 4082 2062 4139 2100
rect 4082 2028 4094 2062
rect 4128 2028 4139 2062
rect 4082 1990 4139 2028
rect 4169 2092 4201 2100
rect 4235 2092 4251 2126
rect 4169 2036 4251 2092
rect 4169 2002 4183 2036
rect 4217 2002 4251 2036
rect 4169 1990 4251 2002
rect 4281 1990 4329 2138
rect 4359 2118 4468 2138
rect 4359 2084 4396 2118
rect 4430 2084 4468 2118
rect 4359 1990 4468 2084
rect 4498 1990 4660 2138
rect 4690 2100 4803 2138
rect 4690 2066 4730 2100
rect 4764 2066 4803 2100
rect 4690 1990 4803 2066
rect 4833 2126 4890 2138
rect 4833 2092 4844 2126
rect 4878 2092 4890 2126
rect 4833 2036 4890 2092
rect 4833 2002 4844 2036
rect 4878 2002 4890 2036
rect 4833 1990 4890 2002
rect 4949 2126 5006 2138
rect 4949 2092 4961 2126
rect 4995 2092 5006 2126
rect 4949 2036 5006 2092
rect 4949 2002 4961 2036
rect 4995 2002 5006 2036
rect 4949 1990 5006 2002
rect 5036 2126 5092 2138
rect 5036 2092 5047 2126
rect 5081 2092 5092 2126
rect 5036 2036 5092 2092
rect 5036 2002 5047 2036
rect 5081 2002 5092 2036
rect 5036 1990 5092 2002
rect 5122 2126 5179 2138
rect 5122 2092 5133 2126
rect 5167 2092 5179 2126
rect 5122 2036 5179 2092
rect 5122 2002 5133 2036
rect 5167 2002 5179 2036
rect 5122 1990 5179 2002
rect 6189 2164 6247 2176
rect 6189 2130 6201 2164
rect 6235 2130 6247 2164
rect 6189 2114 6247 2130
rect 6477 2128 6539 2140
rect 5431 2076 5488 2093
rect 5431 2042 5443 2076
rect 5477 2042 5488 2076
rect 5431 2009 5488 2042
rect 5518 2009 5566 2093
rect 5596 2071 5732 2093
rect 5596 2037 5607 2071
rect 5641 2037 5687 2071
rect 5721 2037 5732 2071
rect 5596 2009 5732 2037
rect 5762 2009 5810 2093
rect 5840 2077 5946 2093
rect 5840 2043 5851 2077
rect 5885 2043 5946 2077
rect 5840 2009 5946 2043
rect 5976 2066 6033 2093
rect 5976 2032 5987 2066
rect 6021 2032 6033 2066
rect 5976 2009 6033 2032
rect 6087 2012 6144 2114
rect 6087 1978 6099 2012
rect 6133 1978 6144 2012
rect 6087 1966 6144 1978
rect 6174 1966 6312 2114
rect 6342 2077 6399 2114
rect 6342 2043 6353 2077
rect 6387 2043 6399 2077
rect 6342 2009 6399 2043
rect 6342 1975 6353 2009
rect 6387 1975 6399 2009
rect 6477 2094 6491 2128
rect 6525 2094 6539 2128
rect 6477 2087 6539 2094
rect 6872 2127 6949 2139
rect 7739 2160 7806 2172
rect 7739 2130 7755 2160
rect 6872 2093 6893 2127
rect 6927 2093 6949 2127
rect 6872 2087 6949 2093
rect 7316 2087 7366 2130
rect 6477 2003 6554 2087
rect 6584 2003 6626 2087
rect 6656 2062 6717 2087
rect 6656 2028 6672 2062
rect 6706 2028 6717 2062
rect 6656 2003 6717 2028
rect 6747 2067 6818 2087
rect 6747 2033 6772 2067
rect 6806 2033 6818 2067
rect 6747 2003 6818 2033
rect 6342 1966 6399 1975
rect 6872 1977 6964 2087
rect 6994 2057 7050 2087
rect 6994 2023 7005 2057
rect 7039 2023 7050 2057
rect 6994 1977 7050 2023
rect 7080 2075 7171 2087
rect 7080 2041 7115 2075
rect 7149 2041 7171 2075
rect 7080 1977 7171 2041
rect 7201 2075 7271 2087
rect 7201 2041 7226 2075
rect 7260 2041 7271 2075
rect 7201 1977 7271 2041
rect 7301 2020 7366 2087
rect 7396 2092 7616 2130
rect 7396 2058 7407 2092
rect 7441 2058 7489 2092
rect 7523 2058 7571 2092
rect 7605 2058 7616 2092
rect 7396 2046 7616 2058
rect 7646 2046 7694 2130
rect 7724 2126 7755 2130
rect 7789 2138 7806 2160
rect 8056 2147 8114 2159
rect 8056 2138 8068 2147
rect 7789 2126 7821 2138
rect 7724 2046 7821 2126
rect 7396 2020 7446 2046
rect 7301 1977 7351 2020
rect 7771 1990 7821 2046
rect 7851 2126 7925 2138
rect 7851 2092 7871 2126
rect 7905 2092 7925 2126
rect 7851 1990 7925 2092
rect 7955 2074 8011 2138
rect 7955 2040 7966 2074
rect 8000 2040 8011 2074
rect 7955 1990 8011 2040
rect 8041 2113 8068 2138
rect 8102 2113 8114 2147
rect 8041 1990 8114 2113
rect 8377 2126 8430 2138
rect 8377 2092 8385 2126
rect 8419 2092 8430 2126
rect 8377 2036 8430 2092
rect 8377 2032 8385 2036
rect 8168 1995 8224 2032
rect 8168 1961 8179 1995
rect 8213 1961 8224 1995
rect 8168 1948 8224 1961
rect 8254 2002 8385 2032
rect 8419 2002 8430 2036
rect 8254 1990 8430 2002
rect 8460 2126 8516 2138
rect 8460 2092 8471 2126
rect 8505 2092 8516 2126
rect 8460 2036 8516 2092
rect 8460 2002 8471 2036
rect 8505 2002 8516 2036
rect 8460 1990 8516 2002
rect 8546 2126 8608 2138
rect 8546 2092 8557 2126
rect 8591 2092 8608 2126
rect 8777 2126 8848 2138
rect 8777 2118 8789 2126
rect 8546 2036 8608 2092
rect 8546 2002 8557 2036
rect 8591 2002 8608 2036
rect 8546 1990 8608 2002
rect 8671 2100 8728 2118
rect 8671 2066 8683 2100
rect 8717 2066 8728 2100
rect 8671 2032 8728 2066
rect 8671 1998 8683 2032
rect 8717 1998 8728 2032
rect 8671 1990 8728 1998
rect 8758 2092 8789 2118
rect 8823 2092 8848 2126
rect 8758 2052 8848 2092
rect 8758 2018 8789 2052
rect 8823 2018 8848 2052
rect 8758 1990 8848 2018
rect 8878 2126 8934 2138
rect 8878 2092 8889 2126
rect 8923 2092 8934 2126
rect 8878 2052 8934 2092
rect 8878 2018 8889 2052
rect 8923 2018 8934 2052
rect 8878 1990 8934 2018
rect 8964 2126 9020 2138
rect 8964 2092 8975 2126
rect 9009 2092 9020 2126
rect 8964 2036 9020 2092
rect 8964 2002 8975 2036
rect 9009 2002 9020 2036
rect 8964 1990 9020 2002
rect 9074 2130 9212 2138
rect 9074 2096 9090 2130
rect 9124 2096 9162 2130
rect 9196 2096 9212 2130
rect 9074 1990 9212 2096
rect 9266 2126 9323 2138
rect 9266 2092 9278 2126
rect 9312 2092 9323 2126
rect 9266 2036 9323 2092
rect 9266 2002 9278 2036
rect 9312 2002 9323 2036
rect 9266 1990 9323 2002
rect 9353 2104 9409 2138
rect 9353 2070 9364 2104
rect 9398 2070 9409 2104
rect 9353 1990 9409 2070
rect 9439 2126 9495 2138
rect 9439 2092 9450 2126
rect 9484 2092 9495 2126
rect 9439 2036 9495 2092
rect 9439 2002 9450 2036
rect 9484 2002 9495 2036
rect 9439 1990 9495 2002
rect 9525 2104 9581 2138
rect 9525 2070 9536 2104
rect 9570 2070 9581 2104
rect 9525 1990 9581 2070
rect 9611 2126 9675 2138
rect 9611 2092 9622 2126
rect 9656 2092 9675 2126
rect 9611 2036 9675 2092
rect 9611 2002 9622 2036
rect 9656 2002 9675 2036
rect 9611 1990 9675 2002
rect 9705 2072 9767 2138
rect 9705 2038 9722 2072
rect 9756 2038 9767 2072
rect 9705 1990 9767 2038
rect 9797 2104 9867 2138
rect 9797 2070 9822 2104
rect 9856 2070 9867 2104
rect 9797 1990 9867 2070
rect 9897 2072 9980 2138
rect 9897 2038 9926 2072
rect 9960 2038 9980 2072
rect 9897 1990 9980 2038
rect 10010 2104 10076 2138
rect 10010 2070 10030 2104
rect 10064 2070 10076 2104
rect 10010 1990 10076 2070
rect 8254 1948 8304 1990
rect 3580 1090 3651 1102
rect 3580 1056 3592 1090
rect 3626 1056 3651 1090
rect 3580 1000 3651 1056
rect 3580 966 3592 1000
rect 3626 966 3651 1000
rect 3580 954 3651 966
rect 3681 1090 3738 1102
rect 3681 1056 3692 1090
rect 3726 1056 3738 1090
rect 3681 1000 3738 1056
rect 4949 1082 5006 1102
rect 4949 1048 4961 1082
rect 4995 1048 5006 1082
rect 3681 966 3692 1000
rect 3726 966 3738 1000
rect 3681 954 3738 966
rect 4949 1000 5006 1048
rect 4949 966 4961 1000
rect 4995 966 5006 1000
rect 4949 954 5006 966
rect 5036 954 5084 1102
rect 5114 1082 5171 1102
rect 5114 1048 5125 1082
rect 5159 1048 5171 1082
rect 5114 1000 5171 1048
rect 5114 966 5125 1000
rect 5159 966 5171 1000
rect 5114 954 5171 966
rect 6087 1114 6144 1126
rect 5431 1050 5488 1083
rect 5431 1016 5443 1050
rect 5477 1016 5488 1050
rect 5431 999 5488 1016
rect 5518 999 5566 1083
rect 5596 1055 5732 1083
rect 5596 1021 5607 1055
rect 5641 1021 5687 1055
rect 5721 1021 5732 1055
rect 5596 999 5732 1021
rect 5762 999 5810 1083
rect 5840 1049 5946 1083
rect 5840 1015 5851 1049
rect 5885 1015 5946 1049
rect 5840 999 5946 1015
rect 5976 1060 6033 1083
rect 5976 1026 5987 1060
rect 6021 1026 6033 1060
rect 5976 999 6033 1026
rect 6087 1080 6099 1114
rect 6133 1080 6144 1114
rect 6087 978 6144 1080
rect 6174 978 6312 1126
rect 6342 1117 6399 1126
rect 6342 1083 6353 1117
rect 6387 1083 6399 1117
rect 6342 1049 6399 1083
rect 6342 1015 6353 1049
rect 6387 1015 6399 1049
rect 6342 978 6399 1015
rect 6477 1005 6554 1089
rect 6584 1005 6626 1089
rect 6656 1064 6717 1089
rect 6656 1030 6672 1064
rect 6706 1030 6717 1064
rect 6656 1005 6717 1030
rect 6747 1059 6818 1089
rect 6747 1025 6772 1059
rect 6806 1025 6818 1059
rect 6747 1005 6818 1025
rect 6872 1005 6964 1115
rect 6994 1069 7050 1115
rect 6994 1035 7005 1069
rect 7039 1035 7050 1069
rect 6994 1005 7050 1035
rect 7080 1051 7171 1115
rect 7080 1017 7115 1051
rect 7149 1017 7171 1051
rect 7080 1005 7171 1017
rect 7201 1051 7271 1115
rect 7201 1017 7226 1051
rect 7260 1017 7271 1051
rect 7201 1005 7271 1017
rect 7301 1072 7351 1115
rect 7301 1005 7366 1072
rect 6477 998 6539 1005
rect 6189 962 6247 978
rect 6189 928 6201 962
rect 6235 928 6247 962
rect 6189 916 6247 928
rect 6477 964 6491 998
rect 6525 964 6539 998
rect 6477 952 6539 964
rect 6872 999 6949 1005
rect 6872 965 6893 999
rect 6927 965 6949 999
rect 6872 953 6949 965
rect 7316 962 7366 1005
rect 7396 1046 7446 1072
rect 8168 1131 8224 1144
rect 7771 1046 7821 1102
rect 7396 1034 7616 1046
rect 7396 1000 7407 1034
rect 7441 1000 7489 1034
rect 7523 1000 7571 1034
rect 7605 1000 7616 1034
rect 7396 962 7616 1000
rect 7646 962 7694 1046
rect 7724 966 7821 1046
rect 7724 962 7755 966
rect 7739 932 7755 962
rect 7789 954 7821 966
rect 7851 1000 7925 1102
rect 7851 966 7871 1000
rect 7905 966 7925 1000
rect 7851 954 7925 966
rect 7955 1052 8011 1102
rect 7955 1018 7966 1052
rect 8000 1018 8011 1052
rect 7955 954 8011 1018
rect 8041 979 8114 1102
rect 8168 1097 8179 1131
rect 8213 1097 8224 1131
rect 8168 1060 8224 1097
rect 8254 1102 8304 1144
rect 9266 1115 9323 1127
rect 8254 1090 8430 1102
rect 8254 1060 8385 1090
rect 8377 1056 8385 1060
rect 8419 1056 8430 1090
rect 8041 954 8068 979
rect 7789 932 7806 954
rect 7739 920 7806 932
rect 8056 945 8068 954
rect 8102 945 8114 979
rect 8377 1000 8430 1056
rect 8377 966 8385 1000
rect 8419 966 8430 1000
rect 8377 954 8430 966
rect 8460 1090 8516 1102
rect 8460 1056 8471 1090
rect 8505 1056 8516 1090
rect 8460 1000 8516 1056
rect 8460 966 8471 1000
rect 8505 966 8516 1000
rect 8460 954 8516 966
rect 8546 1090 8608 1102
rect 8546 1056 8557 1090
rect 8591 1056 8608 1090
rect 8546 1000 8608 1056
rect 8546 966 8557 1000
rect 8591 966 8608 1000
rect 8671 1094 8728 1102
rect 8671 1060 8683 1094
rect 8717 1060 8728 1094
rect 8671 1026 8728 1060
rect 8671 992 8683 1026
rect 8717 992 8728 1026
rect 8671 974 8728 992
rect 8758 1074 8848 1102
rect 8758 1040 8789 1074
rect 8823 1040 8848 1074
rect 8758 1000 8848 1040
rect 8758 974 8789 1000
rect 8546 954 8608 966
rect 8056 933 8114 945
rect 8777 966 8789 974
rect 8823 966 8848 1000
rect 8777 954 8848 966
rect 8878 1074 8934 1102
rect 8878 1040 8889 1074
rect 8923 1040 8934 1074
rect 8878 1000 8934 1040
rect 8878 966 8889 1000
rect 8923 966 8934 1000
rect 8878 954 8934 966
rect 8964 1090 9020 1102
rect 8964 1056 8975 1090
rect 9009 1056 9020 1090
rect 8964 1000 9020 1056
rect 8964 966 8975 1000
rect 9009 966 9020 1000
rect 8964 954 9020 966
rect 9074 996 9212 1102
rect 9266 1081 9278 1115
rect 9312 1081 9323 1115
rect 9266 1045 9323 1081
rect 9266 1011 9278 1045
rect 9312 1011 9323 1045
rect 9266 999 9323 1011
rect 9353 1048 9413 1127
rect 9353 1014 9368 1048
rect 9402 1014 9413 1048
rect 9353 999 9413 1014
rect 9443 1119 9508 1127
rect 9443 1085 9454 1119
rect 9488 1085 9508 1119
rect 9443 1041 9508 1085
rect 9443 1007 9454 1041
rect 9488 1007 9508 1041
rect 9443 999 9508 1007
rect 9538 1109 9599 1127
rect 9538 1075 9554 1109
rect 9588 1075 9599 1109
rect 9538 1041 9599 1075
rect 9538 1007 9554 1041
rect 9588 1007 9599 1041
rect 9538 999 9599 1007
rect 9629 1115 9701 1127
rect 9629 1081 9656 1115
rect 9690 1081 9701 1115
rect 9629 1037 9701 1081
rect 9629 1003 9656 1037
rect 9690 1003 9701 1037
rect 9629 999 9701 1003
rect 9074 962 9090 996
rect 9124 962 9162 996
rect 9196 962 9212 996
rect 9074 954 9212 962
rect 9644 979 9701 999
rect 9731 1099 9817 1127
rect 9731 1065 9758 1099
rect 9792 1065 9817 1099
rect 9731 1025 9817 1065
rect 9731 991 9758 1025
rect 9792 991 9817 1025
rect 9731 979 9817 991
rect 9847 1031 9903 1127
rect 9847 997 9858 1031
rect 9892 997 9903 1031
rect 9847 979 9903 997
rect 9933 1115 9989 1127
rect 9933 1081 9944 1115
rect 9978 1081 9989 1115
rect 9933 1025 9989 1081
rect 9933 991 9944 1025
rect 9978 991 9989 1025
rect 9933 979 9989 991
rect 10019 1115 10076 1127
rect 10019 1081 10030 1115
rect 10064 1081 10076 1115
rect 10019 1025 10076 1081
rect 10019 991 10030 1025
rect 10064 991 10076 1025
rect 10019 979 10076 991
rect 3806 570 3864 582
rect 3806 194 3818 570
rect 3852 194 3864 570
rect 3806 182 3864 194
rect 3894 570 3952 582
rect 3894 194 3906 570
rect 3940 194 3952 570
rect 3894 182 3952 194
rect 10446 1296 10504 1308
rect 10446 320 10458 1296
rect 10492 320 10504 1296
rect 10446 308 10504 320
rect 10904 1296 10962 1308
rect 10904 320 10916 1296
rect 10950 320 10962 1296
rect 10904 308 10962 320
rect 11362 1296 11420 1308
rect 11362 320 11374 1296
rect 11408 320 11420 1296
rect 11362 308 11420 320
rect 11820 1296 11878 1308
rect 11820 320 11832 1296
rect 11866 320 11878 1296
rect 11820 308 11878 320
rect 12278 1296 12336 1308
rect 12278 320 12290 1296
rect 12324 320 12336 1296
rect 12278 308 12336 320
rect 12736 1296 12794 1308
rect 12736 320 12748 1296
rect 12782 320 12794 1296
rect 12736 308 12794 320
rect 13194 1296 13252 1308
rect 13194 320 13206 1296
rect 13240 320 13252 1296
rect 13194 308 13252 320
rect 13652 1296 13710 1308
rect 13652 320 13664 1296
rect 13698 320 13710 1296
rect 13652 308 13710 320
rect 13880 1296 13938 1308
rect 13880 320 13892 1296
rect 13926 320 13938 1296
rect 13880 308 13938 320
rect 13968 1296 14026 1308
rect 13968 320 13980 1296
rect 14014 320 14026 1296
rect 13968 308 14026 320
rect 14196 1296 14254 1308
rect 14196 320 14208 1296
rect 14242 320 14254 1296
rect 14196 308 14254 320
rect 14284 1296 14342 1308
rect 14284 320 14296 1296
rect 14330 320 14342 1296
rect 14284 308 14342 320
rect 15540 901 15940 913
rect 15540 867 15552 901
rect 15928 867 15940 901
rect 15540 855 15940 867
rect 15540 813 15940 825
rect 15540 779 15552 813
rect 15928 779 15940 813
rect 15540 767 15940 779
rect 16254 901 16654 913
rect 16254 867 16266 901
rect 16642 867 16654 901
rect 16254 855 16654 867
rect 16254 813 16654 825
rect 16254 779 16266 813
rect 16642 779 16654 813
rect 16254 767 16654 779
rect 16968 901 17368 913
rect 16968 867 16980 901
rect 17356 867 17368 901
rect 16968 855 17368 867
rect 16968 813 17368 825
rect 16968 779 16980 813
rect 17356 779 17368 813
rect 16968 767 17368 779
rect 17682 901 18082 913
rect 17682 867 17694 901
rect 18070 867 18082 901
rect 17682 855 18082 867
rect 17682 813 18082 825
rect 17682 779 17694 813
rect 18070 779 18082 813
rect 17682 767 18082 779
rect 18396 901 18796 913
rect 18396 867 18408 901
rect 18784 867 18796 901
rect 18396 855 18796 867
rect 18396 813 18796 825
rect 18396 779 18408 813
rect 18784 779 18796 813
rect 18396 767 18796 779
rect 19110 901 19510 913
rect 19110 867 19122 901
rect 19498 867 19510 901
rect 19110 855 19510 867
rect 19110 813 19510 825
rect 19110 779 19122 813
rect 19498 779 19510 813
rect 19110 767 19510 779
rect 19824 901 20224 913
rect 19824 867 19836 901
rect 20212 867 20224 901
rect 19824 855 20224 867
rect 19824 813 20224 825
rect 19824 779 19836 813
rect 20212 779 20224 813
rect 19824 767 20224 779
rect 20538 901 20938 913
rect 20538 867 20550 901
rect 20926 867 20938 901
rect 20538 855 20938 867
rect 20538 813 20938 825
rect 20538 779 20550 813
rect 20926 779 20938 813
rect 20538 767 20938 779
rect 21252 901 21652 913
rect 21252 867 21264 901
rect 21640 867 21652 901
rect 21252 855 21652 867
rect 21252 813 21652 825
rect 21252 779 21264 813
rect 21640 779 21652 813
rect 21252 767 21652 779
rect 21966 901 22366 913
rect 21966 867 21978 901
rect 22354 867 22366 901
rect 21966 855 22366 867
rect 21966 813 22366 825
rect 21966 779 21978 813
rect 22354 779 22366 813
rect 21966 767 22366 779
rect 22680 901 23080 913
rect 22680 867 22692 901
rect 23068 867 23080 901
rect 22680 855 23080 867
rect 22680 813 23080 825
rect 22680 779 22692 813
rect 23068 779 23080 813
rect 22680 767 23080 779
rect 23394 901 23794 913
rect 23394 867 23406 901
rect 23782 867 23794 901
rect 23394 855 23794 867
rect 23394 813 23794 825
rect 23394 779 23406 813
rect 23782 779 23794 813
rect 23394 767 23794 779
rect 24108 901 24508 913
rect 24108 867 24120 901
rect 24496 867 24508 901
rect 24108 855 24508 867
rect 24108 813 24508 825
rect 24108 779 24120 813
rect 24496 779 24508 813
rect 24108 767 24508 779
rect 24822 901 25222 913
rect 24822 867 24834 901
rect 25210 867 25222 901
rect 24822 855 25222 867
rect 24822 813 25222 825
rect 24822 779 24834 813
rect 25210 779 25222 813
rect 24822 767 25222 779
rect 25536 901 25936 913
rect 25536 867 25548 901
rect 25924 867 25936 901
rect 25536 855 25936 867
rect 25536 813 25936 825
rect 25536 779 25548 813
rect 25924 779 25936 813
rect 25536 767 25936 779
rect 26250 901 26650 913
rect 26250 867 26262 901
rect 26638 867 26650 901
rect 26250 855 26650 867
rect 26250 813 26650 825
rect 26250 779 26262 813
rect 26638 779 26650 813
rect 26250 767 26650 779
rect 26964 901 27364 913
rect 26964 867 26976 901
rect 27352 867 27364 901
rect 26964 855 27364 867
rect 26964 813 27364 825
rect 26964 779 26976 813
rect 27352 779 27364 813
rect 26964 767 27364 779
rect 27678 901 28078 913
rect 27678 867 27690 901
rect 28066 867 28078 901
rect 27678 855 28078 867
rect 27678 813 28078 825
rect 27678 779 27690 813
rect 28066 779 28078 813
rect 27678 767 28078 779
rect 28392 901 28792 913
rect 28392 867 28404 901
rect 28780 867 28792 901
rect 28392 855 28792 867
rect 28392 813 28792 825
rect 28392 779 28404 813
rect 28780 779 28792 813
rect 28392 767 28792 779
rect 29106 901 29506 913
rect 29106 867 29118 901
rect 29494 867 29506 901
rect 29106 855 29506 867
rect 29106 813 29506 825
rect 29106 779 29118 813
rect 29494 779 29506 813
rect 29106 767 29506 779
rect 29820 901 30220 913
rect 29820 867 29832 901
rect 30208 867 30220 901
rect 29820 855 30220 867
rect 29820 813 30220 825
rect 29820 779 29832 813
rect 30208 779 30220 813
rect 29820 767 30220 779
rect 30534 901 30934 913
rect 30534 867 30546 901
rect 30922 867 30934 901
rect 30534 855 30934 867
rect 30534 813 30934 825
rect 30534 779 30546 813
rect 30922 779 30934 813
rect 30534 767 30934 779
rect 31248 901 31648 913
rect 31248 867 31260 901
rect 31636 867 31648 901
rect 31248 855 31648 867
rect 31248 813 31648 825
rect 31248 779 31260 813
rect 31636 779 31648 813
rect 31248 767 31648 779
rect 31962 901 32362 913
rect 31962 867 31974 901
rect 32350 867 32362 901
rect 31962 855 32362 867
rect 31962 813 32362 825
rect 31962 779 31974 813
rect 32350 779 32362 813
rect 31962 767 32362 779
rect 32676 901 33076 913
rect 32676 867 32688 901
rect 33064 867 33076 901
rect 32676 855 33076 867
rect 32676 813 33076 825
rect 32676 779 32688 813
rect 33064 779 33076 813
rect 32676 767 33076 779
rect 33390 901 33790 913
rect 33390 867 33402 901
rect 33778 867 33790 901
rect 33390 855 33790 867
rect 33390 813 33790 825
rect 33390 779 33402 813
rect 33778 779 33790 813
rect 33390 767 33790 779
rect 34104 901 34504 913
rect 34104 867 34116 901
rect 34492 867 34504 901
rect 34104 855 34504 867
rect 34104 813 34504 825
rect 34104 779 34116 813
rect 34492 779 34504 813
rect 34104 767 34504 779
rect 34818 901 35218 913
rect 34818 867 34830 901
rect 35206 867 35218 901
rect 34818 855 35218 867
rect 34818 813 35218 825
rect 34818 779 34830 813
rect 35206 779 35218 813
rect 34818 767 35218 779
rect 35532 901 35932 913
rect 35532 867 35544 901
rect 35920 867 35932 901
rect 35532 855 35932 867
rect 35532 813 35932 825
rect 35532 779 35544 813
rect 35920 779 35932 813
rect 35532 767 35932 779
rect 36246 901 36646 913
rect 36246 867 36258 901
rect 36634 867 36646 901
rect 36246 855 36646 867
rect 36246 813 36646 825
rect 36246 779 36258 813
rect 36634 779 36646 813
rect 36246 767 36646 779
rect 36960 901 37360 913
rect 36960 867 36972 901
rect 37348 867 37360 901
rect 36960 855 37360 867
rect 36960 813 37360 825
rect 36960 779 36972 813
rect 37348 779 37360 813
rect 36960 767 37360 779
rect 37674 901 38074 913
rect 37674 867 37686 901
rect 38062 867 38074 901
rect 37674 855 38074 867
rect 37674 813 38074 825
rect 37674 779 37686 813
rect 38062 779 38074 813
rect 37674 767 38074 779
rect 38388 901 38788 913
rect 38388 867 38400 901
rect 38776 867 38788 901
rect 38388 855 38788 867
rect 38388 813 38788 825
rect 38388 779 38400 813
rect 38776 779 38788 813
rect 38388 767 38788 779
rect 3806 -144 3864 -132
rect 3806 -520 3818 -144
rect 3852 -520 3864 -144
rect 3806 -532 3864 -520
rect 3894 -144 3952 -132
rect 3894 -520 3906 -144
rect 3940 -520 3952 -144
rect 3894 -532 3952 -520
rect 15540 83 15940 95
rect 15540 49 15552 83
rect 15928 49 15940 83
rect 15540 37 15940 49
rect 15540 -5 15940 7
rect 15540 -39 15552 -5
rect 15928 -39 15940 -5
rect 15540 -51 15940 -39
rect 16254 83 16654 95
rect 16254 49 16266 83
rect 16642 49 16654 83
rect 16254 37 16654 49
rect 16254 -5 16654 7
rect 16254 -39 16266 -5
rect 16642 -39 16654 -5
rect 16254 -51 16654 -39
rect 16968 83 17368 95
rect 16968 49 16980 83
rect 17356 49 17368 83
rect 16968 37 17368 49
rect 16968 -5 17368 7
rect 16968 -39 16980 -5
rect 17356 -39 17368 -5
rect 16968 -51 17368 -39
rect 17682 83 18082 95
rect 17682 49 17694 83
rect 18070 49 18082 83
rect 17682 37 18082 49
rect 17682 -5 18082 7
rect 17682 -39 17694 -5
rect 18070 -39 18082 -5
rect 17682 -51 18082 -39
rect 18396 83 18796 95
rect 18396 49 18408 83
rect 18784 49 18796 83
rect 18396 37 18796 49
rect 18396 -5 18796 7
rect 18396 -39 18408 -5
rect 18784 -39 18796 -5
rect 18396 -51 18796 -39
rect 19110 83 19510 95
rect 19110 49 19122 83
rect 19498 49 19510 83
rect 19110 37 19510 49
rect 19110 -5 19510 7
rect 19110 -39 19122 -5
rect 19498 -39 19510 -5
rect 19110 -51 19510 -39
rect 19824 83 20224 95
rect 19824 49 19836 83
rect 20212 49 20224 83
rect 19824 37 20224 49
rect 19824 -5 20224 7
rect 19824 -39 19836 -5
rect 20212 -39 20224 -5
rect 19824 -51 20224 -39
rect 20538 83 20938 95
rect 20538 49 20550 83
rect 20926 49 20938 83
rect 20538 37 20938 49
rect 20538 -5 20938 7
rect 20538 -39 20550 -5
rect 20926 -39 20938 -5
rect 20538 -51 20938 -39
rect 21252 83 21652 95
rect 21252 49 21264 83
rect 21640 49 21652 83
rect 21252 37 21652 49
rect 21252 -5 21652 7
rect 21252 -39 21264 -5
rect 21640 -39 21652 -5
rect 21252 -51 21652 -39
rect 21966 83 22366 95
rect 21966 49 21978 83
rect 22354 49 22366 83
rect 21966 37 22366 49
rect 21966 -5 22366 7
rect 21966 -39 21978 -5
rect 22354 -39 22366 -5
rect 21966 -51 22366 -39
rect 22680 83 23080 95
rect 22680 49 22692 83
rect 23068 49 23080 83
rect 22680 37 23080 49
rect 22680 -5 23080 7
rect 22680 -39 22692 -5
rect 23068 -39 23080 -5
rect 22680 -51 23080 -39
rect 23394 83 23794 95
rect 23394 49 23406 83
rect 23782 49 23794 83
rect 23394 37 23794 49
rect 23394 -5 23794 7
rect 23394 -39 23406 -5
rect 23782 -39 23794 -5
rect 23394 -51 23794 -39
rect 24108 83 24508 95
rect 24108 49 24120 83
rect 24496 49 24508 83
rect 24108 37 24508 49
rect 24108 -5 24508 7
rect 24108 -39 24120 -5
rect 24496 -39 24508 -5
rect 24108 -51 24508 -39
rect 24822 83 25222 95
rect 24822 49 24834 83
rect 25210 49 25222 83
rect 24822 37 25222 49
rect 24822 -5 25222 7
rect 24822 -39 24834 -5
rect 25210 -39 25222 -5
rect 24822 -51 25222 -39
rect 25536 83 25936 95
rect 25536 49 25548 83
rect 25924 49 25936 83
rect 25536 37 25936 49
rect 25536 -5 25936 7
rect 25536 -39 25548 -5
rect 25924 -39 25936 -5
rect 25536 -51 25936 -39
rect 26250 83 26650 95
rect 26250 49 26262 83
rect 26638 49 26650 83
rect 26250 37 26650 49
rect 26250 -5 26650 7
rect 26250 -39 26262 -5
rect 26638 -39 26650 -5
rect 26250 -51 26650 -39
rect 26964 83 27364 95
rect 26964 49 26976 83
rect 27352 49 27364 83
rect 26964 37 27364 49
rect 26964 -5 27364 7
rect 26964 -39 26976 -5
rect 27352 -39 27364 -5
rect 26964 -51 27364 -39
rect 27678 83 28078 95
rect 27678 49 27690 83
rect 28066 49 28078 83
rect 27678 37 28078 49
rect 27678 -5 28078 7
rect 27678 -39 27690 -5
rect 28066 -39 28078 -5
rect 27678 -51 28078 -39
rect 28392 83 28792 95
rect 28392 49 28404 83
rect 28780 49 28792 83
rect 28392 37 28792 49
rect 28392 -5 28792 7
rect 28392 -39 28404 -5
rect 28780 -39 28792 -5
rect 28392 -51 28792 -39
rect 29106 83 29506 95
rect 29106 49 29118 83
rect 29494 49 29506 83
rect 29106 37 29506 49
rect 29106 -5 29506 7
rect 29106 -39 29118 -5
rect 29494 -39 29506 -5
rect 29106 -51 29506 -39
rect 29820 83 30220 95
rect 29820 49 29832 83
rect 30208 49 30220 83
rect 29820 37 30220 49
rect 29820 -5 30220 7
rect 29820 -39 29832 -5
rect 30208 -39 30220 -5
rect 29820 -51 30220 -39
rect 30534 83 30934 95
rect 30534 49 30546 83
rect 30922 49 30934 83
rect 30534 37 30934 49
rect 30534 -5 30934 7
rect 30534 -39 30546 -5
rect 30922 -39 30934 -5
rect 30534 -51 30934 -39
rect 31248 83 31648 95
rect 31248 49 31260 83
rect 31636 49 31648 83
rect 31248 37 31648 49
rect 31248 -5 31648 7
rect 31248 -39 31260 -5
rect 31636 -39 31648 -5
rect 31248 -51 31648 -39
rect 31962 83 32362 95
rect 31962 49 31974 83
rect 32350 49 32362 83
rect 31962 37 32362 49
rect 31962 -5 32362 7
rect 31962 -39 31974 -5
rect 32350 -39 32362 -5
rect 31962 -51 32362 -39
rect 32676 83 33076 95
rect 32676 49 32688 83
rect 33064 49 33076 83
rect 32676 37 33076 49
rect 32676 -5 33076 7
rect 32676 -39 32688 -5
rect 33064 -39 33076 -5
rect 32676 -51 33076 -39
rect 33390 83 33790 95
rect 33390 49 33402 83
rect 33778 49 33790 83
rect 33390 37 33790 49
rect 33390 -5 33790 7
rect 33390 -39 33402 -5
rect 33778 -39 33790 -5
rect 33390 -51 33790 -39
rect 34104 83 34504 95
rect 34104 49 34116 83
rect 34492 49 34504 83
rect 34104 37 34504 49
rect 34104 -5 34504 7
rect 34104 -39 34116 -5
rect 34492 -39 34504 -5
rect 34104 -51 34504 -39
rect 34818 83 35218 95
rect 34818 49 34830 83
rect 35206 49 35218 83
rect 34818 37 35218 49
rect 34818 -5 35218 7
rect 34818 -39 34830 -5
rect 35206 -39 35218 -5
rect 34818 -51 35218 -39
rect 35532 83 35932 95
rect 35532 49 35544 83
rect 35920 49 35932 83
rect 35532 37 35932 49
rect 35532 -5 35932 7
rect 35532 -39 35544 -5
rect 35920 -39 35932 -5
rect 35532 -51 35932 -39
rect 36246 83 36646 95
rect 36246 49 36258 83
rect 36634 49 36646 83
rect 36246 37 36646 49
rect 36246 -5 36646 7
rect 36246 -39 36258 -5
rect 36634 -39 36646 -5
rect 36246 -51 36646 -39
rect 36960 83 37360 95
rect 36960 49 36972 83
rect 37348 49 37360 83
rect 36960 37 37360 49
rect 36960 -5 37360 7
rect 36960 -39 36972 -5
rect 37348 -39 37360 -5
rect 36960 -51 37360 -39
rect 37674 83 38074 95
rect 37674 49 37686 83
rect 38062 49 38074 83
rect 37674 37 38074 49
rect 37674 -5 38074 7
rect 37674 -39 37686 -5
rect 38062 -39 38074 -5
rect 37674 -51 38074 -39
rect 38388 83 38788 95
rect 38388 49 38400 83
rect 38776 49 38788 83
rect 38388 37 38788 49
rect 38388 -5 38788 7
rect 38388 -39 38400 -5
rect 38776 -39 38788 -5
rect 38388 -51 38788 -39
rect 10615 -804 10745 -796
rect 10615 -838 10627 -804
rect 10661 -838 10695 -804
rect 10729 -838 10745 -804
rect 10615 -848 10745 -838
rect 10615 -888 10745 -878
rect 10615 -922 10627 -888
rect 10661 -922 10695 -888
rect 10729 -922 10745 -888
rect 10615 -930 10745 -922
rect 5847 -4388 5905 -4376
rect 5847 -6364 5859 -4388
rect 5893 -6364 5905 -4388
rect 5847 -6376 5905 -6364
rect 5965 -4388 6023 -4376
rect 5965 -6364 5977 -4388
rect 6011 -6364 6023 -4388
rect 5965 -6376 6023 -6364
rect 6083 -4388 6141 -4376
rect 6083 -6364 6095 -4388
rect 6129 -6364 6141 -4388
rect 6083 -6376 6141 -6364
rect 6201 -4388 6259 -4376
rect 6201 -6364 6213 -4388
rect 6247 -6364 6259 -4388
rect 6201 -6376 6259 -6364
rect 6319 -4388 6377 -4376
rect 6319 -6364 6331 -4388
rect 6365 -6364 6377 -4388
rect 6319 -6376 6377 -6364
rect 6437 -4388 6495 -4376
rect 6437 -6364 6449 -4388
rect 6483 -6364 6495 -4388
rect 6437 -6376 6495 -6364
rect 6555 -4388 6613 -4376
rect 6555 -6364 6567 -4388
rect 6601 -6364 6613 -4388
rect 6555 -6376 6613 -6364
rect 7055 -3272 7113 -3260
rect 7055 -5248 7067 -3272
rect 7101 -5248 7113 -3272
rect 7055 -5260 7113 -5248
rect 7513 -3272 7571 -3260
rect 7513 -5248 7525 -3272
rect 7559 -5248 7571 -3272
rect 7513 -5260 7571 -5248
rect 7971 -3272 8029 -3260
rect 7971 -5248 7983 -3272
rect 8017 -5248 8029 -3272
rect 7971 -5260 8029 -5248
rect 8429 -3272 8487 -3260
rect 8429 -5248 8441 -3272
rect 8475 -5248 8487 -3272
rect 8429 -5260 8487 -5248
rect 8887 -3272 8945 -3260
rect 8887 -5248 8899 -3272
rect 8933 -5248 8945 -3272
rect 8887 -5260 8945 -5248
rect 10852 -3484 11352 -3472
rect 10852 -3518 10864 -3484
rect 11340 -3518 11352 -3484
rect 10852 -3534 11352 -3518
rect 10852 -3580 11352 -3564
rect 10852 -3614 10864 -3580
rect 11340 -3614 11352 -3580
rect 10852 -3630 11352 -3614
rect 10852 -3676 11352 -3660
rect 10852 -3710 10864 -3676
rect 11340 -3710 11352 -3676
rect 10852 -3726 11352 -3710
rect 10852 -3772 11352 -3756
rect 10852 -3806 10864 -3772
rect 11340 -3806 11352 -3772
rect 10852 -3822 11352 -3806
rect 10852 -3868 11352 -3852
rect 10852 -3902 10864 -3868
rect 11340 -3902 11352 -3868
rect 10852 -3914 11352 -3902
rect 7011 -5712 7073 -5700
rect 7011 -6188 7023 -5712
rect 7057 -6188 7073 -5712
rect 7011 -6200 7073 -6188
rect 7103 -5712 7169 -5700
rect 7103 -6188 7119 -5712
rect 7153 -6188 7169 -5712
rect 7103 -6200 7169 -6188
rect 7199 -5712 7265 -5700
rect 7199 -6188 7215 -5712
rect 7249 -6188 7265 -5712
rect 7199 -6200 7265 -6188
rect 7295 -5712 7361 -5700
rect 7295 -6188 7311 -5712
rect 7345 -6188 7361 -5712
rect 7295 -6200 7361 -6188
rect 7391 -5712 7457 -5700
rect 7391 -6188 7407 -5712
rect 7441 -6188 7457 -5712
rect 7391 -6200 7457 -6188
rect 7487 -5712 7553 -5700
rect 7487 -6188 7503 -5712
rect 7537 -6188 7553 -5712
rect 7487 -6200 7553 -6188
rect 7583 -5712 7649 -5700
rect 7583 -6188 7599 -5712
rect 7633 -6188 7649 -5712
rect 7583 -6200 7649 -6188
rect 7679 -5712 7745 -5700
rect 7679 -6188 7695 -5712
rect 7729 -6188 7745 -5712
rect 7679 -6200 7745 -6188
rect 7775 -5712 7841 -5700
rect 7775 -6188 7791 -5712
rect 7825 -6188 7841 -5712
rect 7775 -6200 7841 -6188
rect 7871 -5712 7937 -5700
rect 7871 -6188 7887 -5712
rect 7921 -6188 7937 -5712
rect 7871 -6200 7937 -6188
rect 7967 -5712 8033 -5700
rect 7967 -6188 7983 -5712
rect 8017 -6188 8033 -5712
rect 7967 -6200 8033 -6188
rect 8063 -5712 8129 -5700
rect 8063 -6188 8079 -5712
rect 8113 -6188 8129 -5712
rect 8063 -6200 8129 -6188
rect 8159 -5712 8225 -5700
rect 8159 -6188 8175 -5712
rect 8209 -6188 8225 -5712
rect 8159 -6200 8225 -6188
rect 8255 -5712 8321 -5700
rect 8255 -6188 8271 -5712
rect 8305 -6188 8321 -5712
rect 8255 -6200 8321 -6188
rect 8351 -5712 8417 -5700
rect 8351 -6188 8367 -5712
rect 8401 -6188 8417 -5712
rect 8351 -6200 8417 -6188
rect 8447 -5712 8513 -5700
rect 8447 -6188 8463 -5712
rect 8497 -6188 8513 -5712
rect 8447 -6200 8513 -6188
rect 8543 -5712 8609 -5700
rect 8543 -6188 8559 -5712
rect 8593 -6188 8609 -5712
rect 8543 -6200 8609 -6188
rect 8639 -5712 8705 -5700
rect 8639 -6188 8655 -5712
rect 8689 -6188 8705 -5712
rect 8639 -6200 8705 -6188
rect 8735 -5712 8801 -5700
rect 8735 -6188 8751 -5712
rect 8785 -6188 8801 -5712
rect 8735 -6200 8801 -6188
rect 8831 -5712 8897 -5700
rect 8831 -6188 8847 -5712
rect 8881 -6188 8897 -5712
rect 8831 -6200 8897 -6188
rect 8927 -5712 8989 -5700
rect 8927 -6188 8943 -5712
rect 8977 -6188 8989 -5712
rect 8927 -6200 8989 -6188
rect 9388 -4388 9446 -4376
rect 9388 -6364 9400 -4388
rect 9434 -6364 9446 -4388
rect 9388 -6376 9446 -6364
rect 9506 -4388 9564 -4376
rect 9506 -6364 9518 -4388
rect 9552 -6364 9564 -4388
rect 9506 -6376 9564 -6364
rect 9624 -4388 9682 -4376
rect 9624 -6364 9636 -4388
rect 9670 -6364 9682 -4388
rect 9624 -6376 9682 -6364
rect 9742 -4388 9800 -4376
rect 9742 -6364 9754 -4388
rect 9788 -6364 9800 -4388
rect 9742 -6376 9800 -6364
rect 9860 -4388 9918 -4376
rect 9860 -6364 9872 -4388
rect 9906 -6364 9918 -4388
rect 9860 -6376 9918 -6364
rect 9978 -4388 10036 -4376
rect 9978 -6364 9990 -4388
rect 10024 -6364 10036 -4388
rect 9978 -6376 10036 -6364
rect 10096 -4388 10154 -4376
rect 10096 -6364 10108 -4388
rect 10142 -6364 10154 -4388
rect 10096 -6376 10154 -6364
<< pdiff >>
rect 6083 12273 6141 12285
rect 6083 10297 6095 12273
rect 6129 10297 6141 12273
rect 6083 10285 6141 10297
rect 6201 12273 6259 12285
rect 6201 10297 6213 12273
rect 6247 10297 6259 12273
rect 6201 10285 6259 10297
rect 6319 12273 6377 12285
rect 6319 10297 6331 12273
rect 6365 10297 6377 12273
rect 6319 10285 6377 10297
rect 6437 12273 6495 12285
rect 6437 10297 6449 12273
rect 6483 10297 6495 12273
rect 6437 10285 6495 10297
rect 6555 12273 6613 12285
rect 6555 10297 6567 12273
rect 6601 10297 6613 12273
rect 6555 10285 6613 10297
rect 6673 12273 6731 12285
rect 6673 10297 6685 12273
rect 6719 10297 6731 12273
rect 6673 10285 6731 10297
rect 6791 12273 6849 12285
rect 6791 10297 6803 12273
rect 6837 10297 6849 12273
rect 6791 10285 6849 10297
rect 6909 12273 6967 12285
rect 6909 10297 6921 12273
rect 6955 10297 6967 12273
rect 6909 10285 6967 10297
rect 7027 12273 7085 12285
rect 7027 10297 7039 12273
rect 7073 10297 7085 12273
rect 7027 10285 7085 10297
rect 7145 12273 7203 12285
rect 7145 10297 7157 12273
rect 7191 10297 7203 12273
rect 7145 10285 7203 10297
rect 7263 12273 7321 12285
rect 7263 10297 7275 12273
rect 7309 10297 7321 12273
rect 7263 10285 7321 10297
rect 7381 12273 7439 12285
rect 7381 10297 7393 12273
rect 7427 10297 7439 12273
rect 7381 10285 7439 10297
rect 7499 12273 7557 12285
rect 7499 10297 7511 12273
rect 7545 10297 7557 12273
rect 7499 10285 7557 10297
rect 7617 12273 7675 12285
rect 7617 10297 7629 12273
rect 7663 10297 7675 12273
rect 7617 10285 7675 10297
rect 7735 12273 7793 12285
rect 7735 10297 7747 12273
rect 7781 10297 7793 12273
rect 7735 10285 7793 10297
rect 7853 12273 7911 12285
rect 7853 10297 7865 12273
rect 7899 10297 7911 12273
rect 7853 10285 7911 10297
rect 7971 12273 8029 12285
rect 7971 10297 7983 12273
rect 8017 10297 8029 12273
rect 7971 10285 8029 10297
rect 8089 12273 8147 12285
rect 8089 10297 8101 12273
rect 8135 10297 8147 12273
rect 8089 10285 8147 10297
rect 8207 12273 8265 12285
rect 8207 10297 8219 12273
rect 8253 10297 8265 12273
rect 8207 10285 8265 10297
rect 8325 12273 8383 12285
rect 8325 10297 8337 12273
rect 8371 10297 8383 12273
rect 8325 10285 8383 10297
rect 8443 12273 8501 12285
rect 8443 10297 8455 12273
rect 8489 10297 8501 12273
rect 8443 10285 8501 10297
rect 8561 12273 8619 12285
rect 8561 10297 8573 12273
rect 8607 10297 8619 12273
rect 8561 10285 8619 10297
rect 8679 12273 8737 12285
rect 8679 10297 8691 12273
rect 8725 10297 8737 12273
rect 8679 10285 8737 10297
rect 8797 12273 8855 12285
rect 8797 10297 8809 12273
rect 8843 10297 8855 12273
rect 8797 10285 8855 10297
rect 8915 12273 8973 12285
rect 8915 10297 8927 12273
rect 8961 10297 8973 12273
rect 8915 10285 8973 10297
rect 9033 12273 9091 12285
rect 9033 10297 9045 12273
rect 9079 10297 9091 12273
rect 9033 10285 9091 10297
rect 9151 12273 9209 12285
rect 9151 10297 9163 12273
rect 9197 10297 9209 12273
rect 9151 10285 9209 10297
rect 9269 12273 9327 12285
rect 9269 10297 9281 12273
rect 9315 10297 9327 12273
rect 9269 10285 9327 10297
rect 9387 12273 9445 12285
rect 9387 10297 9399 12273
rect 9433 10297 9445 12273
rect 9387 10285 9445 10297
rect 9505 12273 9563 12285
rect 9505 10297 9517 12273
rect 9551 10297 9563 12273
rect 9505 10285 9563 10297
rect 9623 12273 9681 12285
rect 9623 10297 9635 12273
rect 9669 10297 9681 12273
rect 9623 10285 9681 10297
rect 9741 12273 9799 12285
rect 9741 10297 9753 12273
rect 9787 10297 9799 12273
rect 9741 10285 9799 10297
rect 9859 12273 9917 12285
rect 9859 10297 9871 12273
rect 9905 10297 9917 12273
rect 9859 10285 9917 10297
rect 2428 2792 2497 2804
rect 2428 2758 2440 2792
rect 2474 2758 2497 2792
rect 2428 2722 2497 2758
rect 2428 2688 2440 2722
rect 2474 2688 2497 2722
rect 2428 2652 2497 2688
rect 2428 2618 2440 2652
rect 2474 2618 2497 2652
rect 2428 2580 2497 2618
rect 2527 2792 2586 2804
rect 2527 2758 2540 2792
rect 2574 2758 2586 2792
rect 2527 2709 2586 2758
rect 2527 2675 2540 2709
rect 2574 2675 2586 2709
rect 2527 2626 2586 2675
rect 3794 2792 3851 2804
rect 3794 2758 3804 2792
rect 3838 2758 3851 2792
rect 3794 2709 3851 2758
rect 3794 2675 3804 2709
rect 3838 2675 3851 2709
rect 2527 2592 2540 2626
rect 2574 2592 2586 2626
rect 2527 2580 2586 2592
rect 3794 2626 3851 2675
rect 3794 2592 3804 2626
rect 3838 2592 3851 2626
rect 3794 2580 3851 2592
rect 3881 2792 3941 2804
rect 3881 2758 3894 2792
rect 3928 2758 3941 2792
rect 3881 2709 3941 2758
rect 3881 2675 3894 2709
rect 3928 2675 3941 2709
rect 3881 2626 3941 2675
rect 3881 2592 3894 2626
rect 3928 2592 3941 2626
rect 3881 2580 3941 2592
rect 3971 2792 4028 2804
rect 3971 2758 3984 2792
rect 4018 2758 4028 2792
rect 3971 2709 4028 2758
rect 3971 2675 3984 2709
rect 4018 2675 4028 2709
rect 3971 2626 4028 2675
rect 3971 2592 3984 2626
rect 4018 2592 4028 2626
rect 4082 2792 4137 2804
rect 4082 2758 4090 2792
rect 4124 2758 4137 2792
rect 4082 2721 4137 2758
rect 4082 2687 4090 2721
rect 4124 2687 4137 2721
rect 4082 2650 4137 2687
rect 4082 2616 4090 2650
rect 4124 2616 4137 2650
rect 4082 2604 4137 2616
rect 4337 2792 4392 2804
rect 4337 2758 4348 2792
rect 4382 2758 4392 2792
rect 4337 2721 4392 2758
rect 4337 2687 4348 2721
rect 4382 2687 4392 2721
rect 4337 2650 4392 2687
rect 4337 2616 4348 2650
rect 4382 2616 4392 2650
rect 4337 2604 4392 2616
rect 4592 2792 4649 2804
rect 4592 2758 4603 2792
rect 4637 2758 4649 2792
rect 4592 2721 4649 2758
rect 4592 2687 4603 2721
rect 4637 2687 4649 2721
rect 4592 2650 4649 2687
rect 4592 2616 4603 2650
rect 4637 2616 4649 2650
rect 5426 2792 5481 2804
rect 5426 2758 5434 2792
rect 5468 2758 5481 2792
rect 5426 2721 5481 2758
rect 5426 2687 5434 2721
rect 5468 2687 5481 2721
rect 5426 2650 5481 2687
rect 4592 2604 4649 2616
rect 5426 2616 5434 2650
rect 5468 2616 5481 2650
rect 5426 2604 5481 2616
rect 5681 2792 5736 2804
rect 5681 2758 5692 2792
rect 5726 2758 5736 2792
rect 5681 2721 5736 2758
rect 5681 2687 5692 2721
rect 5726 2687 5736 2721
rect 5681 2650 5736 2687
rect 5681 2616 5692 2650
rect 5726 2616 5736 2650
rect 5681 2604 5736 2616
rect 5936 2792 5993 2804
rect 5936 2758 5947 2792
rect 5981 2758 5993 2792
rect 5936 2721 5993 2758
rect 5936 2687 5947 2721
rect 5981 2687 5993 2721
rect 5936 2650 5993 2687
rect 5936 2616 5947 2650
rect 5981 2616 5993 2650
rect 5936 2604 5993 2616
rect 6098 2792 6153 2804
rect 6098 2758 6106 2792
rect 6140 2758 6153 2792
rect 6098 2721 6153 2758
rect 6098 2687 6106 2721
rect 6140 2687 6153 2721
rect 6098 2650 6153 2687
rect 6098 2616 6106 2650
rect 6140 2616 6153 2650
rect 6098 2604 6153 2616
rect 6353 2792 6408 2804
rect 6353 2758 6364 2792
rect 6398 2758 6408 2792
rect 6353 2721 6408 2758
rect 6353 2687 6364 2721
rect 6398 2687 6408 2721
rect 6353 2650 6408 2687
rect 6353 2616 6364 2650
rect 6398 2616 6408 2650
rect 6353 2604 6408 2616
rect 6608 2792 6665 2804
rect 6608 2758 6619 2792
rect 6653 2758 6665 2792
rect 6608 2721 6665 2758
rect 6608 2687 6619 2721
rect 6653 2687 6665 2721
rect 6608 2650 6665 2687
rect 6608 2616 6619 2650
rect 6653 2616 6665 2650
rect 6608 2604 6665 2616
rect 6770 2792 6825 2804
rect 6770 2758 6778 2792
rect 6812 2758 6825 2792
rect 6770 2721 6825 2758
rect 6770 2687 6778 2721
rect 6812 2687 6825 2721
rect 6770 2650 6825 2687
rect 6770 2616 6778 2650
rect 6812 2616 6825 2650
rect 6770 2604 6825 2616
rect 7025 2792 7080 2804
rect 7025 2758 7036 2792
rect 7070 2758 7080 2792
rect 7025 2721 7080 2758
rect 7025 2687 7036 2721
rect 7070 2687 7080 2721
rect 7025 2650 7080 2687
rect 7025 2616 7036 2650
rect 7070 2616 7080 2650
rect 7025 2604 7080 2616
rect 7280 2792 7337 2804
rect 7280 2758 7291 2792
rect 7325 2758 7337 2792
rect 7280 2721 7337 2758
rect 7280 2687 7291 2721
rect 7325 2687 7337 2721
rect 7280 2650 7337 2687
rect 7280 2616 7291 2650
rect 7325 2616 7337 2650
rect 7280 2604 7337 2616
rect 8114 2792 8169 2804
rect 8114 2758 8122 2792
rect 8156 2758 8169 2792
rect 8114 2721 8169 2758
rect 8114 2687 8122 2721
rect 8156 2687 8169 2721
rect 8114 2650 8169 2687
rect 8114 2616 8122 2650
rect 8156 2616 8169 2650
rect 8114 2604 8169 2616
rect 8369 2792 8424 2804
rect 8369 2758 8380 2792
rect 8414 2758 8424 2792
rect 8369 2721 8424 2758
rect 8369 2687 8380 2721
rect 8414 2687 8424 2721
rect 8369 2650 8424 2687
rect 8369 2616 8380 2650
rect 8414 2616 8424 2650
rect 8369 2604 8424 2616
rect 8624 2792 8681 2804
rect 8624 2758 8635 2792
rect 8669 2758 8681 2792
rect 8624 2721 8681 2758
rect 8624 2687 8635 2721
rect 8669 2687 8681 2721
rect 8624 2650 8681 2687
rect 8624 2616 8635 2650
rect 8669 2616 8681 2650
rect 8624 2604 8681 2616
rect 8786 2792 8841 2804
rect 8786 2758 8794 2792
rect 8828 2758 8841 2792
rect 8786 2721 8841 2758
rect 8786 2687 8794 2721
rect 8828 2687 8841 2721
rect 8786 2650 8841 2687
rect 8786 2616 8794 2650
rect 8828 2616 8841 2650
rect 8786 2604 8841 2616
rect 9041 2792 9096 2804
rect 9041 2758 9052 2792
rect 9086 2758 9096 2792
rect 9041 2721 9096 2758
rect 9041 2687 9052 2721
rect 9086 2687 9096 2721
rect 9041 2650 9096 2687
rect 9041 2616 9052 2650
rect 9086 2616 9096 2650
rect 9041 2604 9096 2616
rect 9296 2792 9353 2804
rect 9296 2758 9307 2792
rect 9341 2758 9353 2792
rect 9296 2721 9353 2758
rect 9296 2687 9307 2721
rect 9341 2687 9353 2721
rect 9296 2650 9353 2687
rect 9296 2616 9307 2650
rect 9341 2616 9353 2650
rect 9296 2604 9353 2616
rect 9458 2792 9513 2804
rect 9458 2758 9466 2792
rect 9500 2758 9513 2792
rect 9458 2721 9513 2758
rect 9458 2687 9466 2721
rect 9500 2687 9513 2721
rect 9458 2650 9513 2687
rect 9458 2616 9466 2650
rect 9500 2616 9513 2650
rect 9458 2604 9513 2616
rect 9713 2792 9770 2804
rect 9713 2758 9724 2792
rect 9758 2758 9770 2792
rect 9713 2721 9770 2758
rect 9713 2687 9724 2721
rect 9758 2687 9770 2721
rect 9713 2650 9770 2687
rect 9713 2616 9724 2650
rect 9758 2616 9770 2650
rect 9713 2604 9770 2616
rect 3971 2580 4028 2592
rect 2428 1806 2497 1844
rect 2428 1772 2440 1806
rect 2474 1772 2497 1806
rect 2428 1736 2497 1772
rect 2428 1702 2440 1736
rect 2474 1702 2497 1736
rect 2428 1666 2497 1702
rect 2428 1632 2440 1666
rect 2474 1632 2497 1666
rect 2428 1620 2497 1632
rect 2527 1832 2586 1844
rect 2527 1798 2540 1832
rect 2574 1798 2586 1832
rect 2527 1749 2586 1798
rect 3794 1832 3851 1844
rect 3794 1798 3804 1832
rect 3838 1798 3851 1832
rect 2527 1715 2540 1749
rect 2574 1715 2586 1749
rect 2527 1666 2586 1715
rect 2527 1632 2540 1666
rect 2574 1632 2586 1666
rect 2527 1620 2586 1632
rect 3794 1749 3851 1798
rect 3794 1715 3804 1749
rect 3838 1715 3851 1749
rect 3794 1666 3851 1715
rect 3794 1632 3804 1666
rect 3838 1632 3851 1666
rect 3794 1620 3851 1632
rect 3881 1832 3941 1844
rect 3881 1798 3894 1832
rect 3928 1798 3941 1832
rect 3881 1749 3941 1798
rect 3881 1715 3894 1749
rect 3928 1715 3941 1749
rect 3881 1666 3941 1715
rect 3881 1632 3894 1666
rect 3928 1632 3941 1666
rect 3881 1620 3941 1632
rect 3971 1832 4028 1844
rect 3971 1798 3984 1832
rect 4018 1798 4028 1832
rect 3971 1749 4028 1798
rect 3971 1715 3984 1749
rect 4018 1715 4028 1749
rect 3971 1666 4028 1715
rect 4082 1817 4141 1844
rect 4082 1783 4094 1817
rect 4128 1783 4141 1817
rect 4082 1722 4141 1783
rect 4082 1688 4094 1722
rect 4128 1688 4141 1722
rect 4082 1676 4141 1688
rect 4171 1727 4248 1844
rect 4171 1693 4201 1727
rect 4235 1693 4248 1727
rect 4171 1676 4248 1693
rect 3971 1632 3984 1666
rect 4018 1632 4028 1666
rect 4189 1644 4248 1676
rect 4278 1644 4441 1844
rect 4471 1832 4549 1844
rect 4471 1798 4484 1832
rect 4518 1798 4549 1832
rect 4471 1715 4549 1798
rect 4471 1681 4484 1715
rect 4518 1681 4549 1715
rect 4471 1644 4549 1681
rect 4579 1644 4663 1844
rect 4693 1832 4787 1844
rect 4693 1798 4730 1832
rect 4764 1798 4787 1832
rect 4693 1749 4787 1798
rect 4693 1715 4730 1749
rect 4764 1715 4787 1749
rect 4693 1666 4787 1715
rect 4693 1644 4730 1666
rect 3971 1620 4028 1632
rect 4718 1632 4730 1644
rect 4764 1632 4787 1666
rect 4718 1620 4787 1632
rect 4817 1832 4876 1844
rect 4817 1798 4830 1832
rect 4864 1798 4876 1832
rect 4817 1749 4876 1798
rect 4817 1715 4830 1749
rect 4864 1715 4876 1749
rect 4817 1666 4876 1715
rect 4817 1632 4830 1666
rect 4864 1632 4876 1666
rect 4817 1620 4876 1632
rect 4946 1806 5003 1844
rect 4946 1772 4956 1806
rect 4990 1772 5003 1806
rect 4946 1736 5003 1772
rect 4946 1702 4956 1736
rect 4990 1702 5003 1736
rect 4946 1666 5003 1702
rect 4946 1632 4956 1666
rect 4990 1632 5003 1666
rect 4946 1620 5003 1632
rect 5033 1832 5093 1844
rect 5033 1798 5046 1832
rect 5080 1798 5093 1832
rect 5033 1749 5093 1798
rect 5033 1715 5046 1749
rect 5080 1715 5093 1749
rect 5033 1666 5093 1715
rect 5033 1632 5046 1666
rect 5080 1632 5093 1666
rect 5033 1620 5093 1632
rect 5123 1832 5180 1844
rect 5123 1798 5136 1832
rect 5170 1798 5180 1832
rect 5123 1749 5180 1798
rect 5123 1715 5136 1749
rect 5170 1715 5180 1749
rect 5123 1666 5180 1715
rect 5123 1632 5136 1666
rect 5170 1632 5180 1666
rect 5123 1620 5180 1632
rect 6088 1806 6147 1844
rect 6088 1772 6100 1806
rect 6134 1772 6147 1806
rect 5426 1735 5485 1748
rect 5426 1701 5438 1735
rect 5472 1701 5485 1735
rect 5426 1666 5485 1701
rect 5426 1632 5438 1666
rect 5472 1632 5485 1666
rect 5426 1620 5485 1632
rect 5515 1667 5575 1748
rect 5515 1633 5528 1667
rect 5562 1633 5575 1667
rect 5515 1620 5575 1633
rect 5605 1620 5653 1748
rect 5683 1726 5743 1748
rect 5683 1692 5696 1726
rect 5730 1692 5743 1726
rect 5683 1620 5743 1692
rect 5773 1736 5832 1748
rect 5773 1702 5786 1736
rect 5820 1702 5832 1736
rect 5773 1666 5832 1702
rect 5773 1632 5786 1666
rect 5820 1632 5832 1666
rect 5773 1620 5832 1632
rect 5886 1736 5945 1748
rect 5886 1702 5898 1736
rect 5932 1702 5945 1736
rect 5886 1666 5945 1702
rect 5886 1632 5898 1666
rect 5932 1632 5945 1666
rect 5886 1620 5945 1632
rect 5975 1736 6034 1748
rect 5975 1702 5988 1736
rect 6022 1702 6034 1736
rect 5975 1666 6034 1702
rect 5975 1632 5988 1666
rect 6022 1632 6034 1666
rect 5975 1620 6034 1632
rect 6088 1736 6147 1772
rect 6088 1702 6100 1736
rect 6134 1702 6147 1736
rect 6088 1666 6147 1702
rect 6088 1632 6100 1666
rect 6134 1632 6147 1666
rect 6088 1620 6147 1632
rect 6177 1744 6237 1844
rect 6177 1710 6190 1744
rect 6224 1710 6237 1744
rect 6177 1666 6237 1710
rect 6177 1632 6190 1666
rect 6224 1632 6237 1666
rect 6177 1620 6237 1632
rect 6267 1828 6326 1844
rect 6267 1794 6280 1828
rect 6314 1794 6326 1828
rect 6267 1747 6326 1794
rect 6267 1713 6280 1747
rect 6314 1713 6326 1747
rect 6267 1666 6326 1713
rect 6267 1632 6280 1666
rect 6314 1632 6326 1666
rect 6380 1718 6439 1748
rect 6380 1684 6392 1718
rect 6426 1684 6439 1718
rect 6380 1664 6439 1684
rect 6469 1664 6523 1748
rect 6553 1726 6630 1748
rect 6553 1692 6583 1726
rect 6617 1692 6630 1726
rect 6553 1664 6630 1692
rect 6267 1620 6326 1632
rect 6571 1620 6630 1664
rect 6660 1726 6729 1748
rect 6660 1692 6683 1726
rect 6717 1692 6729 1726
rect 6660 1620 6729 1692
rect 6783 1666 6961 1788
rect 6783 1632 6795 1666
rect 6829 1632 6914 1666
rect 6948 1632 6961 1666
rect 6783 1620 6961 1632
rect 6991 1620 7045 1788
rect 7075 1703 7153 1788
rect 7075 1669 7088 1703
rect 7122 1669 7153 1703
rect 7075 1620 7153 1669
rect 7183 1776 7242 1788
rect 7183 1742 7196 1776
rect 7230 1742 7242 1776
rect 7183 1666 7242 1742
rect 7183 1632 7196 1666
rect 7230 1632 7242 1666
rect 7183 1620 7242 1632
rect 7296 1738 7355 1788
rect 7296 1704 7308 1738
rect 7342 1704 7355 1738
rect 7296 1666 7355 1704
rect 7296 1632 7308 1666
rect 7342 1632 7355 1666
rect 7296 1620 7355 1632
rect 7385 1620 7433 1788
rect 7463 1776 7522 1788
rect 7463 1742 7476 1776
rect 7510 1742 7522 1776
rect 7463 1704 7522 1742
rect 7764 1744 7823 1820
rect 7764 1710 7776 1744
rect 7810 1710 7823 1744
rect 7463 1666 7540 1704
rect 7463 1632 7476 1666
rect 7510 1632 7540 1666
rect 7463 1620 7540 1632
rect 7570 1620 7618 1704
rect 7648 1671 7707 1704
rect 7648 1637 7661 1671
rect 7695 1637 7707 1671
rect 7648 1620 7707 1637
rect 7764 1666 7823 1710
rect 7764 1632 7776 1666
rect 7810 1632 7823 1666
rect 7764 1620 7823 1632
rect 7853 1671 7925 1820
rect 7853 1637 7876 1671
rect 7910 1637 7925 1671
rect 7853 1620 7925 1637
rect 7955 1620 8009 1820
rect 8039 1784 8098 1820
rect 8394 1813 8447 1844
rect 8039 1750 8052 1784
rect 8086 1750 8098 1784
rect 8039 1666 8098 1750
rect 8152 1795 8211 1813
rect 8152 1761 8164 1795
rect 8198 1761 8211 1795
rect 8152 1685 8211 1761
rect 8241 1799 8447 1813
rect 8241 1765 8383 1799
rect 8417 1765 8447 1799
rect 8241 1717 8447 1765
rect 8241 1685 8383 1717
rect 8039 1632 8052 1666
rect 8086 1632 8098 1666
rect 8259 1683 8383 1685
rect 8417 1683 8447 1717
rect 8039 1620 8098 1632
rect 8259 1627 8447 1683
rect 8259 1593 8271 1627
rect 8305 1593 8383 1627
rect 8417 1620 8447 1627
rect 8477 1832 8537 1844
rect 8477 1798 8490 1832
rect 8524 1798 8537 1832
rect 8477 1749 8537 1798
rect 8477 1715 8490 1749
rect 8524 1715 8537 1749
rect 8477 1666 8537 1715
rect 8477 1632 8490 1666
rect 8524 1632 8537 1666
rect 8477 1620 8537 1632
rect 8567 1806 8624 1844
rect 8788 1828 8841 1844
rect 8567 1772 8580 1806
rect 8614 1772 8624 1806
rect 8567 1736 8624 1772
rect 8567 1702 8580 1736
rect 8614 1702 8624 1736
rect 8567 1666 8624 1702
rect 8567 1632 8580 1666
rect 8614 1632 8624 1666
rect 8567 1620 8624 1632
rect 8678 1816 8736 1828
rect 8678 1782 8689 1816
rect 8723 1782 8736 1816
rect 8678 1745 8736 1782
rect 8678 1711 8689 1745
rect 8723 1711 8736 1745
rect 8678 1674 8736 1711
rect 8678 1640 8689 1674
rect 8723 1640 8736 1674
rect 8678 1628 8736 1640
rect 8766 1820 8841 1828
rect 8766 1786 8794 1820
rect 8828 1786 8841 1820
rect 8766 1748 8841 1786
rect 8766 1714 8794 1748
rect 8828 1714 8841 1748
rect 8766 1670 8841 1714
rect 8766 1636 8794 1670
rect 8828 1636 8841 1670
rect 8766 1628 8841 1636
rect 8417 1593 8429 1620
rect 8784 1620 8841 1628
rect 8871 1832 8931 1844
rect 8871 1798 8884 1832
rect 8918 1798 8931 1832
rect 8871 1749 8931 1798
rect 8871 1715 8884 1749
rect 8918 1715 8931 1749
rect 8871 1666 8931 1715
rect 8871 1632 8884 1666
rect 8918 1632 8931 1666
rect 8871 1620 8931 1632
rect 8961 1832 9020 1844
rect 8961 1798 8974 1832
rect 9008 1798 9020 1832
rect 8961 1749 9020 1798
rect 8961 1715 8974 1749
rect 9008 1715 9020 1749
rect 8961 1666 9020 1715
rect 8961 1632 8974 1666
rect 9008 1632 9020 1666
rect 8961 1620 9020 1632
rect 9074 1662 9212 1844
rect 9074 1628 9090 1662
rect 9124 1628 9162 1662
rect 9196 1628 9212 1662
rect 9074 1620 9212 1628
rect 9266 1826 9326 1844
rect 9266 1792 9278 1826
rect 9312 1792 9326 1826
rect 9266 1746 9326 1792
rect 9266 1712 9278 1746
rect 9312 1712 9326 1746
rect 9266 1666 9326 1712
rect 9266 1632 9278 1666
rect 9312 1632 9326 1666
rect 9266 1620 9326 1632
rect 9356 1806 9578 1844
rect 9356 1772 9369 1806
rect 9403 1772 9449 1806
rect 9483 1772 9531 1806
rect 9565 1772 9578 1806
rect 9356 1735 9578 1772
rect 9356 1701 9369 1735
rect 9403 1701 9449 1735
rect 9483 1701 9531 1735
rect 9565 1701 9578 1735
rect 9356 1666 9578 1701
rect 9356 1632 9369 1666
rect 9403 1632 9449 1666
rect 9483 1632 9531 1666
rect 9565 1632 9578 1666
rect 9356 1620 9578 1632
rect 9608 1745 9678 1844
rect 9608 1711 9621 1745
rect 9655 1711 9678 1745
rect 9608 1666 9678 1711
rect 9608 1632 9621 1666
rect 9655 1632 9678 1666
rect 9608 1620 9678 1632
rect 9708 1806 9977 1844
rect 9708 1772 9721 1806
rect 9755 1772 9790 1806
rect 9824 1772 9861 1806
rect 9895 1772 9930 1806
rect 9964 1772 9977 1806
rect 9708 1735 9977 1772
rect 9708 1701 9721 1735
rect 9755 1701 9790 1735
rect 9824 1701 9861 1735
rect 9895 1701 9930 1735
rect 9964 1701 9977 1735
rect 9708 1666 9977 1701
rect 9708 1632 9721 1666
rect 9755 1632 9790 1666
rect 9824 1632 9861 1666
rect 9895 1632 9930 1666
rect 9964 1632 9977 1666
rect 9708 1620 9977 1632
rect 10007 1745 10076 1844
rect 10007 1711 10030 1745
rect 10064 1711 10076 1745
rect 10007 1666 10076 1711
rect 10007 1632 10030 1666
rect 10064 1632 10076 1666
rect 10007 1620 10076 1632
rect 8259 1581 8429 1593
rect 11362 3725 11420 3737
rect 11362 1749 11374 3725
rect 11408 1749 11420 3725
rect 11362 1737 11420 1749
rect 11820 3725 11878 3737
rect 11820 1749 11832 3725
rect 11866 1749 11878 3725
rect 11820 1737 11878 1749
rect 12278 3725 12336 3737
rect 12278 1749 12290 3725
rect 12324 1749 12336 3725
rect 12278 1737 12336 1749
rect 12736 3725 12794 3737
rect 12736 1749 12748 3725
rect 12782 1749 12794 3725
rect 12736 1737 12794 1749
rect 13194 3725 13252 3737
rect 13194 1749 13206 3725
rect 13240 1749 13252 3725
rect 13194 1737 13252 1749
rect 13652 3725 13710 3737
rect 13652 1749 13664 3725
rect 13698 1749 13710 3725
rect 13652 1737 13710 1749
rect 13880 3725 13938 3737
rect 13880 1749 13892 3725
rect 13926 1749 13938 3725
rect 13880 1737 13938 1749
rect 13968 3725 14026 3737
rect 13968 1749 13980 3725
rect 14014 1749 14026 3725
rect 13968 1737 14026 1749
rect 14196 3725 14254 3737
rect 14196 1749 14208 3725
rect 14242 1749 14254 3725
rect 14196 1737 14254 1749
rect 14284 3725 14342 3737
rect 14284 1749 14296 3725
rect 14330 1749 14342 3725
rect 14284 1737 14342 1749
rect 8259 1499 8429 1511
rect 3580 1460 3649 1472
rect 3580 1426 3592 1460
rect 3626 1426 3649 1460
rect 3580 1390 3649 1426
rect 3580 1356 3592 1390
rect 3626 1356 3649 1390
rect 3580 1320 3649 1356
rect 3580 1286 3592 1320
rect 3626 1286 3649 1320
rect 3580 1248 3649 1286
rect 3679 1460 3738 1472
rect 3679 1426 3692 1460
rect 3726 1426 3738 1460
rect 3679 1377 3738 1426
rect 3679 1343 3692 1377
rect 3726 1343 3738 1377
rect 3679 1294 3738 1343
rect 4946 1460 5003 1472
rect 4946 1426 4956 1460
rect 4990 1426 5003 1460
rect 4946 1377 5003 1426
rect 4946 1343 4956 1377
rect 4990 1343 5003 1377
rect 3679 1260 3692 1294
rect 3726 1260 3738 1294
rect 3679 1248 3738 1260
rect 4946 1294 5003 1343
rect 4946 1260 4956 1294
rect 4990 1260 5003 1294
rect 4946 1248 5003 1260
rect 5033 1460 5093 1472
rect 5033 1426 5046 1460
rect 5080 1426 5093 1460
rect 5033 1377 5093 1426
rect 5033 1343 5046 1377
rect 5080 1343 5093 1377
rect 5033 1294 5093 1343
rect 5033 1260 5046 1294
rect 5080 1260 5093 1294
rect 5033 1248 5093 1260
rect 5123 1460 5180 1472
rect 5123 1426 5136 1460
rect 5170 1426 5180 1460
rect 5123 1377 5180 1426
rect 5123 1343 5136 1377
rect 5170 1343 5180 1377
rect 5123 1294 5180 1343
rect 5426 1460 5485 1472
rect 5426 1426 5438 1460
rect 5472 1426 5485 1460
rect 5426 1391 5485 1426
rect 5426 1357 5438 1391
rect 5472 1357 5485 1391
rect 5426 1344 5485 1357
rect 5515 1459 5575 1472
rect 5515 1425 5528 1459
rect 5562 1425 5575 1459
rect 5515 1344 5575 1425
rect 5605 1344 5653 1472
rect 5683 1400 5743 1472
rect 5683 1366 5696 1400
rect 5730 1366 5743 1400
rect 5683 1344 5743 1366
rect 5773 1460 5832 1472
rect 5773 1426 5786 1460
rect 5820 1426 5832 1460
rect 5773 1390 5832 1426
rect 5773 1356 5786 1390
rect 5820 1356 5832 1390
rect 5773 1344 5832 1356
rect 5886 1460 5945 1472
rect 5886 1426 5898 1460
rect 5932 1426 5945 1460
rect 5886 1390 5945 1426
rect 5886 1356 5898 1390
rect 5932 1356 5945 1390
rect 5886 1344 5945 1356
rect 5975 1460 6034 1472
rect 5975 1426 5988 1460
rect 6022 1426 6034 1460
rect 5975 1390 6034 1426
rect 5975 1356 5988 1390
rect 6022 1356 6034 1390
rect 5975 1344 6034 1356
rect 6088 1460 6147 1472
rect 6088 1426 6100 1460
rect 6134 1426 6147 1460
rect 6088 1390 6147 1426
rect 6088 1356 6100 1390
rect 6134 1356 6147 1390
rect 5123 1260 5136 1294
rect 5170 1260 5180 1294
rect 5123 1248 5180 1260
rect 6088 1320 6147 1356
rect 6088 1286 6100 1320
rect 6134 1286 6147 1320
rect 6088 1248 6147 1286
rect 6177 1460 6237 1472
rect 6177 1426 6190 1460
rect 6224 1426 6237 1460
rect 6177 1382 6237 1426
rect 6177 1348 6190 1382
rect 6224 1348 6237 1382
rect 6177 1248 6237 1348
rect 6267 1460 6326 1472
rect 6267 1426 6280 1460
rect 6314 1426 6326 1460
rect 6571 1428 6630 1472
rect 6267 1379 6326 1426
rect 6267 1345 6280 1379
rect 6314 1345 6326 1379
rect 6267 1298 6326 1345
rect 6380 1408 6439 1428
rect 6380 1374 6392 1408
rect 6426 1374 6439 1408
rect 6380 1344 6439 1374
rect 6469 1344 6523 1428
rect 6553 1400 6630 1428
rect 6553 1366 6583 1400
rect 6617 1366 6630 1400
rect 6553 1344 6630 1366
rect 6660 1400 6729 1472
rect 6660 1366 6683 1400
rect 6717 1366 6729 1400
rect 6660 1344 6729 1366
rect 6783 1460 6961 1472
rect 6783 1426 6795 1460
rect 6829 1426 6914 1460
rect 6948 1426 6961 1460
rect 6267 1264 6280 1298
rect 6314 1264 6326 1298
rect 6267 1248 6326 1264
rect 6783 1304 6961 1426
rect 6991 1304 7045 1472
rect 7075 1423 7153 1472
rect 7075 1389 7088 1423
rect 7122 1389 7153 1423
rect 7075 1304 7153 1389
rect 7183 1460 7242 1472
rect 7183 1426 7196 1460
rect 7230 1426 7242 1460
rect 7183 1350 7242 1426
rect 7183 1316 7196 1350
rect 7230 1316 7242 1350
rect 7183 1304 7242 1316
rect 7296 1460 7355 1472
rect 7296 1426 7308 1460
rect 7342 1426 7355 1460
rect 7296 1388 7355 1426
rect 7296 1354 7308 1388
rect 7342 1354 7355 1388
rect 7296 1304 7355 1354
rect 7385 1304 7433 1472
rect 7463 1460 7540 1472
rect 7463 1426 7476 1460
rect 7510 1426 7540 1460
rect 7463 1388 7540 1426
rect 7570 1388 7618 1472
rect 7648 1455 7707 1472
rect 7648 1421 7661 1455
rect 7695 1421 7707 1455
rect 7648 1388 7707 1421
rect 7764 1460 7823 1472
rect 7764 1426 7776 1460
rect 7810 1426 7823 1460
rect 7463 1350 7522 1388
rect 7764 1382 7823 1426
rect 7463 1316 7476 1350
rect 7510 1316 7522 1350
rect 7463 1304 7522 1316
rect 7764 1348 7776 1382
rect 7810 1348 7823 1382
rect 7764 1272 7823 1348
rect 7853 1455 7925 1472
rect 7853 1421 7876 1455
rect 7910 1421 7925 1455
rect 7853 1272 7925 1421
rect 7955 1272 8009 1472
rect 8039 1460 8098 1472
rect 8039 1426 8052 1460
rect 8086 1426 8098 1460
rect 8259 1465 8271 1499
rect 8305 1465 8383 1499
rect 8417 1472 8429 1499
rect 8417 1465 8447 1472
rect 8039 1342 8098 1426
rect 8259 1409 8447 1465
rect 8259 1407 8383 1409
rect 8039 1308 8052 1342
rect 8086 1308 8098 1342
rect 8039 1272 8098 1308
rect 8152 1331 8211 1407
rect 8152 1297 8164 1331
rect 8198 1297 8211 1331
rect 8152 1279 8211 1297
rect 8241 1375 8383 1407
rect 8417 1375 8447 1409
rect 8241 1327 8447 1375
rect 8241 1293 8383 1327
rect 8417 1293 8447 1327
rect 8241 1279 8447 1293
rect 8394 1248 8447 1279
rect 8477 1460 8537 1472
rect 8477 1426 8490 1460
rect 8524 1426 8537 1460
rect 8477 1377 8537 1426
rect 8477 1343 8490 1377
rect 8524 1343 8537 1377
rect 8477 1294 8537 1343
rect 8477 1260 8490 1294
rect 8524 1260 8537 1294
rect 8477 1248 8537 1260
rect 8567 1460 8624 1472
rect 8784 1464 8841 1472
rect 8567 1426 8580 1460
rect 8614 1426 8624 1460
rect 8567 1390 8624 1426
rect 8567 1356 8580 1390
rect 8614 1356 8624 1390
rect 8567 1320 8624 1356
rect 8567 1286 8580 1320
rect 8614 1286 8624 1320
rect 8567 1248 8624 1286
rect 8678 1452 8736 1464
rect 8678 1418 8689 1452
rect 8723 1418 8736 1452
rect 8678 1381 8736 1418
rect 8678 1347 8689 1381
rect 8723 1347 8736 1381
rect 8678 1310 8736 1347
rect 8678 1276 8689 1310
rect 8723 1276 8736 1310
rect 8678 1264 8736 1276
rect 8766 1456 8841 1464
rect 8766 1422 8794 1456
rect 8828 1422 8841 1456
rect 8766 1378 8841 1422
rect 8766 1344 8794 1378
rect 8828 1344 8841 1378
rect 8766 1306 8841 1344
rect 8766 1272 8794 1306
rect 8828 1272 8841 1306
rect 8766 1264 8841 1272
rect 8788 1248 8841 1264
rect 8871 1460 8931 1472
rect 8871 1426 8884 1460
rect 8918 1426 8931 1460
rect 8871 1377 8931 1426
rect 8871 1343 8884 1377
rect 8918 1343 8931 1377
rect 8871 1294 8931 1343
rect 8871 1260 8884 1294
rect 8918 1260 8931 1294
rect 8871 1248 8931 1260
rect 8961 1460 9020 1472
rect 8961 1426 8974 1460
rect 9008 1426 9020 1460
rect 8961 1377 9020 1426
rect 8961 1343 8974 1377
rect 9008 1343 9020 1377
rect 8961 1294 9020 1343
rect 8961 1260 8974 1294
rect 9008 1260 9020 1294
rect 8961 1248 9020 1260
rect 9074 1464 9212 1472
rect 9074 1430 9090 1464
rect 9124 1430 9162 1464
rect 9196 1430 9212 1464
rect 9654 1460 9713 1472
rect 9654 1457 9666 1460
rect 9074 1248 9212 1430
rect 9267 1445 9326 1457
rect 9267 1411 9279 1445
rect 9313 1411 9326 1445
rect 9267 1335 9326 1411
rect 9267 1301 9279 1335
rect 9313 1301 9326 1335
rect 9267 1289 9326 1301
rect 9356 1445 9416 1457
rect 9356 1411 9369 1445
rect 9403 1411 9416 1445
rect 9356 1335 9416 1411
rect 9356 1301 9369 1335
rect 9403 1301 9416 1335
rect 9356 1289 9416 1301
rect 9446 1448 9511 1457
rect 9446 1414 9459 1448
rect 9493 1414 9511 1448
rect 9446 1380 9511 1414
rect 9446 1346 9459 1380
rect 9493 1346 9511 1380
rect 9446 1289 9511 1346
rect 9541 1445 9606 1457
rect 9541 1411 9559 1445
rect 9593 1411 9606 1445
rect 9541 1335 9606 1411
rect 9541 1301 9559 1335
rect 9593 1301 9606 1335
rect 9541 1289 9606 1301
rect 9636 1426 9666 1457
rect 9700 1426 9713 1460
rect 9636 1388 9713 1426
rect 9636 1354 9666 1388
rect 9700 1354 9713 1388
rect 9636 1289 9713 1354
rect 9660 1248 9713 1289
rect 9743 1460 9807 1472
rect 9743 1426 9760 1460
rect 9794 1426 9807 1460
rect 9743 1379 9807 1426
rect 9743 1345 9760 1379
rect 9794 1345 9807 1379
rect 9743 1299 9807 1345
rect 9743 1265 9760 1299
rect 9794 1265 9807 1299
rect 9743 1248 9807 1265
rect 9837 1460 9897 1472
rect 9837 1426 9850 1460
rect 9884 1426 9897 1460
rect 9837 1367 9897 1426
rect 9837 1333 9850 1367
rect 9884 1333 9897 1367
rect 9837 1248 9897 1333
rect 9927 1460 9987 1472
rect 9927 1426 9940 1460
rect 9974 1426 9987 1460
rect 9927 1379 9987 1426
rect 9927 1345 9940 1379
rect 9974 1345 9987 1379
rect 9927 1299 9987 1345
rect 9927 1265 9940 1299
rect 9974 1265 9987 1299
rect 9927 1248 9987 1265
rect 10017 1460 10076 1472
rect 10017 1426 10030 1460
rect 10064 1426 10076 1460
rect 10017 1377 10076 1426
rect 10017 1343 10030 1377
rect 10064 1343 10076 1377
rect 10017 1294 10076 1343
rect 10017 1260 10030 1294
rect 10064 1260 10076 1294
rect 10017 1248 10076 1260
rect 10295 -804 10495 -796
rect 10295 -838 10307 -804
rect 10341 -838 10375 -804
rect 10409 -838 10443 -804
rect 10477 -838 10495 -804
rect 10295 -848 10495 -838
rect 10295 -888 10495 -878
rect 10295 -922 10307 -888
rect 10341 -922 10375 -888
rect 10409 -922 10443 -888
rect 10477 -922 10495 -888
rect 10295 -930 10495 -922
rect 6083 -6897 6141 -6885
rect 6083 -8873 6095 -6897
rect 6129 -8873 6141 -6897
rect 6083 -8885 6141 -8873
rect 6201 -6897 6259 -6885
rect 6201 -8873 6213 -6897
rect 6247 -8873 6259 -6897
rect 6201 -8885 6259 -8873
rect 6319 -6897 6377 -6885
rect 6319 -8873 6331 -6897
rect 6365 -8873 6377 -6897
rect 6319 -8885 6377 -8873
rect 6437 -6897 6495 -6885
rect 6437 -8873 6449 -6897
rect 6483 -8873 6495 -6897
rect 6437 -8885 6495 -8873
rect 6555 -6897 6613 -6885
rect 6555 -8873 6567 -6897
rect 6601 -8873 6613 -6897
rect 6555 -8885 6613 -8873
rect 6673 -6897 6731 -6885
rect 6673 -8873 6685 -6897
rect 6719 -8873 6731 -6897
rect 6673 -8885 6731 -8873
rect 6791 -6897 6849 -6885
rect 6791 -8873 6803 -6897
rect 6837 -8873 6849 -6897
rect 6791 -8885 6849 -8873
rect 6909 -6897 6967 -6885
rect 6909 -8873 6921 -6897
rect 6955 -8873 6967 -6897
rect 6909 -8885 6967 -8873
rect 7027 -6897 7085 -6885
rect 7027 -8873 7039 -6897
rect 7073 -8873 7085 -6897
rect 7027 -8885 7085 -8873
rect 7145 -6897 7203 -6885
rect 7145 -8873 7157 -6897
rect 7191 -8873 7203 -6897
rect 7145 -8885 7203 -8873
rect 7263 -6897 7321 -6885
rect 7263 -8873 7275 -6897
rect 7309 -8873 7321 -6897
rect 7263 -8885 7321 -8873
rect 7381 -6897 7439 -6885
rect 7381 -8873 7393 -6897
rect 7427 -8873 7439 -6897
rect 7381 -8885 7439 -8873
rect 7499 -6897 7557 -6885
rect 7499 -8873 7511 -6897
rect 7545 -8873 7557 -6897
rect 7499 -8885 7557 -8873
rect 7617 -6897 7675 -6885
rect 7617 -8873 7629 -6897
rect 7663 -8873 7675 -6897
rect 7617 -8885 7675 -8873
rect 7735 -6897 7793 -6885
rect 7735 -8873 7747 -6897
rect 7781 -8873 7793 -6897
rect 7735 -8885 7793 -8873
rect 7853 -6897 7911 -6885
rect 7853 -8873 7865 -6897
rect 7899 -8873 7911 -6897
rect 7853 -8885 7911 -8873
rect 7971 -6897 8029 -6885
rect 7971 -8873 7983 -6897
rect 8017 -8873 8029 -6897
rect 7971 -8885 8029 -8873
rect 8089 -6897 8147 -6885
rect 8089 -8873 8101 -6897
rect 8135 -8873 8147 -6897
rect 8089 -8885 8147 -8873
rect 8207 -6897 8265 -6885
rect 8207 -8873 8219 -6897
rect 8253 -8873 8265 -6897
rect 8207 -8885 8265 -8873
rect 8325 -6897 8383 -6885
rect 8325 -8873 8337 -6897
rect 8371 -8873 8383 -6897
rect 8325 -8885 8383 -8873
rect 8443 -6897 8501 -6885
rect 8443 -8873 8455 -6897
rect 8489 -8873 8501 -6897
rect 8443 -8885 8501 -8873
rect 8561 -6897 8619 -6885
rect 8561 -8873 8573 -6897
rect 8607 -8873 8619 -6897
rect 8561 -8885 8619 -8873
rect 8679 -6897 8737 -6885
rect 8679 -8873 8691 -6897
rect 8725 -8873 8737 -6897
rect 8679 -8885 8737 -8873
rect 8797 -6897 8855 -6885
rect 8797 -8873 8809 -6897
rect 8843 -8873 8855 -6897
rect 8797 -8885 8855 -8873
rect 8915 -6897 8973 -6885
rect 8915 -8873 8927 -6897
rect 8961 -8873 8973 -6897
rect 8915 -8885 8973 -8873
rect 9033 -6897 9091 -6885
rect 9033 -8873 9045 -6897
rect 9079 -8873 9091 -6897
rect 9033 -8885 9091 -8873
rect 9151 -6897 9209 -6885
rect 9151 -8873 9163 -6897
rect 9197 -8873 9209 -6897
rect 9151 -8885 9209 -8873
rect 9269 -6897 9327 -6885
rect 9269 -8873 9281 -6897
rect 9315 -8873 9327 -6897
rect 9269 -8885 9327 -8873
rect 9387 -6897 9445 -6885
rect 9387 -8873 9399 -6897
rect 9433 -8873 9445 -6897
rect 9387 -8885 9445 -8873
rect 9505 -6897 9563 -6885
rect 9505 -8873 9517 -6897
rect 9551 -8873 9563 -6897
rect 9505 -8885 9563 -8873
rect 9623 -6897 9681 -6885
rect 9623 -8873 9635 -6897
rect 9669 -8873 9681 -6897
rect 9623 -8885 9681 -8873
rect 9741 -6897 9799 -6885
rect 9741 -8873 9753 -6897
rect 9787 -8873 9799 -6897
rect 9741 -8885 9799 -8873
rect 9859 -6897 9917 -6885
rect 9859 -8873 9871 -6897
rect 9905 -8873 9917 -6897
rect 9859 -8885 9917 -8873
<< ndiffc >>
rect 5859 7788 5893 9764
rect 5977 7788 6011 9764
rect 6095 7788 6129 9764
rect 6213 7788 6247 9764
rect 6331 7788 6365 9764
rect 6449 7788 6483 9764
rect 6567 7788 6601 9764
rect 7023 9112 7057 9588
rect 7119 9112 7153 9588
rect 7215 9112 7249 9588
rect 7311 9112 7345 9588
rect 7407 9112 7441 9588
rect 7503 9112 7537 9588
rect 7599 9112 7633 9588
rect 7695 9112 7729 9588
rect 7791 9112 7825 9588
rect 7887 9112 7921 9588
rect 7983 9112 8017 9588
rect 8079 9112 8113 9588
rect 8175 9112 8209 9588
rect 8271 9112 8305 9588
rect 8367 9112 8401 9588
rect 8463 9112 8497 9588
rect 8559 9112 8593 9588
rect 8655 9112 8689 9588
rect 8751 9112 8785 9588
rect 8847 9112 8881 9588
rect 8943 9112 8977 9588
rect 7067 6672 7101 8648
rect 7525 6672 7559 8648
rect 7983 6672 8017 8648
rect 8441 6672 8475 8648
rect 8899 6672 8933 8648
rect 9400 7788 9434 9764
rect 9518 7788 9552 9764
rect 9636 7788 9670 9764
rect 9754 7788 9788 9764
rect 9872 7788 9906 9764
rect 9990 7788 10024 9764
rect 10108 7788 10142 9764
rect 10864 7268 11340 7302
rect 10864 7172 11340 7206
rect 10864 7076 11340 7110
rect 10864 6980 11340 7014
rect 10864 6884 11340 6918
rect 3469 3964 3503 4340
rect 3557 3964 3591 4340
rect 3469 3250 3503 3626
rect 3557 3250 3591 3626
rect 4251 3964 4285 4340
rect 4339 3964 4373 4340
rect 4251 3250 4285 3626
rect 4339 3250 4373 3626
rect 2440 2388 2474 2422
rect 2440 2298 2474 2332
rect 2540 2388 2574 2422
rect 3809 2380 3843 2414
rect 2540 2298 2574 2332
rect 3809 2298 3843 2332
rect 3973 2380 4007 2414
rect 3973 2298 4007 2332
rect 4105 2323 4139 2357
rect 4361 2323 4395 2357
rect 4617 2323 4651 2357
rect 5449 2323 5483 2357
rect 5705 2323 5739 2357
rect 5961 2323 5995 2357
rect 6121 2323 6155 2357
rect 6377 2323 6411 2357
rect 6633 2323 6667 2357
rect 6793 2323 6827 2357
rect 7049 2323 7083 2357
rect 7305 2323 7339 2357
rect 8137 2323 8171 2357
rect 8393 2323 8427 2357
rect 8649 2323 8683 2357
rect 8809 2323 8843 2357
rect 9065 2323 9099 2357
rect 9321 2323 9355 2357
rect 9481 2323 9515 2357
rect 9737 2323 9771 2357
rect 2440 2092 2474 2126
rect 2440 2002 2474 2036
rect 2540 2092 2574 2126
rect 3809 2092 3843 2126
rect 2540 2002 2574 2036
rect 3809 2010 3843 2044
rect 3973 2092 4007 2126
rect 3973 2010 4007 2044
rect 4094 2028 4128 2062
rect 4201 2092 4235 2126
rect 4183 2002 4217 2036
rect 4396 2084 4430 2118
rect 4730 2066 4764 2100
rect 4844 2092 4878 2126
rect 4844 2002 4878 2036
rect 4961 2092 4995 2126
rect 4961 2002 4995 2036
rect 5047 2092 5081 2126
rect 5047 2002 5081 2036
rect 5133 2092 5167 2126
rect 5133 2002 5167 2036
rect 6201 2130 6235 2164
rect 5443 2042 5477 2076
rect 5607 2037 5641 2071
rect 5687 2037 5721 2071
rect 5851 2043 5885 2077
rect 5987 2032 6021 2066
rect 6099 1978 6133 2012
rect 6353 2043 6387 2077
rect 6353 1975 6387 2009
rect 6491 2094 6525 2128
rect 6893 2093 6927 2127
rect 6672 2028 6706 2062
rect 6772 2033 6806 2067
rect 7005 2023 7039 2057
rect 7115 2041 7149 2075
rect 7226 2041 7260 2075
rect 7407 2058 7441 2092
rect 7489 2058 7523 2092
rect 7571 2058 7605 2092
rect 7755 2126 7789 2160
rect 7871 2092 7905 2126
rect 7966 2040 8000 2074
rect 8068 2113 8102 2147
rect 8385 2092 8419 2126
rect 8179 1961 8213 1995
rect 8385 2002 8419 2036
rect 8471 2092 8505 2126
rect 8471 2002 8505 2036
rect 8557 2092 8591 2126
rect 8557 2002 8591 2036
rect 8683 2066 8717 2100
rect 8683 1998 8717 2032
rect 8789 2092 8823 2126
rect 8789 2018 8823 2052
rect 8889 2092 8923 2126
rect 8889 2018 8923 2052
rect 8975 2092 9009 2126
rect 8975 2002 9009 2036
rect 9090 2096 9124 2130
rect 9162 2096 9196 2130
rect 9278 2092 9312 2126
rect 9278 2002 9312 2036
rect 9364 2070 9398 2104
rect 9450 2092 9484 2126
rect 9450 2002 9484 2036
rect 9536 2070 9570 2104
rect 9622 2092 9656 2126
rect 9622 2002 9656 2036
rect 9722 2038 9756 2072
rect 9822 2070 9856 2104
rect 9926 2038 9960 2072
rect 10030 2070 10064 2104
rect 3592 1056 3626 1090
rect 3592 966 3626 1000
rect 3692 1056 3726 1090
rect 4961 1048 4995 1082
rect 3692 966 3726 1000
rect 4961 966 4995 1000
rect 5125 1048 5159 1082
rect 5125 966 5159 1000
rect 5443 1016 5477 1050
rect 5607 1021 5641 1055
rect 5687 1021 5721 1055
rect 5851 1015 5885 1049
rect 5987 1026 6021 1060
rect 6099 1080 6133 1114
rect 6353 1083 6387 1117
rect 6353 1015 6387 1049
rect 6672 1030 6706 1064
rect 6772 1025 6806 1059
rect 7005 1035 7039 1069
rect 7115 1017 7149 1051
rect 7226 1017 7260 1051
rect 6201 928 6235 962
rect 6491 964 6525 998
rect 6893 965 6927 999
rect 7407 1000 7441 1034
rect 7489 1000 7523 1034
rect 7571 1000 7605 1034
rect 7755 932 7789 966
rect 7871 966 7905 1000
rect 7966 1018 8000 1052
rect 8179 1097 8213 1131
rect 8385 1056 8419 1090
rect 8068 945 8102 979
rect 8385 966 8419 1000
rect 8471 1056 8505 1090
rect 8471 966 8505 1000
rect 8557 1056 8591 1090
rect 8557 966 8591 1000
rect 8683 1060 8717 1094
rect 8683 992 8717 1026
rect 8789 1040 8823 1074
rect 8789 966 8823 1000
rect 8889 1040 8923 1074
rect 8889 966 8923 1000
rect 8975 1056 9009 1090
rect 8975 966 9009 1000
rect 9278 1081 9312 1115
rect 9278 1011 9312 1045
rect 9368 1014 9402 1048
rect 9454 1085 9488 1119
rect 9454 1007 9488 1041
rect 9554 1075 9588 1109
rect 9554 1007 9588 1041
rect 9656 1081 9690 1115
rect 9656 1003 9690 1037
rect 9090 962 9124 996
rect 9162 962 9196 996
rect 9758 1065 9792 1099
rect 9758 991 9792 1025
rect 9858 997 9892 1031
rect 9944 1081 9978 1115
rect 9944 991 9978 1025
rect 10030 1081 10064 1115
rect 10030 991 10064 1025
rect 3818 194 3852 570
rect 3906 194 3940 570
rect 10458 320 10492 1296
rect 10916 320 10950 1296
rect 11374 320 11408 1296
rect 11832 320 11866 1296
rect 12290 320 12324 1296
rect 12748 320 12782 1296
rect 13206 320 13240 1296
rect 13664 320 13698 1296
rect 13892 320 13926 1296
rect 13980 320 14014 1296
rect 14208 320 14242 1296
rect 14296 320 14330 1296
rect 15552 867 15928 901
rect 15552 779 15928 813
rect 16266 867 16642 901
rect 16266 779 16642 813
rect 16980 867 17356 901
rect 16980 779 17356 813
rect 17694 867 18070 901
rect 17694 779 18070 813
rect 18408 867 18784 901
rect 18408 779 18784 813
rect 19122 867 19498 901
rect 19122 779 19498 813
rect 19836 867 20212 901
rect 19836 779 20212 813
rect 20550 867 20926 901
rect 20550 779 20926 813
rect 21264 867 21640 901
rect 21264 779 21640 813
rect 21978 867 22354 901
rect 21978 779 22354 813
rect 22692 867 23068 901
rect 22692 779 23068 813
rect 23406 867 23782 901
rect 23406 779 23782 813
rect 24120 867 24496 901
rect 24120 779 24496 813
rect 24834 867 25210 901
rect 24834 779 25210 813
rect 25548 867 25924 901
rect 25548 779 25924 813
rect 26262 867 26638 901
rect 26262 779 26638 813
rect 26976 867 27352 901
rect 26976 779 27352 813
rect 27690 867 28066 901
rect 27690 779 28066 813
rect 28404 867 28780 901
rect 28404 779 28780 813
rect 29118 867 29494 901
rect 29118 779 29494 813
rect 29832 867 30208 901
rect 29832 779 30208 813
rect 30546 867 30922 901
rect 30546 779 30922 813
rect 31260 867 31636 901
rect 31260 779 31636 813
rect 31974 867 32350 901
rect 31974 779 32350 813
rect 32688 867 33064 901
rect 32688 779 33064 813
rect 33402 867 33778 901
rect 33402 779 33778 813
rect 34116 867 34492 901
rect 34116 779 34492 813
rect 34830 867 35206 901
rect 34830 779 35206 813
rect 35544 867 35920 901
rect 35544 779 35920 813
rect 36258 867 36634 901
rect 36258 779 36634 813
rect 36972 867 37348 901
rect 36972 779 37348 813
rect 37686 867 38062 901
rect 37686 779 38062 813
rect 38400 867 38776 901
rect 38400 779 38776 813
rect 3818 -520 3852 -144
rect 3906 -520 3940 -144
rect 15552 49 15928 83
rect 15552 -39 15928 -5
rect 16266 49 16642 83
rect 16266 -39 16642 -5
rect 16980 49 17356 83
rect 16980 -39 17356 -5
rect 17694 49 18070 83
rect 17694 -39 18070 -5
rect 18408 49 18784 83
rect 18408 -39 18784 -5
rect 19122 49 19498 83
rect 19122 -39 19498 -5
rect 19836 49 20212 83
rect 19836 -39 20212 -5
rect 20550 49 20926 83
rect 20550 -39 20926 -5
rect 21264 49 21640 83
rect 21264 -39 21640 -5
rect 21978 49 22354 83
rect 21978 -39 22354 -5
rect 22692 49 23068 83
rect 22692 -39 23068 -5
rect 23406 49 23782 83
rect 23406 -39 23782 -5
rect 24120 49 24496 83
rect 24120 -39 24496 -5
rect 24834 49 25210 83
rect 24834 -39 25210 -5
rect 25548 49 25924 83
rect 25548 -39 25924 -5
rect 26262 49 26638 83
rect 26262 -39 26638 -5
rect 26976 49 27352 83
rect 26976 -39 27352 -5
rect 27690 49 28066 83
rect 27690 -39 28066 -5
rect 28404 49 28780 83
rect 28404 -39 28780 -5
rect 29118 49 29494 83
rect 29118 -39 29494 -5
rect 29832 49 30208 83
rect 29832 -39 30208 -5
rect 30546 49 30922 83
rect 30546 -39 30922 -5
rect 31260 49 31636 83
rect 31260 -39 31636 -5
rect 31974 49 32350 83
rect 31974 -39 32350 -5
rect 32688 49 33064 83
rect 32688 -39 33064 -5
rect 33402 49 33778 83
rect 33402 -39 33778 -5
rect 34116 49 34492 83
rect 34116 -39 34492 -5
rect 34830 49 35206 83
rect 34830 -39 35206 -5
rect 35544 49 35920 83
rect 35544 -39 35920 -5
rect 36258 49 36634 83
rect 36258 -39 36634 -5
rect 36972 49 37348 83
rect 36972 -39 37348 -5
rect 37686 49 38062 83
rect 37686 -39 38062 -5
rect 38400 49 38776 83
rect 38400 -39 38776 -5
rect 10627 -838 10661 -804
rect 10695 -838 10729 -804
rect 10627 -922 10661 -888
rect 10695 -922 10729 -888
rect 5859 -6364 5893 -4388
rect 5977 -6364 6011 -4388
rect 6095 -6364 6129 -4388
rect 6213 -6364 6247 -4388
rect 6331 -6364 6365 -4388
rect 6449 -6364 6483 -4388
rect 6567 -6364 6601 -4388
rect 7067 -5248 7101 -3272
rect 7525 -5248 7559 -3272
rect 7983 -5248 8017 -3272
rect 8441 -5248 8475 -3272
rect 8899 -5248 8933 -3272
rect 10864 -3518 11340 -3484
rect 10864 -3614 11340 -3580
rect 10864 -3710 11340 -3676
rect 10864 -3806 11340 -3772
rect 10864 -3902 11340 -3868
rect 7023 -6188 7057 -5712
rect 7119 -6188 7153 -5712
rect 7215 -6188 7249 -5712
rect 7311 -6188 7345 -5712
rect 7407 -6188 7441 -5712
rect 7503 -6188 7537 -5712
rect 7599 -6188 7633 -5712
rect 7695 -6188 7729 -5712
rect 7791 -6188 7825 -5712
rect 7887 -6188 7921 -5712
rect 7983 -6188 8017 -5712
rect 8079 -6188 8113 -5712
rect 8175 -6188 8209 -5712
rect 8271 -6188 8305 -5712
rect 8367 -6188 8401 -5712
rect 8463 -6188 8497 -5712
rect 8559 -6188 8593 -5712
rect 8655 -6188 8689 -5712
rect 8751 -6188 8785 -5712
rect 8847 -6188 8881 -5712
rect 8943 -6188 8977 -5712
rect 9400 -6364 9434 -4388
rect 9518 -6364 9552 -4388
rect 9636 -6364 9670 -4388
rect 9754 -6364 9788 -4388
rect 9872 -6364 9906 -4388
rect 9990 -6364 10024 -4388
rect 10108 -6364 10142 -4388
<< pdiffc >>
rect 6095 10297 6129 12273
rect 6213 10297 6247 12273
rect 6331 10297 6365 12273
rect 6449 10297 6483 12273
rect 6567 10297 6601 12273
rect 6685 10297 6719 12273
rect 6803 10297 6837 12273
rect 6921 10297 6955 12273
rect 7039 10297 7073 12273
rect 7157 10297 7191 12273
rect 7275 10297 7309 12273
rect 7393 10297 7427 12273
rect 7511 10297 7545 12273
rect 7629 10297 7663 12273
rect 7747 10297 7781 12273
rect 7865 10297 7899 12273
rect 7983 10297 8017 12273
rect 8101 10297 8135 12273
rect 8219 10297 8253 12273
rect 8337 10297 8371 12273
rect 8455 10297 8489 12273
rect 8573 10297 8607 12273
rect 8691 10297 8725 12273
rect 8809 10297 8843 12273
rect 8927 10297 8961 12273
rect 9045 10297 9079 12273
rect 9163 10297 9197 12273
rect 9281 10297 9315 12273
rect 9399 10297 9433 12273
rect 9517 10297 9551 12273
rect 9635 10297 9669 12273
rect 9753 10297 9787 12273
rect 9871 10297 9905 12273
rect 2440 2758 2474 2792
rect 2440 2688 2474 2722
rect 2440 2618 2474 2652
rect 2540 2758 2574 2792
rect 2540 2675 2574 2709
rect 3804 2758 3838 2792
rect 3804 2675 3838 2709
rect 2540 2592 2574 2626
rect 3804 2592 3838 2626
rect 3894 2758 3928 2792
rect 3894 2675 3928 2709
rect 3894 2592 3928 2626
rect 3984 2758 4018 2792
rect 3984 2675 4018 2709
rect 3984 2592 4018 2626
rect 4090 2758 4124 2792
rect 4090 2687 4124 2721
rect 4090 2616 4124 2650
rect 4348 2758 4382 2792
rect 4348 2687 4382 2721
rect 4348 2616 4382 2650
rect 4603 2758 4637 2792
rect 4603 2687 4637 2721
rect 4603 2616 4637 2650
rect 5434 2758 5468 2792
rect 5434 2687 5468 2721
rect 5434 2616 5468 2650
rect 5692 2758 5726 2792
rect 5692 2687 5726 2721
rect 5692 2616 5726 2650
rect 5947 2758 5981 2792
rect 5947 2687 5981 2721
rect 5947 2616 5981 2650
rect 6106 2758 6140 2792
rect 6106 2687 6140 2721
rect 6106 2616 6140 2650
rect 6364 2758 6398 2792
rect 6364 2687 6398 2721
rect 6364 2616 6398 2650
rect 6619 2758 6653 2792
rect 6619 2687 6653 2721
rect 6619 2616 6653 2650
rect 6778 2758 6812 2792
rect 6778 2687 6812 2721
rect 6778 2616 6812 2650
rect 7036 2758 7070 2792
rect 7036 2687 7070 2721
rect 7036 2616 7070 2650
rect 7291 2758 7325 2792
rect 7291 2687 7325 2721
rect 7291 2616 7325 2650
rect 8122 2758 8156 2792
rect 8122 2687 8156 2721
rect 8122 2616 8156 2650
rect 8380 2758 8414 2792
rect 8380 2687 8414 2721
rect 8380 2616 8414 2650
rect 8635 2758 8669 2792
rect 8635 2687 8669 2721
rect 8635 2616 8669 2650
rect 8794 2758 8828 2792
rect 8794 2687 8828 2721
rect 8794 2616 8828 2650
rect 9052 2758 9086 2792
rect 9052 2687 9086 2721
rect 9052 2616 9086 2650
rect 9307 2758 9341 2792
rect 9307 2687 9341 2721
rect 9307 2616 9341 2650
rect 9466 2758 9500 2792
rect 9466 2687 9500 2721
rect 9466 2616 9500 2650
rect 9724 2758 9758 2792
rect 9724 2687 9758 2721
rect 9724 2616 9758 2650
rect 2440 1772 2474 1806
rect 2440 1702 2474 1736
rect 2440 1632 2474 1666
rect 2540 1798 2574 1832
rect 3804 1798 3838 1832
rect 2540 1715 2574 1749
rect 2540 1632 2574 1666
rect 3804 1715 3838 1749
rect 3804 1632 3838 1666
rect 3894 1798 3928 1832
rect 3894 1715 3928 1749
rect 3894 1632 3928 1666
rect 3984 1798 4018 1832
rect 3984 1715 4018 1749
rect 4094 1783 4128 1817
rect 4094 1688 4128 1722
rect 4201 1693 4235 1727
rect 3984 1632 4018 1666
rect 4484 1798 4518 1832
rect 4484 1681 4518 1715
rect 4730 1798 4764 1832
rect 4730 1715 4764 1749
rect 4730 1632 4764 1666
rect 4830 1798 4864 1832
rect 4830 1715 4864 1749
rect 4830 1632 4864 1666
rect 4956 1772 4990 1806
rect 4956 1702 4990 1736
rect 4956 1632 4990 1666
rect 5046 1798 5080 1832
rect 5046 1715 5080 1749
rect 5046 1632 5080 1666
rect 5136 1798 5170 1832
rect 5136 1715 5170 1749
rect 5136 1632 5170 1666
rect 6100 1772 6134 1806
rect 5438 1701 5472 1735
rect 5438 1632 5472 1666
rect 5528 1633 5562 1667
rect 5696 1692 5730 1726
rect 5786 1702 5820 1736
rect 5786 1632 5820 1666
rect 5898 1702 5932 1736
rect 5898 1632 5932 1666
rect 5988 1702 6022 1736
rect 5988 1632 6022 1666
rect 6100 1702 6134 1736
rect 6100 1632 6134 1666
rect 6190 1710 6224 1744
rect 6190 1632 6224 1666
rect 6280 1794 6314 1828
rect 6280 1713 6314 1747
rect 6280 1632 6314 1666
rect 6392 1684 6426 1718
rect 6583 1692 6617 1726
rect 6683 1692 6717 1726
rect 6795 1632 6829 1666
rect 6914 1632 6948 1666
rect 7088 1669 7122 1703
rect 7196 1742 7230 1776
rect 7196 1632 7230 1666
rect 7308 1704 7342 1738
rect 7308 1632 7342 1666
rect 7476 1742 7510 1776
rect 7776 1710 7810 1744
rect 7476 1632 7510 1666
rect 7661 1637 7695 1671
rect 7776 1632 7810 1666
rect 7876 1637 7910 1671
rect 8052 1750 8086 1784
rect 8164 1761 8198 1795
rect 8383 1765 8417 1799
rect 8052 1632 8086 1666
rect 8383 1683 8417 1717
rect 8271 1593 8305 1627
rect 8383 1593 8417 1627
rect 8490 1798 8524 1832
rect 8490 1715 8524 1749
rect 8490 1632 8524 1666
rect 8580 1772 8614 1806
rect 8580 1702 8614 1736
rect 8580 1632 8614 1666
rect 8689 1782 8723 1816
rect 8689 1711 8723 1745
rect 8689 1640 8723 1674
rect 8794 1786 8828 1820
rect 8794 1714 8828 1748
rect 8794 1636 8828 1670
rect 8884 1798 8918 1832
rect 8884 1715 8918 1749
rect 8884 1632 8918 1666
rect 8974 1798 9008 1832
rect 8974 1715 9008 1749
rect 8974 1632 9008 1666
rect 9090 1628 9124 1662
rect 9162 1628 9196 1662
rect 9278 1792 9312 1826
rect 9278 1712 9312 1746
rect 9278 1632 9312 1666
rect 9369 1772 9403 1806
rect 9449 1772 9483 1806
rect 9531 1772 9565 1806
rect 9369 1701 9403 1735
rect 9449 1701 9483 1735
rect 9531 1701 9565 1735
rect 9369 1632 9403 1666
rect 9449 1632 9483 1666
rect 9531 1632 9565 1666
rect 9621 1711 9655 1745
rect 9621 1632 9655 1666
rect 9721 1772 9755 1806
rect 9790 1772 9824 1806
rect 9861 1772 9895 1806
rect 9930 1772 9964 1806
rect 9721 1701 9755 1735
rect 9790 1701 9824 1735
rect 9861 1701 9895 1735
rect 9930 1701 9964 1735
rect 9721 1632 9755 1666
rect 9790 1632 9824 1666
rect 9861 1632 9895 1666
rect 9930 1632 9964 1666
rect 10030 1711 10064 1745
rect 10030 1632 10064 1666
rect 11374 1749 11408 3725
rect 11832 1749 11866 3725
rect 12290 1749 12324 3725
rect 12748 1749 12782 3725
rect 13206 1749 13240 3725
rect 13664 1749 13698 3725
rect 13892 1749 13926 3725
rect 13980 1749 14014 3725
rect 14208 1749 14242 3725
rect 14296 1749 14330 3725
rect 3592 1426 3626 1460
rect 3592 1356 3626 1390
rect 3592 1286 3626 1320
rect 3692 1426 3726 1460
rect 3692 1343 3726 1377
rect 4956 1426 4990 1460
rect 4956 1343 4990 1377
rect 3692 1260 3726 1294
rect 4956 1260 4990 1294
rect 5046 1426 5080 1460
rect 5046 1343 5080 1377
rect 5046 1260 5080 1294
rect 5136 1426 5170 1460
rect 5136 1343 5170 1377
rect 5438 1426 5472 1460
rect 5438 1357 5472 1391
rect 5528 1425 5562 1459
rect 5696 1366 5730 1400
rect 5786 1426 5820 1460
rect 5786 1356 5820 1390
rect 5898 1426 5932 1460
rect 5898 1356 5932 1390
rect 5988 1426 6022 1460
rect 5988 1356 6022 1390
rect 6100 1426 6134 1460
rect 6100 1356 6134 1390
rect 5136 1260 5170 1294
rect 6100 1286 6134 1320
rect 6190 1426 6224 1460
rect 6190 1348 6224 1382
rect 6280 1426 6314 1460
rect 6280 1345 6314 1379
rect 6392 1374 6426 1408
rect 6583 1366 6617 1400
rect 6683 1366 6717 1400
rect 6795 1426 6829 1460
rect 6914 1426 6948 1460
rect 6280 1264 6314 1298
rect 7088 1389 7122 1423
rect 7196 1426 7230 1460
rect 7196 1316 7230 1350
rect 7308 1426 7342 1460
rect 7308 1354 7342 1388
rect 7476 1426 7510 1460
rect 7661 1421 7695 1455
rect 7776 1426 7810 1460
rect 7476 1316 7510 1350
rect 7776 1348 7810 1382
rect 7876 1421 7910 1455
rect 8052 1426 8086 1460
rect 8271 1465 8305 1499
rect 8383 1465 8417 1499
rect 8052 1308 8086 1342
rect 8164 1297 8198 1331
rect 8383 1375 8417 1409
rect 8383 1293 8417 1327
rect 8490 1426 8524 1460
rect 8490 1343 8524 1377
rect 8490 1260 8524 1294
rect 8580 1426 8614 1460
rect 8580 1356 8614 1390
rect 8580 1286 8614 1320
rect 8689 1418 8723 1452
rect 8689 1347 8723 1381
rect 8689 1276 8723 1310
rect 8794 1422 8828 1456
rect 8794 1344 8828 1378
rect 8794 1272 8828 1306
rect 8884 1426 8918 1460
rect 8884 1343 8918 1377
rect 8884 1260 8918 1294
rect 8974 1426 9008 1460
rect 8974 1343 9008 1377
rect 8974 1260 9008 1294
rect 9090 1430 9124 1464
rect 9162 1430 9196 1464
rect 9279 1411 9313 1445
rect 9279 1301 9313 1335
rect 9369 1411 9403 1445
rect 9369 1301 9403 1335
rect 9459 1414 9493 1448
rect 9459 1346 9493 1380
rect 9559 1411 9593 1445
rect 9559 1301 9593 1335
rect 9666 1426 9700 1460
rect 9666 1354 9700 1388
rect 9760 1426 9794 1460
rect 9760 1345 9794 1379
rect 9760 1265 9794 1299
rect 9850 1426 9884 1460
rect 9850 1333 9884 1367
rect 9940 1426 9974 1460
rect 9940 1345 9974 1379
rect 9940 1265 9974 1299
rect 10030 1426 10064 1460
rect 10030 1343 10064 1377
rect 10030 1260 10064 1294
rect 10307 -838 10341 -804
rect 10375 -838 10409 -804
rect 10443 -838 10477 -804
rect 10307 -922 10341 -888
rect 10375 -922 10409 -888
rect 10443 -922 10477 -888
rect 6095 -8873 6129 -6897
rect 6213 -8873 6247 -6897
rect 6331 -8873 6365 -6897
rect 6449 -8873 6483 -6897
rect 6567 -8873 6601 -6897
rect 6685 -8873 6719 -6897
rect 6803 -8873 6837 -6897
rect 6921 -8873 6955 -6897
rect 7039 -8873 7073 -6897
rect 7157 -8873 7191 -6897
rect 7275 -8873 7309 -6897
rect 7393 -8873 7427 -6897
rect 7511 -8873 7545 -6897
rect 7629 -8873 7663 -6897
rect 7747 -8873 7781 -6897
rect 7865 -8873 7899 -6897
rect 7983 -8873 8017 -6897
rect 8101 -8873 8135 -6897
rect 8219 -8873 8253 -6897
rect 8337 -8873 8371 -6897
rect 8455 -8873 8489 -6897
rect 8573 -8873 8607 -6897
rect 8691 -8873 8725 -6897
rect 8809 -8873 8843 -6897
rect 8927 -8873 8961 -6897
rect 9045 -8873 9079 -6897
rect 9163 -8873 9197 -6897
rect 9281 -8873 9315 -6897
rect 9399 -8873 9433 -6897
rect 9517 -8873 9551 -6897
rect 9635 -8873 9669 -6897
rect 9753 -8873 9787 -6897
rect 9871 -8873 9905 -6897
<< psubdiff >>
rect 5745 9916 5841 9950
rect 6619 9916 6715 9950
rect 5745 9854 5779 9916
rect 5042 9548 5138 9582
rect 5578 9548 5674 9582
rect 5042 9486 5076 9548
rect 5640 9486 5674 9548
rect 5042 8320 5076 8382
rect 5640 8320 5674 8382
rect 5042 8286 5138 8320
rect 5578 8286 5674 8320
rect 6681 9854 6715 9916
rect 5745 7636 5779 7698
rect 9286 9916 9382 9950
rect 10160 9916 10256 9950
rect 9286 9854 9320 9916
rect 6909 9740 7005 9774
rect 8995 9740 9091 9774
rect 6909 9678 6943 9740
rect 9057 9678 9091 9740
rect 6909 8960 6943 9022
rect 9057 8960 9091 9022
rect 6909 8926 7005 8960
rect 8995 8926 9091 8960
rect 6681 7636 6715 7698
rect 5745 7602 5841 7636
rect 6619 7602 6715 7636
rect 6953 8800 7049 8834
rect 8951 8800 9047 8834
rect 6953 8738 6987 8800
rect 9013 8738 9047 8800
rect 6953 6520 6987 6582
rect 10222 9854 10256 9916
rect 9286 7636 9320 7698
rect 10222 7636 10256 7698
rect 9286 7602 9382 7636
rect 10160 7602 10256 7636
rect 9013 6520 9047 6582
rect 6953 6486 7049 6520
rect 8951 6486 9047 6520
rect 10678 7382 10774 7416
rect 11430 7382 11526 7416
rect 10678 7320 10712 7382
rect 11492 7320 11526 7382
rect 10678 6388 10712 6470
rect 11492 6388 11526 6470
rect 10678 6354 10774 6388
rect 11430 6354 11526 6388
rect 3355 4492 3451 4526
rect 3609 4492 3705 4526
rect 3355 4430 3389 4492
rect 3671 4430 3705 4492
rect 3355 3812 3389 3874
rect 3671 3812 3705 3874
rect 3355 3778 3451 3812
rect 3609 3778 3705 3812
rect 3355 3716 3389 3778
rect 3671 3716 3705 3778
rect 3355 3098 3389 3160
rect 3671 3098 3705 3160
rect 3355 3064 3451 3098
rect 3609 3064 3705 3098
rect 4137 4492 4233 4526
rect 4391 4492 4487 4526
rect 4137 4430 4171 4492
rect 4453 4430 4487 4492
rect 4137 3812 4171 3874
rect 4453 3812 4487 3874
rect 4137 3778 4233 3812
rect 4391 3778 4487 3812
rect 4137 3716 4171 3778
rect 4453 3716 4487 3778
rect 4137 3098 4171 3160
rect 4453 3098 4487 3160
rect 4137 3064 4233 3098
rect 4391 3064 4487 3098
rect 2070 2417 2104 2441
rect 2070 2334 2104 2383
rect 2070 2276 2104 2300
rect 10692 2716 10788 2750
rect 11092 2716 11188 2750
rect 10692 2654 10726 2716
rect 5238 2417 5368 2441
rect 5272 2383 5334 2417
rect 5238 2334 5368 2383
rect 9846 2417 9880 2441
rect 5272 2300 5334 2334
rect 5238 2276 5368 2300
rect 9846 2334 9880 2383
rect 9846 2276 9880 2300
rect 10134 2417 10168 2441
rect 10134 2334 10168 2383
rect 10134 2276 10168 2300
rect 2070 2124 2104 2148
rect 2070 2041 2104 2090
rect 2070 1983 2104 2007
rect 5238 2124 5368 2148
rect 5272 2090 5334 2124
rect 5238 2041 5368 2090
rect 5272 2007 5334 2041
rect 5238 1983 5368 2007
rect 10134 2124 10168 2148
rect 10134 2041 10168 2090
rect 10134 1983 10168 2007
rect 11154 2654 11188 2716
rect 10692 1588 10726 1650
rect 11154 1588 11188 1650
rect 10692 1554 10788 1588
rect 11092 1554 11188 1588
rect 3222 1085 3256 1109
rect 1796 1051 1830 1075
rect 1796 970 1830 1017
rect 2072 1051 2106 1075
rect 2072 970 2106 1017
rect 2164 1051 2198 1075
rect 2164 970 2198 1017
rect 2440 1051 2474 1075
rect 2440 970 2474 1017
rect 2532 1051 2566 1075
rect 2532 970 2566 1017
rect 2808 1051 2842 1075
rect 2808 970 2842 1017
rect 3222 1002 3256 1051
rect 3222 944 3256 968
rect 5238 1085 5368 1109
rect 5272 1051 5334 1085
rect 5238 1002 5368 1051
rect 5272 968 5334 1002
rect 5238 944 5368 968
rect 10344 1448 10440 1482
rect 13716 1448 13874 1482
rect 14032 1448 14190 1482
rect 14348 1448 14444 1482
rect 10344 1386 10378 1448
rect 10134 1085 10168 1109
rect 10134 1002 10168 1051
rect 10134 944 10168 968
rect 3704 722 3800 756
rect 3958 722 4054 756
rect 3704 660 3738 722
rect 4020 660 4054 722
rect 3704 42 3738 104
rect 13778 1386 13812 1448
rect 10344 168 10378 230
rect 14094 1386 14128 1448
rect 13778 168 13812 230
rect 14410 1386 14444 1448
rect 14094 168 14128 230
rect 39233 1141 39329 1175
rect 40361 1141 40457 1175
rect 39233 1079 39267 1141
rect 15366 981 15462 1015
rect 16018 981 16176 1015
rect 16732 981 16890 1015
rect 17446 981 17604 1015
rect 18160 981 18318 1015
rect 18874 981 19032 1015
rect 19588 981 19746 1015
rect 20302 981 20460 1015
rect 21016 981 21174 1015
rect 21730 981 21888 1015
rect 22444 981 22602 1015
rect 23158 981 23316 1015
rect 23872 981 24030 1015
rect 24586 981 24744 1015
rect 25300 981 25458 1015
rect 26014 981 26172 1015
rect 26728 981 26886 1015
rect 27442 981 27600 1015
rect 28156 981 28314 1015
rect 28870 981 29028 1015
rect 29584 981 29742 1015
rect 30298 981 30456 1015
rect 31012 981 31170 1015
rect 31726 981 31884 1015
rect 32440 981 32598 1015
rect 33154 981 33312 1015
rect 33868 981 34026 1015
rect 34582 981 34740 1015
rect 35296 981 35454 1015
rect 36010 981 36168 1015
rect 36724 981 36882 1015
rect 37438 981 37596 1015
rect 38152 981 38310 1015
rect 38866 981 38962 1015
rect 15366 919 15400 981
rect 16080 919 16114 981
rect 15366 699 15400 761
rect 16794 919 16828 981
rect 16080 699 16114 761
rect 17508 919 17542 981
rect 16794 699 16828 761
rect 18222 919 18256 981
rect 17508 699 17542 761
rect 18936 919 18970 981
rect 18222 699 18256 761
rect 19650 919 19684 981
rect 18936 699 18970 761
rect 20364 919 20398 981
rect 19650 699 19684 761
rect 21078 919 21112 981
rect 20364 699 20398 761
rect 21792 919 21826 981
rect 21078 699 21112 761
rect 22506 919 22540 981
rect 21792 699 21826 761
rect 23220 919 23254 981
rect 22506 699 22540 761
rect 23934 919 23968 981
rect 23220 699 23254 761
rect 24648 919 24682 981
rect 23934 699 23968 761
rect 25362 919 25396 981
rect 24648 699 24682 761
rect 26076 919 26110 981
rect 25362 699 25396 761
rect 26790 919 26824 981
rect 26076 699 26110 761
rect 27504 919 27538 981
rect 26790 699 26824 761
rect 28218 919 28252 981
rect 27504 699 27538 761
rect 28932 919 28966 981
rect 28218 699 28252 761
rect 29646 919 29680 981
rect 28932 699 28966 761
rect 30360 919 30394 981
rect 29646 699 29680 761
rect 31074 919 31108 981
rect 30360 699 30394 761
rect 31788 919 31822 981
rect 31074 699 31108 761
rect 32502 919 32536 981
rect 31788 699 31822 761
rect 33216 919 33250 981
rect 32502 699 32536 761
rect 33930 919 33964 981
rect 33216 699 33250 761
rect 34644 919 34678 981
rect 33930 699 33964 761
rect 35358 919 35392 981
rect 34644 699 34678 761
rect 36072 919 36106 981
rect 35358 699 35392 761
rect 36786 919 36820 981
rect 36072 699 36106 761
rect 37500 919 37534 981
rect 36786 699 36820 761
rect 38214 919 38248 981
rect 37500 699 37534 761
rect 38928 919 38962 981
rect 38214 699 38248 761
rect 38928 699 38962 761
rect 15366 665 15462 699
rect 16018 665 16176 699
rect 16732 665 16890 699
rect 17446 665 17604 699
rect 18160 665 18318 699
rect 18874 665 19032 699
rect 19588 665 19746 699
rect 20302 665 20460 699
rect 21016 665 21174 699
rect 21730 665 21888 699
rect 22444 665 22602 699
rect 23158 665 23316 699
rect 23872 665 24030 699
rect 24586 665 24744 699
rect 25300 665 25458 699
rect 26014 665 26172 699
rect 26728 665 26886 699
rect 27442 665 27600 699
rect 28156 665 28314 699
rect 28870 665 29028 699
rect 29584 665 29742 699
rect 30298 665 30456 699
rect 31012 665 31170 699
rect 31726 665 31884 699
rect 32440 665 32598 699
rect 33154 665 33312 699
rect 33868 665 34026 699
rect 34582 665 34740 699
rect 35296 665 35454 699
rect 36010 665 36168 699
rect 36724 665 36882 699
rect 37438 665 37596 699
rect 38152 665 38310 699
rect 38866 665 38962 699
rect 14410 168 14444 230
rect 10344 134 10440 168
rect 13716 134 13874 168
rect 14032 134 14190 168
rect 14348 134 14444 168
rect 15366 163 15462 197
rect 16018 163 16176 197
rect 16732 163 16890 197
rect 17446 163 17604 197
rect 18160 163 18318 197
rect 18874 163 19032 197
rect 19588 163 19746 197
rect 20302 163 20460 197
rect 21016 163 21174 197
rect 21730 163 21888 197
rect 22444 163 22602 197
rect 23158 163 23316 197
rect 23872 163 24030 197
rect 24586 163 24744 197
rect 25300 163 25458 197
rect 26014 163 26172 197
rect 26728 163 26886 197
rect 27442 163 27600 197
rect 28156 163 28314 197
rect 28870 163 29028 197
rect 29584 163 29742 197
rect 30298 163 30456 197
rect 31012 163 31170 197
rect 31726 163 31884 197
rect 32440 163 32598 197
rect 33154 163 33312 197
rect 33868 163 34026 197
rect 34582 163 34740 197
rect 35296 163 35454 197
rect 36010 163 36168 197
rect 36724 163 36882 197
rect 37438 163 37596 197
rect 38152 163 38310 197
rect 38866 163 38962 197
rect 4020 42 4054 104
rect 3704 8 3800 42
rect 3958 8 4054 42
rect 3704 -54 3738 8
rect 4020 -54 4054 8
rect 3704 -672 3738 -610
rect 15366 101 15400 163
rect 16080 101 16114 163
rect 15366 -119 15400 -57
rect 16794 101 16828 163
rect 16080 -119 16114 -57
rect 17508 101 17542 163
rect 16794 -119 16828 -57
rect 18222 101 18256 163
rect 17508 -119 17542 -57
rect 18936 101 18970 163
rect 18222 -119 18256 -57
rect 19650 101 19684 163
rect 18936 -119 18970 -57
rect 20364 101 20398 163
rect 19650 -119 19684 -57
rect 21078 101 21112 163
rect 20364 -119 20398 -57
rect 21792 101 21826 163
rect 21078 -119 21112 -57
rect 22506 101 22540 163
rect 21792 -119 21826 -57
rect 23220 101 23254 163
rect 22506 -119 22540 -57
rect 23934 101 23968 163
rect 23220 -119 23254 -57
rect 24648 101 24682 163
rect 23934 -119 23968 -57
rect 25362 101 25396 163
rect 24648 -119 24682 -57
rect 26076 101 26110 163
rect 25362 -119 25396 -57
rect 26790 101 26824 163
rect 26076 -119 26110 -57
rect 27504 101 27538 163
rect 26790 -119 26824 -57
rect 28218 101 28252 163
rect 27504 -119 27538 -57
rect 28932 101 28966 163
rect 28218 -119 28252 -57
rect 29646 101 29680 163
rect 28932 -119 28966 -57
rect 30360 101 30394 163
rect 29646 -119 29680 -57
rect 31074 101 31108 163
rect 30360 -119 30394 -57
rect 31788 101 31822 163
rect 31074 -119 31108 -57
rect 32502 101 32536 163
rect 31788 -119 31822 -57
rect 33216 101 33250 163
rect 32502 -119 32536 -57
rect 33930 101 33964 163
rect 33216 -119 33250 -57
rect 34644 101 34678 163
rect 33930 -119 33964 -57
rect 35358 101 35392 163
rect 34644 -119 34678 -57
rect 36072 101 36106 163
rect 35358 -119 35392 -57
rect 36786 101 36820 163
rect 36072 -119 36106 -57
rect 37500 101 37534 163
rect 36786 -119 36820 -57
rect 38214 101 38248 163
rect 37500 -119 37534 -57
rect 38928 101 38962 163
rect 38214 -119 38248 -57
rect 38928 -119 38962 -57
rect 15366 -153 15462 -119
rect 16018 -153 16176 -119
rect 16732 -153 16890 -119
rect 17446 -153 17604 -119
rect 18160 -153 18318 -119
rect 18874 -153 19032 -119
rect 19588 -153 19746 -119
rect 20302 -153 20460 -119
rect 21016 -153 21174 -119
rect 21730 -153 21888 -119
rect 22444 -153 22602 -119
rect 23158 -153 23316 -119
rect 23872 -153 24030 -119
rect 24586 -153 24744 -119
rect 25300 -153 25458 -119
rect 26014 -153 26172 -119
rect 26728 -153 26886 -119
rect 27442 -153 27600 -119
rect 28156 -153 28314 -119
rect 28870 -153 29028 -119
rect 29584 -153 29742 -119
rect 30298 -153 30456 -119
rect 31012 -153 31170 -119
rect 31726 -153 31884 -119
rect 32440 -153 32598 -119
rect 33154 -153 33312 -119
rect 33868 -153 34026 -119
rect 34582 -153 34740 -119
rect 35296 -153 35454 -119
rect 36010 -153 36168 -119
rect 36724 -153 36882 -119
rect 37438 -153 37596 -119
rect 38152 -153 38310 -119
rect 38866 -153 38962 -119
rect 40423 1079 40457 1141
rect 39233 -283 39267 -221
rect 40423 -283 40457 -221
rect 39233 -317 39329 -283
rect 40361 -317 40457 -283
rect 10623 -417 10647 -383
rect 10681 -417 10728 -383
rect 4020 -672 4054 -610
rect 3704 -706 3800 -672
rect 3958 -706 4054 -672
rect 10623 -693 10647 -659
rect 10681 -693 10728 -659
rect 10623 -1061 10647 -1027
rect 10681 -1061 10728 -1027
rect 10623 -1337 10647 -1303
rect 10681 -1337 10728 -1303
rect 10678 -2988 10774 -2954
rect 11430 -2988 11526 -2954
rect 10678 -3070 10712 -2988
rect 6953 -3120 7049 -3086
rect 8951 -3120 9047 -3086
rect 6953 -3182 6987 -3120
rect 5745 -4236 5841 -4202
rect 6619 -4236 6715 -4202
rect 5745 -4298 5779 -4236
rect 5042 -4920 5138 -4886
rect 5578 -4920 5674 -4886
rect 5042 -4982 5076 -4920
rect 5640 -4982 5674 -4920
rect 5042 -6148 5076 -6086
rect 5640 -6148 5674 -6086
rect 5042 -6182 5138 -6148
rect 5578 -6182 5674 -6148
rect 6681 -4298 6715 -4236
rect 5745 -6516 5779 -6454
rect 9013 -3182 9047 -3120
rect 6953 -5400 6987 -5338
rect 11492 -3070 11526 -2988
rect 10678 -3982 10712 -3920
rect 11492 -3982 11526 -3920
rect 10678 -4016 10774 -3982
rect 11430 -4016 11526 -3982
rect 9013 -5400 9047 -5338
rect 6953 -5434 7049 -5400
rect 8951 -5434 9047 -5400
rect 9286 -4236 9382 -4202
rect 10160 -4236 10256 -4202
rect 9286 -4298 9320 -4236
rect 6909 -5560 7005 -5526
rect 8995 -5560 9091 -5526
rect 6909 -5622 6943 -5560
rect 9057 -5622 9091 -5560
rect 6909 -6340 6943 -6278
rect 9057 -6340 9091 -6278
rect 6909 -6374 7005 -6340
rect 8995 -6374 9091 -6340
rect 6681 -6516 6715 -6454
rect 5745 -6550 5841 -6516
rect 6619 -6550 6715 -6516
rect 10222 -4298 10256 -4236
rect 9286 -6516 9320 -6454
rect 10222 -6516 10256 -6454
rect 9286 -6550 9382 -6516
rect 10160 -6550 10256 -6516
<< nsubdiff >>
rect 5981 12434 6077 12468
rect 9923 12434 10019 12468
rect 5981 12372 6015 12434
rect 9985 12372 10019 12434
rect 5981 10136 6015 10198
rect 9985 10136 10019 10198
rect 5981 10102 6077 10136
rect 9923 10102 10019 10136
rect 11260 3886 11356 3920
rect 13716 3886 13874 3920
rect 14032 3886 14190 3920
rect 14348 3886 14444 3920
rect 11260 3824 11294 3886
rect 2070 2790 2104 2814
rect 2070 2704 2104 2756
rect 2070 2646 2104 2670
rect 5238 2790 5368 2814
rect 5272 2756 5334 2790
rect 5238 2704 5368 2756
rect 5272 2670 5334 2704
rect 5238 2646 5368 2670
rect 9846 2790 9880 2814
rect 9846 2704 9880 2756
rect 9846 2646 9880 2670
rect 10134 2790 10168 2814
rect 10134 2704 10168 2756
rect 10134 2646 10168 2670
rect 2070 1754 2104 1778
rect 2070 1668 2104 1720
rect 2070 1610 2104 1634
rect 5238 1754 5368 1778
rect 5272 1720 5334 1754
rect 5238 1668 5368 1720
rect 5272 1634 5334 1668
rect 5238 1610 5368 1634
rect 10134 1754 10168 1778
rect 10134 1668 10168 1720
rect 10134 1610 10168 1634
rect 13778 3824 13812 3886
rect 11260 1588 11294 1650
rect 14094 3824 14128 3886
rect 13778 1588 13812 1650
rect 14410 3824 14444 3886
rect 14094 1588 14128 1650
rect 14410 1588 14444 1650
rect 11260 1554 11356 1588
rect 13716 1554 13874 1588
rect 14032 1554 14190 1588
rect 14348 1554 14444 1588
rect 3222 1458 3256 1482
rect 1796 1362 1830 1386
rect 1796 1269 1830 1328
rect 1796 1211 1830 1235
rect 2072 1362 2106 1386
rect 2072 1269 2106 1328
rect 2072 1211 2106 1235
rect 2164 1362 2198 1386
rect 2164 1269 2198 1328
rect 2164 1211 2198 1235
rect 2440 1362 2474 1386
rect 2440 1269 2474 1328
rect 2440 1211 2474 1235
rect 2532 1362 2566 1386
rect 2532 1269 2566 1328
rect 2532 1211 2566 1235
rect 2808 1362 2842 1386
rect 2808 1269 2842 1328
rect 3222 1372 3256 1424
rect 3222 1314 3256 1338
rect 2808 1211 2842 1235
rect 5238 1458 5368 1482
rect 5272 1424 5334 1458
rect 5238 1372 5368 1424
rect 5272 1338 5334 1372
rect 5238 1314 5368 1338
rect 10134 1458 10168 1482
rect 10134 1372 10168 1424
rect 10134 1314 10168 1338
rect 10312 -417 10336 -383
rect 10370 -417 10429 -383
rect 10463 -417 10487 -383
rect 10312 -693 10336 -659
rect 10370 -693 10429 -659
rect 10463 -693 10487 -659
rect 10312 -1061 10336 -1027
rect 10370 -1061 10429 -1027
rect 10463 -1061 10487 -1027
rect 10312 -1337 10336 -1303
rect 10370 -1337 10429 -1303
rect 10463 -1337 10487 -1303
rect 5981 -6736 6077 -6702
rect 9923 -6736 10019 -6702
rect 5981 -6798 6015 -6736
rect 9985 -6798 10019 -6736
rect 5981 -9034 6015 -8972
rect 9985 -9034 10019 -8972
rect 5981 -9068 6077 -9034
rect 9923 -9068 10019 -9034
<< psubdiffcont >>
rect 5841 9916 6619 9950
rect 5138 9548 5578 9582
rect 5042 8382 5076 9486
rect 5640 8382 5674 9486
rect 5138 8286 5578 8320
rect 5745 7698 5779 9854
rect 6681 7698 6715 9854
rect 9382 9916 10160 9950
rect 7005 9740 8995 9774
rect 6909 9022 6943 9678
rect 9057 9022 9091 9678
rect 7005 8926 8995 8960
rect 5841 7602 6619 7636
rect 7049 8800 8951 8834
rect 6953 6582 6987 8738
rect 9013 6582 9047 8738
rect 9286 7698 9320 9854
rect 10222 7698 10256 9854
rect 9382 7602 10160 7636
rect 7049 6486 8951 6520
rect 10774 7382 11430 7416
rect 10678 6470 10712 7320
rect 11492 6470 11526 7320
rect 10774 6354 11430 6388
rect 3451 4492 3609 4526
rect 3355 3874 3389 4430
rect 3671 3874 3705 4430
rect 3451 3778 3609 3812
rect 3355 3160 3389 3716
rect 3671 3160 3705 3716
rect 3451 3064 3609 3098
rect 4233 4492 4391 4526
rect 4137 3874 4171 4430
rect 4453 3874 4487 4430
rect 4233 3778 4391 3812
rect 4137 3160 4171 3716
rect 4453 3160 4487 3716
rect 4233 3064 4391 3098
rect 2070 2383 2104 2417
rect 2070 2300 2104 2334
rect 10788 2716 11092 2750
rect 5238 2383 5272 2417
rect 5334 2383 5368 2417
rect 9846 2383 9880 2417
rect 5238 2300 5272 2334
rect 5334 2300 5368 2334
rect 9846 2300 9880 2334
rect 10134 2383 10168 2417
rect 10134 2300 10168 2334
rect 2070 2090 2104 2124
rect 2070 2007 2104 2041
rect 5238 2090 5272 2124
rect 5334 2090 5368 2124
rect 5238 2007 5272 2041
rect 5334 2007 5368 2041
rect 10134 2090 10168 2124
rect 10134 2007 10168 2041
rect 10692 1650 10726 2654
rect 11154 1650 11188 2654
rect 10788 1554 11092 1588
rect 1796 1017 1830 1051
rect 2072 1017 2106 1051
rect 2164 1017 2198 1051
rect 2440 1017 2474 1051
rect 2532 1017 2566 1051
rect 2808 1017 2842 1051
rect 3222 1051 3256 1085
rect 3222 968 3256 1002
rect 5238 1051 5272 1085
rect 5334 1051 5368 1085
rect 5238 968 5272 1002
rect 5334 968 5368 1002
rect 10440 1448 13716 1482
rect 13874 1448 14032 1482
rect 14190 1448 14348 1482
rect 10134 1051 10168 1085
rect 10134 968 10168 1002
rect 3800 722 3958 756
rect 3704 104 3738 660
rect 4020 104 4054 660
rect 10344 230 10378 1386
rect 13778 230 13812 1386
rect 14094 230 14128 1386
rect 14410 230 14444 1386
rect 39329 1141 40361 1175
rect 15462 981 16018 1015
rect 16176 981 16732 1015
rect 16890 981 17446 1015
rect 17604 981 18160 1015
rect 18318 981 18874 1015
rect 19032 981 19588 1015
rect 19746 981 20302 1015
rect 20460 981 21016 1015
rect 21174 981 21730 1015
rect 21888 981 22444 1015
rect 22602 981 23158 1015
rect 23316 981 23872 1015
rect 24030 981 24586 1015
rect 24744 981 25300 1015
rect 25458 981 26014 1015
rect 26172 981 26728 1015
rect 26886 981 27442 1015
rect 27600 981 28156 1015
rect 28314 981 28870 1015
rect 29028 981 29584 1015
rect 29742 981 30298 1015
rect 30456 981 31012 1015
rect 31170 981 31726 1015
rect 31884 981 32440 1015
rect 32598 981 33154 1015
rect 33312 981 33868 1015
rect 34026 981 34582 1015
rect 34740 981 35296 1015
rect 35454 981 36010 1015
rect 36168 981 36724 1015
rect 36882 981 37438 1015
rect 37596 981 38152 1015
rect 38310 981 38866 1015
rect 15366 761 15400 919
rect 16080 761 16114 919
rect 16794 761 16828 919
rect 17508 761 17542 919
rect 18222 761 18256 919
rect 18936 761 18970 919
rect 19650 761 19684 919
rect 20364 761 20398 919
rect 21078 761 21112 919
rect 21792 761 21826 919
rect 22506 761 22540 919
rect 23220 761 23254 919
rect 23934 761 23968 919
rect 24648 761 24682 919
rect 25362 761 25396 919
rect 26076 761 26110 919
rect 26790 761 26824 919
rect 27504 761 27538 919
rect 28218 761 28252 919
rect 28932 761 28966 919
rect 29646 761 29680 919
rect 30360 761 30394 919
rect 31074 761 31108 919
rect 31788 761 31822 919
rect 32502 761 32536 919
rect 33216 761 33250 919
rect 33930 761 33964 919
rect 34644 761 34678 919
rect 35358 761 35392 919
rect 36072 761 36106 919
rect 36786 761 36820 919
rect 37500 761 37534 919
rect 38214 761 38248 919
rect 38928 761 38962 919
rect 15462 665 16018 699
rect 16176 665 16732 699
rect 16890 665 17446 699
rect 17604 665 18160 699
rect 18318 665 18874 699
rect 19032 665 19588 699
rect 19746 665 20302 699
rect 20460 665 21016 699
rect 21174 665 21730 699
rect 21888 665 22444 699
rect 22602 665 23158 699
rect 23316 665 23872 699
rect 24030 665 24586 699
rect 24744 665 25300 699
rect 25458 665 26014 699
rect 26172 665 26728 699
rect 26886 665 27442 699
rect 27600 665 28156 699
rect 28314 665 28870 699
rect 29028 665 29584 699
rect 29742 665 30298 699
rect 30456 665 31012 699
rect 31170 665 31726 699
rect 31884 665 32440 699
rect 32598 665 33154 699
rect 33312 665 33868 699
rect 34026 665 34582 699
rect 34740 665 35296 699
rect 35454 665 36010 699
rect 36168 665 36724 699
rect 36882 665 37438 699
rect 37596 665 38152 699
rect 38310 665 38866 699
rect 10440 134 13716 168
rect 13874 134 14032 168
rect 14190 134 14348 168
rect 15462 163 16018 197
rect 16176 163 16732 197
rect 16890 163 17446 197
rect 17604 163 18160 197
rect 18318 163 18874 197
rect 19032 163 19588 197
rect 19746 163 20302 197
rect 20460 163 21016 197
rect 21174 163 21730 197
rect 21888 163 22444 197
rect 22602 163 23158 197
rect 23316 163 23872 197
rect 24030 163 24586 197
rect 24744 163 25300 197
rect 25458 163 26014 197
rect 26172 163 26728 197
rect 26886 163 27442 197
rect 27600 163 28156 197
rect 28314 163 28870 197
rect 29028 163 29584 197
rect 29742 163 30298 197
rect 30456 163 31012 197
rect 31170 163 31726 197
rect 31884 163 32440 197
rect 32598 163 33154 197
rect 33312 163 33868 197
rect 34026 163 34582 197
rect 34740 163 35296 197
rect 35454 163 36010 197
rect 36168 163 36724 197
rect 36882 163 37438 197
rect 37596 163 38152 197
rect 38310 163 38866 197
rect 3800 8 3958 42
rect 3704 -610 3738 -54
rect 4020 -610 4054 -54
rect 15366 -57 15400 101
rect 16080 -57 16114 101
rect 16794 -57 16828 101
rect 17508 -57 17542 101
rect 18222 -57 18256 101
rect 18936 -57 18970 101
rect 19650 -57 19684 101
rect 20364 -57 20398 101
rect 21078 -57 21112 101
rect 21792 -57 21826 101
rect 22506 -57 22540 101
rect 23220 -57 23254 101
rect 23934 -57 23968 101
rect 24648 -57 24682 101
rect 25362 -57 25396 101
rect 26076 -57 26110 101
rect 26790 -57 26824 101
rect 27504 -57 27538 101
rect 28218 -57 28252 101
rect 28932 -57 28966 101
rect 29646 -57 29680 101
rect 30360 -57 30394 101
rect 31074 -57 31108 101
rect 31788 -57 31822 101
rect 32502 -57 32536 101
rect 33216 -57 33250 101
rect 33930 -57 33964 101
rect 34644 -57 34678 101
rect 35358 -57 35392 101
rect 36072 -57 36106 101
rect 36786 -57 36820 101
rect 37500 -57 37534 101
rect 38214 -57 38248 101
rect 38928 -57 38962 101
rect 15462 -153 16018 -119
rect 16176 -153 16732 -119
rect 16890 -153 17446 -119
rect 17604 -153 18160 -119
rect 18318 -153 18874 -119
rect 19032 -153 19588 -119
rect 19746 -153 20302 -119
rect 20460 -153 21016 -119
rect 21174 -153 21730 -119
rect 21888 -153 22444 -119
rect 22602 -153 23158 -119
rect 23316 -153 23872 -119
rect 24030 -153 24586 -119
rect 24744 -153 25300 -119
rect 25458 -153 26014 -119
rect 26172 -153 26728 -119
rect 26886 -153 27442 -119
rect 27600 -153 28156 -119
rect 28314 -153 28870 -119
rect 29028 -153 29584 -119
rect 29742 -153 30298 -119
rect 30456 -153 31012 -119
rect 31170 -153 31726 -119
rect 31884 -153 32440 -119
rect 32598 -153 33154 -119
rect 33312 -153 33868 -119
rect 34026 -153 34582 -119
rect 34740 -153 35296 -119
rect 35454 -153 36010 -119
rect 36168 -153 36724 -119
rect 36882 -153 37438 -119
rect 37596 -153 38152 -119
rect 38310 -153 38866 -119
rect 39233 -221 39267 1079
rect 40423 -221 40457 1079
rect 39329 -317 40361 -283
rect 10647 -417 10681 -383
rect 3800 -706 3958 -672
rect 10647 -693 10681 -659
rect 10647 -1061 10681 -1027
rect 10647 -1337 10681 -1303
rect 10774 -2988 11430 -2954
rect 7049 -3120 8951 -3086
rect 5841 -4236 6619 -4202
rect 5138 -4920 5578 -4886
rect 5042 -6086 5076 -4982
rect 5640 -6086 5674 -4982
rect 5138 -6182 5578 -6148
rect 5745 -6454 5779 -4298
rect 6681 -6454 6715 -4298
rect 6953 -5338 6987 -3182
rect 9013 -5338 9047 -3182
rect 10678 -3920 10712 -3070
rect 11492 -3920 11526 -3070
rect 10774 -4016 11430 -3982
rect 7049 -5434 8951 -5400
rect 9382 -4236 10160 -4202
rect 7005 -5560 8995 -5526
rect 6909 -6278 6943 -5622
rect 9057 -6278 9091 -5622
rect 7005 -6374 8995 -6340
rect 5841 -6550 6619 -6516
rect 9286 -6454 9320 -4298
rect 10222 -6454 10256 -4298
rect 9382 -6550 10160 -6516
<< nsubdiffcont >>
rect 6077 12434 9923 12468
rect 5981 10198 6015 12372
rect 9985 10198 10019 12372
rect 6077 10102 9923 10136
rect 11356 3886 13716 3920
rect 13874 3886 14032 3920
rect 14190 3886 14348 3920
rect 2070 2756 2104 2790
rect 2070 2670 2104 2704
rect 5238 2756 5272 2790
rect 5334 2756 5368 2790
rect 5238 2670 5272 2704
rect 5334 2670 5368 2704
rect 9846 2756 9880 2790
rect 9846 2670 9880 2704
rect 10134 2756 10168 2790
rect 10134 2670 10168 2704
rect 2070 1720 2104 1754
rect 2070 1634 2104 1668
rect 5238 1720 5272 1754
rect 5334 1720 5368 1754
rect 5238 1634 5272 1668
rect 5334 1634 5368 1668
rect 10134 1720 10168 1754
rect 10134 1634 10168 1668
rect 11260 1650 11294 3824
rect 13778 1650 13812 3824
rect 14094 1650 14128 3824
rect 14410 1650 14444 3824
rect 11356 1554 13716 1588
rect 13874 1554 14032 1588
rect 14190 1554 14348 1588
rect 3222 1424 3256 1458
rect 1796 1328 1830 1362
rect 1796 1235 1830 1269
rect 2072 1328 2106 1362
rect 2072 1235 2106 1269
rect 2164 1328 2198 1362
rect 2164 1235 2198 1269
rect 2440 1328 2474 1362
rect 2440 1235 2474 1269
rect 2532 1328 2566 1362
rect 2532 1235 2566 1269
rect 2808 1328 2842 1362
rect 3222 1338 3256 1372
rect 2808 1235 2842 1269
rect 5238 1424 5272 1458
rect 5334 1424 5368 1458
rect 5238 1338 5272 1372
rect 5334 1338 5368 1372
rect 10134 1424 10168 1458
rect 10134 1338 10168 1372
rect 10336 -417 10370 -383
rect 10429 -417 10463 -383
rect 10336 -693 10370 -659
rect 10429 -693 10463 -659
rect 10336 -1061 10370 -1027
rect 10429 -1061 10463 -1027
rect 10336 -1337 10370 -1303
rect 10429 -1337 10463 -1303
rect 6077 -6736 9923 -6702
rect 5981 -8972 6015 -6798
rect 9985 -8972 10019 -6798
rect 6077 -9068 9923 -9034
<< poly >>
rect 6138 12366 6204 12382
rect 6138 12332 6154 12366
rect 6188 12332 6204 12366
rect 6138 12316 6204 12332
rect 6256 12366 6322 12382
rect 6256 12332 6272 12366
rect 6306 12332 6322 12366
rect 6256 12316 6322 12332
rect 6374 12366 6440 12382
rect 6374 12332 6390 12366
rect 6424 12332 6440 12366
rect 6374 12316 6440 12332
rect 6492 12366 6558 12382
rect 6492 12332 6508 12366
rect 6542 12332 6558 12366
rect 6492 12316 6558 12332
rect 6610 12366 6676 12382
rect 6610 12332 6626 12366
rect 6660 12332 6676 12366
rect 6610 12316 6676 12332
rect 6728 12366 6794 12382
rect 6728 12332 6744 12366
rect 6778 12332 6794 12366
rect 6728 12316 6794 12332
rect 6846 12366 6912 12382
rect 6846 12332 6862 12366
rect 6896 12332 6912 12366
rect 6846 12316 6912 12332
rect 6964 12366 7030 12382
rect 6964 12332 6980 12366
rect 7014 12332 7030 12366
rect 6964 12316 7030 12332
rect 7082 12366 7148 12382
rect 7082 12332 7098 12366
rect 7132 12332 7148 12366
rect 7082 12316 7148 12332
rect 7200 12366 7266 12382
rect 7200 12332 7216 12366
rect 7250 12332 7266 12366
rect 7200 12316 7266 12332
rect 7318 12366 7384 12382
rect 7318 12332 7334 12366
rect 7368 12332 7384 12366
rect 7318 12316 7384 12332
rect 7436 12366 7502 12382
rect 7436 12332 7452 12366
rect 7486 12332 7502 12366
rect 7436 12316 7502 12332
rect 7554 12316 7620 12382
rect 7672 12316 7738 12382
rect 7790 12316 7856 12382
rect 7908 12316 7974 12382
rect 8026 12316 8092 12382
rect 8144 12316 8210 12382
rect 8262 12316 8328 12382
rect 8380 12316 8446 12382
rect 8498 12366 8564 12382
rect 8498 12332 8514 12366
rect 8548 12332 8564 12366
rect 8498 12316 8564 12332
rect 8616 12366 8682 12382
rect 8616 12332 8632 12366
rect 8666 12332 8682 12366
rect 8616 12316 8682 12332
rect 8734 12366 8800 12382
rect 8734 12332 8750 12366
rect 8784 12332 8800 12366
rect 8734 12316 8800 12332
rect 8852 12366 8918 12382
rect 8852 12332 8868 12366
rect 8902 12332 8918 12366
rect 8852 12316 8918 12332
rect 8970 12366 9036 12382
rect 8970 12332 8986 12366
rect 9020 12332 9036 12366
rect 8970 12316 9036 12332
rect 9088 12366 9154 12382
rect 9088 12332 9104 12366
rect 9138 12332 9154 12366
rect 9088 12316 9154 12332
rect 9206 12366 9272 12382
rect 9206 12332 9222 12366
rect 9256 12332 9272 12366
rect 9206 12316 9272 12332
rect 9324 12366 9390 12382
rect 9324 12332 9340 12366
rect 9374 12332 9390 12366
rect 9324 12316 9390 12332
rect 9442 12366 9508 12382
rect 9442 12332 9458 12366
rect 9492 12332 9508 12366
rect 9442 12316 9508 12332
rect 9560 12366 9626 12382
rect 9560 12332 9576 12366
rect 9610 12332 9626 12366
rect 9560 12316 9626 12332
rect 9678 12366 9744 12382
rect 9678 12332 9694 12366
rect 9728 12332 9744 12366
rect 9678 12316 9744 12332
rect 9796 12366 9862 12382
rect 9796 12332 9812 12366
rect 9846 12332 9862 12366
rect 9796 12316 9862 12332
rect 6141 12285 6201 12316
rect 6259 12285 6319 12316
rect 6377 12285 6437 12316
rect 6495 12285 6555 12316
rect 6613 12285 6673 12316
rect 6731 12285 6791 12316
rect 6849 12285 6909 12316
rect 6967 12285 7027 12316
rect 7085 12285 7145 12316
rect 7203 12285 7263 12316
rect 7321 12285 7381 12316
rect 7439 12285 7499 12316
rect 7557 12285 7617 12316
rect 7675 12285 7735 12316
rect 7793 12285 7853 12316
rect 7911 12285 7971 12316
rect 8029 12285 8089 12316
rect 8147 12285 8207 12316
rect 8265 12285 8325 12316
rect 8383 12285 8443 12316
rect 8501 12285 8561 12316
rect 8619 12285 8679 12316
rect 8737 12285 8797 12316
rect 8855 12285 8915 12316
rect 8973 12285 9033 12316
rect 9091 12285 9151 12316
rect 9209 12285 9269 12316
rect 9327 12285 9387 12316
rect 9445 12285 9505 12316
rect 9563 12285 9623 12316
rect 9681 12285 9741 12316
rect 9799 12285 9859 12316
rect 6141 10254 6201 10285
rect 6259 10254 6319 10285
rect 6377 10254 6437 10285
rect 6495 10254 6555 10285
rect 6613 10254 6673 10285
rect 6731 10254 6791 10285
rect 6849 10254 6909 10285
rect 6967 10254 7027 10285
rect 7085 10254 7145 10285
rect 7203 10254 7263 10285
rect 7321 10254 7381 10285
rect 7439 10254 7499 10285
rect 7557 10254 7617 10285
rect 7675 10254 7735 10285
rect 7793 10254 7853 10285
rect 7911 10254 7971 10285
rect 8029 10254 8089 10285
rect 8147 10254 8207 10285
rect 8265 10254 8325 10285
rect 8383 10254 8443 10285
rect 8501 10254 8561 10285
rect 8619 10254 8679 10285
rect 8737 10254 8797 10285
rect 8855 10254 8915 10285
rect 8973 10254 9033 10285
rect 9091 10254 9151 10285
rect 9209 10254 9269 10285
rect 9327 10254 9387 10285
rect 9445 10254 9505 10285
rect 9563 10254 9623 10285
rect 9681 10254 9741 10285
rect 9799 10254 9859 10285
rect 6138 10238 6204 10254
rect 6138 10204 6154 10238
rect 6188 10204 6204 10238
rect 6138 10188 6204 10204
rect 6256 10238 6322 10254
rect 6256 10204 6272 10238
rect 6306 10204 6322 10238
rect 6256 10188 6322 10204
rect 6374 10238 6440 10254
rect 6374 10204 6390 10238
rect 6424 10204 6440 10238
rect 6374 10188 6440 10204
rect 6492 10238 6558 10254
rect 6492 10204 6508 10238
rect 6542 10204 6558 10238
rect 6492 10188 6558 10204
rect 6610 10238 6676 10254
rect 6610 10204 6626 10238
rect 6660 10204 6676 10238
rect 6610 10188 6676 10204
rect 6728 10238 6794 10254
rect 6728 10204 6744 10238
rect 6778 10204 6794 10238
rect 6728 10188 6794 10204
rect 6846 10238 6912 10254
rect 6846 10204 6862 10238
rect 6896 10204 6912 10238
rect 6846 10188 6912 10204
rect 6964 10238 7030 10254
rect 6964 10204 6980 10238
rect 7014 10204 7030 10238
rect 6964 10188 7030 10204
rect 7082 10238 7148 10254
rect 7082 10204 7098 10238
rect 7132 10204 7148 10238
rect 7082 10188 7148 10204
rect 7200 10238 7266 10254
rect 7200 10204 7216 10238
rect 7250 10204 7266 10238
rect 7200 10188 7266 10204
rect 7318 10238 7384 10254
rect 7318 10204 7334 10238
rect 7368 10204 7384 10238
rect 7318 10188 7384 10204
rect 7436 10238 7502 10254
rect 7436 10204 7452 10238
rect 7486 10204 7502 10238
rect 7436 10188 7502 10204
rect 7554 10238 7620 10254
rect 7554 10204 7570 10238
rect 7604 10204 7620 10238
rect 7554 10188 7620 10204
rect 7672 10238 7738 10254
rect 7672 10204 7688 10238
rect 7722 10204 7738 10238
rect 7672 10188 7738 10204
rect 7790 10238 7856 10254
rect 7790 10204 7806 10238
rect 7840 10204 7856 10238
rect 7790 10188 7856 10204
rect 7908 10238 7974 10254
rect 7908 10204 7924 10238
rect 7958 10204 7974 10238
rect 7908 10188 7974 10204
rect 8026 10238 8092 10254
rect 8026 10204 8042 10238
rect 8076 10204 8092 10238
rect 8026 10188 8092 10204
rect 8144 10238 8210 10254
rect 8144 10204 8160 10238
rect 8194 10204 8210 10238
rect 8144 10188 8210 10204
rect 8262 10238 8328 10254
rect 8262 10204 8278 10238
rect 8312 10204 8328 10238
rect 8262 10188 8328 10204
rect 8380 10238 8446 10254
rect 8380 10204 8396 10238
rect 8430 10204 8446 10238
rect 8380 10188 8446 10204
rect 8498 10238 8564 10254
rect 8498 10204 8514 10238
rect 8548 10204 8564 10238
rect 8498 10188 8564 10204
rect 8616 10238 8682 10254
rect 8616 10204 8632 10238
rect 8666 10204 8682 10238
rect 8616 10188 8682 10204
rect 8734 10238 8800 10254
rect 8734 10204 8750 10238
rect 8784 10204 8800 10238
rect 8734 10188 8800 10204
rect 8852 10238 8918 10254
rect 8852 10204 8868 10238
rect 8902 10204 8918 10238
rect 8852 10188 8918 10204
rect 8970 10238 9036 10254
rect 8970 10204 8986 10238
rect 9020 10204 9036 10238
rect 8970 10188 9036 10204
rect 9088 10238 9154 10254
rect 9088 10204 9104 10238
rect 9138 10204 9154 10238
rect 9088 10188 9154 10204
rect 9206 10238 9272 10254
rect 9206 10204 9222 10238
rect 9256 10204 9272 10238
rect 9206 10188 9272 10204
rect 9324 10238 9390 10254
rect 9324 10204 9340 10238
rect 9374 10204 9390 10238
rect 9324 10188 9390 10204
rect 9442 10238 9508 10254
rect 9442 10204 9458 10238
rect 9492 10204 9508 10238
rect 9442 10188 9508 10204
rect 9560 10238 9626 10254
rect 9560 10204 9576 10238
rect 9610 10204 9626 10238
rect 9560 10188 9626 10204
rect 9678 10238 9744 10254
rect 9678 10204 9694 10238
rect 9728 10204 9744 10238
rect 9678 10188 9744 10204
rect 9796 10238 9862 10254
rect 9796 10204 9812 10238
rect 9846 10204 9862 10238
rect 9796 10188 9862 10204
rect 5902 9848 5968 9864
rect 5902 9814 5918 9848
rect 5952 9814 5968 9848
rect 5902 9798 5968 9814
rect 6020 9848 6086 9864
rect 6020 9814 6036 9848
rect 6070 9814 6086 9848
rect 6020 9798 6086 9814
rect 6138 9848 6204 9864
rect 6138 9814 6154 9848
rect 6188 9814 6204 9848
rect 6138 9798 6204 9814
rect 6256 9848 6322 9864
rect 6256 9814 6272 9848
rect 6306 9814 6322 9848
rect 6256 9798 6322 9814
rect 6374 9848 6440 9864
rect 6374 9814 6390 9848
rect 6424 9814 6440 9848
rect 6374 9798 6440 9814
rect 6492 9848 6558 9864
rect 6492 9814 6508 9848
rect 6542 9814 6558 9848
rect 6492 9798 6558 9814
rect 5905 9776 5965 9798
rect 6023 9776 6083 9798
rect 6141 9776 6201 9798
rect 6259 9776 6319 9798
rect 6377 9776 6437 9798
rect 6495 9776 6555 9798
rect 5905 7754 5965 7776
rect 6023 7754 6083 7776
rect 6141 7754 6201 7776
rect 6259 7754 6319 7776
rect 6377 7754 6437 7776
rect 6495 7754 6555 7776
rect 5902 7738 5968 7754
rect 5902 7704 5918 7738
rect 5952 7704 5968 7738
rect 5902 7688 5968 7704
rect 6020 7738 6086 7754
rect 6020 7704 6036 7738
rect 6070 7704 6086 7738
rect 6020 7688 6086 7704
rect 6138 7738 6204 7754
rect 6138 7704 6154 7738
rect 6188 7704 6204 7738
rect 6138 7688 6204 7704
rect 6256 7738 6322 7754
rect 6256 7704 6272 7738
rect 6306 7704 6322 7738
rect 6256 7688 6322 7704
rect 6374 7738 6440 7754
rect 6374 7704 6390 7738
rect 6424 7704 6440 7738
rect 6374 7688 6440 7704
rect 6492 7738 6558 7754
rect 6492 7704 6508 7738
rect 6542 7704 6558 7738
rect 6492 7688 6558 7704
rect 7073 9676 7199 9704
rect 7073 9642 7119 9676
rect 7153 9642 7199 9676
rect 7073 9626 7199 9642
rect 8801 9676 8927 9704
rect 8801 9642 8847 9676
rect 8881 9642 8927 9676
rect 8801 9626 8927 9642
rect 7073 9600 7103 9626
rect 7169 9600 7199 9626
rect 7265 9600 7295 9626
rect 7361 9600 7391 9626
rect 7457 9600 7487 9626
rect 7553 9600 7583 9626
rect 7649 9600 7679 9626
rect 7745 9600 7775 9626
rect 7841 9600 7871 9626
rect 7937 9600 7967 9626
rect 8033 9600 8063 9626
rect 8129 9600 8159 9626
rect 8225 9600 8255 9626
rect 8321 9600 8351 9626
rect 8417 9600 8447 9626
rect 8513 9600 8543 9626
rect 8609 9600 8639 9626
rect 8705 9600 8735 9626
rect 8801 9600 8831 9626
rect 8897 9600 8927 9626
rect 7073 9074 7103 9100
rect 7169 9074 7199 9100
rect 7265 9078 7295 9100
rect 7361 9078 7391 9100
rect 7265 9050 7391 9078
rect 7265 9016 7311 9050
rect 7345 9016 7391 9050
rect 7265 9000 7391 9016
rect 7457 9078 7487 9100
rect 7553 9078 7583 9100
rect 7457 9050 7583 9078
rect 7457 9016 7503 9050
rect 7537 9016 7583 9050
rect 7457 9000 7583 9016
rect 7649 9078 7679 9100
rect 7745 9078 7775 9100
rect 7649 9050 7775 9078
rect 7649 9016 7695 9050
rect 7729 9016 7775 9050
rect 7649 9000 7775 9016
rect 7841 9078 7871 9100
rect 7937 9078 7967 9100
rect 7841 9050 7967 9078
rect 7841 9016 7887 9050
rect 7921 9016 7967 9050
rect 7841 9000 7967 9016
rect 8033 9078 8063 9100
rect 8129 9078 8159 9100
rect 8033 9050 8159 9078
rect 8033 9016 8079 9050
rect 8113 9016 8159 9050
rect 8033 9000 8159 9016
rect 8225 9078 8255 9100
rect 8321 9078 8351 9100
rect 8225 9050 8351 9078
rect 8225 9016 8271 9050
rect 8305 9016 8351 9050
rect 8225 9000 8351 9016
rect 8417 9078 8447 9100
rect 8513 9078 8543 9100
rect 8417 9050 8543 9078
rect 8417 9016 8463 9050
rect 8497 9016 8543 9050
rect 8417 9000 8543 9016
rect 8609 9078 8639 9100
rect 8705 9078 8735 9100
rect 8609 9050 8735 9078
rect 8801 9074 8831 9100
rect 8897 9074 8927 9100
rect 8609 9016 8655 9050
rect 8689 9016 8735 9050
rect 8609 9000 8735 9016
rect 7113 8732 7513 8748
rect 7113 8698 7129 8732
rect 7497 8698 7513 8732
rect 7113 8660 7513 8698
rect 7571 8732 7971 8748
rect 7571 8698 7587 8732
rect 7955 8698 7971 8732
rect 7571 8660 7971 8698
rect 8029 8732 8429 8748
rect 8029 8698 8045 8732
rect 8413 8698 8429 8732
rect 8029 8660 8429 8698
rect 8487 8732 8887 8748
rect 8487 8698 8503 8732
rect 8871 8698 8887 8732
rect 8487 8660 8887 8698
rect 7113 6622 7513 6660
rect 7113 6588 7129 6622
rect 7497 6588 7513 6622
rect 7113 6572 7513 6588
rect 7571 6622 7971 6660
rect 7571 6588 7587 6622
rect 7955 6588 7971 6622
rect 7571 6572 7971 6588
rect 8029 6622 8429 6660
rect 8029 6588 8045 6622
rect 8413 6588 8429 6622
rect 8029 6572 8429 6588
rect 8487 6622 8887 6660
rect 8487 6588 8503 6622
rect 8871 6588 8887 6622
rect 8487 6572 8887 6588
rect 9443 9848 9509 9864
rect 9443 9814 9459 9848
rect 9493 9814 9509 9848
rect 9443 9798 9509 9814
rect 9561 9848 9627 9864
rect 9561 9814 9577 9848
rect 9611 9814 9627 9848
rect 9561 9798 9627 9814
rect 9679 9848 9745 9864
rect 9679 9814 9695 9848
rect 9729 9814 9745 9848
rect 9679 9798 9745 9814
rect 9797 9848 9863 9864
rect 9797 9814 9813 9848
rect 9847 9814 9863 9848
rect 9797 9798 9863 9814
rect 9915 9848 9981 9864
rect 9915 9814 9931 9848
rect 9965 9814 9981 9848
rect 9915 9798 9981 9814
rect 10033 9848 10099 9864
rect 10033 9814 10049 9848
rect 10083 9814 10099 9848
rect 10033 9798 10099 9814
rect 9446 9776 9506 9798
rect 9564 9776 9624 9798
rect 9682 9776 9742 9798
rect 9800 9776 9860 9798
rect 9918 9776 9978 9798
rect 10036 9776 10096 9798
rect 9446 7754 9506 7776
rect 9564 7754 9624 7776
rect 9682 7754 9742 7776
rect 9800 7754 9860 7776
rect 9918 7754 9978 7776
rect 10036 7754 10096 7776
rect 9443 7738 9509 7754
rect 9443 7704 9459 7738
rect 9493 7704 9509 7738
rect 9443 7688 9509 7704
rect 9561 7738 9627 7754
rect 9561 7704 9577 7738
rect 9611 7704 9627 7738
rect 9561 7688 9627 7704
rect 9679 7738 9745 7754
rect 9679 7704 9695 7738
rect 9729 7704 9745 7738
rect 9679 7688 9745 7704
rect 9797 7738 9863 7754
rect 9797 7704 9813 7738
rect 9847 7704 9863 7738
rect 9797 7688 9863 7704
rect 9915 7738 9981 7754
rect 9915 7704 9931 7738
rect 9965 7704 9981 7738
rect 9915 7688 9981 7704
rect 10033 7738 10099 7754
rect 10033 7704 10049 7738
rect 10083 7704 10099 7738
rect 10033 7688 10099 7704
rect 10826 7222 10852 7252
rect 11352 7236 11440 7252
rect 11352 7222 11390 7236
rect 11374 7202 11390 7222
rect 11424 7202 11440 7236
rect 11374 7156 11440 7202
rect 10826 7126 10852 7156
rect 11352 7126 11440 7156
rect 10826 7030 10852 7060
rect 11352 7044 11440 7060
rect 11352 7030 11390 7044
rect 11374 7010 11390 7030
rect 11424 7010 11440 7044
rect 11374 6964 11440 7010
rect 10826 6934 10852 6964
rect 11352 6934 11440 6964
rect 3497 4374 3563 4440
rect 3515 4352 3545 4374
rect 3515 3930 3545 3952
rect 3497 3914 3563 3930
rect 3497 3880 3513 3914
rect 3547 3880 3563 3914
rect 3497 3864 3563 3880
rect 3497 3660 3563 3726
rect 3515 3638 3545 3660
rect 3515 3216 3545 3238
rect 3497 3200 3563 3216
rect 3497 3166 3513 3200
rect 3547 3166 3563 3200
rect 3497 3150 3563 3166
rect 4279 4374 4345 4440
rect 4297 4352 4327 4374
rect 4297 3930 4327 3952
rect 4279 3914 4345 3930
rect 4279 3880 4295 3914
rect 4329 3880 4345 3914
rect 4279 3864 4345 3880
rect 4279 3660 4345 3726
rect 4297 3638 4327 3660
rect 4297 3216 4327 3238
rect 4279 3200 4345 3216
rect 4279 3166 4295 3200
rect 4329 3166 4345 3200
rect 4279 3150 4345 3166
rect 2497 2804 2527 2830
rect 3851 2804 3881 2830
rect 3941 2804 3971 2830
rect 4137 2804 4337 2830
rect 4392 2804 4592 2830
rect 2497 2565 2527 2580
rect 2494 2538 2530 2565
rect 2356 2531 2530 2538
rect 2354 2522 2530 2531
rect 2354 2488 2372 2522
rect 2406 2488 2440 2522
rect 2474 2488 2530 2522
rect 2354 2479 2530 2488
rect 2356 2472 2530 2479
rect 2499 2434 2529 2472
rect 5481 2804 5681 2830
rect 5736 2804 5936 2830
rect 6153 2804 6353 2830
rect 6408 2804 6608 2830
rect 6825 2804 7025 2830
rect 7080 2804 7280 2830
rect 8169 2804 8369 2830
rect 8424 2804 8624 2830
rect 8841 2804 9041 2830
rect 9096 2804 9296 2830
rect 9513 2804 9713 2830
rect 3851 2565 3881 2580
rect 3941 2565 3971 2580
rect 4137 2578 4337 2604
rect 4392 2578 4592 2604
rect 3848 2522 3884 2565
rect 3938 2522 3974 2565
rect 3788 2506 3884 2522
rect 3788 2472 3804 2506
rect 3838 2472 3884 2506
rect 3788 2456 3884 2472
rect 3854 2434 3884 2456
rect 3932 2506 4034 2522
rect 3932 2472 3984 2506
rect 4018 2472 4034 2506
rect 3932 2456 4034 2472
rect 4137 2513 4203 2578
rect 4137 2479 4153 2513
rect 4187 2479 4203 2513
rect 4137 2463 4203 2479
rect 4284 2512 4471 2528
rect 4284 2478 4300 2512
rect 4334 2478 4421 2512
rect 4455 2478 4471 2512
rect 3932 2434 3962 2456
rect 4284 2450 4471 2478
rect 4526 2513 4592 2578
rect 4526 2479 4542 2513
rect 4576 2479 4592 2513
rect 4526 2463 4592 2479
rect 5481 2578 5681 2604
rect 5736 2578 5936 2604
rect 5481 2513 5547 2578
rect 5481 2479 5497 2513
rect 5531 2479 5547 2513
rect 5481 2463 5547 2479
rect 5628 2512 5815 2528
rect 5628 2478 5644 2512
rect 5678 2478 5765 2512
rect 5799 2478 5815 2512
rect 4284 2421 4350 2450
rect 4150 2381 4350 2421
rect 4406 2421 4471 2450
rect 5628 2450 5815 2478
rect 5870 2513 5936 2578
rect 5870 2479 5886 2513
rect 5920 2479 5936 2513
rect 5870 2463 5936 2479
rect 6153 2578 6353 2604
rect 6408 2578 6608 2604
rect 6153 2513 6219 2578
rect 6153 2479 6169 2513
rect 6203 2479 6219 2513
rect 6153 2463 6219 2479
rect 6300 2512 6487 2528
rect 6300 2478 6316 2512
rect 6350 2478 6437 2512
rect 6471 2478 6487 2512
rect 4406 2381 4606 2421
rect 5628 2421 5694 2450
rect 5494 2381 5694 2421
rect 5750 2421 5815 2450
rect 6300 2450 6487 2478
rect 6542 2513 6608 2578
rect 6542 2479 6558 2513
rect 6592 2479 6608 2513
rect 6542 2463 6608 2479
rect 6825 2578 7025 2604
rect 7080 2578 7280 2604
rect 6825 2513 6891 2578
rect 6825 2479 6841 2513
rect 6875 2479 6891 2513
rect 6825 2463 6891 2479
rect 6972 2512 7159 2528
rect 6972 2478 6988 2512
rect 7022 2478 7109 2512
rect 7143 2478 7159 2512
rect 6300 2421 6366 2450
rect 5750 2381 5950 2421
rect 6166 2381 6366 2421
rect 6422 2421 6487 2450
rect 6972 2450 7159 2478
rect 7214 2513 7280 2578
rect 7214 2479 7230 2513
rect 7264 2479 7280 2513
rect 7214 2463 7280 2479
rect 8169 2578 8369 2604
rect 8424 2578 8624 2604
rect 8169 2513 8235 2578
rect 8169 2479 8185 2513
rect 8219 2479 8235 2513
rect 8169 2463 8235 2479
rect 8316 2512 8503 2528
rect 8316 2478 8332 2512
rect 8366 2478 8453 2512
rect 8487 2478 8503 2512
rect 6972 2421 7038 2450
rect 6422 2381 6622 2421
rect 6838 2381 7038 2421
rect 7094 2421 7159 2450
rect 8316 2450 8503 2478
rect 8558 2513 8624 2578
rect 8558 2479 8574 2513
rect 8608 2479 8624 2513
rect 8558 2463 8624 2479
rect 8841 2578 9041 2604
rect 9096 2578 9296 2604
rect 8841 2513 8907 2578
rect 8841 2479 8857 2513
rect 8891 2479 8907 2513
rect 8841 2463 8907 2479
rect 8988 2512 9175 2528
rect 8988 2478 9004 2512
rect 9038 2478 9125 2512
rect 9159 2478 9175 2512
rect 8316 2421 8382 2450
rect 7094 2381 7294 2421
rect 8182 2381 8382 2421
rect 8438 2421 8503 2450
rect 8988 2450 9175 2478
rect 9230 2513 9296 2578
rect 9230 2479 9246 2513
rect 9280 2479 9296 2513
rect 9230 2463 9296 2479
rect 9513 2578 9713 2604
rect 9513 2513 9579 2578
rect 9513 2479 9529 2513
rect 9563 2479 9579 2513
rect 9513 2463 9579 2479
rect 9660 2512 9726 2528
rect 9660 2478 9676 2512
rect 9710 2478 9726 2512
rect 8988 2421 9054 2450
rect 8438 2381 8638 2421
rect 8854 2381 9054 2421
rect 9110 2421 9175 2450
rect 9660 2421 9726 2478
rect 9110 2381 9310 2421
rect 9526 2381 9726 2421
rect 2499 2260 2529 2286
rect 3854 2260 3884 2286
rect 3932 2260 3962 2286
rect 4150 2259 4350 2297
rect 4406 2259 4606 2297
rect 5494 2259 5694 2297
rect 5750 2259 5950 2297
rect 6166 2259 6366 2297
rect 6422 2259 6622 2297
rect 6838 2259 7038 2297
rect 7094 2259 7294 2297
rect 8182 2259 8382 2297
rect 8438 2259 8638 2297
rect 8854 2259 9054 2297
rect 9110 2259 9310 2297
rect 9526 2259 9726 2297
rect 2499 2138 2529 2164
rect 3854 2138 3884 2164
rect 3932 2138 3962 2164
rect 4251 2138 4281 2164
rect 4329 2138 4359 2164
rect 4468 2138 4498 2164
rect 4660 2138 4690 2164
rect 4803 2138 4833 2164
rect 5006 2138 5036 2164
rect 5092 2138 5122 2164
rect 5566 2161 5976 2191
rect 2499 1952 2529 1990
rect 2356 1945 2530 1952
rect 2354 1936 2530 1945
rect 2354 1902 2372 1936
rect 2406 1902 2440 1936
rect 2474 1902 2530 1936
rect 2354 1893 2530 1902
rect 2356 1886 2530 1893
rect 2494 1859 2530 1886
rect 2497 1844 2527 1859
rect 4139 2100 4169 2126
rect 5488 2093 5518 2119
rect 5566 2093 5596 2161
rect 5732 2093 5762 2119
rect 5810 2093 5840 2119
rect 5946 2093 5976 2161
rect 6144 2114 6174 2140
rect 6312 2161 7396 2191
rect 6312 2114 6342 2161
rect 3854 1968 3884 1990
rect 3788 1952 3884 1968
rect 3788 1918 3804 1952
rect 3838 1918 3884 1952
rect 3788 1902 3884 1918
rect 3932 1968 3962 1990
rect 3932 1952 4034 1968
rect 3932 1918 3984 1952
rect 4018 1918 4034 1952
rect 4139 1942 4169 1990
rect 4251 1942 4281 1990
rect 4329 1968 4359 1990
rect 4468 1968 4498 1990
rect 3932 1902 4034 1918
rect 4138 1926 4281 1942
rect 3848 1859 3884 1902
rect 3938 1859 3974 1902
rect 4138 1892 4172 1926
rect 4206 1892 4281 1926
rect 4324 1952 4390 1968
rect 4324 1918 4340 1952
rect 4374 1918 4390 1952
rect 4324 1902 4390 1918
rect 4432 1952 4498 1968
rect 4432 1918 4448 1952
rect 4482 1918 4498 1952
rect 4432 1902 4498 1918
rect 4546 1952 4612 1968
rect 4546 1918 4562 1952
rect 4596 1918 4612 1952
rect 4546 1902 4612 1918
rect 4660 1948 4690 1990
rect 4803 1952 4833 1990
rect 5006 1952 5036 1990
rect 5092 1952 5122 1990
rect 5488 1987 5518 2009
rect 5566 1987 5596 2009
rect 5443 1971 5518 1987
rect 4660 1932 4726 1948
rect 4138 1876 4281 1892
rect 4138 1859 4174 1876
rect 4245 1859 4281 1876
rect 4438 1859 4474 1902
rect 4546 1859 4582 1902
rect 4660 1898 4676 1932
rect 4710 1898 4726 1932
rect 4660 1882 4726 1898
rect 4768 1936 4834 1952
rect 4768 1902 4784 1936
rect 4818 1902 4834 1936
rect 4768 1886 4834 1902
rect 4940 1936 5126 1952
rect 4940 1902 4956 1936
rect 4990 1922 5126 1936
rect 4990 1902 5036 1922
rect 4940 1886 5036 1902
rect 4660 1859 4696 1882
rect 4784 1859 4820 1886
rect 5000 1859 5036 1886
rect 5090 1859 5126 1922
rect 5443 1937 5459 1971
rect 5493 1937 5518 1971
rect 5443 1903 5518 1937
rect 5443 1869 5459 1903
rect 5493 1869 5518 1903
rect 3851 1844 3881 1859
rect 3941 1844 3971 1859
rect 4141 1844 4171 1859
rect 4248 1844 4278 1859
rect 4441 1844 4471 1859
rect 4549 1844 4579 1859
rect 4663 1844 4693 1859
rect 4787 1844 4817 1859
rect 5003 1844 5033 1859
rect 5093 1844 5123 1859
rect 4141 1650 4171 1676
rect 2497 1594 2527 1620
rect 3851 1594 3881 1620
rect 3941 1594 3971 1620
rect 4248 1618 4278 1644
rect 4441 1618 4471 1644
rect 4549 1618 4579 1644
rect 4663 1618 4693 1644
rect 5443 1835 5518 1869
rect 5560 1971 5626 1987
rect 5560 1937 5576 1971
rect 5610 1937 5626 1971
rect 5560 1903 5626 1937
rect 5732 1920 5762 2009
rect 5560 1869 5576 1903
rect 5610 1869 5626 1903
rect 5560 1853 5626 1869
rect 5668 1904 5762 1920
rect 5668 1870 5712 1904
rect 5746 1870 5762 1904
rect 5668 1854 5762 1870
rect 5810 1880 5840 2009
rect 5946 1994 5976 2009
rect 5946 1964 6064 1994
rect 6554 2087 6584 2113
rect 6626 2087 6656 2161
rect 7366 2130 7396 2161
rect 7616 2130 7646 2156
rect 7694 2130 7724 2156
rect 6717 2087 6747 2113
rect 6964 2087 6994 2113
rect 7050 2087 7080 2113
rect 7171 2087 7201 2113
rect 7271 2087 7301 2113
rect 6554 1988 6584 2003
rect 5920 1900 5986 1916
rect 5920 1880 5936 1900
rect 5810 1866 5936 1880
rect 5970 1866 5986 1900
rect 5443 1801 5459 1835
rect 5493 1801 5518 1835
rect 5443 1785 5518 1801
rect 5482 1763 5518 1785
rect 5572 1763 5608 1853
rect 5668 1805 5698 1854
rect 5650 1775 5698 1805
rect 5810 1850 5986 1866
rect 5810 1802 5840 1850
rect 6034 1802 6064 1964
rect 6144 1942 6174 1966
rect 6312 1944 6342 1966
rect 6112 1926 6180 1942
rect 6112 1892 6128 1926
rect 6162 1892 6180 1926
rect 6112 1876 6180 1892
rect 6222 1928 6342 1944
rect 6222 1894 6238 1928
rect 6272 1894 6342 1928
rect 6222 1878 6342 1894
rect 6440 1958 6584 1988
rect 6144 1859 6180 1876
rect 6234 1859 6270 1878
rect 6147 1844 6177 1859
rect 6237 1844 6267 1859
rect 6440 1846 6470 1958
rect 6518 1894 6584 1910
rect 6518 1860 6534 1894
rect 6568 1860 6584 1894
rect 5650 1763 5686 1775
rect 5740 1772 5840 1802
rect 5942 1772 6064 1802
rect 5740 1763 5776 1772
rect 5942 1763 5978 1772
rect 5485 1748 5515 1763
rect 5575 1748 5605 1763
rect 5653 1748 5683 1763
rect 5743 1748 5773 1763
rect 5945 1748 5975 1763
rect 4787 1594 4817 1620
rect 5003 1594 5033 1620
rect 5093 1594 5123 1620
rect 6406 1830 6472 1846
rect 6518 1844 6584 1860
rect 6406 1796 6422 1830
rect 6456 1796 6472 1830
rect 6406 1780 6472 1796
rect 6436 1763 6472 1780
rect 6520 1763 6556 1844
rect 6626 1793 6656 2003
rect 6717 1907 6747 2003
rect 7821 2138 7851 2164
rect 7925 2138 7955 2164
rect 8011 2138 8041 2164
rect 7366 2005 7396 2020
rect 6964 1955 6994 1977
rect 7050 1955 7080 1977
rect 6806 1939 6994 1955
rect 6698 1891 6764 1907
rect 6698 1857 6714 1891
rect 6748 1857 6764 1891
rect 6698 1841 6764 1857
rect 6806 1905 6822 1939
rect 6856 1925 6994 1939
rect 6856 1905 6872 1925
rect 6806 1871 6872 1905
rect 6806 1837 6822 1871
rect 6856 1837 6872 1871
rect 6806 1821 6872 1837
rect 6958 1803 6994 1925
rect 7042 1939 7108 1955
rect 7042 1905 7058 1939
rect 7092 1905 7108 1939
rect 7171 1922 7201 1977
rect 7042 1871 7108 1905
rect 7042 1837 7058 1871
rect 7092 1837 7108 1871
rect 7042 1821 7108 1837
rect 7150 1906 7223 1922
rect 7150 1872 7173 1906
rect 7207 1872 7223 1906
rect 7150 1856 7223 1872
rect 7271 1896 7301 1977
rect 7366 1975 7568 2005
rect 7430 1911 7496 1927
rect 7271 1880 7388 1896
rect 7042 1803 7078 1821
rect 7150 1803 7186 1856
rect 7271 1846 7338 1880
rect 7372 1846 7388 1880
rect 7271 1830 7388 1846
rect 7352 1803 7388 1830
rect 7430 1877 7446 1911
rect 7480 1877 7496 1911
rect 7430 1861 7496 1877
rect 7430 1803 7466 1861
rect 7538 1813 7568 1975
rect 7616 1959 7646 2046
rect 7694 2031 7724 2046
rect 7694 2001 7748 2031
rect 7610 1943 7676 1959
rect 7610 1909 7626 1943
rect 7660 1909 7676 1943
rect 7610 1893 7676 1909
rect 6626 1763 6663 1793
rect 6961 1788 6991 1803
rect 7045 1788 7075 1803
rect 7153 1788 7183 1803
rect 7355 1788 7385 1803
rect 7433 1788 7463 1803
rect 6439 1748 6469 1763
rect 6523 1748 6553 1763
rect 6630 1748 6660 1763
rect 6439 1638 6469 1664
rect 6523 1638 6553 1664
rect 7537 1719 7573 1813
rect 7718 1802 7748 2001
rect 8430 2138 8460 2164
rect 8516 2138 8546 2164
rect 8224 2032 8254 2058
rect 7821 1968 7851 1990
rect 7925 1968 7955 1990
rect 7790 1952 7856 1968
rect 7790 1918 7806 1952
rect 7840 1918 7856 1952
rect 7790 1902 7856 1918
rect 7898 1952 7964 1968
rect 7898 1918 7914 1952
rect 7948 1918 7964 1952
rect 8011 1918 8041 1990
rect 8728 2118 8758 2144
rect 8848 2138 8878 2164
rect 8934 2138 8964 2164
rect 9323 2138 9353 2164
rect 9409 2138 9439 2164
rect 9495 2138 9525 2164
rect 9581 2138 9611 2164
rect 9675 2138 9705 2164
rect 9767 2138 9797 2164
rect 9867 2138 9897 2164
rect 9980 2138 10010 2164
rect 7898 1902 7964 1918
rect 8006 1902 8072 1918
rect 8224 1911 8254 1948
rect 8430 1942 8460 1990
rect 8516 1942 8546 1990
rect 8728 1942 8758 1990
rect 8848 1968 8878 1990
rect 8934 1968 8964 1990
rect 8806 1952 8964 1968
rect 8430 1926 8764 1942
rect 7820 1835 7856 1902
rect 7922 1835 7958 1902
rect 8006 1868 8022 1902
rect 8056 1868 8072 1902
rect 8006 1852 8072 1868
rect 8188 1895 8254 1911
rect 8188 1861 8204 1895
rect 8238 1861 8254 1895
rect 8006 1835 8042 1852
rect 8188 1845 8254 1861
rect 8296 1910 8764 1926
rect 8296 1876 8312 1910
rect 8346 1883 8764 1910
rect 8806 1918 8822 1952
rect 8856 1918 8964 1952
rect 8806 1902 8964 1918
rect 8346 1876 8362 1883
rect 8296 1860 8362 1876
rect 8444 1859 8480 1883
rect 8534 1859 8570 1883
rect 8733 1882 8764 1883
rect 7823 1820 7853 1835
rect 7925 1820 7955 1835
rect 8009 1820 8039 1835
rect 8208 1828 8244 1845
rect 8447 1844 8477 1859
rect 8537 1844 8567 1859
rect 7615 1786 7748 1802
rect 7615 1752 7631 1786
rect 7665 1772 7748 1786
rect 7665 1752 7681 1772
rect 7615 1736 7681 1752
rect 7615 1719 7651 1736
rect 7540 1704 7570 1719
rect 7618 1704 7648 1719
rect 8211 1813 8241 1828
rect 8211 1659 8241 1685
rect 5485 1594 5515 1620
rect 5575 1594 5605 1620
rect 5653 1594 5683 1620
rect 5743 1594 5773 1620
rect 5945 1594 5975 1620
rect 6147 1594 6177 1620
rect 6237 1594 6267 1620
rect 6630 1594 6660 1620
rect 6961 1594 6991 1620
rect 7045 1594 7075 1620
rect 7153 1594 7183 1620
rect 7355 1594 7385 1620
rect 7433 1594 7463 1620
rect 7540 1594 7570 1620
rect 7618 1594 7648 1620
rect 7823 1594 7853 1620
rect 7925 1594 7955 1620
rect 8009 1594 8039 1620
rect 8733 1843 8769 1882
rect 8838 1859 8874 1902
rect 8928 1859 8964 1902
rect 9323 1942 9353 1990
rect 9409 1942 9439 1990
rect 9495 1942 9525 1990
rect 9581 1942 9611 1990
rect 9323 1926 9611 1942
rect 9323 1892 9357 1926
rect 9391 1892 9425 1926
rect 9459 1892 9493 1926
rect 9527 1892 9561 1926
rect 9595 1892 9611 1926
rect 9323 1876 9611 1892
rect 9323 1859 9359 1876
rect 9575 1859 9611 1876
rect 9675 1942 9705 1990
rect 9767 1942 9797 1990
rect 9867 1942 9897 1990
rect 9980 1942 10010 1990
rect 9675 1926 10010 1942
rect 9675 1892 9744 1926
rect 9778 1892 9812 1926
rect 9846 1892 9880 1926
rect 9914 1892 9948 1926
rect 9982 1892 10010 1926
rect 9675 1876 10010 1892
rect 9675 1859 9711 1876
rect 9974 1859 10010 1876
rect 8841 1844 8871 1859
rect 8931 1844 8961 1859
rect 9326 1844 9356 1859
rect 9578 1844 9608 1859
rect 9678 1844 9708 1859
rect 9977 1844 10007 1859
rect 8736 1828 8766 1843
rect 8447 1594 8477 1620
rect 8537 1594 8567 1620
rect 8736 1602 8766 1628
rect 8841 1594 8871 1620
rect 8931 1594 8961 1620
rect 9326 1594 9356 1620
rect 9578 1594 9608 1620
rect 9678 1594 9708 1620
rect 9977 1594 10007 1620
rect 11420 3818 11820 3834
rect 11420 3784 11436 3818
rect 11804 3784 11820 3818
rect 11420 3737 11820 3784
rect 11878 3818 12278 3834
rect 11878 3784 11894 3818
rect 12262 3784 12278 3818
rect 11878 3737 12278 3784
rect 12336 3818 12736 3834
rect 12336 3784 12352 3818
rect 12720 3784 12736 3818
rect 12336 3737 12736 3784
rect 12794 3818 13194 3834
rect 12794 3784 12810 3818
rect 13178 3784 13194 3818
rect 12794 3737 13194 3784
rect 13252 3818 13652 3834
rect 13252 3784 13268 3818
rect 13636 3784 13652 3818
rect 13252 3737 13652 3784
rect 11420 1690 11820 1737
rect 11420 1656 11436 1690
rect 11804 1656 11820 1690
rect 11420 1640 11820 1656
rect 11878 1690 12278 1737
rect 11878 1656 11894 1690
rect 12262 1656 12278 1690
rect 11878 1640 12278 1656
rect 12336 1690 12736 1737
rect 12336 1656 12352 1690
rect 12720 1656 12736 1690
rect 12336 1640 12736 1656
rect 12794 1690 13194 1737
rect 12794 1656 12810 1690
rect 13178 1656 13194 1690
rect 12794 1640 13194 1656
rect 13252 1690 13652 1737
rect 13252 1656 13268 1690
rect 13636 1656 13652 1690
rect 13252 1640 13652 1656
rect 13920 3768 13986 3834
rect 13938 3737 13968 3768
rect 13938 1706 13968 1737
rect 13920 1690 13986 1706
rect 13920 1656 13936 1690
rect 13970 1656 13986 1690
rect 13920 1640 13986 1656
rect 14236 3768 14302 3834
rect 14254 3737 14284 3768
rect 14254 1706 14284 1737
rect 14236 1690 14302 1706
rect 14236 1656 14252 1690
rect 14286 1656 14302 1690
rect 14236 1640 14302 1656
rect 3649 1472 3679 1498
rect 5003 1472 5033 1498
rect 5093 1472 5123 1498
rect 3649 1233 3679 1248
rect 3646 1206 3682 1233
rect 3508 1199 3682 1206
rect 3506 1190 3682 1199
rect 3506 1156 3524 1190
rect 3558 1156 3592 1190
rect 3626 1156 3682 1190
rect 3506 1147 3682 1156
rect 3508 1140 3682 1147
rect 3651 1102 3681 1140
rect 5485 1472 5515 1498
rect 5575 1472 5605 1498
rect 5653 1472 5683 1498
rect 5743 1472 5773 1498
rect 5945 1472 5975 1498
rect 6147 1472 6177 1498
rect 6237 1472 6267 1498
rect 6630 1472 6660 1498
rect 6961 1472 6991 1498
rect 7045 1472 7075 1498
rect 7153 1472 7183 1498
rect 7355 1472 7385 1498
rect 7433 1472 7463 1498
rect 7540 1472 7570 1498
rect 7618 1472 7648 1498
rect 7823 1472 7853 1498
rect 7925 1472 7955 1498
rect 8009 1472 8039 1498
rect 5485 1329 5515 1344
rect 5575 1329 5605 1344
rect 5653 1329 5683 1344
rect 5743 1329 5773 1344
rect 5945 1329 5975 1344
rect 5482 1307 5518 1329
rect 5443 1291 5518 1307
rect 5443 1257 5459 1291
rect 5493 1257 5518 1291
rect 5003 1233 5033 1248
rect 5093 1233 5123 1248
rect 5000 1190 5036 1233
rect 5090 1190 5126 1233
rect 5443 1223 5518 1257
rect 5572 1239 5608 1329
rect 5650 1317 5686 1329
rect 5740 1320 5776 1329
rect 5942 1320 5978 1329
rect 5650 1287 5698 1317
rect 5740 1290 5840 1320
rect 5942 1290 6064 1320
rect 4940 1174 5036 1190
rect 4940 1140 4956 1174
rect 4990 1140 5036 1174
rect 4940 1124 5036 1140
rect 5006 1102 5036 1124
rect 5084 1174 5186 1190
rect 5084 1140 5136 1174
rect 5170 1140 5186 1174
rect 5084 1124 5186 1140
rect 5443 1189 5459 1223
rect 5493 1189 5518 1223
rect 5443 1155 5518 1189
rect 5084 1102 5114 1124
rect 5443 1121 5459 1155
rect 5493 1121 5518 1155
rect 5443 1105 5518 1121
rect 5560 1223 5626 1239
rect 5560 1189 5576 1223
rect 5610 1189 5626 1223
rect 5560 1155 5626 1189
rect 5668 1238 5698 1287
rect 5810 1242 5840 1290
rect 5668 1222 5762 1238
rect 5668 1188 5712 1222
rect 5746 1188 5762 1222
rect 5668 1172 5762 1188
rect 5560 1121 5576 1155
rect 5610 1121 5626 1155
rect 5560 1105 5626 1121
rect 5488 1083 5518 1105
rect 5566 1083 5596 1105
rect 5732 1083 5762 1172
rect 5810 1226 5986 1242
rect 5810 1212 5936 1226
rect 5810 1083 5840 1212
rect 5920 1192 5936 1212
rect 5970 1192 5986 1226
rect 5920 1176 5986 1192
rect 6034 1128 6064 1290
rect 6439 1428 6469 1454
rect 6523 1428 6553 1454
rect 6439 1329 6469 1344
rect 6523 1329 6553 1344
rect 6630 1329 6660 1344
rect 6436 1312 6472 1329
rect 6406 1296 6472 1312
rect 6406 1262 6422 1296
rect 6456 1262 6472 1296
rect 6147 1233 6177 1248
rect 6237 1233 6267 1248
rect 6406 1246 6472 1262
rect 6520 1248 6556 1329
rect 6626 1299 6663 1329
rect 7540 1373 7570 1388
rect 7618 1373 7648 1388
rect 6144 1216 6180 1233
rect 6112 1200 6180 1216
rect 6234 1214 6270 1233
rect 6112 1166 6128 1200
rect 6162 1166 6180 1200
rect 6112 1150 6180 1166
rect 6222 1198 6342 1214
rect 6222 1164 6238 1198
rect 6272 1164 6342 1198
rect 5946 1098 6064 1128
rect 6144 1126 6174 1150
rect 6222 1148 6342 1164
rect 6312 1126 6342 1148
rect 6440 1134 6470 1246
rect 6518 1232 6584 1248
rect 6518 1198 6534 1232
rect 6568 1198 6584 1232
rect 6518 1182 6584 1198
rect 5946 1083 5976 1098
rect 5488 973 5518 999
rect 3651 928 3681 954
rect 5006 928 5036 954
rect 5084 928 5114 954
rect 5566 931 5596 999
rect 5732 973 5762 999
rect 5810 973 5840 999
rect 5946 931 5976 999
rect 6440 1104 6584 1134
rect 6554 1089 6584 1104
rect 6626 1089 6656 1299
rect 6961 1289 6991 1304
rect 7045 1289 7075 1304
rect 7153 1289 7183 1304
rect 7355 1289 7385 1304
rect 7433 1289 7463 1304
rect 6806 1255 6872 1271
rect 6698 1235 6764 1251
rect 6698 1201 6714 1235
rect 6748 1201 6764 1235
rect 6698 1185 6764 1201
rect 6806 1221 6822 1255
rect 6856 1221 6872 1255
rect 6806 1187 6872 1221
rect 6717 1089 6747 1185
rect 6806 1153 6822 1187
rect 6856 1167 6872 1187
rect 6958 1167 6994 1289
rect 6856 1153 6994 1167
rect 6806 1137 6994 1153
rect 7042 1271 7078 1289
rect 7042 1255 7108 1271
rect 7042 1221 7058 1255
rect 7092 1221 7108 1255
rect 7042 1187 7108 1221
rect 7042 1153 7058 1187
rect 7092 1153 7108 1187
rect 7150 1236 7186 1289
rect 7352 1262 7388 1289
rect 7271 1246 7388 1262
rect 7150 1220 7223 1236
rect 7150 1186 7173 1220
rect 7207 1186 7223 1220
rect 7150 1170 7223 1186
rect 7271 1212 7338 1246
rect 7372 1212 7388 1246
rect 7271 1196 7388 1212
rect 7430 1231 7466 1289
rect 7537 1279 7573 1373
rect 7615 1356 7651 1373
rect 7615 1340 7681 1356
rect 7615 1306 7631 1340
rect 7665 1320 7681 1340
rect 7665 1306 7748 1320
rect 7615 1290 7748 1306
rect 7430 1215 7496 1231
rect 7042 1137 7108 1153
rect 6964 1115 6994 1137
rect 7050 1115 7080 1137
rect 7171 1115 7201 1170
rect 7271 1115 7301 1196
rect 7430 1181 7446 1215
rect 7480 1181 7496 1215
rect 7430 1165 7496 1181
rect 7538 1117 7568 1279
rect 7610 1183 7676 1199
rect 7610 1149 7626 1183
rect 7660 1149 7676 1183
rect 7610 1133 7676 1149
rect 7366 1087 7568 1117
rect 7366 1072 7396 1087
rect 6144 952 6174 978
rect 5566 901 5976 931
rect 6312 931 6342 978
rect 6554 979 6584 1005
rect 6626 931 6656 1005
rect 6717 979 6747 1005
rect 6964 979 6994 1005
rect 7050 979 7080 1005
rect 7171 979 7201 1005
rect 7271 979 7301 1005
rect 7616 1046 7646 1133
rect 7718 1091 7748 1290
rect 8447 1472 8477 1498
rect 8537 1472 8567 1498
rect 8211 1407 8241 1433
rect 7823 1257 7853 1272
rect 7925 1257 7955 1272
rect 8009 1257 8039 1272
rect 8211 1264 8241 1279
rect 7820 1190 7856 1257
rect 7922 1190 7958 1257
rect 8006 1240 8042 1257
rect 8208 1247 8244 1264
rect 8736 1464 8766 1490
rect 8841 1472 8871 1498
rect 8931 1472 8961 1498
rect 8736 1249 8766 1264
rect 8006 1224 8072 1240
rect 8006 1190 8022 1224
rect 8056 1190 8072 1224
rect 7790 1174 7856 1190
rect 7790 1140 7806 1174
rect 7840 1140 7856 1174
rect 7790 1124 7856 1140
rect 7898 1174 7964 1190
rect 8006 1174 8072 1190
rect 8188 1231 8254 1247
rect 8447 1233 8477 1248
rect 8537 1233 8567 1248
rect 8188 1197 8204 1231
rect 8238 1197 8254 1231
rect 8188 1181 8254 1197
rect 7898 1140 7914 1174
rect 7948 1140 7964 1174
rect 7898 1124 7964 1140
rect 7821 1102 7851 1124
rect 7925 1102 7955 1124
rect 8011 1102 8041 1174
rect 8224 1144 8254 1181
rect 8296 1216 8362 1232
rect 8296 1182 8312 1216
rect 8346 1209 8362 1216
rect 8444 1209 8480 1233
rect 8534 1209 8570 1233
rect 8733 1210 8769 1249
rect 9326 1457 9356 1483
rect 9416 1457 9446 1483
rect 9511 1457 9541 1483
rect 9606 1457 9636 1483
rect 9713 1472 9743 1498
rect 9807 1472 9837 1498
rect 9897 1472 9927 1498
rect 9987 1472 10017 1498
rect 9326 1274 9356 1289
rect 9416 1274 9446 1289
rect 9511 1274 9541 1289
rect 9606 1274 9636 1289
rect 8841 1233 8871 1248
rect 8931 1233 8961 1248
rect 8733 1209 8764 1210
rect 8346 1182 8764 1209
rect 8838 1190 8874 1233
rect 8928 1190 8964 1233
rect 8296 1166 8764 1182
rect 8430 1150 8764 1166
rect 8806 1174 8964 1190
rect 7694 1061 7748 1091
rect 7694 1046 7724 1061
rect 7366 931 7396 962
rect 7616 936 7646 962
rect 7694 936 7724 962
rect 6312 901 7396 931
rect 8430 1102 8460 1150
rect 8516 1102 8546 1150
rect 8728 1102 8758 1150
rect 8806 1140 8822 1174
rect 8856 1140 8964 1174
rect 8806 1124 8964 1140
rect 9323 1142 9359 1274
rect 9413 1263 9449 1274
rect 9508 1263 9544 1274
rect 9413 1220 9544 1263
rect 9413 1186 9468 1220
rect 9502 1186 9544 1220
rect 9603 1215 9639 1274
rect 9713 1233 9743 1248
rect 9807 1233 9837 1248
rect 9897 1233 9927 1248
rect 9987 1233 10017 1248
rect 9710 1215 9746 1233
rect 9804 1215 9840 1233
rect 9894 1215 9930 1233
rect 9984 1215 10020 1233
rect 9413 1170 9544 1186
rect 9586 1199 9652 1215
rect 9323 1127 9353 1142
rect 9413 1127 9443 1170
rect 9508 1127 9538 1170
rect 9586 1165 9602 1199
rect 9636 1165 9652 1199
rect 9586 1149 9652 1165
rect 9700 1199 10020 1215
rect 9700 1165 9716 1199
rect 9750 1165 9784 1199
rect 9818 1165 9852 1199
rect 9886 1165 10020 1199
rect 9700 1149 10020 1165
rect 9599 1127 9629 1149
rect 9701 1127 9731 1149
rect 9817 1127 9847 1149
rect 9903 1127 9933 1149
rect 9989 1127 10019 1149
rect 8848 1102 8878 1124
rect 8934 1102 8964 1124
rect 8224 1034 8254 1060
rect 7821 928 7851 954
rect 7925 928 7955 954
rect 8011 928 8041 954
rect 8430 928 8460 954
rect 8516 928 8546 954
rect 8728 948 8758 974
rect 8848 928 8878 954
rect 8934 928 8964 954
rect 9323 931 9353 999
rect 9413 973 9443 999
rect 9508 973 9538 999
rect 9599 931 9629 999
rect 9701 953 9731 979
rect 9817 953 9847 979
rect 9903 953 9933 979
rect 9989 953 10019 979
rect 9323 901 9629 931
rect 3846 604 3912 670
rect 3864 582 3894 604
rect 3864 160 3894 182
rect 3846 144 3912 160
rect 3846 110 3862 144
rect 3896 110 3912 144
rect 3846 94 3912 110
rect 10504 1380 10904 1396
rect 10504 1346 10520 1380
rect 10888 1346 10904 1380
rect 10504 1308 10904 1346
rect 10962 1380 11362 1396
rect 10962 1346 10978 1380
rect 11346 1346 11362 1380
rect 10962 1308 11362 1346
rect 11420 1380 11820 1396
rect 11420 1346 11436 1380
rect 11804 1346 11820 1380
rect 11420 1308 11820 1346
rect 11878 1380 12278 1396
rect 11878 1346 11894 1380
rect 12262 1346 12278 1380
rect 11878 1308 12278 1346
rect 12336 1380 12736 1396
rect 12336 1346 12352 1380
rect 12720 1346 12736 1380
rect 12336 1308 12736 1346
rect 12794 1380 13194 1396
rect 12794 1346 12810 1380
rect 13178 1346 13194 1380
rect 12794 1308 13194 1346
rect 13252 1380 13652 1396
rect 13252 1346 13268 1380
rect 13636 1346 13652 1380
rect 13252 1308 13652 1346
rect 10504 270 10904 308
rect 10504 236 10520 270
rect 10888 236 10904 270
rect 10504 220 10904 236
rect 10962 270 11362 308
rect 10962 236 10978 270
rect 11346 236 11362 270
rect 10962 220 11362 236
rect 11420 270 11820 308
rect 11420 236 11436 270
rect 11804 236 11820 270
rect 11420 220 11820 236
rect 11878 270 12278 308
rect 11878 236 11894 270
rect 12262 236 12278 270
rect 11878 220 12278 236
rect 12336 270 12736 308
rect 12336 236 12352 270
rect 12720 236 12736 270
rect 12336 220 12736 236
rect 12794 270 13194 308
rect 12794 236 12810 270
rect 13178 236 13194 270
rect 12794 220 13194 236
rect 13252 270 13652 308
rect 13252 236 13268 270
rect 13636 236 13652 270
rect 13252 220 13652 236
rect 13920 1380 13986 1396
rect 13920 1346 13936 1380
rect 13970 1346 13986 1380
rect 13920 1330 13986 1346
rect 13938 1308 13968 1330
rect 13938 286 13968 308
rect 13920 220 13986 286
rect 14236 1380 14302 1396
rect 14236 1346 14252 1380
rect 14286 1346 14302 1380
rect 14236 1330 14302 1346
rect 14254 1308 14284 1330
rect 14254 286 14284 308
rect 14236 220 14302 286
rect 15452 855 15518 873
rect 15962 857 16028 873
rect 15962 855 15978 857
rect 15452 825 15540 855
rect 15940 825 15978 855
rect 15452 807 15518 825
rect 15962 823 15978 825
rect 16012 823 16028 857
rect 15962 807 16028 823
rect 16166 855 16232 873
rect 16676 857 16742 873
rect 16676 855 16692 857
rect 16166 825 16254 855
rect 16654 825 16692 855
rect 16166 807 16232 825
rect 16676 823 16692 825
rect 16726 823 16742 857
rect 16676 807 16742 823
rect 16880 855 16946 873
rect 17390 857 17456 873
rect 17390 855 17406 857
rect 16880 825 16968 855
rect 17368 825 17406 855
rect 16880 807 16946 825
rect 17390 823 17406 825
rect 17440 823 17456 857
rect 17390 807 17456 823
rect 17594 855 17660 873
rect 18104 857 18170 873
rect 18104 855 18120 857
rect 17594 825 17682 855
rect 18082 825 18120 855
rect 17594 807 17660 825
rect 18104 823 18120 825
rect 18154 823 18170 857
rect 18104 807 18170 823
rect 18308 855 18374 873
rect 18818 857 18884 873
rect 18818 855 18834 857
rect 18308 825 18396 855
rect 18796 825 18834 855
rect 18308 807 18374 825
rect 18818 823 18834 825
rect 18868 823 18884 857
rect 18818 807 18884 823
rect 19022 855 19088 873
rect 19532 857 19598 873
rect 19532 855 19548 857
rect 19022 825 19110 855
rect 19510 825 19548 855
rect 19022 807 19088 825
rect 19532 823 19548 825
rect 19582 823 19598 857
rect 19532 807 19598 823
rect 19736 855 19802 873
rect 20246 857 20312 873
rect 20246 855 20262 857
rect 19736 825 19824 855
rect 20224 825 20262 855
rect 19736 807 19802 825
rect 20246 823 20262 825
rect 20296 823 20312 857
rect 20246 807 20312 823
rect 20450 855 20516 873
rect 20960 857 21026 873
rect 20960 855 20976 857
rect 20450 825 20538 855
rect 20938 825 20976 855
rect 20450 807 20516 825
rect 20960 823 20976 825
rect 21010 823 21026 857
rect 20960 807 21026 823
rect 21164 855 21230 873
rect 21674 857 21740 873
rect 21674 855 21690 857
rect 21164 825 21252 855
rect 21652 825 21690 855
rect 21164 807 21230 825
rect 21674 823 21690 825
rect 21724 823 21740 857
rect 21674 807 21740 823
rect 21878 855 21944 873
rect 22388 857 22454 873
rect 22388 855 22404 857
rect 21878 825 21966 855
rect 22366 825 22404 855
rect 21878 807 21944 825
rect 22388 823 22404 825
rect 22438 823 22454 857
rect 22388 807 22454 823
rect 22592 855 22658 873
rect 23102 857 23168 873
rect 23102 855 23118 857
rect 22592 825 22680 855
rect 23080 825 23118 855
rect 22592 807 22658 825
rect 23102 823 23118 825
rect 23152 823 23168 857
rect 23102 807 23168 823
rect 23306 855 23372 873
rect 23816 857 23882 873
rect 23816 855 23832 857
rect 23306 825 23394 855
rect 23794 825 23832 855
rect 23306 807 23372 825
rect 23816 823 23832 825
rect 23866 823 23882 857
rect 23816 807 23882 823
rect 24020 855 24086 873
rect 24530 857 24596 873
rect 24530 855 24546 857
rect 24020 825 24108 855
rect 24508 825 24546 855
rect 24020 807 24086 825
rect 24530 823 24546 825
rect 24580 823 24596 857
rect 24530 807 24596 823
rect 24734 855 24800 873
rect 25244 857 25310 873
rect 25244 855 25260 857
rect 24734 825 24822 855
rect 25222 825 25260 855
rect 24734 807 24800 825
rect 25244 823 25260 825
rect 25294 823 25310 857
rect 25244 807 25310 823
rect 25448 855 25514 873
rect 25958 857 26024 873
rect 25958 855 25974 857
rect 25448 825 25536 855
rect 25936 825 25974 855
rect 25448 807 25514 825
rect 25958 823 25974 825
rect 26008 823 26024 857
rect 25958 807 26024 823
rect 26162 855 26228 873
rect 26672 857 26738 873
rect 26672 855 26688 857
rect 26162 825 26250 855
rect 26650 825 26688 855
rect 26162 807 26228 825
rect 26672 823 26688 825
rect 26722 823 26738 857
rect 26672 807 26738 823
rect 26876 855 26942 873
rect 27386 857 27452 873
rect 27386 855 27402 857
rect 26876 825 26964 855
rect 27364 825 27402 855
rect 26876 807 26942 825
rect 27386 823 27402 825
rect 27436 823 27452 857
rect 27386 807 27452 823
rect 27590 855 27656 873
rect 28100 857 28166 873
rect 28100 855 28116 857
rect 27590 825 27678 855
rect 28078 825 28116 855
rect 27590 807 27656 825
rect 28100 823 28116 825
rect 28150 823 28166 857
rect 28100 807 28166 823
rect 28304 855 28370 873
rect 28814 857 28880 873
rect 28814 855 28830 857
rect 28304 825 28392 855
rect 28792 825 28830 855
rect 28304 807 28370 825
rect 28814 823 28830 825
rect 28864 823 28880 857
rect 28814 807 28880 823
rect 29018 855 29084 873
rect 29528 857 29594 873
rect 29528 855 29544 857
rect 29018 825 29106 855
rect 29506 825 29544 855
rect 29018 807 29084 825
rect 29528 823 29544 825
rect 29578 823 29594 857
rect 29528 807 29594 823
rect 29732 855 29798 873
rect 30242 857 30308 873
rect 30242 855 30258 857
rect 29732 825 29820 855
rect 30220 825 30258 855
rect 29732 807 29798 825
rect 30242 823 30258 825
rect 30292 823 30308 857
rect 30242 807 30308 823
rect 30446 855 30512 873
rect 30956 857 31022 873
rect 30956 855 30972 857
rect 30446 825 30534 855
rect 30934 825 30972 855
rect 30446 807 30512 825
rect 30956 823 30972 825
rect 31006 823 31022 857
rect 30956 807 31022 823
rect 31160 855 31226 873
rect 31670 857 31736 873
rect 31670 855 31686 857
rect 31160 825 31248 855
rect 31648 825 31686 855
rect 31160 807 31226 825
rect 31670 823 31686 825
rect 31720 823 31736 857
rect 31670 807 31736 823
rect 31874 855 31940 873
rect 32384 857 32450 873
rect 32384 855 32400 857
rect 31874 825 31962 855
rect 32362 825 32400 855
rect 31874 807 31940 825
rect 32384 823 32400 825
rect 32434 823 32450 857
rect 32384 807 32450 823
rect 32588 855 32654 873
rect 33098 857 33164 873
rect 33098 855 33114 857
rect 32588 825 32676 855
rect 33076 825 33114 855
rect 32588 807 32654 825
rect 33098 823 33114 825
rect 33148 823 33164 857
rect 33098 807 33164 823
rect 33302 855 33368 873
rect 33812 857 33878 873
rect 33812 855 33828 857
rect 33302 825 33390 855
rect 33790 825 33828 855
rect 33302 807 33368 825
rect 33812 823 33828 825
rect 33862 823 33878 857
rect 33812 807 33878 823
rect 34016 855 34082 873
rect 34526 857 34592 873
rect 34526 855 34542 857
rect 34016 825 34104 855
rect 34504 825 34542 855
rect 34016 807 34082 825
rect 34526 823 34542 825
rect 34576 823 34592 857
rect 34526 807 34592 823
rect 34730 855 34796 873
rect 35240 857 35306 873
rect 35240 855 35256 857
rect 34730 825 34818 855
rect 35218 825 35256 855
rect 34730 807 34796 825
rect 35240 823 35256 825
rect 35290 823 35306 857
rect 35240 807 35306 823
rect 35444 855 35510 873
rect 35954 857 36020 873
rect 35954 855 35970 857
rect 35444 825 35532 855
rect 35932 825 35970 855
rect 35444 807 35510 825
rect 35954 823 35970 825
rect 36004 823 36020 857
rect 35954 807 36020 823
rect 36158 855 36224 873
rect 36668 857 36734 873
rect 36668 855 36684 857
rect 36158 825 36246 855
rect 36646 825 36684 855
rect 36158 807 36224 825
rect 36668 823 36684 825
rect 36718 823 36734 857
rect 36668 807 36734 823
rect 36872 855 36938 873
rect 37382 857 37448 873
rect 37382 855 37398 857
rect 36872 825 36960 855
rect 37360 825 37398 855
rect 36872 807 36938 825
rect 37382 823 37398 825
rect 37432 823 37448 857
rect 37382 807 37448 823
rect 37586 855 37652 873
rect 38096 857 38162 873
rect 38096 855 38112 857
rect 37586 825 37674 855
rect 38074 825 38112 855
rect 37586 807 37652 825
rect 38096 823 38112 825
rect 38146 823 38162 857
rect 38096 807 38162 823
rect 38300 855 38366 873
rect 38810 857 38876 873
rect 38810 855 38826 857
rect 38300 825 38388 855
rect 38788 825 38826 855
rect 38300 807 38366 825
rect 38810 823 38826 825
rect 38860 823 38876 857
rect 38810 807 38876 823
rect 3846 -110 3912 -44
rect 3864 -132 3894 -110
rect 3864 -554 3894 -532
rect 3846 -570 3912 -554
rect 3846 -604 3862 -570
rect 3896 -604 3912 -570
rect 3846 -620 3912 -604
rect 15452 37 15518 55
rect 15962 39 16028 55
rect 15962 37 15978 39
rect 15452 7 15540 37
rect 15940 7 15978 37
rect 15452 -11 15518 7
rect 15962 5 15978 7
rect 16012 5 16028 39
rect 15962 -11 16028 5
rect 16166 37 16232 55
rect 16676 39 16742 55
rect 16676 37 16692 39
rect 16166 7 16254 37
rect 16654 7 16692 37
rect 16166 -11 16232 7
rect 16676 5 16692 7
rect 16726 5 16742 39
rect 16676 -11 16742 5
rect 16880 37 16946 55
rect 17390 39 17456 55
rect 17390 37 17406 39
rect 16880 7 16968 37
rect 17368 7 17406 37
rect 16880 -11 16946 7
rect 17390 5 17406 7
rect 17440 5 17456 39
rect 17390 -11 17456 5
rect 17594 37 17660 55
rect 18104 39 18170 55
rect 18104 37 18120 39
rect 17594 7 17682 37
rect 18082 7 18120 37
rect 17594 -11 17660 7
rect 18104 5 18120 7
rect 18154 5 18170 39
rect 18104 -11 18170 5
rect 18308 37 18374 55
rect 18818 39 18884 55
rect 18818 37 18834 39
rect 18308 7 18396 37
rect 18796 7 18834 37
rect 18308 -11 18374 7
rect 18818 5 18834 7
rect 18868 5 18884 39
rect 18818 -11 18884 5
rect 19022 37 19088 55
rect 19532 39 19598 55
rect 19532 37 19548 39
rect 19022 7 19110 37
rect 19510 7 19548 37
rect 19022 -11 19088 7
rect 19532 5 19548 7
rect 19582 5 19598 39
rect 19532 -11 19598 5
rect 19736 37 19802 55
rect 20246 39 20312 55
rect 20246 37 20262 39
rect 19736 7 19824 37
rect 20224 7 20262 37
rect 19736 -11 19802 7
rect 20246 5 20262 7
rect 20296 5 20312 39
rect 20246 -11 20312 5
rect 20450 37 20516 55
rect 20960 39 21026 55
rect 20960 37 20976 39
rect 20450 7 20538 37
rect 20938 7 20976 37
rect 20450 -11 20516 7
rect 20960 5 20976 7
rect 21010 5 21026 39
rect 20960 -11 21026 5
rect 21164 37 21230 55
rect 21674 39 21740 55
rect 21674 37 21690 39
rect 21164 7 21252 37
rect 21652 7 21690 37
rect 21164 -11 21230 7
rect 21674 5 21690 7
rect 21724 5 21740 39
rect 21674 -11 21740 5
rect 21878 37 21944 55
rect 22388 39 22454 55
rect 22388 37 22404 39
rect 21878 7 21966 37
rect 22366 7 22404 37
rect 21878 -11 21944 7
rect 22388 5 22404 7
rect 22438 5 22454 39
rect 22388 -11 22454 5
rect 22592 37 22658 55
rect 23102 39 23168 55
rect 23102 37 23118 39
rect 22592 7 22680 37
rect 23080 7 23118 37
rect 22592 -11 22658 7
rect 23102 5 23118 7
rect 23152 5 23168 39
rect 23102 -11 23168 5
rect 23306 37 23372 55
rect 23816 39 23882 55
rect 23816 37 23832 39
rect 23306 7 23394 37
rect 23794 7 23832 37
rect 23306 -11 23372 7
rect 23816 5 23832 7
rect 23866 5 23882 39
rect 23816 -11 23882 5
rect 24020 37 24086 55
rect 24530 39 24596 55
rect 24530 37 24546 39
rect 24020 7 24108 37
rect 24508 7 24546 37
rect 24020 -11 24086 7
rect 24530 5 24546 7
rect 24580 5 24596 39
rect 24530 -11 24596 5
rect 24734 37 24800 55
rect 25244 39 25310 55
rect 25244 37 25260 39
rect 24734 7 24822 37
rect 25222 7 25260 37
rect 24734 -11 24800 7
rect 25244 5 25260 7
rect 25294 5 25310 39
rect 25244 -11 25310 5
rect 25448 37 25514 55
rect 25958 39 26024 55
rect 25958 37 25974 39
rect 25448 7 25536 37
rect 25936 7 25974 37
rect 25448 -11 25514 7
rect 25958 5 25974 7
rect 26008 5 26024 39
rect 25958 -11 26024 5
rect 26162 37 26228 55
rect 26672 39 26738 55
rect 26672 37 26688 39
rect 26162 7 26250 37
rect 26650 7 26688 37
rect 26162 -11 26228 7
rect 26672 5 26688 7
rect 26722 5 26738 39
rect 26672 -11 26738 5
rect 26876 37 26942 55
rect 27386 39 27452 55
rect 27386 37 27402 39
rect 26876 7 26964 37
rect 27364 7 27402 37
rect 26876 -11 26942 7
rect 27386 5 27402 7
rect 27436 5 27452 39
rect 27386 -11 27452 5
rect 27590 37 27656 55
rect 28100 39 28166 55
rect 28100 37 28116 39
rect 27590 7 27678 37
rect 28078 7 28116 37
rect 27590 -11 27656 7
rect 28100 5 28116 7
rect 28150 5 28166 39
rect 28100 -11 28166 5
rect 28304 37 28370 55
rect 28814 39 28880 55
rect 28814 37 28830 39
rect 28304 7 28392 37
rect 28792 7 28830 37
rect 28304 -11 28370 7
rect 28814 5 28830 7
rect 28864 5 28880 39
rect 28814 -11 28880 5
rect 29018 37 29084 55
rect 29528 39 29594 55
rect 29528 37 29544 39
rect 29018 7 29106 37
rect 29506 7 29544 37
rect 29018 -11 29084 7
rect 29528 5 29544 7
rect 29578 5 29594 39
rect 29528 -11 29594 5
rect 29732 37 29798 55
rect 30242 39 30308 55
rect 30242 37 30258 39
rect 29732 7 29820 37
rect 30220 7 30258 37
rect 29732 -11 29798 7
rect 30242 5 30258 7
rect 30292 5 30308 39
rect 30242 -11 30308 5
rect 30446 37 30512 55
rect 30956 39 31022 55
rect 30956 37 30972 39
rect 30446 7 30534 37
rect 30934 7 30972 37
rect 30446 -11 30512 7
rect 30956 5 30972 7
rect 31006 5 31022 39
rect 30956 -11 31022 5
rect 31160 37 31226 55
rect 31670 39 31736 55
rect 31670 37 31686 39
rect 31160 7 31248 37
rect 31648 7 31686 37
rect 31160 -11 31226 7
rect 31670 5 31686 7
rect 31720 5 31736 39
rect 31670 -11 31736 5
rect 31874 37 31940 55
rect 32384 39 32450 55
rect 32384 37 32400 39
rect 31874 7 31962 37
rect 32362 7 32400 37
rect 31874 -11 31940 7
rect 32384 5 32400 7
rect 32434 5 32450 39
rect 32384 -11 32450 5
rect 32588 37 32654 55
rect 33098 39 33164 55
rect 33098 37 33114 39
rect 32588 7 32676 37
rect 33076 7 33114 37
rect 32588 -11 32654 7
rect 33098 5 33114 7
rect 33148 5 33164 39
rect 33098 -11 33164 5
rect 33302 37 33368 55
rect 33812 39 33878 55
rect 33812 37 33828 39
rect 33302 7 33390 37
rect 33790 7 33828 37
rect 33302 -11 33368 7
rect 33812 5 33828 7
rect 33862 5 33878 39
rect 33812 -11 33878 5
rect 34016 37 34082 55
rect 34526 39 34592 55
rect 34526 37 34542 39
rect 34016 7 34104 37
rect 34504 7 34542 37
rect 34016 -11 34082 7
rect 34526 5 34542 7
rect 34576 5 34592 39
rect 34526 -11 34592 5
rect 34730 37 34796 55
rect 35240 39 35306 55
rect 35240 37 35256 39
rect 34730 7 34818 37
rect 35218 7 35256 37
rect 34730 -11 34796 7
rect 35240 5 35256 7
rect 35290 5 35306 39
rect 35240 -11 35306 5
rect 35444 37 35510 55
rect 35954 39 36020 55
rect 35954 37 35970 39
rect 35444 7 35532 37
rect 35932 7 35970 37
rect 35444 -11 35510 7
rect 35954 5 35970 7
rect 36004 5 36020 39
rect 35954 -11 36020 5
rect 36158 37 36224 55
rect 36668 39 36734 55
rect 36668 37 36684 39
rect 36158 7 36246 37
rect 36646 7 36684 37
rect 36158 -11 36224 7
rect 36668 5 36684 7
rect 36718 5 36734 39
rect 36668 -11 36734 5
rect 36872 37 36938 55
rect 37382 39 37448 55
rect 37382 37 37398 39
rect 36872 7 36960 37
rect 37360 7 37398 37
rect 36872 -11 36938 7
rect 37382 5 37398 7
rect 37432 5 37448 39
rect 37382 -11 37448 5
rect 37586 37 37652 55
rect 38096 39 38162 55
rect 38096 37 38112 39
rect 37586 7 37674 37
rect 38074 7 38112 37
rect 37586 -11 37652 7
rect 38096 5 38112 7
rect 38146 5 38162 39
rect 38096 -11 38162 5
rect 38300 37 38366 55
rect 38810 39 38876 55
rect 38810 37 38826 39
rect 38300 7 38388 37
rect 38788 7 38826 37
rect 38300 -11 38366 7
rect 38810 5 38826 7
rect 38860 5 38876 39
rect 38810 -11 38876 5
rect 10269 -878 10295 -848
rect 10495 -878 10615 -848
rect 10745 -878 10771 -848
rect 10527 -884 10593 -878
rect 10527 -918 10543 -884
rect 10577 -918 10593 -884
rect 10527 -934 10593 -918
rect 5902 -4304 5968 -4288
rect 5902 -4338 5918 -4304
rect 5952 -4338 5968 -4304
rect 5902 -4354 5968 -4338
rect 6020 -4304 6086 -4288
rect 6020 -4338 6036 -4304
rect 6070 -4338 6086 -4304
rect 6020 -4354 6086 -4338
rect 6138 -4304 6204 -4288
rect 6138 -4338 6154 -4304
rect 6188 -4338 6204 -4304
rect 6138 -4354 6204 -4338
rect 6256 -4304 6322 -4288
rect 6256 -4338 6272 -4304
rect 6306 -4338 6322 -4304
rect 6256 -4354 6322 -4338
rect 6374 -4304 6440 -4288
rect 6374 -4338 6390 -4304
rect 6424 -4338 6440 -4304
rect 6374 -4354 6440 -4338
rect 6492 -4304 6558 -4288
rect 6492 -4338 6508 -4304
rect 6542 -4338 6558 -4304
rect 6492 -4354 6558 -4338
rect 5905 -4376 5965 -4354
rect 6023 -4376 6083 -4354
rect 6141 -4376 6201 -4354
rect 6259 -4376 6319 -4354
rect 6377 -4376 6437 -4354
rect 6495 -4376 6555 -4354
rect 5905 -6398 5965 -6376
rect 6023 -6398 6083 -6376
rect 6141 -6398 6201 -6376
rect 6259 -6398 6319 -6376
rect 6377 -6398 6437 -6376
rect 6495 -6398 6555 -6376
rect 5902 -6414 5968 -6398
rect 5902 -6448 5918 -6414
rect 5952 -6448 5968 -6414
rect 5902 -6464 5968 -6448
rect 6020 -6414 6086 -6398
rect 6020 -6448 6036 -6414
rect 6070 -6448 6086 -6414
rect 6020 -6464 6086 -6448
rect 6138 -6414 6204 -6398
rect 6138 -6448 6154 -6414
rect 6188 -6448 6204 -6414
rect 6138 -6464 6204 -6448
rect 6256 -6414 6322 -6398
rect 6256 -6448 6272 -6414
rect 6306 -6448 6322 -6414
rect 6256 -6464 6322 -6448
rect 6374 -6414 6440 -6398
rect 6374 -6448 6390 -6414
rect 6424 -6448 6440 -6414
rect 6374 -6464 6440 -6448
rect 6492 -6414 6558 -6398
rect 6492 -6448 6508 -6414
rect 6542 -6448 6558 -6414
rect 6492 -6464 6558 -6448
rect 7113 -3188 7513 -3172
rect 7113 -3222 7129 -3188
rect 7497 -3222 7513 -3188
rect 7113 -3260 7513 -3222
rect 7571 -3188 7971 -3172
rect 7571 -3222 7587 -3188
rect 7955 -3222 7971 -3188
rect 7571 -3260 7971 -3222
rect 8029 -3188 8429 -3172
rect 8029 -3222 8045 -3188
rect 8413 -3222 8429 -3188
rect 8029 -3260 8429 -3222
rect 8487 -3188 8887 -3172
rect 8487 -3222 8503 -3188
rect 8871 -3222 8887 -3188
rect 8487 -3260 8887 -3222
rect 7113 -5298 7513 -5260
rect 7113 -5332 7129 -5298
rect 7497 -5332 7513 -5298
rect 7113 -5348 7513 -5332
rect 7571 -5298 7971 -5260
rect 7571 -5332 7587 -5298
rect 7955 -5332 7971 -5298
rect 7571 -5348 7971 -5332
rect 8029 -5298 8429 -5260
rect 8029 -5332 8045 -5298
rect 8413 -5332 8429 -5298
rect 8029 -5348 8429 -5332
rect 8487 -5298 8887 -5260
rect 8487 -5332 8503 -5298
rect 8871 -5332 8887 -5298
rect 8487 -5348 8887 -5332
rect 10826 -3564 10852 -3534
rect 11352 -3564 11440 -3534
rect 11374 -3610 11440 -3564
rect 11374 -3630 11390 -3610
rect 10826 -3660 10852 -3630
rect 11352 -3644 11390 -3630
rect 11424 -3644 11440 -3610
rect 11352 -3660 11440 -3644
rect 10826 -3756 10852 -3726
rect 11352 -3756 11440 -3726
rect 11374 -3802 11440 -3756
rect 11374 -3822 11390 -3802
rect 10826 -3852 10852 -3822
rect 11352 -3836 11390 -3822
rect 11424 -3836 11440 -3802
rect 11352 -3852 11440 -3836
rect 7265 -5616 7391 -5600
rect 7265 -5650 7311 -5616
rect 7345 -5650 7391 -5616
rect 7073 -5700 7103 -5674
rect 7169 -5700 7199 -5674
rect 7265 -5678 7391 -5650
rect 7265 -5700 7295 -5678
rect 7361 -5700 7391 -5678
rect 7457 -5616 7583 -5600
rect 7457 -5650 7503 -5616
rect 7537 -5650 7583 -5616
rect 7457 -5678 7583 -5650
rect 7457 -5700 7487 -5678
rect 7553 -5700 7583 -5678
rect 7649 -5616 7775 -5600
rect 7649 -5650 7695 -5616
rect 7729 -5650 7775 -5616
rect 7649 -5678 7775 -5650
rect 7649 -5700 7679 -5678
rect 7745 -5700 7775 -5678
rect 7841 -5616 7967 -5600
rect 7841 -5650 7887 -5616
rect 7921 -5650 7967 -5616
rect 7841 -5678 7967 -5650
rect 7841 -5700 7871 -5678
rect 7937 -5700 7967 -5678
rect 8033 -5616 8159 -5600
rect 8033 -5650 8079 -5616
rect 8113 -5650 8159 -5616
rect 8033 -5678 8159 -5650
rect 8033 -5700 8063 -5678
rect 8129 -5700 8159 -5678
rect 8225 -5616 8351 -5600
rect 8225 -5650 8271 -5616
rect 8305 -5650 8351 -5616
rect 8225 -5678 8351 -5650
rect 8225 -5700 8255 -5678
rect 8321 -5700 8351 -5678
rect 8417 -5616 8543 -5600
rect 8417 -5650 8463 -5616
rect 8497 -5650 8543 -5616
rect 8417 -5678 8543 -5650
rect 8417 -5700 8447 -5678
rect 8513 -5700 8543 -5678
rect 8609 -5616 8735 -5600
rect 8609 -5650 8655 -5616
rect 8689 -5650 8735 -5616
rect 8609 -5678 8735 -5650
rect 8609 -5700 8639 -5678
rect 8705 -5700 8735 -5678
rect 8801 -5700 8831 -5674
rect 8897 -5700 8927 -5674
rect 7073 -6226 7103 -6200
rect 7169 -6226 7199 -6200
rect 7265 -6226 7295 -6200
rect 7361 -6226 7391 -6200
rect 7457 -6226 7487 -6200
rect 7553 -6226 7583 -6200
rect 7649 -6226 7679 -6200
rect 7745 -6226 7775 -6200
rect 7841 -6226 7871 -6200
rect 7937 -6226 7967 -6200
rect 8033 -6226 8063 -6200
rect 8129 -6226 8159 -6200
rect 8225 -6226 8255 -6200
rect 8321 -6226 8351 -6200
rect 8417 -6226 8447 -6200
rect 8513 -6226 8543 -6200
rect 8609 -6226 8639 -6200
rect 8705 -6226 8735 -6200
rect 8801 -6226 8831 -6200
rect 8897 -6226 8927 -6200
rect 7073 -6242 7199 -6226
rect 7073 -6276 7119 -6242
rect 7153 -6276 7199 -6242
rect 7073 -6304 7199 -6276
rect 8801 -6242 8927 -6226
rect 8801 -6276 8847 -6242
rect 8881 -6276 8927 -6242
rect 8801 -6304 8927 -6276
rect 9443 -4304 9509 -4288
rect 9443 -4338 9459 -4304
rect 9493 -4338 9509 -4304
rect 9443 -4354 9509 -4338
rect 9561 -4304 9627 -4288
rect 9561 -4338 9577 -4304
rect 9611 -4338 9627 -4304
rect 9561 -4354 9627 -4338
rect 9679 -4304 9745 -4288
rect 9679 -4338 9695 -4304
rect 9729 -4338 9745 -4304
rect 9679 -4354 9745 -4338
rect 9797 -4304 9863 -4288
rect 9797 -4338 9813 -4304
rect 9847 -4338 9863 -4304
rect 9797 -4354 9863 -4338
rect 9915 -4304 9981 -4288
rect 9915 -4338 9931 -4304
rect 9965 -4338 9981 -4304
rect 9915 -4354 9981 -4338
rect 10033 -4304 10099 -4288
rect 10033 -4338 10049 -4304
rect 10083 -4338 10099 -4304
rect 10033 -4354 10099 -4338
rect 9446 -4376 9506 -4354
rect 9564 -4376 9624 -4354
rect 9682 -4376 9742 -4354
rect 9800 -4376 9860 -4354
rect 9918 -4376 9978 -4354
rect 10036 -4376 10096 -4354
rect 9446 -6398 9506 -6376
rect 9564 -6398 9624 -6376
rect 9682 -6398 9742 -6376
rect 9800 -6398 9860 -6376
rect 9918 -6398 9978 -6376
rect 10036 -6398 10096 -6376
rect 9443 -6414 9509 -6398
rect 9443 -6448 9459 -6414
rect 9493 -6448 9509 -6414
rect 9443 -6464 9509 -6448
rect 9561 -6414 9627 -6398
rect 9561 -6448 9577 -6414
rect 9611 -6448 9627 -6414
rect 9561 -6464 9627 -6448
rect 9679 -6414 9745 -6398
rect 9679 -6448 9695 -6414
rect 9729 -6448 9745 -6414
rect 9679 -6464 9745 -6448
rect 9797 -6414 9863 -6398
rect 9797 -6448 9813 -6414
rect 9847 -6448 9863 -6414
rect 9797 -6464 9863 -6448
rect 9915 -6414 9981 -6398
rect 9915 -6448 9931 -6414
rect 9965 -6448 9981 -6414
rect 9915 -6464 9981 -6448
rect 10033 -6414 10099 -6398
rect 10033 -6448 10049 -6414
rect 10083 -6448 10099 -6414
rect 10033 -6464 10099 -6448
rect 6138 -6804 6204 -6788
rect 6138 -6838 6154 -6804
rect 6188 -6838 6204 -6804
rect 6138 -6854 6204 -6838
rect 6256 -6804 6322 -6788
rect 6256 -6838 6272 -6804
rect 6306 -6838 6322 -6804
rect 6256 -6854 6322 -6838
rect 6374 -6804 6440 -6788
rect 6374 -6838 6390 -6804
rect 6424 -6838 6440 -6804
rect 6374 -6854 6440 -6838
rect 6492 -6804 6558 -6788
rect 6492 -6838 6508 -6804
rect 6542 -6838 6558 -6804
rect 6492 -6854 6558 -6838
rect 6610 -6804 6676 -6788
rect 6610 -6838 6626 -6804
rect 6660 -6838 6676 -6804
rect 6610 -6854 6676 -6838
rect 6728 -6804 6794 -6788
rect 6728 -6838 6744 -6804
rect 6778 -6838 6794 -6804
rect 6728 -6854 6794 -6838
rect 6846 -6804 6912 -6788
rect 6846 -6838 6862 -6804
rect 6896 -6838 6912 -6804
rect 6846 -6854 6912 -6838
rect 6964 -6804 7030 -6788
rect 6964 -6838 6980 -6804
rect 7014 -6838 7030 -6804
rect 6964 -6854 7030 -6838
rect 7082 -6804 7148 -6788
rect 7082 -6838 7098 -6804
rect 7132 -6838 7148 -6804
rect 7082 -6854 7148 -6838
rect 7200 -6804 7266 -6788
rect 7200 -6838 7216 -6804
rect 7250 -6838 7266 -6804
rect 7200 -6854 7266 -6838
rect 7318 -6804 7384 -6788
rect 7318 -6838 7334 -6804
rect 7368 -6838 7384 -6804
rect 7318 -6854 7384 -6838
rect 7436 -6804 7502 -6788
rect 7436 -6838 7452 -6804
rect 7486 -6838 7502 -6804
rect 7436 -6854 7502 -6838
rect 7554 -6804 7620 -6788
rect 7554 -6838 7570 -6804
rect 7604 -6838 7620 -6804
rect 7554 -6854 7620 -6838
rect 7672 -6804 7738 -6788
rect 7672 -6838 7688 -6804
rect 7722 -6838 7738 -6804
rect 7672 -6854 7738 -6838
rect 7790 -6804 7856 -6788
rect 7790 -6838 7806 -6804
rect 7840 -6838 7856 -6804
rect 7790 -6854 7856 -6838
rect 7908 -6804 7974 -6788
rect 7908 -6838 7924 -6804
rect 7958 -6838 7974 -6804
rect 7908 -6854 7974 -6838
rect 8026 -6804 8092 -6788
rect 8026 -6838 8042 -6804
rect 8076 -6838 8092 -6804
rect 8026 -6854 8092 -6838
rect 8144 -6804 8210 -6788
rect 8144 -6838 8160 -6804
rect 8194 -6838 8210 -6804
rect 8144 -6854 8210 -6838
rect 8262 -6804 8328 -6788
rect 8262 -6838 8278 -6804
rect 8312 -6838 8328 -6804
rect 8262 -6854 8328 -6838
rect 8380 -6804 8446 -6788
rect 8380 -6838 8396 -6804
rect 8430 -6838 8446 -6804
rect 8380 -6854 8446 -6838
rect 8498 -6804 8564 -6788
rect 8498 -6838 8514 -6804
rect 8548 -6838 8564 -6804
rect 8498 -6854 8564 -6838
rect 8616 -6804 8682 -6788
rect 8616 -6838 8632 -6804
rect 8666 -6838 8682 -6804
rect 8616 -6854 8682 -6838
rect 8734 -6804 8800 -6788
rect 8734 -6838 8750 -6804
rect 8784 -6838 8800 -6804
rect 8734 -6854 8800 -6838
rect 8852 -6804 8918 -6788
rect 8852 -6838 8868 -6804
rect 8902 -6838 8918 -6804
rect 8852 -6854 8918 -6838
rect 8970 -6804 9036 -6788
rect 8970 -6838 8986 -6804
rect 9020 -6838 9036 -6804
rect 8970 -6854 9036 -6838
rect 9088 -6804 9154 -6788
rect 9088 -6838 9104 -6804
rect 9138 -6838 9154 -6804
rect 9088 -6854 9154 -6838
rect 9206 -6804 9272 -6788
rect 9206 -6838 9222 -6804
rect 9256 -6838 9272 -6804
rect 9206 -6854 9272 -6838
rect 9324 -6804 9390 -6788
rect 9324 -6838 9340 -6804
rect 9374 -6838 9390 -6804
rect 9324 -6854 9390 -6838
rect 9442 -6804 9508 -6788
rect 9442 -6838 9458 -6804
rect 9492 -6838 9508 -6804
rect 9442 -6854 9508 -6838
rect 9560 -6804 9626 -6788
rect 9560 -6838 9576 -6804
rect 9610 -6838 9626 -6804
rect 9560 -6854 9626 -6838
rect 9678 -6804 9744 -6788
rect 9678 -6838 9694 -6804
rect 9728 -6838 9744 -6804
rect 9678 -6854 9744 -6838
rect 9796 -6804 9862 -6788
rect 9796 -6838 9812 -6804
rect 9846 -6838 9862 -6804
rect 9796 -6854 9862 -6838
rect 6141 -6885 6201 -6854
rect 6259 -6885 6319 -6854
rect 6377 -6885 6437 -6854
rect 6495 -6885 6555 -6854
rect 6613 -6885 6673 -6854
rect 6731 -6885 6791 -6854
rect 6849 -6885 6909 -6854
rect 6967 -6885 7027 -6854
rect 7085 -6885 7145 -6854
rect 7203 -6885 7263 -6854
rect 7321 -6885 7381 -6854
rect 7439 -6885 7499 -6854
rect 7557 -6885 7617 -6854
rect 7675 -6885 7735 -6854
rect 7793 -6885 7853 -6854
rect 7911 -6885 7971 -6854
rect 8029 -6885 8089 -6854
rect 8147 -6885 8207 -6854
rect 8265 -6885 8325 -6854
rect 8383 -6885 8443 -6854
rect 8501 -6885 8561 -6854
rect 8619 -6885 8679 -6854
rect 8737 -6885 8797 -6854
rect 8855 -6885 8915 -6854
rect 8973 -6885 9033 -6854
rect 9091 -6885 9151 -6854
rect 9209 -6885 9269 -6854
rect 9327 -6885 9387 -6854
rect 9445 -6885 9505 -6854
rect 9563 -6885 9623 -6854
rect 9681 -6885 9741 -6854
rect 9799 -6885 9859 -6854
rect 6141 -8916 6201 -8885
rect 6259 -8916 6319 -8885
rect 6377 -8916 6437 -8885
rect 6495 -8916 6555 -8885
rect 6613 -8916 6673 -8885
rect 6731 -8916 6791 -8885
rect 6849 -8916 6909 -8885
rect 6967 -8916 7027 -8885
rect 7085 -8916 7145 -8885
rect 7203 -8916 7263 -8885
rect 7321 -8916 7381 -8885
rect 7439 -8916 7499 -8885
rect 7557 -8916 7617 -8885
rect 7675 -8916 7735 -8885
rect 7793 -8916 7853 -8885
rect 7911 -8916 7971 -8885
rect 8029 -8916 8089 -8885
rect 8147 -8916 8207 -8885
rect 8265 -8916 8325 -8885
rect 8383 -8916 8443 -8885
rect 8501 -8916 8561 -8885
rect 8619 -8916 8679 -8885
rect 8737 -8916 8797 -8885
rect 8855 -8916 8915 -8885
rect 8973 -8916 9033 -8885
rect 9091 -8916 9151 -8885
rect 9209 -8916 9269 -8885
rect 9327 -8916 9387 -8885
rect 9445 -8916 9505 -8885
rect 9563 -8916 9623 -8885
rect 9681 -8916 9741 -8885
rect 9799 -8916 9859 -8885
rect 6138 -8932 6204 -8916
rect 6138 -8966 6154 -8932
rect 6188 -8966 6204 -8932
rect 6138 -8982 6204 -8966
rect 6256 -8932 6322 -8916
rect 6256 -8966 6272 -8932
rect 6306 -8966 6322 -8932
rect 6256 -8982 6322 -8966
rect 6374 -8932 6440 -8916
rect 6374 -8966 6390 -8932
rect 6424 -8966 6440 -8932
rect 6374 -8982 6440 -8966
rect 6492 -8932 6558 -8916
rect 6492 -8966 6508 -8932
rect 6542 -8966 6558 -8932
rect 6492 -8982 6558 -8966
rect 6610 -8932 6676 -8916
rect 6610 -8966 6626 -8932
rect 6660 -8966 6676 -8932
rect 6610 -8982 6676 -8966
rect 6728 -8932 6794 -8916
rect 6728 -8966 6744 -8932
rect 6778 -8966 6794 -8932
rect 6728 -8982 6794 -8966
rect 6846 -8932 6912 -8916
rect 6846 -8966 6862 -8932
rect 6896 -8966 6912 -8932
rect 6846 -8982 6912 -8966
rect 6964 -8932 7030 -8916
rect 6964 -8966 6980 -8932
rect 7014 -8966 7030 -8932
rect 6964 -8982 7030 -8966
rect 7082 -8932 7148 -8916
rect 7082 -8966 7098 -8932
rect 7132 -8966 7148 -8932
rect 7082 -8982 7148 -8966
rect 7200 -8932 7266 -8916
rect 7200 -8966 7216 -8932
rect 7250 -8966 7266 -8932
rect 7200 -8982 7266 -8966
rect 7318 -8932 7384 -8916
rect 7318 -8966 7334 -8932
rect 7368 -8966 7384 -8932
rect 7318 -8982 7384 -8966
rect 7436 -8932 7502 -8916
rect 7436 -8966 7452 -8932
rect 7486 -8966 7502 -8932
rect 7436 -8982 7502 -8966
rect 7554 -8982 7620 -8916
rect 7672 -8982 7738 -8916
rect 7790 -8982 7856 -8916
rect 7908 -8982 7974 -8916
rect 8026 -8982 8092 -8916
rect 8144 -8982 8210 -8916
rect 8262 -8982 8328 -8916
rect 8380 -8982 8446 -8916
rect 8498 -8932 8564 -8916
rect 8498 -8966 8514 -8932
rect 8548 -8966 8564 -8932
rect 8498 -8982 8564 -8966
rect 8616 -8932 8682 -8916
rect 8616 -8966 8632 -8932
rect 8666 -8966 8682 -8932
rect 8616 -8982 8682 -8966
rect 8734 -8932 8800 -8916
rect 8734 -8966 8750 -8932
rect 8784 -8966 8800 -8932
rect 8734 -8982 8800 -8966
rect 8852 -8932 8918 -8916
rect 8852 -8966 8868 -8932
rect 8902 -8966 8918 -8932
rect 8852 -8982 8918 -8966
rect 8970 -8932 9036 -8916
rect 8970 -8966 8986 -8932
rect 9020 -8966 9036 -8932
rect 8970 -8982 9036 -8966
rect 9088 -8932 9154 -8916
rect 9088 -8966 9104 -8932
rect 9138 -8966 9154 -8932
rect 9088 -8982 9154 -8966
rect 9206 -8932 9272 -8916
rect 9206 -8966 9222 -8932
rect 9256 -8966 9272 -8932
rect 9206 -8982 9272 -8966
rect 9324 -8932 9390 -8916
rect 9324 -8966 9340 -8932
rect 9374 -8966 9390 -8932
rect 9324 -8982 9390 -8966
rect 9442 -8932 9508 -8916
rect 9442 -8966 9458 -8932
rect 9492 -8966 9508 -8932
rect 9442 -8982 9508 -8966
rect 9560 -8932 9626 -8916
rect 9560 -8966 9576 -8932
rect 9610 -8966 9626 -8932
rect 9560 -8982 9626 -8966
rect 9678 -8932 9744 -8916
rect 9678 -8966 9694 -8932
rect 9728 -8966 9744 -8932
rect 9678 -8982 9744 -8966
rect 9796 -8932 9862 -8916
rect 9796 -8966 9812 -8932
rect 9846 -8966 9862 -8932
rect 9796 -8982 9862 -8966
<< polycont >>
rect 6154 12332 6188 12366
rect 6272 12332 6306 12366
rect 6390 12332 6424 12366
rect 6508 12332 6542 12366
rect 6626 12332 6660 12366
rect 6744 12332 6778 12366
rect 6862 12332 6896 12366
rect 6980 12332 7014 12366
rect 7098 12332 7132 12366
rect 7216 12332 7250 12366
rect 7334 12332 7368 12366
rect 7452 12332 7486 12366
rect 8514 12332 8548 12366
rect 8632 12332 8666 12366
rect 8750 12332 8784 12366
rect 8868 12332 8902 12366
rect 8986 12332 9020 12366
rect 9104 12332 9138 12366
rect 9222 12332 9256 12366
rect 9340 12332 9374 12366
rect 9458 12332 9492 12366
rect 9576 12332 9610 12366
rect 9694 12332 9728 12366
rect 9812 12332 9846 12366
rect 6154 10204 6188 10238
rect 6272 10204 6306 10238
rect 6390 10204 6424 10238
rect 6508 10204 6542 10238
rect 6626 10204 6660 10238
rect 6744 10204 6778 10238
rect 6862 10204 6896 10238
rect 6980 10204 7014 10238
rect 7098 10204 7132 10238
rect 7216 10204 7250 10238
rect 7334 10204 7368 10238
rect 7452 10204 7486 10238
rect 7570 10204 7604 10238
rect 7688 10204 7722 10238
rect 7806 10204 7840 10238
rect 7924 10204 7958 10238
rect 8042 10204 8076 10238
rect 8160 10204 8194 10238
rect 8278 10204 8312 10238
rect 8396 10204 8430 10238
rect 8514 10204 8548 10238
rect 8632 10204 8666 10238
rect 8750 10204 8784 10238
rect 8868 10204 8902 10238
rect 8986 10204 9020 10238
rect 9104 10204 9138 10238
rect 9222 10204 9256 10238
rect 9340 10204 9374 10238
rect 9458 10204 9492 10238
rect 9576 10204 9610 10238
rect 9694 10204 9728 10238
rect 9812 10204 9846 10238
rect 5918 9814 5952 9848
rect 6036 9814 6070 9848
rect 6154 9814 6188 9848
rect 6272 9814 6306 9848
rect 6390 9814 6424 9848
rect 6508 9814 6542 9848
rect 5918 7704 5952 7738
rect 6036 7704 6070 7738
rect 6154 7704 6188 7738
rect 6272 7704 6306 7738
rect 6390 7704 6424 7738
rect 6508 7704 6542 7738
rect 7119 9642 7153 9676
rect 8847 9642 8881 9676
rect 7311 9016 7345 9050
rect 7503 9016 7537 9050
rect 7695 9016 7729 9050
rect 7887 9016 7921 9050
rect 8079 9016 8113 9050
rect 8271 9016 8305 9050
rect 8463 9016 8497 9050
rect 8655 9016 8689 9050
rect 7129 8698 7497 8732
rect 7587 8698 7955 8732
rect 8045 8698 8413 8732
rect 8503 8698 8871 8732
rect 7129 6588 7497 6622
rect 7587 6588 7955 6622
rect 8045 6588 8413 6622
rect 8503 6588 8871 6622
rect 9459 9814 9493 9848
rect 9577 9814 9611 9848
rect 9695 9814 9729 9848
rect 9813 9814 9847 9848
rect 9931 9814 9965 9848
rect 10049 9814 10083 9848
rect 9459 7704 9493 7738
rect 9577 7704 9611 7738
rect 9695 7704 9729 7738
rect 9813 7704 9847 7738
rect 9931 7704 9965 7738
rect 10049 7704 10083 7738
rect 11390 7202 11424 7236
rect 11390 7010 11424 7044
rect 3513 3880 3547 3914
rect 3513 3166 3547 3200
rect 4295 3880 4329 3914
rect 4295 3166 4329 3200
rect 2372 2488 2406 2522
rect 2440 2488 2474 2522
rect 3804 2472 3838 2506
rect 3984 2472 4018 2506
rect 4153 2479 4187 2513
rect 4300 2478 4334 2512
rect 4421 2478 4455 2512
rect 4542 2479 4576 2513
rect 5497 2479 5531 2513
rect 5644 2478 5678 2512
rect 5765 2478 5799 2512
rect 5886 2479 5920 2513
rect 6169 2479 6203 2513
rect 6316 2478 6350 2512
rect 6437 2478 6471 2512
rect 6558 2479 6592 2513
rect 6841 2479 6875 2513
rect 6988 2478 7022 2512
rect 7109 2478 7143 2512
rect 7230 2479 7264 2513
rect 8185 2479 8219 2513
rect 8332 2478 8366 2512
rect 8453 2478 8487 2512
rect 8574 2479 8608 2513
rect 8857 2479 8891 2513
rect 9004 2478 9038 2512
rect 9125 2478 9159 2512
rect 9246 2479 9280 2513
rect 9529 2479 9563 2513
rect 9676 2478 9710 2512
rect 2372 1902 2406 1936
rect 2440 1902 2474 1936
rect 3804 1918 3838 1952
rect 3984 1918 4018 1952
rect 4172 1892 4206 1926
rect 4340 1918 4374 1952
rect 4448 1918 4482 1952
rect 4562 1918 4596 1952
rect 4676 1898 4710 1932
rect 4784 1902 4818 1936
rect 4956 1902 4990 1936
rect 5459 1937 5493 1971
rect 5459 1869 5493 1903
rect 5576 1937 5610 1971
rect 5576 1869 5610 1903
rect 5712 1870 5746 1904
rect 5936 1866 5970 1900
rect 5459 1801 5493 1835
rect 6128 1892 6162 1926
rect 6238 1894 6272 1928
rect 6534 1860 6568 1894
rect 6422 1796 6456 1830
rect 6714 1857 6748 1891
rect 6822 1905 6856 1939
rect 6822 1837 6856 1871
rect 7058 1905 7092 1939
rect 7058 1837 7092 1871
rect 7173 1872 7207 1906
rect 7338 1846 7372 1880
rect 7446 1877 7480 1911
rect 7626 1909 7660 1943
rect 7806 1918 7840 1952
rect 7914 1918 7948 1952
rect 8022 1868 8056 1902
rect 8204 1861 8238 1895
rect 8312 1876 8346 1910
rect 8822 1918 8856 1952
rect 7631 1752 7665 1786
rect 9357 1892 9391 1926
rect 9425 1892 9459 1926
rect 9493 1892 9527 1926
rect 9561 1892 9595 1926
rect 9744 1892 9778 1926
rect 9812 1892 9846 1926
rect 9880 1892 9914 1926
rect 9948 1892 9982 1926
rect 11436 3784 11804 3818
rect 11894 3784 12262 3818
rect 12352 3784 12720 3818
rect 12810 3784 13178 3818
rect 13268 3784 13636 3818
rect 11436 1656 11804 1690
rect 11894 1656 12262 1690
rect 12352 1656 12720 1690
rect 12810 1656 13178 1690
rect 13268 1656 13636 1690
rect 13936 1656 13970 1690
rect 14252 1656 14286 1690
rect 3524 1156 3558 1190
rect 3592 1156 3626 1190
rect 5459 1257 5493 1291
rect 4956 1140 4990 1174
rect 5136 1140 5170 1174
rect 5459 1189 5493 1223
rect 5459 1121 5493 1155
rect 5576 1189 5610 1223
rect 5712 1188 5746 1222
rect 5576 1121 5610 1155
rect 5936 1192 5970 1226
rect 6422 1262 6456 1296
rect 6128 1166 6162 1200
rect 6238 1164 6272 1198
rect 6534 1198 6568 1232
rect 6714 1201 6748 1235
rect 6822 1221 6856 1255
rect 6822 1153 6856 1187
rect 7058 1221 7092 1255
rect 7058 1153 7092 1187
rect 7173 1186 7207 1220
rect 7338 1212 7372 1246
rect 7631 1306 7665 1340
rect 7446 1181 7480 1215
rect 7626 1149 7660 1183
rect 8022 1190 8056 1224
rect 7806 1140 7840 1174
rect 8204 1197 8238 1231
rect 7914 1140 7948 1174
rect 8312 1182 8346 1216
rect 8822 1140 8856 1174
rect 9468 1186 9502 1220
rect 9602 1165 9636 1199
rect 9716 1165 9750 1199
rect 9784 1165 9818 1199
rect 9852 1165 9886 1199
rect 3862 110 3896 144
rect 10520 1346 10888 1380
rect 10978 1346 11346 1380
rect 11436 1346 11804 1380
rect 11894 1346 12262 1380
rect 12352 1346 12720 1380
rect 12810 1346 13178 1380
rect 13268 1346 13636 1380
rect 10520 236 10888 270
rect 10978 236 11346 270
rect 11436 236 11804 270
rect 11894 236 12262 270
rect 12352 236 12720 270
rect 12810 236 13178 270
rect 13268 236 13636 270
rect 13936 1346 13970 1380
rect 14252 1346 14286 1380
rect 15978 823 16012 857
rect 16692 823 16726 857
rect 17406 823 17440 857
rect 18120 823 18154 857
rect 18834 823 18868 857
rect 19548 823 19582 857
rect 20262 823 20296 857
rect 20976 823 21010 857
rect 21690 823 21724 857
rect 22404 823 22438 857
rect 23118 823 23152 857
rect 23832 823 23866 857
rect 24546 823 24580 857
rect 25260 823 25294 857
rect 25974 823 26008 857
rect 26688 823 26722 857
rect 27402 823 27436 857
rect 28116 823 28150 857
rect 28830 823 28864 857
rect 29544 823 29578 857
rect 30258 823 30292 857
rect 30972 823 31006 857
rect 31686 823 31720 857
rect 32400 823 32434 857
rect 33114 823 33148 857
rect 33828 823 33862 857
rect 34542 823 34576 857
rect 35256 823 35290 857
rect 35970 823 36004 857
rect 36684 823 36718 857
rect 37398 823 37432 857
rect 38112 823 38146 857
rect 38826 823 38860 857
rect 3862 -604 3896 -570
rect 15978 5 16012 39
rect 16692 5 16726 39
rect 17406 5 17440 39
rect 18120 5 18154 39
rect 18834 5 18868 39
rect 19548 5 19582 39
rect 20262 5 20296 39
rect 20976 5 21010 39
rect 21690 5 21724 39
rect 22404 5 22438 39
rect 23118 5 23152 39
rect 23832 5 23866 39
rect 24546 5 24580 39
rect 25260 5 25294 39
rect 25974 5 26008 39
rect 26688 5 26722 39
rect 27402 5 27436 39
rect 28116 5 28150 39
rect 28830 5 28864 39
rect 29544 5 29578 39
rect 30258 5 30292 39
rect 30972 5 31006 39
rect 31686 5 31720 39
rect 32400 5 32434 39
rect 33114 5 33148 39
rect 33828 5 33862 39
rect 34542 5 34576 39
rect 35256 5 35290 39
rect 35970 5 36004 39
rect 36684 5 36718 39
rect 37398 5 37432 39
rect 38112 5 38146 39
rect 38826 5 38860 39
rect 10543 -918 10577 -884
rect 5918 -4338 5952 -4304
rect 6036 -4338 6070 -4304
rect 6154 -4338 6188 -4304
rect 6272 -4338 6306 -4304
rect 6390 -4338 6424 -4304
rect 6508 -4338 6542 -4304
rect 5918 -6448 5952 -6414
rect 6036 -6448 6070 -6414
rect 6154 -6448 6188 -6414
rect 6272 -6448 6306 -6414
rect 6390 -6448 6424 -6414
rect 6508 -6448 6542 -6414
rect 7129 -3222 7497 -3188
rect 7587 -3222 7955 -3188
rect 8045 -3222 8413 -3188
rect 8503 -3222 8871 -3188
rect 7129 -5332 7497 -5298
rect 7587 -5332 7955 -5298
rect 8045 -5332 8413 -5298
rect 8503 -5332 8871 -5298
rect 11390 -3644 11424 -3610
rect 11390 -3836 11424 -3802
rect 7311 -5650 7345 -5616
rect 7503 -5650 7537 -5616
rect 7695 -5650 7729 -5616
rect 7887 -5650 7921 -5616
rect 8079 -5650 8113 -5616
rect 8271 -5650 8305 -5616
rect 8463 -5650 8497 -5616
rect 8655 -5650 8689 -5616
rect 7119 -6276 7153 -6242
rect 8847 -6276 8881 -6242
rect 9459 -4338 9493 -4304
rect 9577 -4338 9611 -4304
rect 9695 -4338 9729 -4304
rect 9813 -4338 9847 -4304
rect 9931 -4338 9965 -4304
rect 10049 -4338 10083 -4304
rect 9459 -6448 9493 -6414
rect 9577 -6448 9611 -6414
rect 9695 -6448 9729 -6414
rect 9813 -6448 9847 -6414
rect 9931 -6448 9965 -6414
rect 10049 -6448 10083 -6414
rect 6154 -6838 6188 -6804
rect 6272 -6838 6306 -6804
rect 6390 -6838 6424 -6804
rect 6508 -6838 6542 -6804
rect 6626 -6838 6660 -6804
rect 6744 -6838 6778 -6804
rect 6862 -6838 6896 -6804
rect 6980 -6838 7014 -6804
rect 7098 -6838 7132 -6804
rect 7216 -6838 7250 -6804
rect 7334 -6838 7368 -6804
rect 7452 -6838 7486 -6804
rect 7570 -6838 7604 -6804
rect 7688 -6838 7722 -6804
rect 7806 -6838 7840 -6804
rect 7924 -6838 7958 -6804
rect 8042 -6838 8076 -6804
rect 8160 -6838 8194 -6804
rect 8278 -6838 8312 -6804
rect 8396 -6838 8430 -6804
rect 8514 -6838 8548 -6804
rect 8632 -6838 8666 -6804
rect 8750 -6838 8784 -6804
rect 8868 -6838 8902 -6804
rect 8986 -6838 9020 -6804
rect 9104 -6838 9138 -6804
rect 9222 -6838 9256 -6804
rect 9340 -6838 9374 -6804
rect 9458 -6838 9492 -6804
rect 9576 -6838 9610 -6804
rect 9694 -6838 9728 -6804
rect 9812 -6838 9846 -6804
rect 6154 -8966 6188 -8932
rect 6272 -8966 6306 -8932
rect 6390 -8966 6424 -8932
rect 6508 -8966 6542 -8932
rect 6626 -8966 6660 -8932
rect 6744 -8966 6778 -8932
rect 6862 -8966 6896 -8932
rect 6980 -8966 7014 -8932
rect 7098 -8966 7132 -8932
rect 7216 -8966 7250 -8932
rect 7334 -8966 7368 -8932
rect 7452 -8966 7486 -8932
rect 8514 -8966 8548 -8932
rect 8632 -8966 8666 -8932
rect 8750 -8966 8784 -8932
rect 8868 -8966 8902 -8932
rect 8986 -8966 9020 -8932
rect 9104 -8966 9138 -8932
rect 9222 -8966 9256 -8932
rect 9340 -8966 9374 -8932
rect 9458 -8966 9492 -8932
rect 9576 -8966 9610 -8932
rect 9694 -8966 9728 -8932
rect 9812 -8966 9846 -8932
<< xpolycontact >>
rect 5172 9020 5310 9452
rect 5406 9020 5544 9452
rect 10964 6696 11396 6766
rect 10964 6530 11396 6600
rect 2691 2347 3123 2629
rect 3223 2347 3655 2629
rect 2691 1795 3123 2077
rect 3223 1795 3655 2077
rect 10822 1684 10892 2116
rect 10988 1684 11058 2116
rect 3843 1015 4275 1297
rect 4375 1015 4807 1297
rect 39363 975 39795 1045
rect 39895 975 40327 1045
rect 39363 809 39795 879
rect 39895 809 40327 879
rect 39363 643 39795 713
rect 39895 643 40327 713
rect 39363 477 39795 547
rect 39895 477 40327 547
rect 39363 311 39795 381
rect 39895 311 40327 381
rect 39363 145 39795 215
rect 39895 145 40327 215
rect 39363 -21 39795 49
rect 39895 -21 40327 49
rect 39363 -187 39795 -117
rect 39895 -187 40327 -117
rect 5172 -6052 5310 -5620
rect 5406 -6052 5544 -5620
rect 10964 -3200 11396 -3130
rect 10964 -3366 11396 -3296
<< ppolyres >>
rect 5172 8554 5310 9020
rect 5406 8554 5544 9020
rect 5172 8416 5544 8554
rect 5172 -5154 5544 -5016
rect 5172 -5620 5310 -5154
rect 5406 -5620 5544 -5154
<< xpolyres >>
rect 10828 6696 10964 6766
rect 10828 6600 10898 6696
rect 10828 6530 10964 6600
rect 3123 2347 3223 2629
rect 3123 1795 3223 2077
rect 10822 2550 11058 2620
rect 10822 2116 10892 2550
rect 10988 2116 11058 2550
rect 4275 1015 4375 1297
rect 39795 975 39895 1045
rect 39795 809 39895 879
rect 39795 643 39895 713
rect 39795 477 39895 547
rect 39795 311 39895 381
rect 39795 145 39895 215
rect 39795 -21 39895 49
rect 39795 -187 39895 -117
rect 10828 -3200 10964 -3130
rect 10828 -3296 10898 -3200
rect 10828 -3366 10964 -3296
<< pdiode >>
rect 1890 1393 2016 1411
rect 1890 1223 1899 1393
rect 2007 1223 2016 1393
rect 2258 1393 2384 1411
rect 1890 1203 2016 1223
rect 2258 1223 2267 1393
rect 2375 1223 2384 1393
rect 2626 1393 2752 1411
rect 2258 1203 2384 1223
rect 2626 1223 2635 1393
rect 2743 1223 2752 1393
rect 2626 1203 2752 1223
rect 10287 -486 10495 -477
rect 10287 -594 10305 -486
rect 10475 -594 10495 -486
rect 10287 -603 10495 -594
rect 10287 -1130 10495 -1121
rect 10287 -1238 10305 -1130
rect 10475 -1238 10495 -1130
rect 10287 -1247 10495 -1238
<< ndiode >>
rect 2162 2454 2300 2462
rect 2162 2420 2174 2454
rect 2208 2420 2254 2454
rect 2288 2420 2300 2454
rect 2162 2386 2300 2420
rect 2162 2352 2174 2386
rect 2208 2352 2254 2386
rect 2288 2352 2300 2386
rect 2162 2318 2300 2352
rect 2162 2284 2174 2318
rect 2208 2284 2254 2318
rect 2288 2284 2300 2318
rect 2162 2276 2300 2284
rect 2162 2140 2300 2148
rect 2162 2106 2174 2140
rect 2208 2106 2254 2140
rect 2288 2106 2300 2140
rect 2162 2072 2300 2106
rect 2162 2038 2174 2072
rect 2208 2038 2254 2072
rect 2288 2038 2300 2072
rect 2162 2004 2300 2038
rect 2162 1970 2174 2004
rect 2208 1970 2254 2004
rect 2288 1970 2300 2004
rect 2162 1962 2300 1970
rect 3314 1122 3452 1130
rect 1890 1065 2016 1083
rect 1890 963 1899 1065
rect 2008 963 2016 1065
rect 2258 1065 2384 1083
rect 1890 945 2016 963
rect 2258 963 2267 1065
rect 2376 963 2384 1065
rect 2626 1065 2752 1083
rect 2258 945 2384 963
rect 2626 963 2635 1065
rect 2744 963 2752 1065
rect 2626 945 2752 963
rect 3314 1088 3326 1122
rect 3360 1088 3406 1122
rect 3440 1088 3452 1122
rect 3314 1054 3452 1088
rect 3314 1020 3326 1054
rect 3360 1020 3406 1054
rect 3440 1020 3452 1054
rect 3314 986 3452 1020
rect 3314 952 3326 986
rect 3360 952 3406 986
rect 3440 952 3452 986
rect 3314 944 3452 952
rect 10615 -486 10753 -477
rect 10615 -595 10633 -486
rect 10735 -595 10753 -486
rect 10615 -603 10753 -595
rect 10615 -1130 10753 -1121
rect 10615 -1239 10633 -1130
rect 10735 -1239 10753 -1130
rect 10615 -1247 10753 -1239
<< pdiodec >>
rect 1899 1223 2007 1393
rect 2267 1223 2375 1393
rect 2635 1223 2743 1393
rect 10305 -594 10475 -486
rect 10305 -1238 10475 -1130
<< ndiodec >>
rect 2174 2420 2208 2454
rect 2254 2420 2288 2454
rect 2174 2352 2208 2386
rect 2254 2352 2288 2386
rect 2174 2284 2208 2318
rect 2254 2284 2288 2318
rect 2174 2106 2208 2140
rect 2254 2106 2288 2140
rect 2174 2038 2208 2072
rect 2254 2038 2288 2072
rect 2174 1970 2208 2004
rect 2254 1970 2288 2004
rect 1899 963 2008 1065
rect 2267 963 2376 1065
rect 2635 963 2744 1065
rect 3326 1088 3360 1122
rect 3406 1088 3440 1122
rect 3326 1020 3360 1054
rect 3406 1020 3440 1054
rect 3326 952 3360 986
rect 3406 952 3440 986
rect 10633 -595 10735 -486
rect 10633 -1239 10735 -1130
<< locali >>
rect 5981 12434 6077 12468
rect 9923 12434 10019 12468
rect 5981 12372 6015 12434
rect 9985 12372 10019 12434
rect 6138 12332 6154 12366
rect 6188 12332 6204 12366
rect 6256 12332 6272 12366
rect 6306 12332 6322 12366
rect 6374 12332 6390 12366
rect 6424 12332 6440 12366
rect 6492 12332 6508 12366
rect 6542 12332 6558 12366
rect 6610 12332 6626 12366
rect 6660 12332 6676 12366
rect 6728 12332 6744 12366
rect 6778 12332 6794 12366
rect 6846 12332 6862 12366
rect 6896 12332 6912 12366
rect 6964 12332 6980 12366
rect 7014 12332 7030 12366
rect 7082 12332 7098 12366
rect 7132 12332 7148 12366
rect 7200 12332 7216 12366
rect 7250 12332 7266 12366
rect 7318 12332 7334 12366
rect 7368 12332 7384 12366
rect 7436 12332 7452 12366
rect 7486 12332 7502 12366
rect 8498 12332 8514 12366
rect 8548 12332 8564 12366
rect 8616 12332 8632 12366
rect 8666 12332 8682 12366
rect 8734 12332 8750 12366
rect 8784 12332 8800 12366
rect 8852 12332 8868 12366
rect 8902 12332 8918 12366
rect 8970 12332 8986 12366
rect 9020 12332 9036 12366
rect 9088 12332 9104 12366
rect 9138 12332 9154 12366
rect 9206 12332 9222 12366
rect 9256 12332 9272 12366
rect 9324 12332 9340 12366
rect 9374 12332 9390 12366
rect 9442 12332 9458 12366
rect 9492 12332 9508 12366
rect 9560 12332 9576 12366
rect 9610 12332 9626 12366
rect 9678 12332 9694 12366
rect 9728 12332 9744 12366
rect 9796 12332 9812 12366
rect 9846 12332 9862 12366
rect 6095 12273 6129 12289
rect 6095 10281 6129 10297
rect 6213 12273 6247 12289
rect 6213 10281 6247 10297
rect 6331 12273 6365 12289
rect 6331 10281 6365 10297
rect 6449 12273 6483 12289
rect 6449 10281 6483 10297
rect 6567 12273 6601 12289
rect 6567 10281 6601 10297
rect 6685 12273 6719 12289
rect 6685 10281 6719 10297
rect 6803 12273 6837 12289
rect 6803 10281 6837 10297
rect 6921 12273 6955 12289
rect 6921 10281 6955 10297
rect 7039 12273 7073 12289
rect 7039 10281 7073 10297
rect 7157 12273 7191 12289
rect 7157 10281 7191 10297
rect 7275 12273 7309 12289
rect 7275 10281 7309 10297
rect 7393 12273 7427 12289
rect 7393 10281 7427 10297
rect 7511 12273 7545 12289
rect 7511 10281 7545 10297
rect 7629 12273 7663 12289
rect 7629 10281 7663 10297
rect 7747 12273 7781 12289
rect 7747 10281 7781 10297
rect 7865 12273 7899 12289
rect 7865 10281 7899 10297
rect 7983 12273 8017 12289
rect 7983 10281 8017 10297
rect 8101 12273 8135 12289
rect 8101 10281 8135 10297
rect 8219 12273 8253 12289
rect 8219 10281 8253 10297
rect 8337 12273 8371 12289
rect 8337 10281 8371 10297
rect 8455 12273 8489 12289
rect 8455 10281 8489 10297
rect 8573 12273 8607 12289
rect 8573 10281 8607 10297
rect 8691 12273 8725 12289
rect 8691 10281 8725 10297
rect 8809 12273 8843 12289
rect 8809 10281 8843 10297
rect 8927 12273 8961 12289
rect 8927 10281 8961 10297
rect 9045 12273 9079 12289
rect 9045 10281 9079 10297
rect 9163 12273 9197 12289
rect 9163 10281 9197 10297
rect 9281 12273 9315 12289
rect 9281 10281 9315 10297
rect 9399 12273 9433 12289
rect 9399 10281 9433 10297
rect 9517 12273 9551 12289
rect 9517 10281 9551 10297
rect 9635 12273 9669 12289
rect 9635 10281 9669 10297
rect 9753 12273 9787 12289
rect 9753 10281 9787 10297
rect 9871 12273 9905 12289
rect 9871 10281 9905 10297
rect 6138 10204 6154 10238
rect 6188 10204 6204 10238
rect 6256 10204 6272 10238
rect 6306 10204 6322 10238
rect 6374 10204 6390 10238
rect 6424 10204 6440 10238
rect 6492 10204 6508 10238
rect 6542 10204 6558 10238
rect 6610 10204 6626 10238
rect 6660 10204 6676 10238
rect 6728 10204 6744 10238
rect 6778 10204 6794 10238
rect 6846 10204 6862 10238
rect 6896 10204 6912 10238
rect 6964 10204 6980 10238
rect 7014 10204 7030 10238
rect 7082 10204 7098 10238
rect 7132 10204 7148 10238
rect 7200 10204 7216 10238
rect 7250 10204 7266 10238
rect 7318 10204 7334 10238
rect 7368 10204 7384 10238
rect 7436 10204 7452 10238
rect 7486 10204 7502 10238
rect 7554 10204 7570 10238
rect 7604 10204 7620 10238
rect 7672 10204 7688 10238
rect 7722 10204 7738 10238
rect 7790 10204 7806 10238
rect 7840 10204 7856 10238
rect 7908 10204 7924 10238
rect 7958 10204 7974 10238
rect 8026 10204 8042 10238
rect 8076 10204 8092 10238
rect 8144 10204 8160 10238
rect 8194 10204 8210 10238
rect 8262 10204 8278 10238
rect 8312 10204 8328 10238
rect 8380 10204 8396 10238
rect 8430 10204 8446 10238
rect 8498 10204 8514 10238
rect 8548 10204 8564 10238
rect 8616 10204 8632 10238
rect 8666 10204 8682 10238
rect 8734 10204 8750 10238
rect 8784 10204 8800 10238
rect 8852 10204 8868 10238
rect 8902 10204 8918 10238
rect 8970 10204 8986 10238
rect 9020 10204 9036 10238
rect 9088 10204 9104 10238
rect 9138 10204 9154 10238
rect 9206 10204 9222 10238
rect 9256 10204 9272 10238
rect 9324 10204 9340 10238
rect 9374 10204 9390 10238
rect 9442 10204 9458 10238
rect 9492 10204 9508 10238
rect 9560 10204 9576 10238
rect 9610 10204 9626 10238
rect 9678 10204 9694 10238
rect 9728 10204 9744 10238
rect 9796 10204 9812 10238
rect 9846 10204 9862 10238
rect 5981 10136 6015 10198
rect 9985 10136 10019 10198
rect 5981 10102 6077 10136
rect 9923 10102 10019 10136
rect 5745 9916 5841 9950
rect 6619 9916 6715 9950
rect 5745 9854 5779 9916
rect 6681 9854 6715 9916
rect 5902 9814 5918 9848
rect 5952 9814 5968 9848
rect 6020 9814 6036 9848
rect 6070 9814 6086 9848
rect 6138 9814 6154 9848
rect 6188 9814 6204 9848
rect 6256 9814 6272 9848
rect 6306 9814 6322 9848
rect 6374 9814 6390 9848
rect 6424 9814 6440 9848
rect 6492 9814 6508 9848
rect 6542 9814 6558 9848
rect 5042 9548 5138 9582
rect 5578 9560 5674 9582
rect 5578 9548 5745 9560
rect 5042 9486 5076 9548
rect 5640 9486 5745 9548
rect 5042 8320 5076 8382
rect 5674 8382 5745 9486
rect 5640 8320 5745 8382
rect 5042 8286 5138 8320
rect 5578 8286 5674 8320
rect 5859 9764 5893 9780
rect 5859 7772 5893 7788
rect 5977 9764 6011 9780
rect 5977 7772 6011 7788
rect 6095 9764 6129 9780
rect 6095 7772 6129 7788
rect 6213 9764 6247 9780
rect 6213 7772 6247 7788
rect 6331 9764 6365 9780
rect 6331 7772 6365 7788
rect 6449 9764 6483 9780
rect 6449 7772 6483 7788
rect 6567 9764 6601 9780
rect 6567 7772 6601 7788
rect 9286 9916 9382 9950
rect 10160 9916 10256 9950
rect 9286 9854 9320 9916
rect 10222 9854 10256 9916
rect 9443 9814 9459 9848
rect 9493 9814 9509 9848
rect 9561 9814 9577 9848
rect 9611 9814 9627 9848
rect 9679 9814 9695 9848
rect 9729 9814 9745 9848
rect 9797 9814 9813 9848
rect 9847 9814 9863 9848
rect 9915 9814 9931 9848
rect 9965 9814 9981 9848
rect 10033 9814 10049 9848
rect 10083 9814 10099 9848
rect 6909 9740 7005 9774
rect 8995 9740 9091 9774
rect 6909 9678 6943 9740
rect 9057 9678 9091 9740
rect 7103 9642 7119 9676
rect 7153 9642 7169 9676
rect 8831 9642 8847 9676
rect 8881 9642 8897 9676
rect 7023 9588 7057 9604
rect 7023 9096 7057 9112
rect 7119 9588 7153 9604
rect 7119 9096 7153 9112
rect 7215 9588 7249 9604
rect 7215 9096 7249 9112
rect 7311 9588 7345 9604
rect 7311 9096 7345 9112
rect 7407 9588 7441 9604
rect 7407 9096 7441 9112
rect 7503 9588 7537 9604
rect 7503 9096 7537 9112
rect 7599 9588 7633 9604
rect 7599 9096 7633 9112
rect 7695 9588 7729 9604
rect 7695 9096 7729 9112
rect 7791 9588 7825 9604
rect 7791 9096 7825 9112
rect 7887 9588 7921 9604
rect 7887 9096 7921 9112
rect 7983 9588 8017 9604
rect 7983 9096 8017 9112
rect 8079 9588 8113 9604
rect 8079 9096 8113 9112
rect 8175 9588 8209 9604
rect 8175 9096 8209 9112
rect 8271 9588 8305 9604
rect 8271 9096 8305 9112
rect 8367 9588 8401 9604
rect 8367 9096 8401 9112
rect 8463 9588 8497 9604
rect 8463 9096 8497 9112
rect 8559 9588 8593 9604
rect 8559 9096 8593 9112
rect 8655 9588 8689 9604
rect 8655 9096 8689 9112
rect 8751 9588 8785 9604
rect 8751 9096 8785 9112
rect 8847 9588 8881 9604
rect 8847 9096 8881 9112
rect 8943 9588 8977 9604
rect 8943 9096 8977 9112
rect 6909 8960 6943 9022
rect 7295 9016 7311 9050
rect 7345 9016 7361 9050
rect 7487 9016 7503 9050
rect 7537 9016 7553 9050
rect 7679 9016 7695 9050
rect 7729 9016 7745 9050
rect 7871 9016 7887 9050
rect 7921 9016 7937 9050
rect 8063 9016 8079 9050
rect 8113 9016 8129 9050
rect 8255 9016 8271 9050
rect 8305 9016 8321 9050
rect 8447 9016 8463 9050
rect 8497 9016 8513 9050
rect 8639 9016 8655 9050
rect 8689 9016 8705 9050
rect 9057 8960 9091 9022
rect 6909 8926 7005 8960
rect 8995 8926 9091 8960
rect 5902 7704 5918 7738
rect 5952 7704 5968 7738
rect 6020 7704 6036 7738
rect 6070 7704 6086 7738
rect 6138 7704 6154 7738
rect 6188 7704 6204 7738
rect 6256 7704 6272 7738
rect 6306 7704 6322 7738
rect 6374 7704 6390 7738
rect 6424 7704 6440 7738
rect 6492 7704 6508 7738
rect 6542 7704 6558 7738
rect 5745 7636 5779 7698
rect 6681 7636 6715 7698
rect 5745 7602 5841 7636
rect 6619 7602 6715 7636
rect 6953 8800 7049 8834
rect 8951 8800 9047 8834
rect 6953 8738 6987 8800
rect 9013 8738 9047 8800
rect 7113 8698 7129 8732
rect 7497 8698 7513 8732
rect 7571 8698 7587 8732
rect 7955 8698 7971 8732
rect 8029 8698 8045 8732
rect 8413 8698 8429 8732
rect 8487 8698 8503 8732
rect 8871 8698 8887 8732
rect 7067 8648 7101 8664
rect 7067 6656 7101 6672
rect 7525 8648 7559 8664
rect 7525 6656 7559 6672
rect 7983 8648 8017 8664
rect 7983 6656 8017 6672
rect 8441 8648 8475 8664
rect 8441 6656 8475 6672
rect 8899 8648 8933 8664
rect 8899 6656 8933 6672
rect 9400 9764 9434 9780
rect 9400 7772 9434 7788
rect 9518 9764 9552 9780
rect 9518 7772 9552 7788
rect 9636 9764 9670 9780
rect 9636 7772 9670 7788
rect 9754 9764 9788 9780
rect 9754 7772 9788 7788
rect 9872 9764 9906 9780
rect 9872 7772 9906 7788
rect 9990 9764 10024 9780
rect 9990 7772 10024 7788
rect 10108 9764 10142 9780
rect 10108 7772 10142 7788
rect 9443 7704 9459 7738
rect 9493 7704 9509 7738
rect 9561 7704 9577 7738
rect 9611 7704 9627 7738
rect 9679 7704 9695 7738
rect 9729 7704 9745 7738
rect 9797 7704 9813 7738
rect 9847 7704 9863 7738
rect 9915 7704 9931 7738
rect 9965 7704 9981 7738
rect 10033 7704 10049 7738
rect 10083 7704 10099 7738
rect 9286 7636 9320 7698
rect 10222 7636 10256 7698
rect 9286 7602 9382 7636
rect 10160 7602 10256 7636
rect 10644 7416 11560 7450
rect 10644 7382 10774 7416
rect 11430 7382 11560 7416
rect 10644 7320 10712 7382
rect 10644 7280 10678 7320
rect 7113 6588 7129 6622
rect 7497 6588 7513 6622
rect 7571 6588 7587 6622
rect 7955 6588 7971 6622
rect 8029 6588 8045 6622
rect 8413 6588 8429 6622
rect 8487 6588 8503 6622
rect 8871 6588 8887 6622
rect 6953 6520 6987 6582
rect 9013 6520 9047 6582
rect 6953 6486 7049 6520
rect 8951 6486 9047 6520
rect 10522 7260 10678 7280
rect 10522 6340 10542 7260
rect 10602 6470 10678 7260
rect 11492 7320 11560 7382
rect 10848 7268 10864 7302
rect 11340 7268 11356 7302
rect 11390 7236 11424 7252
rect 10848 7172 10864 7206
rect 11340 7172 11356 7206
rect 11390 7186 11424 7202
rect 10848 7076 10864 7110
rect 11340 7076 11356 7110
rect 11390 7044 11424 7060
rect 10712 6980 10864 7014
rect 11340 6980 11356 7014
rect 11390 6994 11424 7010
rect 10848 6884 10864 6918
rect 11340 6884 11435 6918
rect 11384 6766 11435 6884
rect 11396 6696 11435 6766
rect 11396 6592 11435 6600
rect 11412 6539 11435 6592
rect 11396 6530 11435 6539
rect 10602 6388 10712 6470
rect 11526 6470 11560 7320
rect 11492 6388 11560 6470
rect 10602 6354 10774 6388
rect 11430 6354 11560 6388
rect 10602 6340 11560 6354
rect 10522 6320 11560 6340
rect 3355 4492 3451 4526
rect 3609 4492 3739 4526
rect 3355 4430 3389 4492
rect 3671 4430 3739 4492
rect 3469 4340 3503 4356
rect 3469 3948 3503 3964
rect 3557 4340 3591 4356
rect 3557 3948 3591 3964
rect 3497 3880 3513 3914
rect 3547 3880 3563 3914
rect 3355 3812 3389 3874
rect 3705 3874 3739 4430
rect 3671 3812 3739 3874
rect 3355 3778 3451 3812
rect 3609 3778 3739 3812
rect 3355 3716 3389 3778
rect 3671 3716 3739 3778
rect 3469 3626 3503 3642
rect 3469 3234 3503 3250
rect 3557 3626 3591 3642
rect 3557 3234 3591 3250
rect 3497 3166 3513 3200
rect 3547 3166 3563 3200
rect 3355 3098 3389 3160
rect 3705 3160 3739 3716
rect 3671 3098 3739 3160
rect 3355 3064 3451 3098
rect 3609 3064 3739 3098
rect 4103 4492 4233 4526
rect 4391 4492 4487 4526
rect 4103 4430 4171 4492
rect 4103 3874 4137 4430
rect 4453 4430 4487 4492
rect 4251 4340 4285 4356
rect 4251 3948 4285 3964
rect 4339 4340 4373 4356
rect 4339 3948 4373 3964
rect 4279 3880 4295 3914
rect 4329 3880 4345 3914
rect 4103 3812 4171 3874
rect 11268 3978 14438 3988
rect 11268 3920 11278 3978
rect 14428 3920 14438 3978
rect 4453 3812 4487 3874
rect 4103 3778 4233 3812
rect 4391 3778 4487 3812
rect 4103 3716 4171 3778
rect 4103 3160 4137 3716
rect 4453 3716 4487 3778
rect 4251 3626 4285 3642
rect 4251 3234 4285 3250
rect 4339 3626 4373 3642
rect 4339 3234 4373 3250
rect 4279 3166 4295 3200
rect 4329 3166 4345 3200
rect 4103 3098 4171 3160
rect 4453 3098 4487 3160
rect 4103 3064 4233 3098
rect 4391 3064 4487 3098
rect 11260 3908 11278 3920
rect 14428 3908 14444 3920
rect 11260 3886 11356 3908
rect 13716 3886 13874 3908
rect 14032 3886 14190 3908
rect 14348 3886 14444 3908
rect 11260 3824 11294 3886
rect 2039 2861 2070 2895
rect 2104 2861 2166 2895
rect 2200 2861 2262 2895
rect 2296 2861 2358 2895
rect 2392 2861 2454 2895
rect 2488 2861 2550 2895
rect 2584 2861 2646 2895
rect 2680 2861 2742 2895
rect 2776 2861 2838 2895
rect 2872 2861 2934 2895
rect 2968 2861 3030 2895
rect 3064 2861 3126 2895
rect 3160 2861 3222 2895
rect 3256 2861 3318 2895
rect 3352 2861 3414 2895
rect 3448 2861 3510 2895
rect 3544 2861 3606 2895
rect 3640 2861 3702 2895
rect 3736 2861 3798 2895
rect 3832 2861 3894 2895
rect 3928 2861 3990 2895
rect 4024 2861 4086 2895
rect 4120 2861 4182 2895
rect 4216 2861 4278 2895
rect 4312 2861 4374 2895
rect 4408 2861 4470 2895
rect 4504 2861 4566 2895
rect 4600 2861 4662 2895
rect 4696 2861 4758 2895
rect 4792 2861 4854 2895
rect 4888 2861 4950 2895
rect 4984 2861 5046 2895
rect 5080 2861 5142 2895
rect 5176 2861 5238 2895
rect 5272 2861 5334 2895
rect 5368 2861 5430 2895
rect 5464 2861 5526 2895
rect 5560 2861 5622 2895
rect 5656 2861 5718 2895
rect 5752 2861 5814 2895
rect 5848 2861 5910 2895
rect 5944 2861 6006 2895
rect 6040 2861 6102 2895
rect 6136 2861 6198 2895
rect 6232 2861 6294 2895
rect 6328 2861 6390 2895
rect 6424 2861 6486 2895
rect 6520 2861 6582 2895
rect 6616 2861 6678 2895
rect 6712 2861 6774 2895
rect 6808 2861 6870 2895
rect 6904 2861 6966 2895
rect 7000 2861 7062 2895
rect 7096 2861 7158 2895
rect 7192 2861 7254 2895
rect 7288 2861 7350 2895
rect 7384 2861 7446 2895
rect 7480 2861 7542 2895
rect 7576 2861 7638 2895
rect 7672 2861 7734 2895
rect 7768 2861 7830 2895
rect 7864 2861 7926 2895
rect 7960 2861 8022 2895
rect 8056 2861 8118 2895
rect 8152 2861 8214 2895
rect 8248 2861 8310 2895
rect 8344 2861 8406 2895
rect 8440 2861 8502 2895
rect 8536 2861 8598 2895
rect 8632 2861 8694 2895
rect 8728 2861 8790 2895
rect 8824 2861 8886 2895
rect 8920 2861 8982 2895
rect 9016 2861 9078 2895
rect 9112 2861 9174 2895
rect 9208 2861 9270 2895
rect 9304 2861 9366 2895
rect 9400 2861 9462 2895
rect 9496 2861 9558 2895
rect 9592 2861 9654 2895
rect 9688 2861 9750 2895
rect 9784 2861 9846 2895
rect 9880 2861 9942 2895
rect 9976 2861 10038 2895
rect 10072 2861 10134 2895
rect 10168 2861 10199 2895
rect 2057 2790 2117 2861
rect 2057 2756 2070 2790
rect 2104 2756 2117 2790
rect 2057 2704 2117 2756
rect 2057 2670 2070 2704
rect 2104 2670 2117 2704
rect 2057 2653 2117 2670
rect 2154 2568 2308 2825
rect 2424 2792 2490 2861
rect 2424 2758 2440 2792
rect 2474 2758 2490 2792
rect 2424 2722 2490 2758
rect 2424 2688 2440 2722
rect 2474 2688 2490 2722
rect 2424 2652 2490 2688
rect 2424 2618 2440 2652
rect 2474 2618 2490 2652
rect 2424 2602 2490 2618
rect 2524 2792 2590 2808
rect 2524 2758 2540 2792
rect 2574 2758 2590 2792
rect 2524 2709 2590 2758
rect 2524 2675 2540 2709
rect 2574 2675 2590 2709
rect 2524 2626 2590 2675
rect 3788 2792 3854 2861
rect 3788 2758 3804 2792
rect 3838 2758 3854 2792
rect 3788 2709 3854 2758
rect 3788 2675 3804 2709
rect 3838 2675 3854 2709
rect 2524 2592 2540 2626
rect 2574 2592 2590 2626
rect 2154 2522 2490 2568
rect 2154 2488 2368 2522
rect 2406 2488 2440 2522
rect 2474 2488 2490 2522
rect 2154 2472 2490 2488
rect 2524 2539 2590 2592
rect 2524 2480 2691 2539
rect 2154 2454 2308 2472
rect 2057 2417 2117 2433
rect 2057 2383 2070 2417
rect 2104 2383 2117 2417
rect 2057 2334 2117 2383
rect 2057 2300 2070 2334
rect 2104 2300 2117 2334
rect 2057 2229 2117 2300
rect 2154 2420 2174 2454
rect 2208 2420 2254 2454
rect 2288 2420 2308 2454
rect 2154 2386 2308 2420
rect 2154 2352 2174 2386
rect 2208 2352 2254 2386
rect 2288 2352 2308 2386
rect 2154 2318 2308 2352
rect 2154 2284 2174 2318
rect 2208 2284 2254 2318
rect 2288 2284 2308 2318
rect 2154 2265 2308 2284
rect 2424 2422 2490 2438
rect 2424 2388 2440 2422
rect 2474 2388 2490 2422
rect 2424 2332 2490 2388
rect 2424 2298 2440 2332
rect 2474 2298 2490 2332
rect 2424 2229 2490 2298
rect 2524 2422 2590 2480
rect 2524 2388 2540 2422
rect 2574 2388 2590 2422
rect 2524 2332 2590 2388
rect 3788 2626 3854 2675
rect 3788 2592 3804 2626
rect 3838 2592 3854 2626
rect 3788 2576 3854 2592
rect 3888 2792 3934 2808
rect 3888 2758 3894 2792
rect 3928 2758 3934 2792
rect 3888 2709 3934 2758
rect 3888 2675 3894 2709
rect 3928 2675 3934 2709
rect 3888 2626 3934 2675
rect 3888 2592 3894 2626
rect 3928 2592 3934 2626
rect 3655 2506 3854 2522
rect 3655 2472 3804 2506
rect 3838 2472 3854 2506
rect 3655 2456 3854 2472
rect 3788 2448 3854 2456
rect 3888 2448 3934 2592
rect 3968 2792 4034 2861
rect 3968 2758 3984 2792
rect 4018 2758 4034 2792
rect 3968 2709 4034 2758
rect 3968 2675 3984 2709
rect 4018 2675 4034 2709
rect 3968 2626 4034 2675
rect 3968 2592 3984 2626
rect 4018 2592 4034 2626
rect 4074 2792 4140 2861
rect 4074 2758 4090 2792
rect 4124 2758 4140 2792
rect 4074 2721 4140 2758
rect 4074 2687 4090 2721
rect 4124 2687 4140 2721
rect 4074 2650 4140 2687
rect 4074 2616 4090 2650
rect 4124 2616 4140 2650
rect 4074 2598 4140 2616
rect 4284 2792 4471 2861
rect 4284 2758 4348 2792
rect 4382 2758 4471 2792
rect 4284 2721 4471 2758
rect 4284 2687 4348 2721
rect 4382 2687 4471 2721
rect 4284 2650 4471 2687
rect 4284 2616 4348 2650
rect 4382 2616 4471 2650
rect 3968 2576 4034 2592
rect 3968 2506 4034 2522
rect 3968 2472 3984 2506
rect 4018 2472 4034 2506
rect 3968 2448 4034 2472
rect 4089 2513 4203 2529
rect 4089 2479 4153 2513
rect 4187 2479 4203 2513
rect 3900 2414 3934 2448
rect 3793 2380 3809 2414
rect 3843 2380 3859 2414
rect 3900 2380 3973 2414
rect 4007 2380 4023 2414
rect 2524 2298 2540 2332
rect 2574 2298 2590 2332
rect 2524 2282 2590 2298
rect 3793 2332 3859 2380
rect 3793 2298 3809 2332
rect 3843 2298 3859 2332
rect 3793 2229 3859 2298
rect 3957 2338 4023 2380
rect 3957 2332 3974 2338
rect 3957 2298 3973 2332
rect 4008 2304 4023 2338
rect 4007 2298 4023 2304
rect 3957 2282 4023 2298
rect 4089 2357 4203 2479
rect 4284 2512 4471 2616
rect 4587 2792 4653 2861
rect 4587 2758 4603 2792
rect 4637 2758 4653 2792
rect 4587 2721 4653 2758
rect 4587 2687 4603 2721
rect 4637 2687 4653 2721
rect 4587 2650 4653 2687
rect 5225 2790 5381 2825
rect 5225 2756 5238 2790
rect 5272 2756 5334 2790
rect 5225 2750 5334 2756
rect 5368 2750 5381 2790
rect 5225 2704 5381 2750
rect 5225 2670 5238 2704
rect 5272 2670 5334 2704
rect 5368 2670 5381 2704
rect 5225 2654 5381 2670
rect 5418 2792 5484 2861
rect 5418 2758 5434 2792
rect 5468 2758 5484 2792
rect 5418 2721 5484 2758
rect 5418 2687 5434 2721
rect 5468 2687 5484 2721
rect 4587 2616 4603 2650
rect 4637 2616 4653 2650
rect 4587 2600 4653 2616
rect 5418 2650 5484 2687
rect 5418 2616 5434 2650
rect 5468 2616 5484 2650
rect 5418 2598 5484 2616
rect 5628 2792 5815 2861
rect 5628 2758 5692 2792
rect 5726 2758 5815 2792
rect 5628 2721 5815 2758
rect 5628 2687 5692 2721
rect 5726 2687 5815 2721
rect 5628 2650 5815 2687
rect 5628 2616 5692 2650
rect 5726 2616 5815 2650
rect 4284 2478 4300 2512
rect 4334 2478 4421 2512
rect 4455 2478 4471 2512
rect 4284 2462 4471 2478
rect 4526 2513 4666 2528
rect 4526 2479 4542 2513
rect 4576 2479 4666 2513
rect 4089 2323 4105 2357
rect 4139 2323 4203 2357
rect 4089 2229 4203 2323
rect 4345 2357 4411 2373
rect 4345 2323 4361 2357
rect 4395 2323 4411 2357
rect 4345 2229 4411 2323
rect 4526 2357 4666 2479
rect 5433 2513 5547 2529
rect 5433 2479 5497 2513
rect 5531 2479 5547 2513
rect 4526 2323 4617 2357
rect 4651 2323 4666 2357
rect 4526 2229 4666 2323
rect 5225 2417 5381 2433
rect 5225 2383 5238 2417
rect 5272 2383 5334 2417
rect 5368 2383 5381 2417
rect 5225 2340 5381 2383
rect 5225 2300 5238 2340
rect 5272 2334 5381 2340
rect 5272 2300 5334 2334
rect 5368 2300 5381 2334
rect 5225 2265 5381 2300
rect 5433 2357 5547 2479
rect 5628 2512 5815 2616
rect 5931 2792 5997 2861
rect 5931 2758 5947 2792
rect 5981 2758 5997 2792
rect 5931 2721 5997 2758
rect 5931 2687 5947 2721
rect 5981 2687 5997 2721
rect 5931 2650 5997 2687
rect 5931 2616 5947 2650
rect 5981 2616 5997 2650
rect 5931 2600 5997 2616
rect 6090 2792 6156 2861
rect 6090 2758 6106 2792
rect 6140 2758 6156 2792
rect 6090 2721 6156 2758
rect 6090 2687 6106 2721
rect 6140 2687 6156 2721
rect 6090 2650 6156 2687
rect 6090 2616 6106 2650
rect 6140 2616 6156 2650
rect 6090 2598 6156 2616
rect 6300 2792 6487 2861
rect 6300 2758 6364 2792
rect 6398 2758 6487 2792
rect 6300 2721 6487 2758
rect 6300 2687 6364 2721
rect 6398 2687 6487 2721
rect 6300 2650 6487 2687
rect 6300 2616 6364 2650
rect 6398 2616 6487 2650
rect 5628 2478 5644 2512
rect 5678 2478 5765 2512
rect 5799 2478 5815 2512
rect 5628 2462 5815 2478
rect 5870 2513 6010 2528
rect 5870 2479 5886 2513
rect 5920 2479 6010 2513
rect 5433 2323 5449 2357
rect 5483 2323 5547 2357
rect 5433 2229 5547 2323
rect 5689 2357 5755 2373
rect 5689 2323 5705 2357
rect 5739 2323 5755 2357
rect 5689 2229 5755 2323
rect 5870 2357 6010 2479
rect 5870 2323 5961 2357
rect 5995 2323 6010 2357
rect 5870 2229 6010 2323
rect 6105 2513 6219 2529
rect 6105 2479 6169 2513
rect 6203 2479 6219 2513
rect 6105 2357 6219 2479
rect 6300 2512 6487 2616
rect 6603 2792 6669 2861
rect 6603 2758 6619 2792
rect 6653 2758 6669 2792
rect 6603 2721 6669 2758
rect 6603 2687 6619 2721
rect 6653 2687 6669 2721
rect 6603 2650 6669 2687
rect 6603 2616 6619 2650
rect 6653 2616 6669 2650
rect 6603 2600 6669 2616
rect 6762 2792 6828 2861
rect 6762 2758 6778 2792
rect 6812 2758 6828 2792
rect 6762 2721 6828 2758
rect 6762 2687 6778 2721
rect 6812 2687 6828 2721
rect 6762 2650 6828 2687
rect 6762 2616 6778 2650
rect 6812 2616 6828 2650
rect 6762 2598 6828 2616
rect 6972 2792 7159 2861
rect 6972 2758 7036 2792
rect 7070 2758 7159 2792
rect 6972 2721 7159 2758
rect 6972 2687 7036 2721
rect 7070 2687 7159 2721
rect 6972 2650 7159 2687
rect 6972 2616 7036 2650
rect 7070 2616 7159 2650
rect 6300 2478 6316 2512
rect 6350 2478 6437 2512
rect 6471 2478 6487 2512
rect 6300 2462 6487 2478
rect 6542 2513 6682 2528
rect 6542 2479 6558 2513
rect 6592 2479 6682 2513
rect 6105 2323 6121 2357
rect 6155 2323 6219 2357
rect 6105 2229 6219 2323
rect 6361 2357 6427 2373
rect 6361 2323 6377 2357
rect 6411 2323 6427 2357
rect 6361 2229 6427 2323
rect 6542 2357 6682 2479
rect 6542 2323 6633 2357
rect 6667 2323 6682 2357
rect 6542 2229 6682 2323
rect 6777 2513 6891 2529
rect 6777 2479 6841 2513
rect 6875 2479 6891 2513
rect 6777 2357 6891 2479
rect 6972 2512 7159 2616
rect 7275 2792 7341 2861
rect 7275 2758 7291 2792
rect 7325 2758 7341 2792
rect 7275 2721 7341 2758
rect 7275 2687 7291 2721
rect 7325 2687 7341 2721
rect 7275 2650 7341 2687
rect 7275 2616 7291 2650
rect 7325 2616 7341 2650
rect 7275 2600 7341 2616
rect 8106 2792 8172 2861
rect 8106 2758 8122 2792
rect 8156 2758 8172 2792
rect 8106 2721 8172 2758
rect 8106 2687 8122 2721
rect 8156 2687 8172 2721
rect 8106 2650 8172 2687
rect 8106 2616 8122 2650
rect 8156 2616 8172 2650
rect 8106 2598 8172 2616
rect 8316 2792 8503 2861
rect 8316 2758 8380 2792
rect 8414 2758 8503 2792
rect 8316 2721 8503 2758
rect 8316 2687 8380 2721
rect 8414 2687 8503 2721
rect 8316 2650 8503 2687
rect 8316 2616 8380 2650
rect 8414 2616 8503 2650
rect 6972 2478 6988 2512
rect 7022 2478 7109 2512
rect 7143 2478 7159 2512
rect 6972 2462 7159 2478
rect 7214 2513 7354 2528
rect 7214 2479 7230 2513
rect 7264 2479 7354 2513
rect 6777 2323 6793 2357
rect 6827 2323 6891 2357
rect 6777 2229 6891 2323
rect 7033 2357 7099 2373
rect 7033 2323 7049 2357
rect 7083 2323 7099 2357
rect 7033 2229 7099 2323
rect 7214 2357 7354 2479
rect 7214 2323 7305 2357
rect 7339 2323 7354 2357
rect 7214 2229 7354 2323
rect 8121 2513 8235 2529
rect 8121 2479 8185 2513
rect 8219 2479 8235 2513
rect 8121 2357 8235 2479
rect 8316 2512 8503 2616
rect 8619 2792 8685 2861
rect 8619 2758 8635 2792
rect 8669 2758 8685 2792
rect 8619 2721 8685 2758
rect 8619 2687 8635 2721
rect 8669 2687 8685 2721
rect 8619 2650 8685 2687
rect 8619 2616 8635 2650
rect 8669 2616 8685 2650
rect 8619 2600 8685 2616
rect 8778 2792 8844 2861
rect 8778 2758 8794 2792
rect 8828 2758 8844 2792
rect 8778 2721 8844 2758
rect 8778 2687 8794 2721
rect 8828 2687 8844 2721
rect 8778 2650 8844 2687
rect 8778 2616 8794 2650
rect 8828 2616 8844 2650
rect 8778 2598 8844 2616
rect 8988 2792 9175 2861
rect 8988 2758 9052 2792
rect 9086 2758 9175 2792
rect 8988 2721 9175 2758
rect 8988 2687 9052 2721
rect 9086 2687 9175 2721
rect 8988 2650 9175 2687
rect 8988 2616 9052 2650
rect 9086 2616 9175 2650
rect 8316 2478 8332 2512
rect 8366 2478 8453 2512
rect 8487 2478 8503 2512
rect 8316 2462 8503 2478
rect 8558 2513 8698 2528
rect 8558 2479 8574 2513
rect 8608 2479 8698 2513
rect 8121 2323 8137 2357
rect 8171 2323 8235 2357
rect 8121 2229 8235 2323
rect 8377 2357 8443 2373
rect 8377 2323 8393 2357
rect 8427 2323 8443 2357
rect 8377 2229 8443 2323
rect 8558 2357 8698 2479
rect 8558 2323 8649 2357
rect 8683 2323 8698 2357
rect 8558 2229 8698 2323
rect 8793 2513 8907 2529
rect 8793 2479 8857 2513
rect 8891 2479 8907 2513
rect 8793 2357 8907 2479
rect 8988 2512 9175 2616
rect 9291 2792 9357 2861
rect 9291 2758 9307 2792
rect 9341 2758 9357 2792
rect 9291 2721 9357 2758
rect 9291 2687 9307 2721
rect 9341 2687 9357 2721
rect 9291 2650 9357 2687
rect 9291 2616 9307 2650
rect 9341 2616 9357 2650
rect 9291 2600 9357 2616
rect 9450 2792 9516 2861
rect 9450 2758 9466 2792
rect 9500 2758 9516 2792
rect 9450 2721 9516 2758
rect 9450 2687 9466 2721
rect 9500 2687 9516 2721
rect 9450 2650 9516 2687
rect 9450 2616 9466 2650
rect 9500 2616 9516 2650
rect 9450 2598 9516 2616
rect 9660 2792 9774 2861
rect 9660 2758 9724 2792
rect 9758 2758 9774 2792
rect 9660 2721 9774 2758
rect 9660 2687 9724 2721
rect 9758 2687 9774 2721
rect 9660 2650 9774 2687
rect 9833 2790 9893 2861
rect 9833 2756 9846 2790
rect 9880 2756 9893 2790
rect 9833 2704 9893 2756
rect 9833 2670 9846 2704
rect 9880 2670 9893 2704
rect 9833 2653 9893 2670
rect 10121 2790 10181 2861
rect 10121 2756 10134 2790
rect 10168 2756 10181 2790
rect 10121 2704 10181 2756
rect 10121 2670 10134 2704
rect 10168 2670 10181 2704
rect 10121 2653 10181 2670
rect 10692 2716 10788 2750
rect 11092 2716 11188 2750
rect 10692 2654 10726 2716
rect 9660 2616 9724 2650
rect 9758 2616 9774 2650
rect 8988 2478 9004 2512
rect 9038 2478 9125 2512
rect 9159 2478 9175 2512
rect 8988 2462 9175 2478
rect 9230 2513 9370 2528
rect 9230 2479 9246 2513
rect 9280 2479 9370 2513
rect 8793 2323 8809 2357
rect 8843 2323 8907 2357
rect 8793 2229 8907 2323
rect 9049 2357 9115 2373
rect 9049 2323 9065 2357
rect 9099 2323 9115 2357
rect 9049 2229 9115 2323
rect 9230 2357 9370 2479
rect 9230 2323 9321 2357
rect 9355 2323 9370 2357
rect 9230 2229 9370 2323
rect 9465 2513 9579 2529
rect 9465 2479 9529 2513
rect 9563 2479 9579 2513
rect 9465 2357 9579 2479
rect 9660 2512 9774 2616
rect 9660 2478 9676 2512
rect 9710 2478 9774 2512
rect 9660 2462 9774 2478
rect 9833 2417 9893 2433
rect 9833 2383 9846 2417
rect 9880 2383 9893 2417
rect 9465 2323 9481 2357
rect 9515 2323 9579 2357
rect 9465 2229 9579 2323
rect 9721 2357 9787 2373
rect 9721 2323 9737 2357
rect 9771 2323 9787 2357
rect 9721 2229 9787 2323
rect 9833 2334 9893 2383
rect 9833 2300 9846 2334
rect 9880 2300 9893 2334
rect 9833 2229 9893 2300
rect 10121 2417 10181 2433
rect 10121 2383 10134 2417
rect 10168 2383 10181 2417
rect 10121 2334 10181 2383
rect 10121 2300 10134 2334
rect 10168 2300 10181 2334
rect 10121 2229 10181 2300
rect 2039 2195 2070 2229
rect 2104 2195 2166 2229
rect 2200 2195 2262 2229
rect 2296 2195 2358 2229
rect 2392 2195 2454 2229
rect 2488 2195 2550 2229
rect 2584 2195 2646 2229
rect 2680 2195 2742 2229
rect 2776 2195 2838 2229
rect 2872 2195 2934 2229
rect 2968 2195 3030 2229
rect 3064 2195 3126 2229
rect 3160 2195 3222 2229
rect 3256 2195 3318 2229
rect 3352 2195 3414 2229
rect 3448 2195 3510 2229
rect 3544 2195 3606 2229
rect 3640 2195 3702 2229
rect 3736 2195 3798 2229
rect 3832 2195 3894 2229
rect 3928 2195 3990 2229
rect 4024 2195 4086 2229
rect 4120 2195 4182 2229
rect 4216 2195 4278 2229
rect 4312 2195 4374 2229
rect 4408 2195 4470 2229
rect 4504 2195 4566 2229
rect 4600 2195 4662 2229
rect 4696 2195 4758 2229
rect 4792 2195 4854 2229
rect 4888 2195 4950 2229
rect 4984 2195 5046 2229
rect 5080 2195 5142 2229
rect 5176 2195 5238 2229
rect 5272 2195 5334 2229
rect 5368 2195 5430 2229
rect 5464 2195 5526 2229
rect 5560 2195 5622 2229
rect 5656 2195 5718 2229
rect 5752 2195 5814 2229
rect 5848 2195 5910 2229
rect 5944 2195 6006 2229
rect 6040 2195 6102 2229
rect 6136 2195 6198 2229
rect 6232 2195 6294 2229
rect 6328 2195 6390 2229
rect 6424 2195 6486 2229
rect 6520 2195 6582 2229
rect 6616 2195 6678 2229
rect 6712 2195 6774 2229
rect 6808 2195 6870 2229
rect 6904 2195 6966 2229
rect 7000 2195 7062 2229
rect 7096 2195 7158 2229
rect 7192 2195 7254 2229
rect 7288 2195 7350 2229
rect 7384 2195 7446 2229
rect 7480 2195 7542 2229
rect 7576 2195 7638 2229
rect 7672 2195 7734 2229
rect 7768 2195 7830 2229
rect 7864 2195 7926 2229
rect 7960 2195 8022 2229
rect 8056 2195 8118 2229
rect 8152 2195 8214 2229
rect 8248 2195 8310 2229
rect 8344 2195 8406 2229
rect 8440 2195 8502 2229
rect 8536 2195 8598 2229
rect 8632 2195 8694 2229
rect 8728 2195 8790 2229
rect 8824 2195 8886 2229
rect 8920 2195 8982 2229
rect 9016 2195 9078 2229
rect 9112 2195 9174 2229
rect 9208 2195 9270 2229
rect 9304 2195 9366 2229
rect 9400 2195 9462 2229
rect 9496 2195 9558 2229
rect 9592 2195 9654 2229
rect 9688 2195 9750 2229
rect 9784 2195 9846 2229
rect 9880 2195 9942 2229
rect 9976 2195 10038 2229
rect 10072 2195 10134 2229
rect 10168 2195 10199 2229
rect 2057 2124 2117 2195
rect 2057 2090 2070 2124
rect 2104 2090 2117 2124
rect 2057 2041 2117 2090
rect 2057 2007 2070 2041
rect 2104 2007 2117 2041
rect 2057 1991 2117 2007
rect 2154 2140 2308 2159
rect 2154 2106 2174 2140
rect 2208 2106 2254 2140
rect 2288 2106 2308 2140
rect 2154 2072 2308 2106
rect 2154 2038 2174 2072
rect 2208 2038 2254 2072
rect 2288 2038 2308 2072
rect 2154 2004 2308 2038
rect 2154 1970 2174 2004
rect 2208 1970 2254 2004
rect 2288 1970 2308 2004
rect 2424 2126 2490 2195
rect 2424 2092 2440 2126
rect 2474 2092 2490 2126
rect 2424 2036 2490 2092
rect 2424 2002 2440 2036
rect 2474 2002 2490 2036
rect 2424 1986 2490 2002
rect 2524 2126 2590 2142
rect 2524 2092 2540 2126
rect 2574 2092 2590 2126
rect 2524 2036 2590 2092
rect 3793 2126 3859 2195
rect 3793 2092 3809 2126
rect 3843 2092 3859 2126
rect 2524 2002 2540 2036
rect 2574 2002 2590 2036
rect 2154 1952 2308 1970
rect 2154 1936 2490 1952
rect 2154 1902 2368 1936
rect 2406 1902 2440 1936
rect 2474 1902 2490 1936
rect 2154 1856 2490 1902
rect 2524 1944 2590 2002
rect 2524 1885 2691 1944
rect 2057 1754 2117 1771
rect 2057 1720 2070 1754
rect 2104 1720 2117 1754
rect 2057 1668 2117 1720
rect 2057 1634 2070 1668
rect 2104 1634 2117 1668
rect 2057 1563 2117 1634
rect 2154 1599 2308 1856
rect 2524 1832 2590 1885
rect 2424 1806 2490 1822
rect 2424 1772 2440 1806
rect 2474 1772 2490 1806
rect 2424 1736 2490 1772
rect 2424 1702 2440 1736
rect 2474 1702 2490 1736
rect 2424 1666 2490 1702
rect 2424 1632 2440 1666
rect 2474 1632 2490 1666
rect 2424 1563 2490 1632
rect 2524 1798 2540 1832
rect 2574 1798 2590 1832
rect 2524 1749 2590 1798
rect 3793 2044 3859 2092
rect 3957 2126 4023 2142
rect 3957 2092 3973 2126
rect 4007 2120 4023 2126
rect 3957 2086 3974 2092
rect 4008 2086 4023 2120
rect 4180 2126 4256 2195
rect 3957 2044 4023 2086
rect 3793 2010 3809 2044
rect 3843 2010 3859 2044
rect 3900 2010 3973 2044
rect 4007 2010 4023 2044
rect 4078 2062 4144 2104
rect 4078 2028 4094 2062
rect 4128 2028 4144 2062
rect 3900 1976 3934 2010
rect 4078 1986 4144 2028
rect 4180 2092 4201 2126
rect 4235 2092 4256 2126
rect 4180 2076 4256 2092
rect 4290 2118 4680 2134
rect 4290 2084 4396 2118
rect 4430 2084 4680 2118
rect 4180 2036 4222 2076
rect 4290 2042 4324 2084
rect 4180 2002 4183 2036
rect 4217 2002 4222 2036
rect 4180 1986 4222 2002
rect 4256 2008 4324 2042
rect 4358 2016 4612 2050
rect 3788 1968 3854 1976
rect 3655 1952 3854 1968
rect 3655 1918 3804 1952
rect 3838 1918 3854 1952
rect 3655 1902 3854 1918
rect 3788 1832 3854 1848
rect 3788 1798 3804 1832
rect 3838 1798 3854 1832
rect 2524 1715 2540 1749
rect 2574 1715 2590 1749
rect 2524 1666 2590 1715
rect 2524 1632 2540 1666
rect 2574 1632 2590 1666
rect 2524 1616 2590 1632
rect 3788 1749 3854 1798
rect 3788 1715 3804 1749
rect 3838 1715 3854 1749
rect 3788 1666 3854 1715
rect 3788 1632 3804 1666
rect 3838 1632 3854 1666
rect 3788 1563 3854 1632
rect 3888 1832 3934 1976
rect 3968 1952 4034 1976
rect 3968 1918 3984 1952
rect 4018 1918 4034 1952
rect 3968 1902 4034 1918
rect 3888 1798 3894 1832
rect 3928 1798 3934 1832
rect 3888 1749 3934 1798
rect 3888 1715 3894 1749
rect 3928 1715 3934 1749
rect 3888 1666 3934 1715
rect 3888 1632 3894 1666
rect 3928 1632 3934 1666
rect 3888 1616 3934 1632
rect 3968 1832 4034 1848
rect 3968 1798 3984 1832
rect 4018 1798 4034 1832
rect 3968 1749 4034 1798
rect 3968 1715 3984 1749
rect 4018 1715 4034 1749
rect 3968 1666 4034 1715
rect 4078 1822 4112 1986
rect 4156 1929 4222 1942
rect 4156 1895 4171 1929
rect 4205 1926 4222 1929
rect 4156 1892 4172 1895
rect 4206 1892 4222 1926
rect 4156 1856 4222 1892
rect 4256 1868 4290 2008
rect 4358 1968 4392 2016
rect 4324 1952 4392 1968
rect 4324 1918 4340 1952
rect 4374 1918 4392 1952
rect 4324 1902 4392 1918
rect 4432 1952 4510 1976
rect 4432 1918 4448 1952
rect 4482 1918 4510 1952
rect 4432 1902 4510 1918
rect 4546 1954 4612 2016
rect 4646 2016 4680 2084
rect 4714 2100 4780 2195
rect 4714 2066 4730 2100
rect 4764 2066 4780 2100
rect 4714 2050 4780 2066
rect 4828 2126 4902 2142
rect 4828 2092 4844 2126
rect 4878 2092 4902 2126
rect 4828 2036 4902 2092
rect 4646 1982 4794 2016
rect 4828 2002 4844 2036
rect 4878 2002 4902 2036
rect 4828 1986 4902 2002
rect 4945 2126 4995 2195
rect 4945 2092 4961 2126
rect 4945 2036 4995 2092
rect 4945 2002 4961 2036
rect 4945 1986 4995 2002
rect 5031 2126 5097 2142
rect 5031 2092 5047 2126
rect 5081 2092 5097 2126
rect 5031 2036 5097 2092
rect 5031 2002 5047 2036
rect 5081 2002 5097 2036
rect 5031 1986 5097 2002
rect 5133 2126 5183 2195
rect 5167 2092 5183 2126
rect 5133 2036 5183 2092
rect 5167 2002 5183 2036
rect 5133 1986 5183 2002
rect 5225 2124 5381 2159
rect 5225 2084 5238 2124
rect 5272 2090 5334 2124
rect 5368 2090 5381 2124
rect 5272 2084 5381 2090
rect 5225 2041 5381 2084
rect 5225 2007 5238 2041
rect 5272 2007 5334 2041
rect 5368 2007 5381 2041
rect 5225 1991 5381 2007
rect 5427 2076 5493 2195
rect 5427 2042 5443 2076
rect 5477 2042 5493 2076
rect 5427 2021 5493 2042
rect 5591 2071 5737 2087
rect 5591 2037 5607 2071
rect 5641 2037 5687 2071
rect 5721 2037 5737 2071
rect 5591 2021 5737 2037
rect 5835 2077 5885 2195
rect 6185 2164 6235 2195
rect 5835 2043 5851 2077
rect 5835 2022 5885 2043
rect 5919 2127 6106 2161
rect 5427 1987 5492 2021
rect 5696 1988 5737 2021
rect 5919 1988 5953 2127
rect 4546 1918 4562 1954
rect 4596 1918 4612 1954
rect 4760 1952 4794 1982
rect 4546 1902 4612 1918
rect 4646 1932 4726 1948
rect 4646 1898 4676 1932
rect 4710 1898 4726 1932
rect 4646 1882 4726 1898
rect 4760 1936 4834 1952
rect 4760 1902 4784 1936
rect 4818 1902 4834 1936
rect 4760 1886 4834 1902
rect 4256 1834 4534 1868
rect 4468 1832 4534 1834
rect 4078 1817 4144 1822
rect 4078 1783 4094 1817
rect 4128 1800 4144 1817
rect 4128 1783 4319 1800
rect 4078 1766 4319 1783
rect 4078 1722 4144 1766
rect 4078 1688 4094 1722
rect 4128 1688 4144 1722
rect 4078 1672 4144 1688
rect 4185 1727 4251 1732
rect 4185 1693 4201 1727
rect 4235 1693 4251 1727
rect 3968 1632 3984 1666
rect 4018 1632 4034 1666
rect 3968 1563 4034 1632
rect 4185 1563 4251 1693
rect 4285 1631 4319 1766
rect 4468 1798 4484 1832
rect 4518 1798 4534 1832
rect 4468 1715 4534 1798
rect 4468 1681 4484 1715
rect 4518 1681 4534 1715
rect 4468 1665 4534 1681
rect 4646 1631 4680 1882
rect 4868 1848 4902 1986
rect 4940 1941 5006 1952
rect 4940 1907 4955 1941
rect 4989 1936 5006 1941
rect 4940 1902 4956 1907
rect 4990 1902 5006 1936
rect 4940 1856 5006 1902
rect 4285 1597 4680 1631
rect 4714 1832 4780 1848
rect 4714 1798 4730 1832
rect 4764 1798 4780 1832
rect 4714 1749 4780 1798
rect 4714 1715 4730 1749
rect 4764 1715 4780 1749
rect 4714 1666 4780 1715
rect 4714 1632 4730 1666
rect 4764 1632 4780 1666
rect 4714 1563 4780 1632
rect 4814 1832 4902 1848
rect 4814 1798 4830 1832
rect 4864 1798 4902 1832
rect 5040 1832 5097 1986
rect 5424 1971 5662 1987
rect 5424 1937 5459 1971
rect 5493 1937 5576 1971
rect 5610 1937 5662 1971
rect 5696 1954 5953 1988
rect 5987 2066 6038 2093
rect 6021 2032 6038 2066
rect 6072 2080 6106 2127
rect 6185 2130 6201 2164
rect 6185 2114 6235 2130
rect 6269 2127 6455 2161
rect 6269 2080 6303 2127
rect 6072 2046 6303 2080
rect 6337 2077 6387 2093
rect 5424 1920 5662 1937
rect 5424 1903 5509 1920
rect 5424 1869 5459 1903
rect 5493 1869 5509 1903
rect 4814 1767 4902 1798
rect 4814 1749 4847 1767
rect 4814 1715 4830 1749
rect 4881 1733 4902 1767
rect 4864 1715 4902 1733
rect 4814 1666 4902 1715
rect 4814 1632 4830 1666
rect 4864 1632 4902 1666
rect 4814 1616 4902 1632
rect 4940 1806 5006 1822
rect 4940 1772 4956 1806
rect 4990 1772 5006 1806
rect 4940 1736 5006 1772
rect 4940 1702 4956 1736
rect 4990 1702 5006 1736
rect 4940 1666 5006 1702
rect 4940 1632 4956 1666
rect 4990 1632 5006 1666
rect 4940 1563 5006 1632
rect 5040 1798 5046 1832
rect 5080 1798 5097 1832
rect 5040 1749 5097 1798
rect 5040 1715 5046 1749
rect 5080 1715 5097 1749
rect 5040 1695 5097 1715
rect 5040 1666 5049 1695
rect 5040 1632 5046 1666
rect 5083 1661 5097 1695
rect 5080 1632 5097 1661
rect 5040 1616 5097 1632
rect 5136 1832 5186 1848
rect 5170 1798 5186 1832
rect 5136 1749 5186 1798
rect 5424 1835 5509 1869
rect 5560 1903 5662 1920
rect 5560 1869 5576 1903
rect 5610 1869 5662 1903
rect 5560 1853 5662 1869
rect 5696 1905 5762 1920
rect 5696 1904 5716 1905
rect 5696 1870 5712 1904
rect 5750 1871 5762 1905
rect 5746 1870 5762 1871
rect 5696 1854 5762 1870
rect 5424 1801 5459 1835
rect 5493 1801 5509 1835
rect 5796 1820 5830 1954
rect 5987 1916 6038 2032
rect 6337 2043 6353 2077
rect 6083 1978 6099 2012
rect 6133 1978 6246 2012
rect 6212 1944 6246 1978
rect 6337 2009 6387 2043
rect 6421 2044 6455 2127
rect 6489 2128 6543 2195
rect 6489 2094 6491 2128
rect 6525 2094 6543 2128
rect 6489 2078 6543 2094
rect 6588 2125 6822 2159
rect 6588 2044 6622 2125
rect 6421 2010 6622 2044
rect 6656 2062 6722 2091
rect 6656 2028 6672 2062
rect 6706 2028 6722 2062
rect 6337 1976 6353 2009
rect 6322 1975 6353 1976
rect 6387 1975 6622 1976
rect 6322 1970 6622 1975
rect 5920 1900 6038 1916
rect 5920 1866 5936 1900
rect 5970 1866 6038 1900
rect 5920 1850 6038 1866
rect 6096 1926 6178 1942
rect 6096 1892 6124 1926
rect 6162 1892 6178 1926
rect 6096 1856 6178 1892
rect 6212 1928 6288 1944
rect 6212 1894 6238 1928
rect 6272 1894 6288 1928
rect 6212 1878 6288 1894
rect 6322 1942 6582 1970
rect 5424 1785 5509 1801
rect 5696 1786 5830 1820
rect 5170 1715 5186 1749
rect 5136 1666 5186 1715
rect 5170 1632 5186 1666
rect 5136 1563 5186 1632
rect 5225 1754 5381 1770
rect 5225 1720 5238 1754
rect 5272 1720 5334 1754
rect 5368 1720 5381 1754
rect 5696 1752 5730 1786
rect 5225 1674 5381 1720
rect 5225 1668 5334 1674
rect 5225 1634 5238 1668
rect 5272 1634 5334 1668
rect 5368 1634 5381 1674
rect 5225 1599 5381 1634
rect 5422 1735 5646 1751
rect 5422 1701 5438 1735
rect 5472 1717 5646 1735
rect 5422 1666 5472 1701
rect 5422 1632 5438 1666
rect 5422 1616 5472 1632
rect 5512 1667 5578 1683
rect 5512 1633 5528 1667
rect 5562 1633 5578 1667
rect 5512 1563 5578 1633
rect 5612 1631 5646 1717
rect 5680 1726 5730 1752
rect 5680 1692 5696 1726
rect 5680 1665 5730 1692
rect 5770 1736 5836 1752
rect 5770 1702 5786 1736
rect 5820 1702 5836 1736
rect 5770 1666 5836 1702
rect 5770 1632 5786 1666
rect 5820 1632 5836 1666
rect 5770 1631 5836 1632
rect 5612 1597 5836 1631
rect 5882 1736 5948 1752
rect 5882 1702 5898 1736
rect 5932 1702 5948 1736
rect 5882 1666 5948 1702
rect 5882 1632 5898 1666
rect 5932 1632 5948 1666
rect 5882 1563 5948 1632
rect 5988 1736 6038 1850
rect 6212 1822 6246 1878
rect 6322 1844 6356 1942
rect 6518 1936 6582 1942
rect 6616 1936 6622 1970
rect 6656 1975 6722 2028
rect 6756 2067 6822 2125
rect 6868 2127 7123 2159
rect 6868 2093 6893 2127
rect 6927 2125 7123 2127
rect 6927 2093 6953 2125
rect 6868 2077 6953 2093
rect 7089 2091 7123 2125
rect 6756 2033 6772 2067
rect 6806 2043 6822 2067
rect 6989 2057 7055 2091
rect 6806 2033 6940 2043
rect 6756 2009 6940 2033
rect 6989 2023 7005 2057
rect 7039 2023 7055 2057
rect 7089 2075 7176 2091
rect 7089 2041 7115 2075
rect 7149 2041 7176 2075
rect 7089 2025 7176 2041
rect 7210 2075 7276 2195
rect 7735 2160 7810 2195
rect 7210 2041 7226 2075
rect 7260 2041 7276 2075
rect 7210 2024 7276 2041
rect 7310 2126 7701 2160
rect 7735 2126 7755 2160
rect 7789 2126 7810 2160
rect 7846 2147 8118 2161
rect 7846 2127 8068 2147
rect 7846 2126 7930 2127
rect 6656 1941 6872 1975
rect 6518 1907 6622 1936
rect 6806 1939 6872 1941
rect 6518 1894 6764 1907
rect 6518 1860 6534 1894
rect 6568 1891 6764 1894
rect 6568 1860 6714 1891
rect 6518 1857 6714 1860
rect 6748 1857 6764 1891
rect 6022 1702 6038 1736
rect 5988 1666 6038 1702
rect 6022 1632 6038 1666
rect 5988 1616 6038 1632
rect 6084 1806 6246 1822
rect 6084 1772 6100 1806
rect 6134 1788 6246 1806
rect 6280 1828 6356 1844
rect 6314 1794 6356 1828
rect 6084 1736 6134 1772
rect 6084 1702 6100 1736
rect 6084 1666 6134 1702
rect 6084 1632 6100 1666
rect 6084 1616 6134 1632
rect 6174 1744 6240 1754
rect 6174 1710 6190 1744
rect 6224 1710 6240 1744
rect 6174 1666 6240 1710
rect 6174 1632 6190 1666
rect 6224 1632 6240 1666
rect 6174 1563 6240 1632
rect 6280 1747 6356 1794
rect 6406 1830 6472 1846
rect 6518 1844 6764 1857
rect 6698 1841 6764 1844
rect 6806 1905 6822 1939
rect 6856 1905 6872 1939
rect 6806 1871 6872 1905
rect 6406 1796 6422 1830
rect 6456 1810 6472 1830
rect 6806 1837 6822 1871
rect 6856 1837 6872 1871
rect 6456 1796 6510 1810
rect 6806 1804 6872 1837
rect 6406 1776 6510 1796
rect 6314 1713 6356 1747
rect 6280 1666 6356 1713
rect 6314 1632 6356 1666
rect 6280 1616 6356 1632
rect 6392 1718 6442 1742
rect 6426 1684 6442 1718
rect 6392 1563 6442 1684
rect 6476 1631 6510 1776
rect 6567 1770 6872 1804
rect 6567 1726 6633 1770
rect 6906 1736 6940 2009
rect 6567 1692 6583 1726
rect 6617 1692 6633 1726
rect 6567 1665 6633 1692
rect 6667 1726 6940 1736
rect 6667 1692 6683 1726
rect 6717 1702 6940 1726
rect 6974 1989 7055 2023
rect 7310 1990 7344 2126
rect 7667 2092 7701 2126
rect 7846 2092 7871 2126
rect 7905 2092 7930 2126
rect 8052 2113 8068 2127
rect 8102 2113 8118 2147
rect 8364 2126 8421 2195
rect 7391 2058 7407 2092
rect 7441 2058 7489 2092
rect 7523 2058 7571 2092
rect 7605 2058 7621 2092
rect 7667 2058 7812 2092
rect 7966 2079 8016 2093
rect 8364 2092 8385 2126
rect 8419 2092 8421 2126
rect 7966 2074 8297 2079
rect 7391 2042 7621 2058
rect 7587 2024 7621 2042
rect 7778 2024 7932 2058
rect 7587 1990 7744 2024
rect 6974 1787 7008 1989
rect 7089 1956 7344 1990
rect 7430 1970 7496 1976
rect 7089 1955 7123 1956
rect 7042 1939 7123 1955
rect 7042 1905 7058 1939
rect 7092 1905 7123 1939
rect 7430 1936 7446 1970
rect 7480 1956 7496 1970
rect 7480 1943 7676 1956
rect 7480 1936 7626 1943
rect 7042 1871 7123 1905
rect 7042 1837 7058 1871
rect 7092 1837 7123 1871
rect 7157 1906 7288 1922
rect 7157 1872 7173 1906
rect 7207 1896 7288 1906
rect 7430 1911 7626 1936
rect 7207 1872 7254 1896
rect 7157 1862 7254 1872
rect 7157 1856 7288 1862
rect 7322 1880 7388 1896
rect 7042 1821 7123 1837
rect 7322 1846 7338 1880
rect 7372 1846 7388 1880
rect 7430 1877 7446 1911
rect 7480 1909 7626 1911
rect 7660 1909 7676 1943
rect 7480 1896 7676 1909
rect 7480 1877 7496 1896
rect 7430 1861 7496 1877
rect 7710 1862 7744 1990
rect 7898 1986 7932 2024
rect 8000 2045 8297 2074
rect 8000 2040 8016 2045
rect 7966 2020 8016 2040
rect 8263 2011 8330 2045
rect 8120 1995 8229 2011
rect 8120 1986 8179 1995
rect 7790 1952 7864 1976
rect 7790 1918 7806 1952
rect 7840 1918 7864 1952
rect 7790 1896 7864 1918
rect 7898 1961 8179 1986
rect 8213 1961 8229 1995
rect 7898 1952 8229 1961
rect 7898 1918 7914 1952
rect 7948 1918 7964 1952
rect 8120 1945 8229 1952
rect 7898 1902 7964 1918
rect 8006 1902 8072 1918
rect 7790 1862 7830 1896
rect 8006 1868 8022 1902
rect 8056 1868 8072 1902
rect 7322 1822 7388 1846
rect 7180 1788 7388 1822
rect 7547 1828 7749 1862
rect 7898 1834 8072 1868
rect 7898 1828 7932 1834
rect 7547 1792 7581 1828
rect 7715 1794 7932 1828
rect 8120 1811 8154 1945
rect 8296 1926 8330 2011
rect 8364 2036 8421 2092
rect 8364 2002 8385 2036
rect 8419 2002 8421 2036
rect 8364 1986 8421 2002
rect 8455 2126 8521 2142
rect 8455 2092 8471 2126
rect 8505 2092 8521 2126
rect 8455 2036 8521 2092
rect 8455 2002 8471 2036
rect 8505 2002 8521 2036
rect 8455 1968 8521 2002
rect 8555 2126 8621 2195
rect 8555 2092 8557 2126
rect 8591 2092 8621 2126
rect 8773 2126 8839 2195
rect 8555 2036 8621 2092
rect 8555 2002 8557 2036
rect 8591 2002 8621 2036
rect 8555 1986 8621 2002
rect 8667 2100 8733 2104
rect 8667 2066 8683 2100
rect 8717 2066 8733 2100
rect 8667 2032 8733 2066
rect 8667 1998 8683 2032
rect 8717 1998 8733 2032
rect 8773 2092 8789 2126
rect 8823 2092 8839 2126
rect 8773 2052 8839 2092
rect 8773 2018 8789 2052
rect 8823 2018 8839 2052
rect 8773 2002 8839 2018
rect 8873 2126 8940 2142
rect 8873 2092 8889 2126
rect 8923 2092 8940 2126
rect 8873 2052 8940 2092
rect 8873 2018 8889 2052
rect 8923 2018 8940 2052
rect 8873 2002 8940 2018
rect 8188 1895 8254 1911
rect 8188 1894 8204 1895
rect 8188 1860 8203 1894
rect 8238 1861 8254 1895
rect 8237 1860 8254 1861
rect 8188 1845 8254 1860
rect 8296 1910 8362 1926
rect 8296 1876 8312 1910
rect 8346 1876 8362 1910
rect 8296 1860 8362 1876
rect 8474 1902 8521 1968
rect 8667 1968 8733 1998
rect 8667 1952 8872 1968
rect 8667 1918 8822 1952
rect 8856 1918 8872 1952
rect 8667 1902 8872 1918
rect 7180 1787 7246 1788
rect 6974 1776 7246 1787
rect 6974 1753 7196 1776
rect 6717 1692 6733 1702
rect 6667 1665 6733 1692
rect 6974 1666 7008 1753
rect 7180 1742 7196 1753
rect 7230 1742 7246 1776
rect 7460 1776 7581 1792
rect 6779 1632 6795 1666
rect 6829 1632 6914 1666
rect 6948 1632 7008 1666
rect 7072 1703 7138 1719
rect 7072 1669 7088 1703
rect 7122 1669 7138 1703
rect 6779 1631 6964 1632
rect 6476 1597 6964 1631
rect 7072 1563 7138 1669
rect 7180 1666 7246 1742
rect 7180 1632 7196 1666
rect 7230 1632 7246 1666
rect 7180 1616 7246 1632
rect 7292 1738 7358 1754
rect 7292 1704 7308 1738
rect 7342 1704 7358 1738
rect 7292 1666 7358 1704
rect 7292 1632 7308 1666
rect 7342 1632 7358 1666
rect 7292 1563 7358 1632
rect 7460 1742 7476 1776
rect 7510 1758 7581 1776
rect 7615 1786 7681 1794
rect 7510 1742 7526 1758
rect 7460 1666 7526 1742
rect 7615 1752 7631 1786
rect 7665 1760 7681 1786
rect 8036 1784 8086 1800
rect 8036 1760 8052 1784
rect 7665 1752 8052 1760
rect 7615 1750 8052 1752
rect 7615 1744 8086 1750
rect 8120 1795 8214 1811
rect 8120 1761 8164 1795
rect 8198 1761 8214 1795
rect 8120 1745 8214 1761
rect 7615 1726 7776 1744
rect 7760 1710 7776 1726
rect 7810 1726 8086 1744
rect 7810 1710 7826 1726
rect 7460 1632 7476 1666
rect 7510 1632 7526 1666
rect 7460 1616 7526 1632
rect 7645 1671 7711 1692
rect 7645 1637 7661 1671
rect 7695 1637 7711 1671
rect 7645 1563 7711 1637
rect 7760 1666 7826 1710
rect 8036 1711 8086 1726
rect 8296 1711 8330 1860
rect 8474 1856 8542 1902
rect 8474 1832 8524 1856
rect 7760 1632 7776 1666
rect 7810 1632 7826 1666
rect 7760 1616 7826 1632
rect 7860 1671 7926 1692
rect 7860 1637 7876 1671
rect 7910 1637 7926 1671
rect 7860 1563 7926 1637
rect 8036 1677 8330 1711
rect 8364 1799 8433 1822
rect 8364 1765 8383 1799
rect 8417 1765 8433 1799
rect 8364 1717 8433 1765
rect 8364 1683 8383 1717
rect 8417 1683 8433 1717
rect 8036 1666 8086 1677
rect 8036 1632 8052 1666
rect 8364 1643 8433 1683
rect 8036 1616 8086 1632
rect 8255 1627 8433 1643
rect 8255 1593 8271 1627
rect 8305 1593 8383 1627
rect 8417 1593 8433 1627
rect 8474 1798 8490 1832
rect 8474 1749 8524 1798
rect 8474 1715 8490 1749
rect 8474 1666 8524 1715
rect 8474 1632 8490 1666
rect 8474 1616 8524 1632
rect 8564 1806 8630 1822
rect 8564 1772 8580 1806
rect 8614 1772 8630 1806
rect 8564 1736 8630 1772
rect 8564 1702 8580 1736
rect 8614 1702 8630 1736
rect 8564 1666 8630 1702
rect 8564 1632 8580 1666
rect 8614 1632 8630 1666
rect 8255 1563 8433 1593
rect 8564 1563 8630 1632
rect 8667 1816 8739 1902
rect 8906 1848 8940 2002
rect 8975 2126 9025 2195
rect 9009 2092 9025 2126
rect 9074 2130 9212 2195
rect 9074 2096 9090 2130
rect 9124 2096 9162 2130
rect 9196 2096 9212 2130
rect 9262 2126 9312 2142
rect 8975 2036 9025 2092
rect 9009 2002 9025 2036
rect 8975 1986 9025 2002
rect 9262 2092 9278 2126
rect 9262 2036 9312 2092
rect 9348 2104 9414 2195
rect 9348 2070 9364 2104
rect 9398 2070 9414 2104
rect 9348 2051 9414 2070
rect 9450 2126 9484 2142
rect 9262 2002 9278 2036
rect 9450 2036 9484 2092
rect 9520 2104 9586 2195
rect 9520 2070 9536 2104
rect 9570 2070 9586 2104
rect 9520 2051 9586 2070
rect 9622 2127 10080 2161
rect 9622 2126 9672 2127
rect 9656 2092 9672 2126
rect 9312 2002 9450 2010
rect 9622 2036 9672 2092
rect 9806 2104 9872 2127
rect 9484 2002 9622 2010
rect 9656 2002 9672 2036
rect 9262 1976 9672 2002
rect 9706 2072 9772 2090
rect 9706 2038 9722 2072
rect 9756 2038 9772 2072
rect 9806 2070 9822 2104
rect 9856 2070 9872 2104
rect 10014 2104 10080 2127
rect 9806 2051 9872 2070
rect 9906 2072 9980 2090
rect 9706 2010 9772 2038
rect 9906 2038 9926 2072
rect 9960 2038 9980 2072
rect 10014 2070 10030 2104
rect 10064 2070 10080 2104
rect 10014 2051 10080 2070
rect 10121 2124 10181 2195
rect 10121 2090 10134 2124
rect 10168 2090 10181 2124
rect 9906 2010 9980 2038
rect 10121 2041 10181 2090
rect 9706 1976 10078 2010
rect 10121 2007 10134 2041
rect 10168 2007 10181 2041
rect 10121 1991 10181 2007
rect 9341 1926 9694 1942
rect 9341 1892 9357 1926
rect 9391 1892 9425 1926
rect 9459 1892 9489 1926
rect 9527 1892 9561 1926
rect 9595 1892 9694 1926
rect 9341 1876 9694 1892
rect 9456 1856 9694 1876
rect 9728 1926 9998 1942
rect 9728 1892 9744 1926
rect 9778 1892 9812 1926
rect 9846 1892 9876 1926
rect 9914 1892 9948 1926
rect 9982 1892 9998 1926
rect 9728 1856 9998 1892
rect 10032 1930 10078 1976
rect 10180 1930 10280 1950
rect 10032 1850 10200 1930
rect 10260 1850 10280 1930
rect 8667 1782 8689 1816
rect 8723 1782 8739 1816
rect 8667 1745 8739 1782
rect 8667 1711 8689 1745
rect 8723 1711 8739 1745
rect 8667 1674 8739 1711
rect 8667 1640 8689 1674
rect 8723 1640 8739 1674
rect 8667 1624 8739 1640
rect 8778 1820 8844 1848
rect 8778 1786 8794 1820
rect 8828 1786 8844 1820
rect 8778 1748 8844 1786
rect 8778 1714 8794 1748
rect 8828 1714 8844 1748
rect 8778 1670 8844 1714
rect 8778 1636 8794 1670
rect 8828 1636 8844 1670
rect 8778 1563 8844 1636
rect 8878 1832 8940 1848
rect 8878 1798 8884 1832
rect 8918 1823 8940 1832
rect 8878 1789 8887 1798
rect 8921 1789 8940 1823
rect 8878 1751 8940 1789
rect 8878 1749 8887 1751
rect 8878 1715 8884 1749
rect 8921 1717 8940 1751
rect 8918 1715 8940 1717
rect 8878 1666 8940 1715
rect 8878 1632 8884 1666
rect 8918 1632 8940 1666
rect 8878 1616 8940 1632
rect 8974 1832 9024 1848
rect 9008 1798 9024 1832
rect 8974 1749 9024 1798
rect 9008 1715 9024 1749
rect 8974 1666 9024 1715
rect 9008 1632 9024 1666
rect 9262 1826 9328 1842
rect 9262 1792 9278 1826
rect 9312 1792 9328 1826
rect 10032 1822 10078 1850
rect 10180 1830 10280 1850
rect 9262 1746 9328 1792
rect 9262 1712 9278 1746
rect 9312 1712 9328 1746
rect 9262 1666 9328 1712
rect 8974 1563 9024 1632
rect 9074 1628 9090 1662
rect 9124 1628 9162 1662
rect 9196 1628 9212 1662
rect 9074 1563 9212 1628
rect 9262 1632 9278 1666
rect 9312 1632 9328 1666
rect 9262 1563 9328 1632
rect 9362 1806 10078 1822
rect 9362 1772 9369 1806
rect 9403 1772 9449 1806
rect 9483 1772 9531 1806
rect 9565 1788 9721 1806
rect 9565 1772 9571 1788
rect 9362 1735 9571 1772
rect 9705 1772 9721 1788
rect 9755 1772 9790 1806
rect 9824 1772 9861 1806
rect 9895 1772 9930 1806
rect 9964 1788 10078 1806
rect 9964 1772 9980 1788
rect 9362 1701 9369 1735
rect 9403 1701 9449 1735
rect 9483 1701 9531 1735
rect 9565 1701 9571 1735
rect 9362 1666 9571 1701
rect 9362 1632 9369 1666
rect 9403 1632 9449 1666
rect 9483 1632 9531 1666
rect 9565 1632 9571 1666
rect 9362 1616 9571 1632
rect 9605 1745 9671 1754
rect 9605 1711 9621 1745
rect 9655 1711 9671 1745
rect 9605 1666 9671 1711
rect 9605 1632 9621 1666
rect 9655 1632 9671 1666
rect 9605 1563 9671 1632
rect 9705 1735 9980 1772
rect 10121 1754 10181 1771
rect 9705 1701 9721 1735
rect 9755 1701 9790 1735
rect 9824 1701 9861 1735
rect 9895 1701 9930 1735
rect 9964 1701 9980 1735
rect 9705 1666 9980 1701
rect 9705 1632 9721 1666
rect 9755 1632 9790 1666
rect 9824 1632 9861 1666
rect 9895 1632 9930 1666
rect 9964 1632 9980 1666
rect 9705 1616 9980 1632
rect 10014 1745 10080 1754
rect 10014 1711 10030 1745
rect 10064 1711 10080 1745
rect 10014 1666 10080 1711
rect 10014 1632 10030 1666
rect 10064 1632 10080 1666
rect 10014 1563 10080 1632
rect 10121 1720 10134 1754
rect 10168 1720 10181 1754
rect 10121 1668 10181 1720
rect 10121 1634 10134 1668
rect 10168 1634 10181 1668
rect 10121 1563 10181 1634
rect 11154 2654 11188 2716
rect 10818 1684 10822 2108
rect 10892 1684 10898 2108
rect 10818 1678 10898 1684
rect 10692 1588 10726 1650
rect 11154 1588 11188 1650
rect 2039 1529 2070 1563
rect 2104 1529 2166 1563
rect 2200 1529 2262 1563
rect 2296 1529 2358 1563
rect 2392 1529 2454 1563
rect 2488 1529 2550 1563
rect 2584 1529 2646 1563
rect 2680 1529 2742 1563
rect 2776 1529 2838 1563
rect 2872 1529 2934 1563
rect 2968 1529 3030 1563
rect 3064 1529 3126 1563
rect 3160 1529 3222 1563
rect 3256 1529 3318 1563
rect 3352 1529 3414 1563
rect 3448 1529 3510 1563
rect 3544 1529 3606 1563
rect 3640 1529 3702 1563
rect 3736 1529 3798 1563
rect 3832 1529 3894 1563
rect 3928 1529 3990 1563
rect 4024 1529 4086 1563
rect 4120 1529 4182 1563
rect 4216 1529 4278 1563
rect 4312 1529 4374 1563
rect 4408 1529 4470 1563
rect 4504 1529 4566 1563
rect 4600 1529 4662 1563
rect 4696 1529 4758 1563
rect 4792 1529 4854 1563
rect 4888 1529 4950 1563
rect 4984 1529 5046 1563
rect 5080 1529 5142 1563
rect 5176 1529 5238 1563
rect 5272 1529 5334 1563
rect 5368 1529 5430 1563
rect 5464 1529 5526 1563
rect 5560 1529 5622 1563
rect 5656 1529 5718 1563
rect 5752 1529 5814 1563
rect 5848 1529 5910 1563
rect 5944 1529 6006 1563
rect 6040 1529 6102 1563
rect 6136 1529 6198 1563
rect 6232 1529 6294 1563
rect 6328 1529 6390 1563
rect 6424 1529 6486 1563
rect 6520 1529 6582 1563
rect 6616 1529 6678 1563
rect 6712 1529 6774 1563
rect 6808 1529 6870 1563
rect 6904 1529 6966 1563
rect 7000 1529 7062 1563
rect 7096 1529 7158 1563
rect 7192 1529 7254 1563
rect 7288 1529 7350 1563
rect 7384 1529 7446 1563
rect 7480 1529 7542 1563
rect 7576 1529 7638 1563
rect 7672 1529 7734 1563
rect 7768 1529 7830 1563
rect 7864 1529 7926 1563
rect 7960 1529 8022 1563
rect 8056 1529 8118 1563
rect 8152 1529 8214 1563
rect 8248 1529 8310 1563
rect 8344 1529 8406 1563
rect 8440 1529 8502 1563
rect 8536 1529 8598 1563
rect 8632 1529 8694 1563
rect 8728 1529 8790 1563
rect 8824 1529 8886 1563
rect 8920 1529 8982 1563
rect 9016 1529 9078 1563
rect 9112 1529 9174 1563
rect 9208 1529 9270 1563
rect 9304 1529 9366 1563
rect 9400 1529 9462 1563
rect 9496 1529 9558 1563
rect 9592 1529 9654 1563
rect 9688 1529 9750 1563
rect 9784 1529 9846 1563
rect 9880 1529 9942 1563
rect 9976 1529 10038 1563
rect 10072 1529 10134 1563
rect 10168 1529 10199 1563
rect 10692 1554 10788 1588
rect 11092 1554 11188 1588
rect 13778 3824 13812 3886
rect 11420 3784 11436 3818
rect 11804 3784 11820 3818
rect 11878 3784 11894 3818
rect 12262 3784 12278 3818
rect 12336 3784 12352 3818
rect 12720 3784 12736 3818
rect 12794 3784 12810 3818
rect 13178 3784 13194 3818
rect 13252 3784 13268 3818
rect 13636 3784 13652 3818
rect 11374 3725 11408 3741
rect 11374 1733 11408 1749
rect 11832 3725 11866 3741
rect 11832 1733 11866 1749
rect 12290 3725 12324 3741
rect 12290 1733 12324 1749
rect 12748 3725 12782 3741
rect 12748 1733 12782 1749
rect 13206 3725 13240 3741
rect 13206 1733 13240 1749
rect 13664 3725 13698 3741
rect 13664 1733 13698 1749
rect 11420 1656 11436 1690
rect 11804 1656 11820 1690
rect 11878 1656 11894 1690
rect 12262 1656 12278 1690
rect 12336 1656 12352 1690
rect 12720 1656 12736 1690
rect 12794 1656 12810 1690
rect 13178 1656 13194 1690
rect 13252 1656 13268 1690
rect 13636 1656 13652 1690
rect 11260 1588 11294 1650
rect 14094 3824 14128 3886
rect 13892 3725 13926 3741
rect 13892 1733 13926 1749
rect 13980 3725 14014 3741
rect 13980 1733 14014 1749
rect 13920 1656 13936 1690
rect 13970 1656 13986 1690
rect 13778 1588 13812 1650
rect 14410 3824 14444 3886
rect 14208 3725 14242 3741
rect 14208 1733 14242 1749
rect 14296 3725 14330 3741
rect 14296 1733 14330 1749
rect 14236 1656 14252 1690
rect 14286 1656 14302 1690
rect 14094 1588 14128 1650
rect 14410 1588 14444 1650
rect 11260 1554 11356 1588
rect 13716 1554 13874 1588
rect 14032 1554 14190 1588
rect 14348 1554 14444 1588
rect 1767 1433 1796 1467
rect 1830 1433 1888 1467
rect 1922 1433 1980 1467
rect 2014 1433 2072 1467
rect 2106 1433 2164 1467
rect 2198 1433 2256 1467
rect 2290 1433 2348 1467
rect 2382 1433 2440 1467
rect 2474 1433 2532 1467
rect 2566 1433 2624 1467
rect 2658 1433 2716 1467
rect 2750 1433 2808 1467
rect 2842 1433 2871 1467
rect 3209 1458 3269 1529
rect 1784 1362 1842 1433
rect 1784 1328 1796 1362
rect 1830 1328 1842 1362
rect 1784 1269 1842 1328
rect 1784 1235 1796 1269
rect 1830 1235 1842 1269
rect 1784 1200 1842 1235
rect 1876 1393 2026 1399
rect 1876 1223 1899 1393
rect 2007 1223 2026 1393
rect 1876 1158 2026 1223
rect 2060 1362 2118 1433
rect 2060 1328 2072 1362
rect 2106 1328 2118 1362
rect 2060 1269 2118 1328
rect 2060 1235 2072 1269
rect 2106 1235 2118 1269
rect 2060 1200 2118 1235
rect 2152 1362 2210 1433
rect 2152 1328 2164 1362
rect 2198 1328 2210 1362
rect 2152 1269 2210 1328
rect 2152 1235 2164 1269
rect 2198 1235 2210 1269
rect 2152 1200 2210 1235
rect 2244 1393 2394 1399
rect 2244 1223 2267 1393
rect 2375 1223 2394 1393
rect 1876 1118 1891 1158
rect 2011 1118 2026 1158
rect 1784 1051 1842 1068
rect 1784 1017 1796 1051
rect 1830 1017 1842 1051
rect 1784 923 1842 1017
rect 1876 1065 2026 1118
rect 2244 1158 2394 1223
rect 2428 1362 2486 1433
rect 2428 1328 2440 1362
rect 2474 1328 2486 1362
rect 2428 1269 2486 1328
rect 2428 1235 2440 1269
rect 2474 1235 2486 1269
rect 2428 1200 2486 1235
rect 2520 1362 2578 1433
rect 2520 1328 2532 1362
rect 2566 1328 2578 1362
rect 2520 1269 2578 1328
rect 2520 1235 2532 1269
rect 2566 1235 2578 1269
rect 2520 1200 2578 1235
rect 2612 1393 2762 1399
rect 2612 1223 2635 1393
rect 2743 1223 2762 1393
rect 2244 1118 2259 1158
rect 2379 1118 2394 1158
rect 1876 963 1899 1065
rect 2008 963 2026 1065
rect 1876 957 2026 963
rect 2060 1051 2118 1068
rect 2060 1017 2072 1051
rect 2106 1017 2118 1051
rect 2060 923 2118 1017
rect 2152 1051 2210 1068
rect 2152 1017 2164 1051
rect 2198 1017 2210 1051
rect 2152 923 2210 1017
rect 2244 1065 2394 1118
rect 2612 1158 2762 1223
rect 2796 1362 2854 1433
rect 2796 1328 2808 1362
rect 2842 1328 2854 1362
rect 2796 1269 2854 1328
rect 3209 1424 3222 1458
rect 3256 1424 3269 1458
rect 3209 1372 3269 1424
rect 3209 1338 3222 1372
rect 3256 1338 3269 1372
rect 3209 1321 3269 1338
rect 2796 1235 2808 1269
rect 2842 1235 2854 1269
rect 2796 1200 2854 1235
rect 3306 1236 3460 1493
rect 3576 1460 3642 1529
rect 3576 1426 3592 1460
rect 3626 1426 3642 1460
rect 3576 1390 3642 1426
rect 3576 1356 3592 1390
rect 3626 1356 3642 1390
rect 3576 1320 3642 1356
rect 3576 1286 3592 1320
rect 3626 1286 3642 1320
rect 3576 1270 3642 1286
rect 3676 1460 3742 1476
rect 3676 1426 3692 1460
rect 3726 1426 3742 1460
rect 3676 1377 3742 1426
rect 3676 1343 3692 1377
rect 3726 1343 3742 1377
rect 3676 1294 3742 1343
rect 4940 1460 5006 1529
rect 4940 1426 4956 1460
rect 4990 1426 5006 1460
rect 4940 1377 5006 1426
rect 4940 1343 4956 1377
rect 4990 1343 5006 1377
rect 3676 1260 3692 1294
rect 3726 1260 3742 1294
rect 2612 1118 2627 1158
rect 2747 1118 2762 1158
rect 2244 963 2267 1065
rect 2376 963 2394 1065
rect 2244 957 2394 963
rect 2428 1051 2486 1068
rect 2428 1017 2440 1051
rect 2474 1017 2486 1051
rect 2428 923 2486 1017
rect 2520 1051 2578 1068
rect 2520 1017 2532 1051
rect 2566 1017 2578 1051
rect 2520 923 2578 1017
rect 2612 1065 2762 1118
rect 3306 1190 3642 1236
rect 3306 1156 3520 1190
rect 3558 1156 3592 1190
rect 3626 1156 3642 1190
rect 3306 1140 3642 1156
rect 3676 1207 3742 1260
rect 3676 1148 3843 1207
rect 3306 1122 3460 1140
rect 3209 1085 3269 1101
rect 2612 963 2635 1065
rect 2744 963 2762 1065
rect 2612 957 2762 963
rect 2796 1051 2854 1068
rect 2796 1017 2808 1051
rect 2842 1017 2854 1051
rect 2796 923 2854 1017
rect 3209 1051 3222 1085
rect 3256 1051 3269 1085
rect 3209 1002 3269 1051
rect 3209 968 3222 1002
rect 3256 968 3269 1002
rect 1767 889 1796 923
rect 1830 889 1888 923
rect 1922 889 1980 923
rect 2014 889 2072 923
rect 2106 889 2164 923
rect 2198 889 2256 923
rect 2290 889 2348 923
rect 2382 889 2440 923
rect 2474 889 2532 923
rect 2566 889 2624 923
rect 2658 889 2716 923
rect 2750 889 2808 923
rect 2842 889 2871 923
rect 3209 897 3269 968
rect 3306 1088 3326 1122
rect 3360 1088 3406 1122
rect 3440 1088 3460 1122
rect 3306 1054 3460 1088
rect 3306 1020 3326 1054
rect 3360 1020 3406 1054
rect 3440 1020 3460 1054
rect 3306 986 3460 1020
rect 3306 952 3326 986
rect 3360 952 3406 986
rect 3440 952 3460 986
rect 3306 933 3460 952
rect 3576 1090 3642 1106
rect 3576 1056 3592 1090
rect 3626 1056 3642 1090
rect 3576 1000 3642 1056
rect 3576 966 3592 1000
rect 3626 966 3642 1000
rect 3576 897 3642 966
rect 3676 1090 3742 1148
rect 3676 1056 3692 1090
rect 3726 1056 3742 1090
rect 3676 1000 3742 1056
rect 4940 1294 5006 1343
rect 4940 1260 4956 1294
rect 4990 1260 5006 1294
rect 4940 1244 5006 1260
rect 5040 1460 5086 1476
rect 5040 1426 5046 1460
rect 5080 1426 5086 1460
rect 5040 1377 5086 1426
rect 5040 1343 5046 1377
rect 5080 1343 5086 1377
rect 5040 1294 5086 1343
rect 5040 1260 5046 1294
rect 5080 1260 5086 1294
rect 4807 1174 5006 1190
rect 4807 1140 4956 1174
rect 4990 1140 5006 1174
rect 4807 1124 5006 1140
rect 4940 1116 5006 1124
rect 5040 1116 5086 1260
rect 5120 1460 5186 1529
rect 5120 1426 5136 1460
rect 5170 1426 5186 1460
rect 5120 1377 5186 1426
rect 5120 1343 5136 1377
rect 5170 1343 5186 1377
rect 5120 1294 5186 1343
rect 5225 1458 5381 1493
rect 5225 1424 5238 1458
rect 5272 1424 5334 1458
rect 5225 1418 5334 1424
rect 5368 1418 5381 1458
rect 5225 1372 5381 1418
rect 5225 1338 5238 1372
rect 5272 1338 5334 1372
rect 5368 1338 5381 1372
rect 5422 1460 5472 1476
rect 5422 1426 5438 1460
rect 5422 1391 5472 1426
rect 5512 1459 5578 1529
rect 5512 1425 5528 1459
rect 5562 1425 5578 1459
rect 5512 1409 5578 1425
rect 5612 1461 5836 1495
rect 5422 1357 5438 1391
rect 5612 1375 5646 1461
rect 5770 1460 5836 1461
rect 5472 1357 5646 1375
rect 5422 1341 5646 1357
rect 5680 1400 5730 1427
rect 5680 1366 5696 1400
rect 5680 1340 5730 1366
rect 5770 1426 5786 1460
rect 5820 1426 5836 1460
rect 5770 1390 5836 1426
rect 5770 1356 5786 1390
rect 5820 1356 5836 1390
rect 5770 1340 5836 1356
rect 5882 1460 5948 1529
rect 5882 1426 5898 1460
rect 5932 1426 5948 1460
rect 5882 1390 5948 1426
rect 5882 1356 5898 1390
rect 5932 1356 5948 1390
rect 5882 1340 5948 1356
rect 5988 1460 6038 1476
rect 6022 1426 6038 1460
rect 5988 1390 6038 1426
rect 6022 1356 6038 1390
rect 5225 1322 5381 1338
rect 5120 1260 5136 1294
rect 5170 1260 5186 1294
rect 5120 1244 5186 1260
rect 5424 1291 5509 1307
rect 5424 1257 5459 1291
rect 5493 1257 5509 1291
rect 5696 1306 5730 1340
rect 5696 1272 5830 1306
rect 5424 1223 5509 1257
rect 5120 1174 5186 1190
rect 5120 1140 5136 1174
rect 5170 1140 5186 1174
rect 5120 1116 5186 1140
rect 5424 1189 5459 1223
rect 5493 1189 5509 1223
rect 5424 1172 5509 1189
rect 5560 1223 5662 1239
rect 5560 1189 5576 1223
rect 5610 1189 5662 1223
rect 5560 1172 5662 1189
rect 5696 1222 5762 1238
rect 5696 1188 5712 1222
rect 5746 1188 5762 1222
rect 5696 1172 5762 1188
rect 5424 1155 5662 1172
rect 5424 1121 5459 1155
rect 5493 1121 5576 1155
rect 5610 1121 5662 1155
rect 5796 1138 5830 1272
rect 5988 1242 6038 1356
rect 6084 1460 6134 1476
rect 6084 1426 6100 1460
rect 6084 1390 6134 1426
rect 6084 1356 6100 1390
rect 6084 1320 6134 1356
rect 6174 1460 6240 1529
rect 6174 1426 6190 1460
rect 6224 1426 6240 1460
rect 6174 1382 6240 1426
rect 6174 1348 6190 1382
rect 6224 1348 6240 1382
rect 6174 1338 6240 1348
rect 6280 1460 6356 1476
rect 6314 1426 6356 1460
rect 6280 1379 6356 1426
rect 6314 1345 6356 1379
rect 6392 1408 6442 1529
rect 6426 1374 6442 1408
rect 6392 1350 6442 1374
rect 6476 1461 6964 1495
rect 6084 1286 6100 1320
rect 6134 1286 6246 1304
rect 6084 1270 6246 1286
rect 5920 1226 6038 1242
rect 5920 1192 5936 1226
rect 5970 1192 6038 1226
rect 5920 1176 6038 1192
rect 5052 1082 5086 1116
rect 5424 1105 5662 1121
rect 5225 1085 5381 1101
rect 4945 1048 4961 1082
rect 4995 1048 5011 1082
rect 5052 1048 5125 1082
rect 5159 1048 5175 1082
rect 3676 966 3692 1000
rect 3726 966 3742 1000
rect 3676 950 3742 966
rect 4945 1000 5011 1048
rect 4945 966 4961 1000
rect 4995 966 5011 1000
rect 4945 897 5011 966
rect 5109 1006 5175 1048
rect 5109 1000 5126 1006
rect 5109 966 5125 1000
rect 5160 972 5175 1006
rect 5159 966 5175 972
rect 5109 950 5175 966
rect 5225 1051 5238 1085
rect 5272 1051 5334 1085
rect 5368 1051 5381 1085
rect 5225 1008 5381 1051
rect 5225 968 5238 1008
rect 5272 1002 5381 1008
rect 5272 968 5334 1002
rect 5368 968 5381 1002
rect 5225 933 5381 968
rect 5427 1050 5493 1105
rect 5696 1104 5953 1138
rect 5696 1071 5737 1104
rect 5427 1016 5443 1050
rect 5477 1016 5493 1050
rect 5427 897 5493 1016
rect 5591 1055 5737 1071
rect 5591 1021 5607 1055
rect 5641 1021 5687 1055
rect 5721 1021 5737 1055
rect 5591 1005 5737 1021
rect 5835 1049 5885 1070
rect 5835 1015 5851 1049
rect 5835 897 5885 1015
rect 5919 965 5953 1104
rect 5987 1060 6038 1176
rect 6096 1200 6178 1236
rect 6096 1166 6128 1200
rect 6162 1166 6178 1200
rect 6096 1150 6178 1166
rect 6212 1214 6246 1270
rect 6280 1298 6356 1345
rect 6476 1316 6510 1461
rect 6779 1460 6964 1461
rect 6314 1264 6356 1298
rect 6280 1248 6356 1264
rect 6212 1198 6288 1214
rect 6212 1164 6238 1198
rect 6272 1164 6288 1198
rect 6212 1148 6288 1164
rect 6322 1150 6356 1248
rect 6406 1296 6510 1316
rect 6406 1262 6422 1296
rect 6456 1282 6510 1296
rect 6567 1400 6633 1427
rect 6567 1366 6583 1400
rect 6617 1366 6633 1400
rect 6567 1322 6633 1366
rect 6667 1400 6733 1427
rect 6779 1426 6795 1460
rect 6829 1426 6914 1460
rect 6948 1426 7008 1460
rect 6667 1366 6683 1400
rect 6717 1390 6733 1400
rect 6717 1366 6940 1390
rect 6667 1356 6940 1366
rect 6567 1288 6872 1322
rect 6456 1262 6472 1282
rect 6406 1246 6472 1262
rect 6806 1255 6872 1288
rect 6698 1248 6764 1251
rect 6518 1235 6764 1248
rect 6518 1232 6714 1235
rect 6518 1198 6534 1232
rect 6568 1201 6714 1232
rect 6748 1201 6764 1235
rect 6568 1198 6764 1201
rect 6518 1185 6764 1198
rect 6806 1221 6822 1255
rect 6856 1221 6872 1255
rect 6806 1187 6872 1221
rect 6518 1156 6622 1185
rect 6518 1150 6582 1156
rect 6212 1114 6246 1148
rect 6322 1122 6582 1150
rect 6616 1122 6622 1156
rect 6806 1153 6822 1187
rect 6856 1153 6872 1187
rect 6806 1151 6872 1153
rect 6322 1117 6622 1122
rect 6322 1116 6353 1117
rect 6083 1080 6099 1114
rect 6133 1080 6246 1114
rect 6337 1083 6353 1116
rect 6387 1116 6622 1117
rect 6656 1117 6872 1151
rect 6021 1026 6038 1060
rect 6337 1049 6387 1083
rect 5987 999 6038 1026
rect 6072 1012 6303 1046
rect 6072 965 6106 1012
rect 5919 931 6106 965
rect 6185 962 6235 978
rect 6185 928 6201 962
rect 6269 965 6303 1012
rect 6337 1015 6353 1049
rect 6337 999 6387 1015
rect 6421 1048 6622 1082
rect 6421 965 6455 1048
rect 6269 931 6455 965
rect 6489 998 6543 1014
rect 6489 964 6491 998
rect 6525 964 6543 998
rect 6185 897 6235 928
rect 6489 897 6543 964
rect 6588 967 6622 1048
rect 6656 1064 6722 1117
rect 6906 1083 6940 1356
rect 6656 1030 6672 1064
rect 6706 1030 6722 1064
rect 6656 1001 6722 1030
rect 6756 1059 6940 1083
rect 6974 1339 7008 1426
rect 7072 1423 7138 1529
rect 7072 1389 7088 1423
rect 7122 1389 7138 1423
rect 7072 1373 7138 1389
rect 7180 1460 7246 1476
rect 7180 1426 7196 1460
rect 7230 1426 7246 1460
rect 7180 1350 7246 1426
rect 7180 1339 7196 1350
rect 6974 1316 7196 1339
rect 7230 1316 7246 1350
rect 7292 1460 7358 1529
rect 7292 1426 7308 1460
rect 7342 1426 7358 1460
rect 7292 1388 7358 1426
rect 7292 1354 7308 1388
rect 7342 1354 7358 1388
rect 7292 1338 7358 1354
rect 7460 1460 7526 1476
rect 7460 1426 7476 1460
rect 7510 1426 7526 1460
rect 7460 1350 7526 1426
rect 7645 1455 7711 1529
rect 7645 1421 7661 1455
rect 7695 1421 7711 1455
rect 7645 1400 7711 1421
rect 7760 1460 7826 1476
rect 7760 1426 7776 1460
rect 7810 1426 7826 1460
rect 7760 1382 7826 1426
rect 7860 1455 7926 1529
rect 8255 1499 8433 1529
rect 7860 1421 7876 1455
rect 7910 1421 7926 1455
rect 7860 1400 7926 1421
rect 8036 1460 8086 1476
rect 8036 1426 8052 1460
rect 8255 1465 8271 1499
rect 8305 1465 8383 1499
rect 8417 1465 8433 1499
rect 8255 1449 8433 1465
rect 8036 1415 8086 1426
rect 7760 1366 7776 1382
rect 6974 1305 7246 1316
rect 6974 1103 7008 1305
rect 7180 1304 7246 1305
rect 7460 1316 7476 1350
rect 7510 1334 7526 1350
rect 7615 1348 7776 1366
rect 7810 1366 7826 1382
rect 8036 1381 8330 1415
rect 8036 1366 8086 1381
rect 7810 1348 8086 1366
rect 7615 1342 8086 1348
rect 7615 1340 8052 1342
rect 7510 1316 7581 1334
rect 7042 1255 7123 1271
rect 7180 1270 7388 1304
rect 7460 1300 7581 1316
rect 7042 1221 7058 1255
rect 7092 1221 7123 1255
rect 7322 1246 7388 1270
rect 7042 1187 7123 1221
rect 7042 1153 7058 1187
rect 7092 1153 7123 1187
rect 7157 1230 7288 1236
rect 7157 1220 7254 1230
rect 7157 1186 7173 1220
rect 7207 1196 7254 1220
rect 7322 1212 7338 1246
rect 7372 1212 7388 1246
rect 7547 1264 7581 1300
rect 7615 1306 7631 1340
rect 7665 1332 8052 1340
rect 7665 1306 7681 1332
rect 7615 1298 7681 1306
rect 8036 1308 8052 1332
rect 7715 1264 7932 1298
rect 8036 1292 8086 1308
rect 8120 1331 8214 1347
rect 8120 1297 8164 1331
rect 8198 1297 8214 1331
rect 7322 1196 7388 1212
rect 7430 1215 7496 1231
rect 7547 1230 7749 1264
rect 7898 1258 7932 1264
rect 8120 1281 8214 1297
rect 7207 1186 7288 1196
rect 7157 1170 7288 1186
rect 7430 1181 7446 1215
rect 7480 1196 7496 1215
rect 7480 1183 7676 1196
rect 7480 1181 7626 1183
rect 7042 1137 7123 1153
rect 7089 1136 7123 1137
rect 7430 1156 7626 1181
rect 6974 1069 7055 1103
rect 7089 1102 7344 1136
rect 7430 1122 7446 1156
rect 7480 1149 7626 1156
rect 7660 1149 7676 1183
rect 7480 1136 7676 1149
rect 7480 1122 7496 1136
rect 7430 1116 7496 1122
rect 7710 1102 7744 1230
rect 7790 1196 7830 1230
rect 7898 1224 8072 1258
rect 7790 1174 7864 1196
rect 8006 1190 8022 1224
rect 8056 1190 8072 1224
rect 7790 1140 7806 1174
rect 7840 1140 7864 1174
rect 7790 1116 7864 1140
rect 7898 1174 7964 1190
rect 8006 1174 8072 1190
rect 7898 1140 7914 1174
rect 7948 1140 7964 1174
rect 8120 1147 8154 1281
rect 8188 1233 8254 1247
rect 8188 1231 8205 1233
rect 8188 1197 8204 1231
rect 8239 1199 8254 1233
rect 8238 1197 8254 1199
rect 8188 1181 8254 1197
rect 8296 1232 8330 1381
rect 8364 1409 8433 1449
rect 8364 1375 8383 1409
rect 8417 1375 8433 1409
rect 8474 1460 8524 1476
rect 8474 1426 8490 1460
rect 8474 1385 8524 1426
rect 8364 1327 8433 1375
rect 8364 1293 8383 1327
rect 8417 1293 8433 1327
rect 8364 1270 8433 1293
rect 8472 1377 8524 1385
rect 8472 1370 8490 1377
rect 8472 1336 8481 1370
rect 8515 1336 8524 1343
rect 8472 1298 8524 1336
rect 8472 1264 8481 1298
rect 8515 1294 8524 1298
rect 8564 1460 8630 1529
rect 8564 1426 8580 1460
rect 8614 1426 8630 1460
rect 8564 1390 8630 1426
rect 8564 1356 8580 1390
rect 8614 1356 8630 1390
rect 8564 1320 8630 1356
rect 8564 1286 8580 1320
rect 8614 1286 8630 1320
rect 8564 1270 8630 1286
rect 8667 1452 8739 1468
rect 8667 1418 8689 1452
rect 8723 1418 8739 1452
rect 8667 1381 8739 1418
rect 8667 1347 8689 1381
rect 8723 1347 8739 1381
rect 8667 1310 8739 1347
rect 8667 1276 8689 1310
rect 8723 1276 8739 1310
rect 8472 1260 8490 1264
rect 8472 1249 8524 1260
rect 8474 1236 8524 1249
rect 8296 1216 8362 1232
rect 8296 1182 8312 1216
rect 8346 1182 8362 1216
rect 8296 1166 8362 1182
rect 8474 1190 8542 1236
rect 8667 1190 8739 1276
rect 8778 1456 8844 1529
rect 8778 1422 8794 1456
rect 8828 1422 8844 1456
rect 8778 1378 8844 1422
rect 8778 1344 8794 1378
rect 8828 1344 8844 1378
rect 8778 1306 8844 1344
rect 8778 1272 8794 1306
rect 8828 1272 8844 1306
rect 8778 1244 8844 1272
rect 8878 1460 8940 1476
rect 8878 1426 8884 1460
rect 8918 1426 8940 1460
rect 8878 1377 8940 1426
rect 8878 1343 8884 1377
rect 8918 1366 8940 1377
rect 8878 1332 8890 1343
rect 8924 1332 8940 1366
rect 8878 1294 8940 1332
rect 8878 1260 8884 1294
rect 8924 1260 8940 1294
rect 8878 1244 8940 1260
rect 8974 1460 9024 1529
rect 9008 1426 9024 1460
rect 9074 1464 9212 1529
rect 9074 1430 9090 1464
rect 9124 1430 9162 1464
rect 9196 1430 9212 1464
rect 9263 1445 9329 1529
rect 8974 1377 9024 1426
rect 9008 1343 9024 1377
rect 8974 1294 9024 1343
rect 9008 1260 9024 1294
rect 9263 1411 9279 1445
rect 9313 1411 9329 1445
rect 9263 1335 9329 1411
rect 9263 1301 9279 1335
rect 9313 1301 9329 1335
rect 9263 1285 9329 1301
rect 9369 1445 9403 1461
rect 9369 1335 9403 1411
rect 9443 1448 9509 1529
rect 9443 1414 9459 1448
rect 9493 1414 9509 1448
rect 9443 1380 9509 1414
rect 9443 1346 9459 1380
rect 9493 1346 9509 1380
rect 9443 1338 9509 1346
rect 9543 1445 9609 1461
rect 9543 1411 9559 1445
rect 9593 1411 9609 1445
rect 9543 1335 9609 1411
rect 9650 1460 9716 1529
rect 9650 1426 9666 1460
rect 9700 1426 9716 1460
rect 9650 1388 9716 1426
rect 9650 1354 9666 1388
rect 9700 1354 9716 1388
rect 9650 1338 9716 1354
rect 9760 1460 9810 1476
rect 9794 1426 9810 1460
rect 9760 1379 9810 1426
rect 9794 1345 9810 1379
rect 9543 1304 9559 1335
rect 9403 1301 9559 1304
rect 9593 1304 9609 1335
rect 9593 1301 9726 1304
rect 8974 1244 9024 1260
rect 9369 1270 9726 1301
rect 8120 1140 8229 1147
rect 7898 1131 8229 1140
rect 6756 1025 6772 1059
rect 6806 1049 6940 1059
rect 6806 1025 6822 1049
rect 6756 967 6822 1025
rect 6989 1035 7005 1069
rect 7039 1035 7055 1069
rect 6588 933 6822 967
rect 6868 999 6953 1015
rect 6989 1001 7055 1035
rect 7089 1051 7176 1067
rect 7089 1017 7115 1051
rect 7149 1017 7176 1051
rect 7089 1001 7176 1017
rect 7210 1051 7276 1068
rect 7210 1017 7226 1051
rect 7260 1017 7276 1051
rect 6868 965 6893 999
rect 6927 967 6953 999
rect 7089 967 7123 1001
rect 6927 965 7123 967
rect 6868 933 7123 965
rect 7210 897 7276 1017
rect 7310 966 7344 1102
rect 7587 1068 7744 1102
rect 7898 1106 8179 1131
rect 7898 1068 7932 1106
rect 8120 1097 8179 1106
rect 8213 1097 8229 1131
rect 8120 1081 8229 1097
rect 8296 1081 8330 1166
rect 8474 1124 8521 1190
rect 7587 1050 7621 1068
rect 7391 1034 7621 1050
rect 7778 1034 7932 1068
rect 7966 1052 8016 1072
rect 7391 1000 7407 1034
rect 7441 1000 7489 1034
rect 7523 1000 7571 1034
rect 7605 1000 7621 1034
rect 7667 1000 7812 1034
rect 8000 1047 8016 1052
rect 8263 1047 8330 1081
rect 8364 1090 8421 1106
rect 8364 1056 8385 1090
rect 8419 1056 8421 1090
rect 8000 1018 8297 1047
rect 7966 1013 8297 1018
rect 7667 966 7701 1000
rect 7846 966 7871 1000
rect 7905 966 7930 1000
rect 7966 999 8016 1013
rect 8364 1000 8421 1056
rect 7310 932 7701 966
rect 7735 932 7755 966
rect 7789 932 7810 966
rect 7735 897 7810 932
rect 7846 965 7930 966
rect 8052 965 8068 979
rect 7846 945 8068 965
rect 8102 945 8118 979
rect 7846 931 8118 945
rect 8364 966 8385 1000
rect 8419 966 8421 1000
rect 8364 897 8421 966
rect 8455 1090 8521 1124
rect 8667 1174 8872 1190
rect 8667 1140 8822 1174
rect 8856 1140 8872 1174
rect 8667 1124 8872 1140
rect 8455 1056 8471 1090
rect 8505 1056 8521 1090
rect 8455 1000 8521 1056
rect 8455 966 8471 1000
rect 8505 966 8521 1000
rect 8455 950 8521 966
rect 8555 1090 8621 1106
rect 8555 1056 8557 1090
rect 8591 1056 8621 1090
rect 8555 1000 8621 1056
rect 8555 966 8557 1000
rect 8591 966 8621 1000
rect 8667 1094 8733 1124
rect 8667 1060 8683 1094
rect 8717 1060 8733 1094
rect 8906 1090 8940 1244
rect 9369 1136 9403 1270
rect 9452 1221 9518 1236
rect 9452 1220 9469 1221
rect 9452 1186 9468 1220
rect 9503 1187 9518 1221
rect 9502 1186 9518 1187
rect 9452 1170 9518 1186
rect 9552 1223 9652 1236
rect 9552 1214 9657 1223
rect 9552 1180 9594 1214
rect 9628 1199 9657 1214
rect 9552 1165 9602 1180
rect 9636 1171 9657 1199
rect 9692 1215 9726 1270
rect 9760 1299 9810 1345
rect 9850 1460 9900 1529
rect 9884 1426 9900 1460
rect 9850 1367 9900 1426
rect 9884 1333 9900 1367
rect 9850 1317 9900 1333
rect 9940 1460 9994 1476
rect 9974 1426 9994 1460
rect 9940 1379 9994 1426
rect 9974 1345 9994 1379
rect 9794 1283 9810 1299
rect 9940 1299 9994 1345
rect 9794 1265 9940 1283
rect 9974 1265 9994 1299
rect 9760 1249 9994 1265
rect 9692 1199 9902 1215
rect 9636 1165 9652 1171
rect 9552 1149 9652 1165
rect 9692 1165 9716 1199
rect 9750 1165 9784 1199
rect 9818 1165 9852 1199
rect 9886 1165 9902 1199
rect 9936 1207 9994 1249
rect 10030 1460 10080 1529
rect 10064 1426 10080 1460
rect 10030 1377 10080 1426
rect 10064 1343 10080 1377
rect 10030 1294 10080 1343
rect 10121 1458 10181 1529
rect 10692 1482 11188 1554
rect 10121 1424 10134 1458
rect 10168 1424 10181 1458
rect 10121 1372 10181 1424
rect 10121 1338 10134 1372
rect 10168 1338 10181 1372
rect 10121 1321 10181 1338
rect 10344 1448 10440 1482
rect 13716 1448 13874 1482
rect 14032 1448 14190 1482
rect 14348 1448 14444 1482
rect 10344 1386 10378 1448
rect 10064 1260 10080 1294
rect 10030 1244 10080 1260
rect 10180 1240 10280 1260
rect 10180 1225 10200 1240
rect 10123 1207 10200 1225
rect 9936 1190 10200 1207
rect 9692 1149 9902 1165
rect 9944 1167 10200 1190
rect 9262 1115 9328 1131
rect 8667 1026 8733 1060
rect 8667 992 8683 1026
rect 8717 992 8733 1026
rect 8667 988 8733 992
rect 8773 1074 8839 1090
rect 8773 1040 8789 1074
rect 8823 1040 8839 1074
rect 8773 1000 8839 1040
rect 8555 897 8621 966
rect 8773 966 8789 1000
rect 8823 966 8839 1000
rect 8773 897 8839 966
rect 8873 1074 8940 1090
rect 8873 1040 8889 1074
rect 8923 1040 8940 1074
rect 8873 1000 8940 1040
rect 8873 966 8889 1000
rect 8923 966 8940 1000
rect 8873 950 8940 966
rect 8975 1090 9025 1106
rect 9009 1056 9025 1090
rect 8975 1000 9025 1056
rect 9009 966 9025 1000
rect 9262 1081 9278 1115
rect 9312 1081 9328 1115
rect 9369 1119 9504 1136
rect 9369 1102 9454 1119
rect 9262 1045 9328 1081
rect 9438 1085 9454 1102
rect 9488 1085 9504 1119
rect 9944 1115 9994 1167
rect 10123 1160 10200 1167
rect 10260 1160 10280 1240
rect 10123 1145 10280 1160
rect 10180 1140 10280 1145
rect 9262 1011 9278 1045
rect 9312 1011 9328 1045
rect 8975 897 9025 966
rect 9074 962 9090 996
rect 9124 962 9162 996
rect 9196 962 9212 996
rect 9074 897 9212 962
rect 9262 897 9328 1011
rect 9368 1048 9402 1068
rect 9368 965 9402 1014
rect 9438 1041 9504 1085
rect 9438 1007 9454 1041
rect 9488 1007 9504 1041
rect 9438 999 9504 1007
rect 9538 1109 9604 1115
rect 9538 1075 9554 1109
rect 9588 1075 9604 1109
rect 9538 1041 9604 1075
rect 9538 1007 9554 1041
rect 9588 1007 9604 1041
rect 9538 965 9604 1007
rect 9368 931 9604 965
rect 9640 1081 9656 1115
rect 9690 1081 9706 1115
rect 9640 1037 9706 1081
rect 9640 1003 9656 1037
rect 9690 1003 9706 1037
rect 9640 897 9706 1003
rect 9758 1099 9944 1115
rect 9792 1081 9944 1099
rect 9978 1081 9994 1115
rect 9792 1065 9808 1081
rect 9758 1025 9808 1065
rect 9792 991 9808 1025
rect 9758 975 9808 991
rect 9842 1031 9908 1047
rect 9842 997 9858 1031
rect 9892 997 9908 1031
rect 9842 897 9908 997
rect 9944 1025 9994 1081
rect 9978 991 9994 1025
rect 9944 975 9994 991
rect 10030 1115 10080 1131
rect 10064 1081 10080 1115
rect 10030 1025 10080 1081
rect 10064 991 10080 1025
rect 10030 897 10080 991
rect 10121 1085 10181 1101
rect 10121 1051 10134 1085
rect 10168 1051 10181 1085
rect 10121 1002 10181 1051
rect 10121 968 10134 1002
rect 10168 968 10181 1002
rect 10121 897 10181 968
rect 3191 863 3222 897
rect 3256 863 3318 897
rect 3352 863 3414 897
rect 3448 863 3510 897
rect 3544 863 3606 897
rect 3640 863 3702 897
rect 3736 863 3798 897
rect 3832 863 3894 897
rect 3928 863 3990 897
rect 4024 863 4086 897
rect 4120 863 4182 897
rect 4216 863 4278 897
rect 4312 863 4374 897
rect 4408 863 4470 897
rect 4504 863 4566 897
rect 4600 863 4662 897
rect 4696 863 4758 897
rect 4792 863 4854 897
rect 4888 863 4950 897
rect 4984 863 5046 897
rect 5080 863 5142 897
rect 5176 863 5238 897
rect 5272 863 5334 897
rect 5368 863 5430 897
rect 5464 863 5526 897
rect 5560 863 5622 897
rect 5656 863 5718 897
rect 5752 863 5814 897
rect 5848 863 5910 897
rect 5944 863 6006 897
rect 6040 863 6102 897
rect 6136 863 6198 897
rect 6232 863 6294 897
rect 6328 863 6390 897
rect 6424 863 6486 897
rect 6520 863 6582 897
rect 6616 863 6678 897
rect 6712 863 6774 897
rect 6808 863 6870 897
rect 6904 863 6966 897
rect 7000 863 7062 897
rect 7096 863 7158 897
rect 7192 863 7254 897
rect 7288 863 7350 897
rect 7384 863 7446 897
rect 7480 863 7542 897
rect 7576 863 7638 897
rect 7672 863 7734 897
rect 7768 863 7830 897
rect 7864 863 7926 897
rect 7960 863 8022 897
rect 8056 863 8118 897
rect 8152 863 8214 897
rect 8248 863 8310 897
rect 8344 863 8406 897
rect 8440 863 8502 897
rect 8536 863 8598 897
rect 8632 863 8694 897
rect 8728 863 8790 897
rect 8824 863 8886 897
rect 8920 863 8982 897
rect 9016 863 9078 897
rect 9112 863 9174 897
rect 9208 863 9270 897
rect 9304 863 9366 897
rect 9400 863 9462 897
rect 9496 863 9558 897
rect 9592 863 9654 897
rect 9688 863 9750 897
rect 9784 863 9846 897
rect 9880 863 9942 897
rect 9976 863 10038 897
rect 10072 863 10134 897
rect 10168 863 10199 897
rect 3670 722 3800 756
rect 3958 722 4054 756
rect 3670 660 3738 722
rect 3670 104 3704 660
rect 4020 660 4054 722
rect 3818 570 3852 586
rect 3818 178 3852 194
rect 3906 570 3940 586
rect 3906 178 3940 194
rect 3846 110 3862 144
rect 3896 110 3912 144
rect 3670 42 3738 104
rect 13778 1386 13812 1448
rect 10504 1346 10520 1380
rect 10888 1346 10904 1380
rect 10962 1346 10978 1380
rect 11346 1346 11362 1380
rect 11420 1346 11436 1380
rect 11804 1346 11820 1380
rect 11878 1346 11894 1380
rect 12262 1346 12278 1380
rect 12336 1346 12352 1380
rect 12720 1346 12736 1380
rect 12794 1346 12810 1380
rect 13178 1346 13194 1380
rect 13252 1346 13268 1380
rect 13636 1346 13652 1380
rect 10458 1296 10492 1312
rect 10458 304 10492 320
rect 10916 1296 10950 1312
rect 10916 304 10950 320
rect 11374 1296 11408 1312
rect 11374 304 11408 320
rect 11832 1296 11866 1312
rect 11832 304 11866 320
rect 12290 1296 12324 1312
rect 12290 304 12324 320
rect 12748 1296 12782 1312
rect 12748 304 12782 320
rect 13206 1296 13240 1312
rect 13206 304 13240 320
rect 13664 1296 13698 1312
rect 13664 304 13698 320
rect 10504 236 10520 270
rect 10888 236 10904 270
rect 10962 236 10978 270
rect 11346 236 11362 270
rect 11420 236 11436 270
rect 11804 236 11820 270
rect 11878 236 11894 270
rect 12262 236 12278 270
rect 12336 236 12352 270
rect 12720 236 12736 270
rect 12794 236 12810 270
rect 13178 236 13194 270
rect 13252 236 13268 270
rect 13636 236 13652 270
rect 10344 168 10378 230
rect 14094 1386 14128 1448
rect 13920 1346 13936 1380
rect 13970 1346 13986 1380
rect 13892 1296 13926 1312
rect 13892 304 13926 320
rect 13980 1296 14014 1312
rect 13980 304 14014 320
rect 13778 168 13812 230
rect 14410 1386 14444 1448
rect 14236 1346 14252 1380
rect 14286 1346 14302 1380
rect 14208 1296 14242 1312
rect 14208 304 14242 320
rect 14296 1296 14330 1312
rect 14296 304 14330 320
rect 14094 168 14128 230
rect 39160 1175 39260 1210
rect 39160 1141 39329 1175
rect 40361 1141 40457 1175
rect 39160 1079 39267 1141
rect 15366 981 15462 1015
rect 16018 981 16176 1015
rect 16732 981 16890 1015
rect 17446 981 17604 1015
rect 18160 981 18318 1015
rect 18874 981 19032 1015
rect 19588 981 19746 1015
rect 20302 981 20460 1015
rect 21016 981 21174 1015
rect 21730 981 21888 1015
rect 22444 981 22602 1015
rect 23158 981 23316 1015
rect 23872 981 24030 1015
rect 24586 981 24744 1015
rect 25300 981 25458 1015
rect 26014 981 26172 1015
rect 26728 981 26886 1015
rect 27442 981 27600 1015
rect 28156 981 28314 1015
rect 28870 981 29028 1015
rect 29584 981 29742 1015
rect 30298 981 30456 1015
rect 31012 981 31170 1015
rect 31726 981 31884 1015
rect 32440 981 32598 1015
rect 33154 981 33312 1015
rect 33868 981 34026 1015
rect 34582 981 34740 1015
rect 35296 981 35454 1015
rect 36010 981 36168 1015
rect 36724 981 36882 1015
rect 37438 981 37596 1015
rect 38152 981 38310 1015
rect 38866 981 38962 1015
rect 15366 919 15400 981
rect 16080 919 16114 981
rect 15536 867 15552 901
rect 15928 867 15944 901
rect 15978 857 16012 873
rect 15536 779 15552 813
rect 15928 779 15944 813
rect 15978 807 16012 823
rect 15366 699 15400 761
rect 16794 919 16828 981
rect 16250 867 16266 901
rect 16642 867 16658 901
rect 16692 857 16726 873
rect 16250 779 16266 813
rect 16642 779 16658 813
rect 16692 807 16726 823
rect 16080 699 16114 761
rect 17508 919 17542 981
rect 16964 867 16980 901
rect 17356 867 17372 901
rect 17406 857 17440 873
rect 16964 779 16980 813
rect 17356 779 17372 813
rect 17406 807 17440 823
rect 16794 699 16828 761
rect 18222 919 18256 981
rect 17678 867 17694 901
rect 18070 867 18086 901
rect 18120 857 18154 873
rect 17678 779 17694 813
rect 18070 779 18086 813
rect 18120 807 18154 823
rect 17508 699 17542 761
rect 18936 919 18970 981
rect 18392 867 18408 901
rect 18784 867 18800 901
rect 18834 857 18868 873
rect 18392 779 18408 813
rect 18784 779 18800 813
rect 18834 807 18868 823
rect 18222 699 18256 761
rect 19650 919 19684 981
rect 19106 867 19122 901
rect 19498 867 19514 901
rect 19548 857 19582 873
rect 19106 779 19122 813
rect 19498 779 19514 813
rect 19548 807 19582 823
rect 18936 699 18970 761
rect 20364 919 20398 981
rect 19820 867 19836 901
rect 20212 867 20228 901
rect 20262 857 20296 873
rect 19820 779 19836 813
rect 20212 779 20228 813
rect 20262 807 20296 823
rect 19650 699 19684 761
rect 21078 919 21112 981
rect 20534 867 20550 901
rect 20926 867 20942 901
rect 20976 857 21010 873
rect 20534 779 20550 813
rect 20926 779 20942 813
rect 20976 807 21010 823
rect 20364 699 20398 761
rect 21792 919 21826 981
rect 21248 867 21264 901
rect 21640 867 21656 901
rect 21690 857 21724 873
rect 21248 779 21264 813
rect 21640 779 21656 813
rect 21690 807 21724 823
rect 21078 699 21112 761
rect 22506 919 22540 981
rect 21962 867 21978 901
rect 22354 867 22370 901
rect 22404 857 22438 873
rect 21962 779 21978 813
rect 22354 779 22370 813
rect 22404 807 22438 823
rect 21792 699 21826 761
rect 23220 919 23254 981
rect 22676 867 22692 901
rect 23068 867 23084 901
rect 23118 857 23152 873
rect 22676 779 22692 813
rect 23068 779 23084 813
rect 23118 807 23152 823
rect 22506 699 22540 761
rect 23934 919 23968 981
rect 23390 867 23406 901
rect 23782 867 23798 901
rect 23832 857 23866 873
rect 23390 779 23406 813
rect 23782 779 23798 813
rect 23832 807 23866 823
rect 23220 699 23254 761
rect 24648 919 24682 981
rect 24104 867 24120 901
rect 24496 867 24512 901
rect 24546 857 24580 873
rect 24104 779 24120 813
rect 24496 779 24512 813
rect 24546 807 24580 823
rect 23934 699 23968 761
rect 25362 919 25396 981
rect 24818 867 24834 901
rect 25210 867 25226 901
rect 25260 857 25294 873
rect 24818 779 24834 813
rect 25210 779 25226 813
rect 25260 807 25294 823
rect 24648 699 24682 761
rect 26076 919 26110 981
rect 25532 867 25548 901
rect 25924 867 25940 901
rect 25974 857 26008 873
rect 25532 779 25548 813
rect 25924 779 25940 813
rect 25974 807 26008 823
rect 25362 699 25396 761
rect 26790 919 26824 981
rect 26246 867 26262 901
rect 26638 867 26654 901
rect 26688 857 26722 873
rect 26246 779 26262 813
rect 26638 779 26654 813
rect 26688 807 26722 823
rect 26076 699 26110 761
rect 27504 919 27538 981
rect 26960 867 26976 901
rect 27352 867 27368 901
rect 27402 857 27436 873
rect 26960 779 26976 813
rect 27352 779 27368 813
rect 27402 807 27436 823
rect 26790 699 26824 761
rect 28218 919 28252 981
rect 27674 867 27690 901
rect 28066 867 28082 901
rect 28116 857 28150 873
rect 27674 779 27690 813
rect 28066 779 28082 813
rect 28116 807 28150 823
rect 27504 699 27538 761
rect 28932 919 28966 981
rect 28388 867 28404 901
rect 28780 867 28796 901
rect 28830 857 28864 873
rect 28388 779 28404 813
rect 28780 779 28796 813
rect 28830 807 28864 823
rect 28218 699 28252 761
rect 29646 919 29680 981
rect 29102 867 29118 901
rect 29494 867 29510 901
rect 29544 857 29578 873
rect 29102 779 29118 813
rect 29494 779 29510 813
rect 29544 807 29578 823
rect 28932 699 28966 761
rect 30360 919 30394 981
rect 29816 867 29832 901
rect 30208 867 30224 901
rect 30258 857 30292 873
rect 29816 779 29832 813
rect 30208 779 30224 813
rect 30258 807 30292 823
rect 29646 699 29680 761
rect 31074 919 31108 981
rect 30530 867 30546 901
rect 30922 867 30938 901
rect 30972 857 31006 873
rect 30530 779 30546 813
rect 30922 779 30938 813
rect 30972 807 31006 823
rect 30360 699 30394 761
rect 31788 919 31822 981
rect 31244 867 31260 901
rect 31636 867 31652 901
rect 31686 857 31720 873
rect 31244 779 31260 813
rect 31636 779 31652 813
rect 31686 807 31720 823
rect 31074 699 31108 761
rect 32502 919 32536 981
rect 31958 867 31974 901
rect 32350 867 32366 901
rect 32400 857 32434 873
rect 31958 779 31974 813
rect 32350 779 32366 813
rect 32400 807 32434 823
rect 31788 699 31822 761
rect 33216 919 33250 981
rect 32672 867 32688 901
rect 33064 867 33080 901
rect 33114 857 33148 873
rect 32672 779 32688 813
rect 33064 779 33080 813
rect 33114 807 33148 823
rect 32502 699 32536 761
rect 33930 919 33964 981
rect 33386 867 33402 901
rect 33778 867 33794 901
rect 33828 857 33862 873
rect 33386 779 33402 813
rect 33778 779 33794 813
rect 33828 807 33862 823
rect 33216 699 33250 761
rect 34644 919 34678 981
rect 34100 867 34116 901
rect 34492 867 34508 901
rect 34542 857 34576 873
rect 34100 779 34116 813
rect 34492 779 34508 813
rect 34542 807 34576 823
rect 33930 699 33964 761
rect 35358 919 35392 981
rect 34814 867 34830 901
rect 35206 867 35222 901
rect 35256 857 35290 873
rect 34814 779 34830 813
rect 35206 779 35222 813
rect 35256 807 35290 823
rect 34644 699 34678 761
rect 36072 919 36106 981
rect 35528 867 35544 901
rect 35920 867 35936 901
rect 35970 857 36004 873
rect 35528 779 35544 813
rect 35920 779 35936 813
rect 35970 807 36004 823
rect 35358 699 35392 761
rect 36786 919 36820 981
rect 36242 867 36258 901
rect 36634 867 36650 901
rect 36684 857 36718 873
rect 36242 779 36258 813
rect 36634 779 36650 813
rect 36684 807 36718 823
rect 36072 699 36106 761
rect 37500 919 37534 981
rect 36956 867 36972 901
rect 37348 867 37364 901
rect 37398 857 37432 873
rect 36956 779 36972 813
rect 37348 779 37364 813
rect 37398 807 37432 823
rect 36786 699 36820 761
rect 38214 919 38248 981
rect 37670 867 37686 901
rect 38062 867 38078 901
rect 38112 857 38146 873
rect 37670 779 37686 813
rect 38062 779 38078 813
rect 38112 807 38146 823
rect 37500 699 37534 761
rect 38928 919 38962 981
rect 38384 867 38400 901
rect 38776 867 38792 901
rect 38826 857 38860 873
rect 38384 779 38400 813
rect 38776 779 38792 813
rect 38826 807 38860 823
rect 38214 699 38248 761
rect 38928 699 38962 761
rect 15366 665 15462 699
rect 16018 665 16176 699
rect 16732 665 16890 699
rect 17446 665 17604 699
rect 18160 665 18318 699
rect 18874 665 19032 699
rect 19588 665 19746 699
rect 20302 665 20460 699
rect 21016 665 21174 699
rect 21730 665 21888 699
rect 22444 665 22602 699
rect 23158 665 23316 699
rect 23872 665 24030 699
rect 24586 665 24744 699
rect 25300 665 25458 699
rect 26014 665 26172 699
rect 26728 665 26886 699
rect 27442 665 27600 699
rect 28156 665 28314 699
rect 28870 665 29028 699
rect 29584 665 29742 699
rect 30298 665 30456 699
rect 31012 665 31170 699
rect 31726 665 31884 699
rect 32440 665 32598 699
rect 33154 665 33312 699
rect 33868 665 34026 699
rect 34582 665 34740 699
rect 35296 665 35454 699
rect 36010 665 36168 699
rect 36724 665 36882 699
rect 37438 665 37596 699
rect 38152 665 38310 699
rect 38866 665 38962 699
rect 15366 631 38962 665
rect 39160 470 39233 1079
rect 40423 1079 40457 1141
rect 39160 380 39170 470
rect 14410 168 14444 230
rect 15366 197 38962 231
rect 10344 158 10440 168
rect 13716 158 13874 168
rect 14032 158 14190 168
rect 14348 158 14448 168
rect 10344 138 10358 158
rect 4020 42 4054 104
rect 10338 78 10358 138
rect 14428 78 14448 158
rect 10338 68 14448 78
rect 15366 163 15462 197
rect 16018 163 16176 197
rect 16732 163 16890 197
rect 17446 163 17604 197
rect 18160 163 18318 197
rect 18874 163 19032 197
rect 19588 163 19746 197
rect 20302 163 20460 197
rect 21016 163 21174 197
rect 21730 163 21888 197
rect 22444 163 22602 197
rect 23158 163 23316 197
rect 23872 163 24030 197
rect 24586 163 24744 197
rect 25300 163 25458 197
rect 26014 163 26172 197
rect 26728 163 26886 197
rect 27442 163 27600 197
rect 28156 163 28314 197
rect 28870 163 29028 197
rect 29584 163 29742 197
rect 30298 163 30456 197
rect 31012 163 31170 197
rect 31726 163 31884 197
rect 32440 163 32598 197
rect 33154 163 33312 197
rect 33868 163 34026 197
rect 34582 163 34740 197
rect 35296 163 35454 197
rect 36010 163 36168 197
rect 36724 163 36882 197
rect 37438 163 37596 197
rect 38152 163 38310 197
rect 38866 163 38962 197
rect 15366 101 15400 163
rect 3670 8 3800 42
rect 3958 8 4054 42
rect 3670 -54 3738 8
rect 3670 -610 3704 -54
rect 4020 -54 4054 8
rect 3818 -144 3852 -128
rect 3818 -536 3852 -520
rect 3906 -144 3940 -128
rect 3906 -536 3940 -520
rect 3846 -604 3862 -570
rect 3896 -604 3912 -570
rect 3670 -672 3738 -610
rect 16080 101 16114 163
rect 15536 49 15552 83
rect 15928 49 15944 83
rect 15978 39 16012 55
rect 15536 -39 15552 -5
rect 15928 -39 15944 -5
rect 15978 -11 16012 5
rect 15366 -119 15400 -57
rect 16794 101 16828 163
rect 16250 49 16266 83
rect 16642 49 16658 83
rect 16692 39 16726 55
rect 16250 -39 16266 -5
rect 16642 -39 16658 -5
rect 16692 -11 16726 5
rect 16080 -119 16114 -57
rect 17508 101 17542 163
rect 16964 49 16980 83
rect 17356 49 17372 83
rect 17406 39 17440 55
rect 16964 -39 16980 -5
rect 17356 -39 17372 -5
rect 17406 -11 17440 5
rect 16794 -119 16828 -57
rect 18222 101 18256 163
rect 17678 49 17694 83
rect 18070 49 18086 83
rect 18120 39 18154 55
rect 17678 -39 17694 -5
rect 18070 -39 18086 -5
rect 18120 -11 18154 5
rect 17508 -119 17542 -57
rect 18936 101 18970 163
rect 18392 49 18408 83
rect 18784 49 18800 83
rect 18834 39 18868 55
rect 18392 -39 18408 -5
rect 18784 -39 18800 -5
rect 18834 -11 18868 5
rect 18222 -119 18256 -57
rect 19650 101 19684 163
rect 19106 49 19122 83
rect 19498 49 19514 83
rect 19548 39 19582 55
rect 19106 -39 19122 -5
rect 19498 -39 19514 -5
rect 19548 -11 19582 5
rect 18936 -119 18970 -57
rect 20364 101 20398 163
rect 19820 49 19836 83
rect 20212 49 20228 83
rect 20262 39 20296 55
rect 19820 -39 19836 -5
rect 20212 -39 20228 -5
rect 20262 -11 20296 5
rect 19650 -119 19684 -57
rect 21078 101 21112 163
rect 20534 49 20550 83
rect 20926 49 20942 83
rect 20976 39 21010 55
rect 20534 -39 20550 -5
rect 20926 -39 20942 -5
rect 20976 -11 21010 5
rect 20364 -119 20398 -57
rect 21792 101 21826 163
rect 21248 49 21264 83
rect 21640 49 21656 83
rect 21690 39 21724 55
rect 21248 -39 21264 -5
rect 21640 -39 21656 -5
rect 21690 -11 21724 5
rect 21078 -119 21112 -57
rect 22506 101 22540 163
rect 21962 49 21978 83
rect 22354 49 22370 83
rect 22404 39 22438 55
rect 21962 -39 21978 -5
rect 22354 -39 22370 -5
rect 22404 -11 22438 5
rect 21792 -119 21826 -57
rect 23220 101 23254 163
rect 22676 49 22692 83
rect 23068 49 23084 83
rect 23118 39 23152 55
rect 22676 -39 22692 -5
rect 23068 -39 23084 -5
rect 23118 -11 23152 5
rect 22506 -119 22540 -57
rect 23934 101 23968 163
rect 23390 49 23406 83
rect 23782 49 23798 83
rect 23832 39 23866 55
rect 23390 -39 23406 -5
rect 23782 -39 23798 -5
rect 23832 -11 23866 5
rect 23220 -119 23254 -57
rect 24648 101 24682 163
rect 24104 49 24120 83
rect 24496 49 24512 83
rect 24546 39 24580 55
rect 24104 -39 24120 -5
rect 24496 -39 24512 -5
rect 24546 -11 24580 5
rect 23934 -119 23968 -57
rect 25362 101 25396 163
rect 24818 49 24834 83
rect 25210 49 25226 83
rect 25260 39 25294 55
rect 24818 -39 24834 -5
rect 25210 -39 25226 -5
rect 25260 -11 25294 5
rect 24648 -119 24682 -57
rect 26076 101 26110 163
rect 25532 49 25548 83
rect 25924 49 25940 83
rect 25974 39 26008 55
rect 25532 -39 25548 -5
rect 25924 -39 25940 -5
rect 25974 -11 26008 5
rect 25362 -119 25396 -57
rect 26790 101 26824 163
rect 26246 49 26262 83
rect 26638 49 26654 83
rect 26688 39 26722 55
rect 26246 -39 26262 -5
rect 26638 -39 26654 -5
rect 26688 -11 26722 5
rect 26076 -119 26110 -57
rect 27504 101 27538 163
rect 26960 49 26976 83
rect 27352 49 27368 83
rect 27402 39 27436 55
rect 26960 -39 26976 -5
rect 27352 -39 27368 -5
rect 27402 -11 27436 5
rect 26790 -119 26824 -57
rect 28218 101 28252 163
rect 27674 49 27690 83
rect 28066 49 28082 83
rect 28116 39 28150 55
rect 27674 -39 27690 -5
rect 28066 -39 28082 -5
rect 28116 -11 28150 5
rect 27504 -119 27538 -57
rect 28932 101 28966 163
rect 28388 49 28404 83
rect 28780 49 28796 83
rect 28830 39 28864 55
rect 28388 -39 28404 -5
rect 28780 -39 28796 -5
rect 28830 -11 28864 5
rect 28218 -119 28252 -57
rect 29646 101 29680 163
rect 29102 49 29118 83
rect 29494 49 29510 83
rect 29544 39 29578 55
rect 29102 -39 29118 -5
rect 29494 -39 29510 -5
rect 29544 -11 29578 5
rect 28932 -119 28966 -57
rect 30360 101 30394 163
rect 29816 49 29832 83
rect 30208 49 30224 83
rect 30258 39 30292 55
rect 29816 -39 29832 -5
rect 30208 -39 30224 -5
rect 30258 -11 30292 5
rect 29646 -119 29680 -57
rect 31074 101 31108 163
rect 30530 49 30546 83
rect 30922 49 30938 83
rect 30972 39 31006 55
rect 30530 -39 30546 -5
rect 30922 -39 30938 -5
rect 30972 -11 31006 5
rect 30360 -119 30394 -57
rect 31788 101 31822 163
rect 31244 49 31260 83
rect 31636 49 31652 83
rect 31686 39 31720 55
rect 31244 -39 31260 -5
rect 31636 -39 31652 -5
rect 31686 -11 31720 5
rect 31074 -119 31108 -57
rect 32502 101 32536 163
rect 31958 49 31974 83
rect 32350 49 32366 83
rect 32400 39 32434 55
rect 31958 -39 31974 -5
rect 32350 -39 32366 -5
rect 32400 -11 32434 5
rect 31788 -119 31822 -57
rect 33216 101 33250 163
rect 32672 49 32688 83
rect 33064 49 33080 83
rect 33114 39 33148 55
rect 32672 -39 32688 -5
rect 33064 -39 33080 -5
rect 33114 -11 33148 5
rect 32502 -119 32536 -57
rect 33930 101 33964 163
rect 33386 49 33402 83
rect 33778 49 33794 83
rect 33828 39 33862 55
rect 33386 -39 33402 -5
rect 33778 -39 33794 -5
rect 33828 -11 33862 5
rect 33216 -119 33250 -57
rect 34644 101 34678 163
rect 34100 49 34116 83
rect 34492 49 34508 83
rect 34542 39 34576 55
rect 34100 -39 34116 -5
rect 34492 -39 34508 -5
rect 34542 -11 34576 5
rect 33930 -119 33964 -57
rect 35358 101 35392 163
rect 34814 49 34830 83
rect 35206 49 35222 83
rect 35256 39 35290 55
rect 34814 -39 34830 -5
rect 35206 -39 35222 -5
rect 35256 -11 35290 5
rect 34644 -119 34678 -57
rect 36072 101 36106 163
rect 35528 49 35544 83
rect 35920 49 35936 83
rect 35970 39 36004 55
rect 35528 -39 35544 -5
rect 35920 -39 35936 -5
rect 35970 -11 36004 5
rect 35358 -119 35392 -57
rect 36786 101 36820 163
rect 36242 49 36258 83
rect 36634 49 36650 83
rect 36684 39 36718 55
rect 36242 -39 36258 -5
rect 36634 -39 36650 -5
rect 36684 -11 36718 5
rect 36072 -119 36106 -57
rect 37500 101 37534 163
rect 36956 49 36972 83
rect 37348 49 37364 83
rect 37398 39 37432 55
rect 36956 -39 36972 -5
rect 37348 -39 37364 -5
rect 37398 -11 37432 5
rect 36786 -119 36820 -57
rect 38214 101 38248 163
rect 37670 49 37686 83
rect 38062 49 38078 83
rect 38112 39 38146 55
rect 37670 -39 37686 -5
rect 38062 -39 38078 -5
rect 38112 -11 38146 5
rect 37500 -119 37534 -57
rect 38928 101 38962 163
rect 38384 49 38400 83
rect 38776 49 38792 83
rect 38826 39 38860 55
rect 38384 -39 38400 -5
rect 38776 -39 38792 -5
rect 38826 -11 38860 5
rect 38214 -119 38248 -57
rect 38928 -119 38962 -57
rect 15366 -153 15462 -119
rect 16018 -153 16176 -119
rect 16732 -153 16890 -119
rect 17446 -153 17604 -119
rect 18160 -153 18318 -119
rect 18874 -153 19032 -119
rect 19588 -153 19746 -119
rect 20302 -153 20460 -119
rect 21016 -153 21174 -119
rect 21730 -153 21888 -119
rect 22444 -153 22602 -119
rect 23158 -153 23316 -119
rect 23872 -153 24030 -119
rect 24586 -153 24744 -119
rect 25300 -153 25458 -119
rect 26014 -153 26172 -119
rect 26728 -153 26886 -119
rect 27442 -153 27600 -119
rect 28156 -153 28314 -119
rect 28870 -153 29028 -119
rect 29584 -153 29742 -119
rect 30298 -153 30456 -119
rect 31012 -153 31170 -119
rect 31726 -153 31884 -119
rect 32440 -153 32598 -119
rect 33154 -153 33312 -119
rect 33868 -153 34026 -119
rect 34582 -153 34740 -119
rect 35296 -153 35454 -119
rect 36010 -153 36168 -119
rect 36724 -153 36882 -119
rect 37438 -153 37596 -119
rect 38152 -153 38310 -119
rect 38866 -153 38962 -119
rect 39160 -221 39233 380
rect 39160 -283 39267 -221
rect 40423 -283 40457 -221
rect 39160 -317 39329 -283
rect 40361 -317 40457 -283
rect 39160 -320 39260 -317
rect 4020 -672 4054 -610
rect 3670 -706 3800 -672
rect 3958 -706 4054 -672
rect 10231 -371 10265 -354
rect 10775 -371 10809 -354
rect 10231 -383 10498 -371
rect 10265 -417 10336 -383
rect 10370 -417 10429 -383
rect 10463 -417 10498 -383
rect 10231 -429 10498 -417
rect 10630 -383 10809 -371
rect 10630 -417 10647 -383
rect 10681 -417 10775 -383
rect 10630 -429 10809 -417
rect 10231 -475 10265 -429
rect 10231 -567 10265 -509
rect 10231 -647 10265 -601
rect 10299 -478 10741 -463
rect 10299 -486 10540 -478
rect 10299 -594 10305 -486
rect 10475 -594 10540 -486
rect 10299 -598 10540 -594
rect 10580 -486 10741 -478
rect 10580 -595 10633 -486
rect 10735 -595 10741 -486
rect 10580 -598 10741 -595
rect 10299 -613 10741 -598
rect 10775 -475 10809 -429
rect 10775 -567 10809 -509
rect 10775 -647 10809 -601
rect 10231 -659 10498 -647
rect 10265 -693 10336 -659
rect 10370 -693 10429 -659
rect 10463 -693 10498 -659
rect 10231 -705 10498 -693
rect 10630 -659 10809 -647
rect 10630 -693 10647 -659
rect 10681 -693 10775 -659
rect 10630 -705 10809 -693
rect 10231 -751 10265 -705
rect 10231 -843 10265 -785
rect 10775 -751 10809 -705
rect 10514 -788 10616 -786
rect 10299 -793 10741 -788
rect 10299 -804 10570 -793
rect 10299 -838 10307 -804
rect 10341 -838 10375 -804
rect 10409 -838 10443 -804
rect 10477 -827 10570 -804
rect 10604 -804 10741 -793
rect 10604 -827 10627 -804
rect 10477 -834 10627 -827
rect 10477 -838 10495 -834
rect 10299 -854 10495 -838
rect 10615 -838 10627 -834
rect 10661 -838 10695 -804
rect 10729 -838 10741 -804
rect 10615 -854 10741 -838
rect 10775 -843 10809 -785
rect 10231 -888 10265 -877
rect 10529 -884 10577 -868
rect 10231 -922 10307 -888
rect 10341 -922 10375 -888
rect 10409 -922 10443 -888
rect 10477 -922 10493 -888
rect 10231 -930 10493 -922
rect 10529 -918 10543 -884
rect 10775 -888 10809 -877
rect 10231 -935 10265 -930
rect 10231 -1015 10265 -969
rect 10529 -980 10577 -918
rect 10611 -922 10627 -888
rect 10661 -922 10695 -888
rect 10729 -922 10809 -888
rect 10611 -934 10809 -922
rect 10231 -1027 10498 -1015
rect 10265 -1061 10336 -1027
rect 10370 -1061 10429 -1027
rect 10463 -1061 10498 -1027
rect 10231 -1073 10498 -1061
rect 10231 -1119 10265 -1073
rect 10540 -1107 10577 -980
rect 10775 -935 10809 -934
rect 10775 -1015 10809 -969
rect 10630 -1027 10809 -1015
rect 10630 -1061 10647 -1027
rect 10681 -1061 10775 -1027
rect 10630 -1073 10809 -1061
rect 10231 -1211 10265 -1153
rect 10231 -1291 10265 -1245
rect 10299 -1122 10741 -1107
rect 10299 -1130 10540 -1122
rect 10299 -1238 10305 -1130
rect 10475 -1238 10540 -1130
rect 10299 -1242 10540 -1238
rect 10580 -1130 10741 -1122
rect 10580 -1239 10633 -1130
rect 10735 -1239 10741 -1130
rect 10580 -1242 10741 -1239
rect 10299 -1257 10741 -1242
rect 10775 -1119 10809 -1073
rect 10775 -1211 10809 -1153
rect 10775 -1291 10809 -1245
rect 10231 -1303 10498 -1291
rect 10265 -1337 10336 -1303
rect 10370 -1337 10429 -1303
rect 10463 -1337 10498 -1303
rect 10231 -1349 10498 -1337
rect 10630 -1303 10809 -1291
rect 10630 -1337 10647 -1303
rect 10681 -1337 10775 -1303
rect 10630 -1349 10809 -1337
rect 10231 -1366 10265 -1349
rect 10775 -1366 10809 -1349
rect 10522 -2940 11560 -2920
rect 6953 -3120 7049 -3086
rect 8951 -3120 9047 -3086
rect 6953 -3182 6987 -3120
rect 9013 -3182 9047 -3120
rect 7113 -3222 7129 -3188
rect 7497 -3222 7513 -3188
rect 7571 -3222 7587 -3188
rect 7955 -3222 7971 -3188
rect 8029 -3222 8045 -3188
rect 8413 -3222 8429 -3188
rect 8487 -3222 8503 -3188
rect 8871 -3222 8887 -3188
rect 5745 -4236 5841 -4202
rect 6619 -4236 6715 -4202
rect 5745 -4298 5779 -4236
rect 6681 -4298 6715 -4236
rect 5902 -4338 5918 -4304
rect 5952 -4338 5968 -4304
rect 6020 -4338 6036 -4304
rect 6070 -4338 6086 -4304
rect 6138 -4338 6154 -4304
rect 6188 -4338 6204 -4304
rect 6256 -4338 6272 -4304
rect 6306 -4338 6322 -4304
rect 6374 -4338 6390 -4304
rect 6424 -4338 6440 -4304
rect 6492 -4338 6508 -4304
rect 6542 -4338 6558 -4304
rect 5042 -4920 5138 -4886
rect 5578 -4920 5674 -4886
rect 5042 -4982 5076 -4920
rect 5640 -4982 5745 -4920
rect 5042 -6148 5076 -6086
rect 5674 -6086 5745 -4982
rect 5640 -6148 5745 -6086
rect 5042 -6182 5138 -6148
rect 5578 -6160 5745 -6148
rect 5578 -6182 5674 -6160
rect 5859 -4388 5893 -4372
rect 5859 -6380 5893 -6364
rect 5977 -4388 6011 -4372
rect 5977 -6380 6011 -6364
rect 6095 -4388 6129 -4372
rect 6095 -6380 6129 -6364
rect 6213 -4388 6247 -4372
rect 6213 -6380 6247 -6364
rect 6331 -4388 6365 -4372
rect 6331 -6380 6365 -6364
rect 6449 -4388 6483 -4372
rect 6449 -6380 6483 -6364
rect 6567 -4388 6601 -4372
rect 6567 -6380 6601 -6364
rect 7067 -3272 7101 -3256
rect 7067 -5264 7101 -5248
rect 7525 -3272 7559 -3256
rect 7525 -5264 7559 -5248
rect 7983 -3272 8017 -3256
rect 7983 -5264 8017 -5248
rect 8441 -3272 8475 -3256
rect 8441 -5264 8475 -5248
rect 8899 -3272 8933 -3256
rect 8899 -5264 8933 -5248
rect 10522 -3860 10542 -2940
rect 10602 -2954 11560 -2940
rect 10602 -2988 10774 -2954
rect 11430 -2988 11560 -2954
rect 10602 -3070 10712 -2988
rect 10602 -3860 10678 -3070
rect 10522 -3880 10678 -3860
rect 10644 -3920 10678 -3880
rect 11492 -3070 11560 -2988
rect 11396 -3139 11435 -3130
rect 11412 -3192 11435 -3139
rect 11396 -3200 11435 -3192
rect 11396 -3366 11435 -3296
rect 11384 -3484 11435 -3366
rect 10848 -3518 10864 -3484
rect 11340 -3518 11435 -3484
rect 10712 -3614 10864 -3580
rect 11340 -3614 11356 -3580
rect 11390 -3610 11424 -3594
rect 11390 -3660 11424 -3644
rect 10848 -3710 10864 -3676
rect 11340 -3710 11356 -3676
rect 10848 -3806 10864 -3772
rect 11340 -3806 11356 -3772
rect 11390 -3802 11424 -3786
rect 11390 -3852 11424 -3836
rect 10848 -3902 10864 -3868
rect 11340 -3902 11356 -3868
rect 10644 -3982 10712 -3920
rect 11526 -3920 11560 -3070
rect 11492 -3982 11560 -3920
rect 10644 -4016 10774 -3982
rect 11430 -4016 11560 -3982
rect 10644 -4050 11560 -4016
rect 7113 -5332 7129 -5298
rect 7497 -5332 7513 -5298
rect 7571 -5332 7587 -5298
rect 7955 -5332 7971 -5298
rect 8029 -5332 8045 -5298
rect 8413 -5332 8429 -5298
rect 8487 -5332 8503 -5298
rect 8871 -5332 8887 -5298
rect 6953 -5400 6987 -5338
rect 9013 -5400 9047 -5338
rect 6953 -5434 7049 -5400
rect 8951 -5434 9047 -5400
rect 9286 -4236 9382 -4202
rect 10160 -4236 10256 -4202
rect 9286 -4298 9320 -4236
rect 10222 -4298 10256 -4236
rect 9443 -4338 9459 -4304
rect 9493 -4338 9509 -4304
rect 9561 -4338 9577 -4304
rect 9611 -4338 9627 -4304
rect 9679 -4338 9695 -4304
rect 9729 -4338 9745 -4304
rect 9797 -4338 9813 -4304
rect 9847 -4338 9863 -4304
rect 9915 -4338 9931 -4304
rect 9965 -4338 9981 -4304
rect 10033 -4338 10049 -4304
rect 10083 -4338 10099 -4304
rect 6909 -5560 7005 -5526
rect 8995 -5560 9091 -5526
rect 6909 -5622 6943 -5560
rect 7295 -5650 7311 -5616
rect 7345 -5650 7361 -5616
rect 7487 -5650 7503 -5616
rect 7537 -5650 7553 -5616
rect 7679 -5650 7695 -5616
rect 7729 -5650 7745 -5616
rect 7871 -5650 7887 -5616
rect 7921 -5650 7937 -5616
rect 8063 -5650 8079 -5616
rect 8113 -5650 8129 -5616
rect 8255 -5650 8271 -5616
rect 8305 -5650 8321 -5616
rect 8447 -5650 8463 -5616
rect 8497 -5650 8513 -5616
rect 8639 -5650 8655 -5616
rect 8689 -5650 8705 -5616
rect 9057 -5622 9091 -5560
rect 7023 -5712 7057 -5696
rect 7023 -6204 7057 -6188
rect 7119 -5712 7153 -5696
rect 7119 -6204 7153 -6188
rect 7215 -5712 7249 -5696
rect 7215 -6204 7249 -6188
rect 7311 -5712 7345 -5696
rect 7311 -6204 7345 -6188
rect 7407 -5712 7441 -5696
rect 7407 -6204 7441 -6188
rect 7503 -5712 7537 -5696
rect 7503 -6204 7537 -6188
rect 7599 -5712 7633 -5696
rect 7599 -6204 7633 -6188
rect 7695 -5712 7729 -5696
rect 7695 -6204 7729 -6188
rect 7791 -5712 7825 -5696
rect 7791 -6204 7825 -6188
rect 7887 -5712 7921 -5696
rect 7887 -6204 7921 -6188
rect 7983 -5712 8017 -5696
rect 7983 -6204 8017 -6188
rect 8079 -5712 8113 -5696
rect 8079 -6204 8113 -6188
rect 8175 -5712 8209 -5696
rect 8175 -6204 8209 -6188
rect 8271 -5712 8305 -5696
rect 8271 -6204 8305 -6188
rect 8367 -5712 8401 -5696
rect 8367 -6204 8401 -6188
rect 8463 -5712 8497 -5696
rect 8463 -6204 8497 -6188
rect 8559 -5712 8593 -5696
rect 8559 -6204 8593 -6188
rect 8655 -5712 8689 -5696
rect 8655 -6204 8689 -6188
rect 8751 -5712 8785 -5696
rect 8751 -6204 8785 -6188
rect 8847 -5712 8881 -5696
rect 8847 -6204 8881 -6188
rect 8943 -5712 8977 -5696
rect 8943 -6204 8977 -6188
rect 7103 -6276 7119 -6242
rect 7153 -6276 7169 -6242
rect 8831 -6276 8847 -6242
rect 8881 -6276 8897 -6242
rect 6909 -6340 6943 -6278
rect 9057 -6340 9091 -6278
rect 6909 -6374 7005 -6340
rect 8995 -6374 9091 -6340
rect 5902 -6448 5918 -6414
rect 5952 -6448 5968 -6414
rect 6020 -6448 6036 -6414
rect 6070 -6448 6086 -6414
rect 6138 -6448 6154 -6414
rect 6188 -6448 6204 -6414
rect 6256 -6448 6272 -6414
rect 6306 -6448 6322 -6414
rect 6374 -6448 6390 -6414
rect 6424 -6448 6440 -6414
rect 6492 -6448 6508 -6414
rect 6542 -6448 6558 -6414
rect 5745 -6516 5779 -6454
rect 6681 -6516 6715 -6454
rect 5745 -6550 5841 -6516
rect 6619 -6550 6715 -6516
rect 9400 -4388 9434 -4372
rect 9400 -6380 9434 -6364
rect 9518 -4388 9552 -4372
rect 9518 -6380 9552 -6364
rect 9636 -4388 9670 -4372
rect 9636 -6380 9670 -6364
rect 9754 -4388 9788 -4372
rect 9754 -6380 9788 -6364
rect 9872 -4388 9906 -4372
rect 9872 -6380 9906 -6364
rect 9990 -4388 10024 -4372
rect 9990 -6380 10024 -6364
rect 10108 -4388 10142 -4372
rect 10108 -6380 10142 -6364
rect 9443 -6448 9459 -6414
rect 9493 -6448 9509 -6414
rect 9561 -6448 9577 -6414
rect 9611 -6448 9627 -6414
rect 9679 -6448 9695 -6414
rect 9729 -6448 9745 -6414
rect 9797 -6448 9813 -6414
rect 9847 -6448 9863 -6414
rect 9915 -6448 9931 -6414
rect 9965 -6448 9981 -6414
rect 10033 -6448 10049 -6414
rect 10083 -6448 10099 -6414
rect 9286 -6516 9320 -6454
rect 10222 -6516 10256 -6454
rect 9286 -6550 9382 -6516
rect 10160 -6550 10256 -6516
rect 5981 -6736 6077 -6702
rect 9923 -6736 10019 -6702
rect 5981 -6798 6015 -6736
rect 9985 -6798 10019 -6736
rect 6138 -6838 6154 -6804
rect 6188 -6838 6204 -6804
rect 6256 -6838 6272 -6804
rect 6306 -6838 6322 -6804
rect 6374 -6838 6390 -6804
rect 6424 -6838 6440 -6804
rect 6492 -6838 6508 -6804
rect 6542 -6838 6558 -6804
rect 6610 -6838 6626 -6804
rect 6660 -6838 6676 -6804
rect 6728 -6838 6744 -6804
rect 6778 -6838 6794 -6804
rect 6846 -6838 6862 -6804
rect 6896 -6838 6912 -6804
rect 6964 -6838 6980 -6804
rect 7014 -6838 7030 -6804
rect 7082 -6838 7098 -6804
rect 7132 -6838 7148 -6804
rect 7200 -6838 7216 -6804
rect 7250 -6838 7266 -6804
rect 7318 -6838 7334 -6804
rect 7368 -6838 7384 -6804
rect 7436 -6838 7452 -6804
rect 7486 -6838 7502 -6804
rect 7554 -6838 7570 -6804
rect 7604 -6838 7620 -6804
rect 7672 -6838 7688 -6804
rect 7722 -6838 7738 -6804
rect 7790 -6838 7806 -6804
rect 7840 -6838 7856 -6804
rect 7908 -6838 7924 -6804
rect 7958 -6838 7974 -6804
rect 8026 -6838 8042 -6804
rect 8076 -6838 8092 -6804
rect 8144 -6838 8160 -6804
rect 8194 -6838 8210 -6804
rect 8262 -6838 8278 -6804
rect 8312 -6838 8328 -6804
rect 8380 -6838 8396 -6804
rect 8430 -6838 8446 -6804
rect 8498 -6838 8514 -6804
rect 8548 -6838 8564 -6804
rect 8616 -6838 8632 -6804
rect 8666 -6838 8682 -6804
rect 8734 -6838 8750 -6804
rect 8784 -6838 8800 -6804
rect 8852 -6838 8868 -6804
rect 8902 -6838 8918 -6804
rect 8970 -6838 8986 -6804
rect 9020 -6838 9036 -6804
rect 9088 -6838 9104 -6804
rect 9138 -6838 9154 -6804
rect 9206 -6838 9222 -6804
rect 9256 -6838 9272 -6804
rect 9324 -6838 9340 -6804
rect 9374 -6838 9390 -6804
rect 9442 -6838 9458 -6804
rect 9492 -6838 9508 -6804
rect 9560 -6838 9576 -6804
rect 9610 -6838 9626 -6804
rect 9678 -6838 9694 -6804
rect 9728 -6838 9744 -6804
rect 9796 -6838 9812 -6804
rect 9846 -6838 9862 -6804
rect 6095 -6897 6129 -6881
rect 6095 -8889 6129 -8873
rect 6213 -6897 6247 -6881
rect 6213 -8889 6247 -8873
rect 6331 -6897 6365 -6881
rect 6331 -8889 6365 -8873
rect 6449 -6897 6483 -6881
rect 6449 -8889 6483 -8873
rect 6567 -6897 6601 -6881
rect 6567 -8889 6601 -8873
rect 6685 -6897 6719 -6881
rect 6685 -8889 6719 -8873
rect 6803 -6897 6837 -6881
rect 6803 -8889 6837 -8873
rect 6921 -6897 6955 -6881
rect 6921 -8889 6955 -8873
rect 7039 -6897 7073 -6881
rect 7039 -8889 7073 -8873
rect 7157 -6897 7191 -6881
rect 7157 -8889 7191 -8873
rect 7275 -6897 7309 -6881
rect 7275 -8889 7309 -8873
rect 7393 -6897 7427 -6881
rect 7393 -8889 7427 -8873
rect 7511 -6897 7545 -6881
rect 7511 -8889 7545 -8873
rect 7629 -6897 7663 -6881
rect 7629 -8889 7663 -8873
rect 7747 -6897 7781 -6881
rect 7747 -8889 7781 -8873
rect 7865 -6897 7899 -6881
rect 7865 -8889 7899 -8873
rect 7983 -6897 8017 -6881
rect 7983 -8889 8017 -8873
rect 8101 -6897 8135 -6881
rect 8101 -8889 8135 -8873
rect 8219 -6897 8253 -6881
rect 8219 -8889 8253 -8873
rect 8337 -6897 8371 -6881
rect 8337 -8889 8371 -8873
rect 8455 -6897 8489 -6881
rect 8455 -8889 8489 -8873
rect 8573 -6897 8607 -6881
rect 8573 -8889 8607 -8873
rect 8691 -6897 8725 -6881
rect 8691 -8889 8725 -8873
rect 8809 -6897 8843 -6881
rect 8809 -8889 8843 -8873
rect 8927 -6897 8961 -6881
rect 8927 -8889 8961 -8873
rect 9045 -6897 9079 -6881
rect 9045 -8889 9079 -8873
rect 9163 -6897 9197 -6881
rect 9163 -8889 9197 -8873
rect 9281 -6897 9315 -6881
rect 9281 -8889 9315 -8873
rect 9399 -6897 9433 -6881
rect 9399 -8889 9433 -8873
rect 9517 -6897 9551 -6881
rect 9517 -8889 9551 -8873
rect 9635 -6897 9669 -6881
rect 9635 -8889 9669 -8873
rect 9753 -6897 9787 -6881
rect 9753 -8889 9787 -8873
rect 9871 -6897 9905 -6881
rect 9871 -8889 9905 -8873
rect 6138 -8966 6154 -8932
rect 6188 -8966 6204 -8932
rect 6256 -8966 6272 -8932
rect 6306 -8966 6322 -8932
rect 6374 -8966 6390 -8932
rect 6424 -8966 6440 -8932
rect 6492 -8966 6508 -8932
rect 6542 -8966 6558 -8932
rect 6610 -8966 6626 -8932
rect 6660 -8966 6676 -8932
rect 6728 -8966 6744 -8932
rect 6778 -8966 6794 -8932
rect 6846 -8966 6862 -8932
rect 6896 -8966 6912 -8932
rect 6964 -8966 6980 -8932
rect 7014 -8966 7030 -8932
rect 7082 -8966 7098 -8932
rect 7132 -8966 7148 -8932
rect 7200 -8966 7216 -8932
rect 7250 -8966 7266 -8932
rect 7318 -8966 7334 -8932
rect 7368 -8966 7384 -8932
rect 7436 -8966 7452 -8932
rect 7486 -8966 7502 -8932
rect 8498 -8966 8514 -8932
rect 8548 -8966 8564 -8932
rect 8616 -8966 8632 -8932
rect 8666 -8966 8682 -8932
rect 8734 -8966 8750 -8932
rect 8784 -8966 8800 -8932
rect 8852 -8966 8868 -8932
rect 8902 -8966 8918 -8932
rect 8970 -8966 8986 -8932
rect 9020 -8966 9036 -8932
rect 9088 -8966 9104 -8932
rect 9138 -8966 9154 -8932
rect 9206 -8966 9222 -8932
rect 9256 -8966 9272 -8932
rect 9324 -8966 9340 -8932
rect 9374 -8966 9390 -8932
rect 9442 -8966 9458 -8932
rect 9492 -8966 9508 -8932
rect 9560 -8966 9576 -8932
rect 9610 -8966 9626 -8932
rect 9678 -8966 9694 -8932
rect 9728 -8966 9744 -8932
rect 9796 -8966 9812 -8932
rect 9846 -8966 9862 -8932
rect 5981 -9034 6015 -8972
rect 9985 -9034 10019 -8972
rect 5981 -9068 6077 -9034
rect 9923 -9068 10019 -9034
<< viali >>
rect 6154 12332 6188 12366
rect 6272 12332 6306 12366
rect 6390 12332 6424 12366
rect 6508 12332 6542 12366
rect 6626 12332 6660 12366
rect 6744 12332 6778 12366
rect 6862 12332 6896 12366
rect 6980 12332 7014 12366
rect 7098 12332 7132 12366
rect 7216 12332 7250 12366
rect 7334 12332 7368 12366
rect 7452 12332 7486 12366
rect 8514 12332 8548 12366
rect 8632 12332 8666 12366
rect 8750 12332 8784 12366
rect 8868 12332 8902 12366
rect 8986 12332 9020 12366
rect 9104 12332 9138 12366
rect 9222 12332 9256 12366
rect 9340 12332 9374 12366
rect 9458 12332 9492 12366
rect 9576 12332 9610 12366
rect 9694 12332 9728 12366
rect 9812 12332 9846 12366
rect 5981 11885 6015 12285
rect 5981 10285 6015 10685
rect 6095 10297 6129 12273
rect 6213 10297 6247 12273
rect 6331 10297 6365 12273
rect 6449 10297 6483 12273
rect 6567 10297 6601 12273
rect 6685 10297 6719 12273
rect 6803 10297 6837 12273
rect 6921 10297 6955 12273
rect 7039 10297 7073 12273
rect 7157 10297 7191 12273
rect 7275 10297 7309 12273
rect 7393 10297 7427 12273
rect 7511 10297 7545 12273
rect 7629 10297 7663 12273
rect 7747 10297 7781 12273
rect 7865 10297 7899 12273
rect 7983 10297 8017 12273
rect 8101 10297 8135 12273
rect 8219 10297 8253 12273
rect 8337 10297 8371 12273
rect 8455 10297 8489 12273
rect 8573 10297 8607 12273
rect 8691 10297 8725 12273
rect 8809 10297 8843 12273
rect 8927 10297 8961 12273
rect 9045 10297 9079 12273
rect 9163 10297 9197 12273
rect 9281 10297 9315 12273
rect 9399 10297 9433 12273
rect 9517 10297 9551 12273
rect 9635 10297 9669 12273
rect 9753 10297 9787 12273
rect 9871 10297 9905 12273
rect 9985 11885 10019 12285
rect 9985 10285 10019 10685
rect 6154 10204 6188 10238
rect 6272 10204 6306 10238
rect 6390 10204 6424 10238
rect 6508 10204 6542 10238
rect 6626 10204 6660 10238
rect 6744 10204 6778 10238
rect 6862 10204 6896 10238
rect 6980 10204 7014 10238
rect 7098 10204 7132 10238
rect 7216 10204 7250 10238
rect 7334 10204 7368 10238
rect 7452 10204 7486 10238
rect 7570 10204 7604 10238
rect 7688 10204 7722 10238
rect 7806 10204 7840 10238
rect 7924 10204 7958 10238
rect 8042 10204 8076 10238
rect 8160 10204 8194 10238
rect 8278 10204 8312 10238
rect 8396 10204 8430 10238
rect 8514 10204 8548 10238
rect 8632 10204 8666 10238
rect 8750 10204 8784 10238
rect 8868 10204 8902 10238
rect 8986 10204 9020 10238
rect 9104 10204 9138 10238
rect 9222 10204 9256 10238
rect 9340 10204 9374 10238
rect 9458 10204 9492 10238
rect 9576 10204 9610 10238
rect 9694 10204 9728 10238
rect 9812 10204 9846 10238
rect 5918 9814 5952 9848
rect 6036 9814 6070 9848
rect 6154 9814 6188 9848
rect 6272 9814 6306 9848
rect 6390 9814 6424 9848
rect 6508 9814 6542 9848
rect 5190 9040 5300 9430
rect 5420 9040 5530 9430
rect 5745 9376 5779 9776
rect 5745 7776 5779 8176
rect 5859 7788 5893 9764
rect 5977 7788 6011 9764
rect 6095 7788 6129 9764
rect 6213 7788 6247 9764
rect 6331 7788 6365 9764
rect 6449 7788 6483 9764
rect 6567 7788 6601 9764
rect 6681 9376 6715 9776
rect 9459 9814 9493 9848
rect 9577 9814 9611 9848
rect 9695 9814 9729 9848
rect 9813 9814 9847 9848
rect 9931 9814 9965 9848
rect 10049 9814 10083 9848
rect 7119 9642 7153 9676
rect 8847 9642 8881 9676
rect 6909 9100 6943 9600
rect 7023 9112 7057 9588
rect 7119 9112 7153 9588
rect 7215 9112 7249 9588
rect 7311 9112 7345 9588
rect 7407 9112 7441 9588
rect 7503 9112 7537 9588
rect 7599 9112 7633 9588
rect 7695 9112 7729 9588
rect 7791 9112 7825 9588
rect 7887 9112 7921 9588
rect 7983 9112 8017 9588
rect 8079 9112 8113 9588
rect 8175 9112 8209 9588
rect 8271 9112 8305 9588
rect 8367 9112 8401 9588
rect 8463 9112 8497 9588
rect 8559 9112 8593 9588
rect 8655 9112 8689 9588
rect 8751 9112 8785 9588
rect 8847 9112 8881 9588
rect 8943 9112 8977 9588
rect 9057 9100 9091 9600
rect 7311 9016 7345 9050
rect 7503 9016 7537 9050
rect 7695 9016 7729 9050
rect 7887 9016 7921 9050
rect 8079 9016 8113 9050
rect 8271 9016 8305 9050
rect 8463 9016 8497 9050
rect 8655 9016 8689 9050
rect 9286 9376 9320 9776
rect 6681 7776 6715 8176
rect 5918 7704 5952 7738
rect 6036 7704 6070 7738
rect 6154 7704 6188 7738
rect 6272 7704 6306 7738
rect 6390 7704 6424 7738
rect 6508 7704 6542 7738
rect 7129 8698 7497 8732
rect 7587 8698 7955 8732
rect 8045 8698 8413 8732
rect 8503 8698 8871 8732
rect 6953 8260 6987 8660
rect 6953 6660 6987 7060
rect 7067 6672 7101 8648
rect 7525 6672 7559 8648
rect 7983 6672 8017 8648
rect 8441 6672 8475 8648
rect 8899 6672 8933 8648
rect 9013 8260 9047 8660
rect 9286 7776 9320 8176
rect 9400 7788 9434 9764
rect 9518 7788 9552 9764
rect 9636 7788 9670 9764
rect 9754 7788 9788 9764
rect 9872 7788 9906 9764
rect 9990 7788 10024 9764
rect 10108 7788 10142 9764
rect 10222 9376 10256 9776
rect 10222 7776 10256 8176
rect 9459 7704 9493 7738
rect 9577 7704 9611 7738
rect 9695 7704 9729 7738
rect 9813 7704 9847 7738
rect 9931 7704 9965 7738
rect 10049 7704 10083 7738
rect 9013 6660 9047 7060
rect 7129 6588 7497 6622
rect 7587 6588 7955 6622
rect 8045 6588 8413 6622
rect 8503 6588 8871 6622
rect 10542 6340 10602 7260
rect 10864 7268 11340 7302
rect 10864 7172 11340 7206
rect 11390 7202 11424 7236
rect 10864 7076 11340 7110
rect 10864 6980 11340 7014
rect 11390 7010 11424 7044
rect 10864 6884 11340 6918
rect 10980 6539 11396 6592
rect 11396 6539 11412 6592
rect 3469 3964 3503 4340
rect 3557 3964 3591 4340
rect 3671 3958 3705 4346
rect 3513 3880 3547 3914
rect 3469 3250 3503 3626
rect 3557 3250 3591 3626
rect 3671 3244 3705 3632
rect 3513 3166 3547 3200
rect 4137 3958 4171 4346
rect 4251 3964 4285 4340
rect 4339 3964 4373 4340
rect 4295 3880 4329 3914
rect 11278 3920 14428 3978
rect 4137 3244 4171 3632
rect 4251 3250 4285 3626
rect 4339 3250 4373 3626
rect 4295 3166 4329 3200
rect 11278 3908 11356 3920
rect 11356 3908 13716 3920
rect 13716 3908 13874 3920
rect 13874 3908 14032 3920
rect 14032 3908 14190 3920
rect 14190 3908 14348 3920
rect 14348 3908 14428 3920
rect 2070 2861 2104 2895
rect 2166 2861 2200 2895
rect 2262 2861 2296 2895
rect 2358 2861 2392 2895
rect 2454 2861 2488 2895
rect 2550 2861 2584 2895
rect 2646 2861 2680 2895
rect 2742 2861 2776 2895
rect 2838 2861 2872 2895
rect 2934 2861 2968 2895
rect 3030 2861 3064 2895
rect 3126 2861 3160 2895
rect 3222 2861 3256 2895
rect 3318 2861 3352 2895
rect 3414 2861 3448 2895
rect 3510 2861 3544 2895
rect 3606 2861 3640 2895
rect 3702 2861 3736 2895
rect 3798 2861 3832 2895
rect 3894 2861 3928 2895
rect 3990 2861 4024 2895
rect 4086 2861 4120 2895
rect 4182 2861 4216 2895
rect 4278 2861 4312 2895
rect 4374 2861 4408 2895
rect 4470 2861 4504 2895
rect 4566 2861 4600 2895
rect 4662 2861 4696 2895
rect 4758 2861 4792 2895
rect 4854 2861 4888 2895
rect 4950 2861 4984 2895
rect 5046 2861 5080 2895
rect 5142 2861 5176 2895
rect 5238 2861 5272 2895
rect 5334 2861 5368 2895
rect 5430 2861 5464 2895
rect 5526 2861 5560 2895
rect 5622 2861 5656 2895
rect 5718 2861 5752 2895
rect 5814 2861 5848 2895
rect 5910 2861 5944 2895
rect 6006 2861 6040 2895
rect 6102 2861 6136 2895
rect 6198 2861 6232 2895
rect 6294 2861 6328 2895
rect 6390 2861 6424 2895
rect 6486 2861 6520 2895
rect 6582 2861 6616 2895
rect 6678 2861 6712 2895
rect 6774 2861 6808 2895
rect 6870 2861 6904 2895
rect 6966 2861 7000 2895
rect 7062 2861 7096 2895
rect 7158 2861 7192 2895
rect 7254 2861 7288 2895
rect 7350 2861 7384 2895
rect 7446 2861 7480 2895
rect 7542 2861 7576 2895
rect 7638 2861 7672 2895
rect 7734 2861 7768 2895
rect 7830 2861 7864 2895
rect 7926 2861 7960 2895
rect 8022 2861 8056 2895
rect 8118 2861 8152 2895
rect 8214 2861 8248 2895
rect 8310 2861 8344 2895
rect 8406 2861 8440 2895
rect 8502 2861 8536 2895
rect 8598 2861 8632 2895
rect 8694 2861 8728 2895
rect 8790 2861 8824 2895
rect 8886 2861 8920 2895
rect 8982 2861 9016 2895
rect 9078 2861 9112 2895
rect 9174 2861 9208 2895
rect 9270 2861 9304 2895
rect 9366 2861 9400 2895
rect 9462 2861 9496 2895
rect 9558 2861 9592 2895
rect 9654 2861 9688 2895
rect 9750 2861 9784 2895
rect 9846 2861 9880 2895
rect 9942 2861 9976 2895
rect 10038 2861 10072 2895
rect 10134 2861 10168 2895
rect 2368 2488 2372 2522
rect 2372 2488 2402 2522
rect 2440 2488 2474 2522
rect 2709 2363 3106 2613
rect 3240 2363 3637 2613
rect 3984 2472 4018 2506
rect 3974 2332 4008 2338
rect 3974 2304 4007 2332
rect 4007 2304 4008 2332
rect 5334 2756 5368 2784
rect 5334 2750 5368 2756
rect 5238 2334 5272 2340
rect 5238 2306 5272 2334
rect 2070 2195 2104 2229
rect 2166 2195 2200 2229
rect 2262 2195 2296 2229
rect 2358 2195 2392 2229
rect 2454 2195 2488 2229
rect 2550 2195 2584 2229
rect 2646 2195 2680 2229
rect 2742 2195 2776 2229
rect 2838 2195 2872 2229
rect 2934 2195 2968 2229
rect 3030 2195 3064 2229
rect 3126 2195 3160 2229
rect 3222 2195 3256 2229
rect 3318 2195 3352 2229
rect 3414 2195 3448 2229
rect 3510 2195 3544 2229
rect 3606 2195 3640 2229
rect 3702 2195 3736 2229
rect 3798 2195 3832 2229
rect 3894 2195 3928 2229
rect 3990 2195 4024 2229
rect 4086 2195 4120 2229
rect 4182 2195 4216 2229
rect 4278 2195 4312 2229
rect 4374 2195 4408 2229
rect 4470 2195 4504 2229
rect 4566 2195 4600 2229
rect 4662 2195 4696 2229
rect 4758 2195 4792 2229
rect 4854 2195 4888 2229
rect 4950 2195 4984 2229
rect 5046 2195 5080 2229
rect 5142 2195 5176 2229
rect 5238 2195 5272 2229
rect 5334 2195 5368 2229
rect 5430 2195 5464 2229
rect 5526 2195 5560 2229
rect 5622 2195 5656 2229
rect 5718 2195 5752 2229
rect 5814 2195 5848 2229
rect 5910 2195 5944 2229
rect 6006 2195 6040 2229
rect 6102 2195 6136 2229
rect 6198 2195 6232 2229
rect 6294 2195 6328 2229
rect 6390 2195 6424 2229
rect 6486 2195 6520 2229
rect 6582 2195 6616 2229
rect 6678 2195 6712 2229
rect 6774 2195 6808 2229
rect 6870 2195 6904 2229
rect 6966 2195 7000 2229
rect 7062 2195 7096 2229
rect 7158 2195 7192 2229
rect 7254 2195 7288 2229
rect 7350 2195 7384 2229
rect 7446 2195 7480 2229
rect 7542 2195 7576 2229
rect 7638 2195 7672 2229
rect 7734 2195 7768 2229
rect 7830 2195 7864 2229
rect 7926 2195 7960 2229
rect 8022 2195 8056 2229
rect 8118 2195 8152 2229
rect 8214 2195 8248 2229
rect 8310 2195 8344 2229
rect 8406 2195 8440 2229
rect 8502 2195 8536 2229
rect 8598 2195 8632 2229
rect 8694 2195 8728 2229
rect 8790 2195 8824 2229
rect 8886 2195 8920 2229
rect 8982 2195 9016 2229
rect 9078 2195 9112 2229
rect 9174 2195 9208 2229
rect 9270 2195 9304 2229
rect 9366 2195 9400 2229
rect 9462 2195 9496 2229
rect 9558 2195 9592 2229
rect 9654 2195 9688 2229
rect 9750 2195 9784 2229
rect 9846 2195 9880 2229
rect 9942 2195 9976 2229
rect 10038 2195 10072 2229
rect 10134 2195 10168 2229
rect 2368 1902 2372 1936
rect 2372 1902 2402 1936
rect 2440 1902 2474 1936
rect 2709 1811 3106 2061
rect 3240 1811 3637 2061
rect 3974 2092 4007 2120
rect 4007 2092 4008 2120
rect 3974 2086 4008 2092
rect 3984 1918 4018 1952
rect 4171 1926 4205 1929
rect 4171 1895 4172 1926
rect 4172 1895 4205 1926
rect 4448 1918 4482 1952
rect 5238 2090 5272 2118
rect 5238 2084 5272 2090
rect 4562 1952 4596 1954
rect 4562 1920 4596 1952
rect 4955 1936 4989 1941
rect 4955 1907 4956 1936
rect 4956 1907 4989 1936
rect 4847 1749 4881 1767
rect 4847 1733 4864 1749
rect 4864 1733 4881 1749
rect 5049 1666 5083 1695
rect 5049 1661 5080 1666
rect 5080 1661 5083 1666
rect 5716 1904 5750 1905
rect 5716 1871 5746 1904
rect 5746 1871 5750 1904
rect 6124 1892 6128 1926
rect 6128 1892 6158 1926
rect 5334 1668 5368 1674
rect 5334 1640 5368 1668
rect 6582 1936 6616 1970
rect 7446 1936 7480 1970
rect 7254 1862 7288 1896
rect 7830 1862 7864 1896
rect 8203 1861 8204 1894
rect 8204 1861 8237 1894
rect 8203 1860 8237 1861
rect 9489 1892 9493 1926
rect 9493 1892 9523 1926
rect 9561 1892 9595 1926
rect 9876 1892 9880 1926
rect 9880 1892 9910 1926
rect 9948 1892 9982 1926
rect 10200 1850 10260 1930
rect 8887 1798 8918 1823
rect 8918 1798 8921 1823
rect 8887 1789 8921 1798
rect 8887 1749 8921 1751
rect 8887 1717 8918 1749
rect 8918 1717 8921 1749
rect 10828 1688 10888 2098
rect 10998 1688 11058 2098
rect 2070 1529 2104 1563
rect 2166 1529 2200 1563
rect 2262 1529 2296 1563
rect 2358 1529 2392 1563
rect 2454 1529 2488 1563
rect 2550 1529 2584 1563
rect 2646 1529 2680 1563
rect 2742 1529 2776 1563
rect 2838 1529 2872 1563
rect 2934 1529 2968 1563
rect 3030 1529 3064 1563
rect 3126 1529 3160 1563
rect 3222 1529 3256 1563
rect 3318 1529 3352 1563
rect 3414 1529 3448 1563
rect 3510 1529 3544 1563
rect 3606 1529 3640 1563
rect 3702 1529 3736 1563
rect 3798 1529 3832 1563
rect 3894 1529 3928 1563
rect 3990 1529 4024 1563
rect 4086 1529 4120 1563
rect 4182 1529 4216 1563
rect 4278 1529 4312 1563
rect 4374 1529 4408 1563
rect 4470 1529 4504 1563
rect 4566 1529 4600 1563
rect 4662 1529 4696 1563
rect 4758 1529 4792 1563
rect 4854 1529 4888 1563
rect 4950 1529 4984 1563
rect 5046 1529 5080 1563
rect 5142 1529 5176 1563
rect 5238 1529 5272 1563
rect 5334 1529 5368 1563
rect 5430 1529 5464 1563
rect 5526 1529 5560 1563
rect 5622 1529 5656 1563
rect 5718 1529 5752 1563
rect 5814 1529 5848 1563
rect 5910 1529 5944 1563
rect 6006 1529 6040 1563
rect 6102 1529 6136 1563
rect 6198 1529 6232 1563
rect 6294 1529 6328 1563
rect 6390 1529 6424 1563
rect 6486 1529 6520 1563
rect 6582 1529 6616 1563
rect 6678 1529 6712 1563
rect 6774 1529 6808 1563
rect 6870 1529 6904 1563
rect 6966 1529 7000 1563
rect 7062 1529 7096 1563
rect 7158 1529 7192 1563
rect 7254 1529 7288 1563
rect 7350 1529 7384 1563
rect 7446 1529 7480 1563
rect 7542 1529 7576 1563
rect 7638 1529 7672 1563
rect 7734 1529 7768 1563
rect 7830 1529 7864 1563
rect 7926 1529 7960 1563
rect 8022 1529 8056 1563
rect 8118 1529 8152 1563
rect 8214 1529 8248 1563
rect 8310 1529 8344 1563
rect 8406 1529 8440 1563
rect 8502 1529 8536 1563
rect 8598 1529 8632 1563
rect 8694 1529 8728 1563
rect 8790 1529 8824 1563
rect 8886 1529 8920 1563
rect 8982 1529 9016 1563
rect 9078 1529 9112 1563
rect 9174 1529 9208 1563
rect 9270 1529 9304 1563
rect 9366 1529 9400 1563
rect 9462 1529 9496 1563
rect 9558 1529 9592 1563
rect 9654 1529 9688 1563
rect 9750 1529 9784 1563
rect 9846 1529 9880 1563
rect 9942 1529 9976 1563
rect 10038 1529 10072 1563
rect 10134 1529 10168 1563
rect 11436 3784 11804 3818
rect 11894 3784 12262 3818
rect 12352 3784 12720 3818
rect 12810 3784 13178 3818
rect 13268 3784 13636 3818
rect 11374 1749 11408 3725
rect 11832 1749 11866 3725
rect 12290 1749 12324 3725
rect 12748 1749 12782 3725
rect 13206 1749 13240 3725
rect 13664 1749 13698 3725
rect 11436 1656 11804 1690
rect 11894 1656 12262 1690
rect 12352 1656 12720 1690
rect 12810 1656 13178 1690
rect 13268 1656 13636 1690
rect 13892 1749 13926 3725
rect 13980 1749 14014 3725
rect 13936 1656 13970 1690
rect 14208 1749 14242 3725
rect 14296 1749 14330 3725
rect 14252 1656 14286 1690
rect 1796 1433 1830 1467
rect 1888 1433 1922 1467
rect 1980 1433 2014 1467
rect 2072 1433 2106 1467
rect 2164 1433 2198 1467
rect 2256 1433 2290 1467
rect 2348 1433 2382 1467
rect 2440 1433 2474 1467
rect 2532 1433 2566 1467
rect 2624 1433 2658 1467
rect 2716 1433 2750 1467
rect 2808 1433 2842 1467
rect 1891 1118 2011 1158
rect 2259 1118 2379 1158
rect 2627 1118 2747 1158
rect 3520 1156 3524 1190
rect 3524 1156 3554 1190
rect 3592 1156 3626 1190
rect 1796 889 1830 923
rect 1888 889 1922 923
rect 1980 889 2014 923
rect 2072 889 2106 923
rect 2164 889 2198 923
rect 2256 889 2290 923
rect 2348 889 2382 923
rect 2440 889 2474 923
rect 2532 889 2566 923
rect 2624 889 2658 923
rect 2716 889 2750 923
rect 2808 889 2842 923
rect 3861 1031 4258 1281
rect 4392 1031 4789 1281
rect 5334 1424 5368 1452
rect 5334 1418 5368 1424
rect 5136 1140 5170 1174
rect 5712 1188 5746 1222
rect 5126 1000 5160 1006
rect 5126 972 5159 1000
rect 5159 972 5160 1000
rect 5238 1002 5272 1008
rect 5238 974 5272 1002
rect 6128 1166 6162 1200
rect 6582 1122 6616 1156
rect 7254 1196 7288 1230
rect 7446 1122 7480 1156
rect 7830 1196 7864 1230
rect 8205 1231 8239 1233
rect 8205 1199 8238 1231
rect 8238 1199 8239 1231
rect 8481 1343 8490 1370
rect 8490 1343 8515 1370
rect 8481 1336 8515 1343
rect 8481 1294 8515 1298
rect 8481 1264 8490 1294
rect 8490 1264 8515 1294
rect 8890 1343 8918 1366
rect 8918 1343 8924 1366
rect 8890 1332 8924 1343
rect 8890 1260 8918 1294
rect 8918 1260 8924 1294
rect 9469 1220 9503 1221
rect 9469 1187 9502 1220
rect 9502 1187 9503 1220
rect 9594 1199 9628 1214
rect 9594 1180 9602 1199
rect 9602 1180 9628 1199
rect 10200 1160 10260 1240
rect 3222 863 3256 897
rect 3318 863 3352 897
rect 3414 863 3448 897
rect 3510 863 3544 897
rect 3606 863 3640 897
rect 3702 863 3736 897
rect 3798 863 3832 897
rect 3894 863 3928 897
rect 3990 863 4024 897
rect 4086 863 4120 897
rect 4182 863 4216 897
rect 4278 863 4312 897
rect 4374 863 4408 897
rect 4470 863 4504 897
rect 4566 863 4600 897
rect 4662 863 4696 897
rect 4758 863 4792 897
rect 4854 863 4888 897
rect 4950 863 4984 897
rect 5046 863 5080 897
rect 5142 863 5176 897
rect 5238 863 5272 897
rect 5334 863 5368 897
rect 5430 863 5464 897
rect 5526 863 5560 897
rect 5622 863 5656 897
rect 5718 863 5752 897
rect 5814 863 5848 897
rect 5910 863 5944 897
rect 6006 863 6040 897
rect 6102 863 6136 897
rect 6198 863 6232 897
rect 6294 863 6328 897
rect 6390 863 6424 897
rect 6486 863 6520 897
rect 6582 863 6616 897
rect 6678 863 6712 897
rect 6774 863 6808 897
rect 6870 863 6904 897
rect 6966 863 7000 897
rect 7062 863 7096 897
rect 7158 863 7192 897
rect 7254 863 7288 897
rect 7350 863 7384 897
rect 7446 863 7480 897
rect 7542 863 7576 897
rect 7638 863 7672 897
rect 7734 863 7768 897
rect 7830 863 7864 897
rect 7926 863 7960 897
rect 8022 863 8056 897
rect 8118 863 8152 897
rect 8214 863 8248 897
rect 8310 863 8344 897
rect 8406 863 8440 897
rect 8502 863 8536 897
rect 8598 863 8632 897
rect 8694 863 8728 897
rect 8790 863 8824 897
rect 8886 863 8920 897
rect 8982 863 9016 897
rect 9078 863 9112 897
rect 9174 863 9208 897
rect 9270 863 9304 897
rect 9366 863 9400 897
rect 9462 863 9496 897
rect 9558 863 9592 897
rect 9654 863 9688 897
rect 9750 863 9784 897
rect 9846 863 9880 897
rect 9942 863 9976 897
rect 10038 863 10072 897
rect 10134 863 10168 897
rect 3704 188 3738 576
rect 3818 194 3852 570
rect 3906 194 3940 570
rect 3862 110 3896 144
rect 10520 1346 10888 1380
rect 10978 1346 11346 1380
rect 11436 1346 11804 1380
rect 11894 1346 12262 1380
rect 12352 1346 12720 1380
rect 12810 1346 13178 1380
rect 13268 1346 13636 1380
rect 10458 320 10492 1296
rect 10916 320 10950 1296
rect 11374 320 11408 1296
rect 11832 320 11866 1296
rect 12290 320 12324 1296
rect 12748 320 12782 1296
rect 13206 320 13240 1296
rect 13664 320 13698 1296
rect 10520 236 10888 270
rect 10978 236 11346 270
rect 11436 236 11804 270
rect 11894 236 12262 270
rect 12352 236 12720 270
rect 12810 236 13178 270
rect 13268 236 13636 270
rect 13936 1346 13970 1380
rect 13892 320 13926 1296
rect 13980 320 14014 1296
rect 14252 1346 14286 1380
rect 14208 320 14242 1296
rect 14296 320 14330 1296
rect 15552 867 15928 901
rect 15978 823 16012 857
rect 15552 779 15928 813
rect 16266 867 16642 901
rect 16692 823 16726 857
rect 16266 779 16642 813
rect 16980 867 17356 901
rect 17406 823 17440 857
rect 16980 779 17356 813
rect 17694 867 18070 901
rect 18120 823 18154 857
rect 17694 779 18070 813
rect 18408 867 18784 901
rect 18834 823 18868 857
rect 18408 779 18784 813
rect 19122 867 19498 901
rect 19548 823 19582 857
rect 19122 779 19498 813
rect 19836 867 20212 901
rect 20262 823 20296 857
rect 19836 779 20212 813
rect 20550 867 20926 901
rect 20976 823 21010 857
rect 20550 779 20926 813
rect 21264 867 21640 901
rect 21690 823 21724 857
rect 21264 779 21640 813
rect 21978 867 22354 901
rect 22404 823 22438 857
rect 21978 779 22354 813
rect 22692 867 23068 901
rect 23118 823 23152 857
rect 22692 779 23068 813
rect 23406 867 23782 901
rect 23832 823 23866 857
rect 23406 779 23782 813
rect 24120 867 24496 901
rect 24546 823 24580 857
rect 24120 779 24496 813
rect 24834 867 25210 901
rect 25260 823 25294 857
rect 24834 779 25210 813
rect 25548 867 25924 901
rect 25974 823 26008 857
rect 25548 779 25924 813
rect 26262 867 26638 901
rect 26688 823 26722 857
rect 26262 779 26638 813
rect 26976 867 27352 901
rect 27402 823 27436 857
rect 26976 779 27352 813
rect 27690 867 28066 901
rect 28116 823 28150 857
rect 27690 779 28066 813
rect 28404 867 28780 901
rect 28830 823 28864 857
rect 28404 779 28780 813
rect 29118 867 29494 901
rect 29544 823 29578 857
rect 29118 779 29494 813
rect 29832 867 30208 901
rect 30258 823 30292 857
rect 29832 779 30208 813
rect 30546 867 30922 901
rect 30972 823 31006 857
rect 30546 779 30922 813
rect 31260 867 31636 901
rect 31686 823 31720 857
rect 31260 779 31636 813
rect 31974 867 32350 901
rect 32400 823 32434 857
rect 31974 779 32350 813
rect 32688 867 33064 901
rect 33114 823 33148 857
rect 32688 779 33064 813
rect 33402 867 33778 901
rect 33828 823 33862 857
rect 33402 779 33778 813
rect 34116 867 34492 901
rect 34542 823 34576 857
rect 34116 779 34492 813
rect 34830 867 35206 901
rect 35256 823 35290 857
rect 34830 779 35206 813
rect 35544 867 35920 901
rect 35970 823 36004 857
rect 35544 779 35920 813
rect 36258 867 36634 901
rect 36684 823 36718 857
rect 36258 779 36634 813
rect 36972 867 37348 901
rect 37398 823 37432 857
rect 36972 779 37348 813
rect 37686 867 38062 901
rect 38112 823 38146 857
rect 37686 779 38062 813
rect 38400 867 38776 901
rect 38826 823 38860 857
rect 38400 779 38776 813
rect 15546 665 15934 699
rect 16260 665 16648 699
rect 16974 665 17362 699
rect 17688 665 18076 699
rect 18402 665 18790 699
rect 19116 665 19504 699
rect 19830 665 20218 699
rect 20544 665 20932 699
rect 21258 665 21646 699
rect 21972 665 22360 699
rect 22686 665 23074 699
rect 23400 665 23788 699
rect 24114 665 24502 699
rect 24828 665 25216 699
rect 25542 665 25930 699
rect 26256 665 26644 699
rect 26970 665 27358 699
rect 27684 665 28072 699
rect 28398 665 28786 699
rect 29112 665 29500 699
rect 29826 665 30214 699
rect 30540 665 30928 699
rect 31254 665 31642 699
rect 31968 665 32356 699
rect 32682 665 33070 699
rect 33396 665 33784 699
rect 34110 665 34498 699
rect 34824 665 35212 699
rect 35538 665 35926 699
rect 36252 665 36640 699
rect 36966 665 37354 699
rect 37680 665 38068 699
rect 38394 665 38782 699
rect 39381 991 39778 1029
rect 39912 991 40309 1029
rect 39381 825 39778 863
rect 39912 825 40309 863
rect 39381 659 39778 697
rect 39912 659 40309 697
rect 39381 493 39778 531
rect 39912 493 40309 531
rect 39170 380 39233 470
rect 39233 380 39250 470
rect 10358 134 10440 158
rect 10440 134 13716 158
rect 13716 134 13874 158
rect 13874 134 14032 158
rect 14032 134 14190 158
rect 14190 134 14348 158
rect 14348 134 14428 158
rect 10358 78 14428 134
rect 15546 163 15934 197
rect 16260 163 16648 197
rect 16974 163 17362 197
rect 17688 163 18076 197
rect 18402 163 18790 197
rect 19116 163 19504 197
rect 19830 163 20218 197
rect 20544 163 20932 197
rect 21258 163 21646 197
rect 21972 163 22360 197
rect 22686 163 23074 197
rect 23400 163 23788 197
rect 24114 163 24502 197
rect 24828 163 25216 197
rect 25542 163 25930 197
rect 26256 163 26644 197
rect 26970 163 27358 197
rect 27684 163 28072 197
rect 28398 163 28786 197
rect 29112 163 29500 197
rect 29826 163 30214 197
rect 30540 163 30928 197
rect 31254 163 31642 197
rect 31968 163 32356 197
rect 32682 163 33070 197
rect 33396 163 33784 197
rect 34110 163 34498 197
rect 34824 163 35212 197
rect 35538 163 35926 197
rect 36252 163 36640 197
rect 36966 163 37354 197
rect 37680 163 38068 197
rect 38394 163 38782 197
rect 3704 -526 3738 -138
rect 3818 -520 3852 -144
rect 3906 -520 3940 -144
rect 3862 -604 3896 -570
rect 15552 49 15928 83
rect 15978 5 16012 39
rect 15552 -39 15928 -5
rect 16266 49 16642 83
rect 16692 5 16726 39
rect 16266 -39 16642 -5
rect 16980 49 17356 83
rect 17406 5 17440 39
rect 16980 -39 17356 -5
rect 17694 49 18070 83
rect 18120 5 18154 39
rect 17694 -39 18070 -5
rect 18408 49 18784 83
rect 18834 5 18868 39
rect 18408 -39 18784 -5
rect 19122 49 19498 83
rect 19548 5 19582 39
rect 19122 -39 19498 -5
rect 19836 49 20212 83
rect 20262 5 20296 39
rect 19836 -39 20212 -5
rect 20550 49 20926 83
rect 20976 5 21010 39
rect 20550 -39 20926 -5
rect 21264 49 21640 83
rect 21690 5 21724 39
rect 21264 -39 21640 -5
rect 21978 49 22354 83
rect 22404 5 22438 39
rect 21978 -39 22354 -5
rect 22692 49 23068 83
rect 23118 5 23152 39
rect 22692 -39 23068 -5
rect 23406 49 23782 83
rect 23832 5 23866 39
rect 23406 -39 23782 -5
rect 24120 49 24496 83
rect 24546 5 24580 39
rect 24120 -39 24496 -5
rect 24834 49 25210 83
rect 25260 5 25294 39
rect 24834 -39 25210 -5
rect 25548 49 25924 83
rect 25974 5 26008 39
rect 25548 -39 25924 -5
rect 26262 49 26638 83
rect 26688 5 26722 39
rect 26262 -39 26638 -5
rect 26976 49 27352 83
rect 27402 5 27436 39
rect 26976 -39 27352 -5
rect 27690 49 28066 83
rect 28116 5 28150 39
rect 27690 -39 28066 -5
rect 28404 49 28780 83
rect 28830 5 28864 39
rect 28404 -39 28780 -5
rect 29118 49 29494 83
rect 29544 5 29578 39
rect 29118 -39 29494 -5
rect 29832 49 30208 83
rect 30258 5 30292 39
rect 29832 -39 30208 -5
rect 30546 49 30922 83
rect 30972 5 31006 39
rect 30546 -39 30922 -5
rect 31260 49 31636 83
rect 31686 5 31720 39
rect 31260 -39 31636 -5
rect 31974 49 32350 83
rect 32400 5 32434 39
rect 31974 -39 32350 -5
rect 32688 49 33064 83
rect 33114 5 33148 39
rect 32688 -39 33064 -5
rect 33402 49 33778 83
rect 33828 5 33862 39
rect 33402 -39 33778 -5
rect 34116 49 34492 83
rect 34542 5 34576 39
rect 34116 -39 34492 -5
rect 34830 49 35206 83
rect 35256 5 35290 39
rect 34830 -39 35206 -5
rect 35544 49 35920 83
rect 35970 5 36004 39
rect 35544 -39 35920 -5
rect 36258 49 36634 83
rect 36684 5 36718 39
rect 36258 -39 36634 -5
rect 36972 49 37348 83
rect 37398 5 37432 39
rect 36972 -39 37348 -5
rect 37686 49 38062 83
rect 38112 5 38146 39
rect 37686 -39 38062 -5
rect 38400 49 38776 83
rect 38826 5 38860 39
rect 38400 -39 38776 -5
rect 39381 327 39778 365
rect 39912 327 40309 365
rect 39381 161 39778 199
rect 39912 161 40309 199
rect 39381 -5 39778 33
rect 39912 -5 40309 33
rect 39381 -171 39778 -133
rect 39912 -171 40309 -133
rect 10231 -417 10265 -383
rect 10775 -417 10809 -383
rect 10231 -509 10265 -475
rect 10231 -601 10265 -567
rect 10540 -598 10580 -478
rect 10775 -509 10809 -475
rect 10775 -601 10809 -567
rect 10231 -693 10265 -659
rect 10775 -693 10809 -659
rect 10231 -785 10265 -751
rect 10775 -785 10809 -751
rect 10231 -877 10265 -843
rect 10570 -827 10604 -793
rect 10775 -877 10809 -843
rect 10231 -969 10265 -935
rect 10231 -1061 10265 -1027
rect 10775 -969 10809 -935
rect 10775 -1061 10809 -1027
rect 10231 -1153 10265 -1119
rect 10231 -1245 10265 -1211
rect 10540 -1242 10580 -1122
rect 10775 -1153 10809 -1119
rect 10775 -1245 10809 -1211
rect 10231 -1337 10265 -1303
rect 10775 -1337 10809 -1303
rect 7129 -3222 7497 -3188
rect 7587 -3222 7955 -3188
rect 8045 -3222 8413 -3188
rect 8503 -3222 8871 -3188
rect 6953 -3660 6987 -3260
rect 5918 -4338 5952 -4304
rect 6036 -4338 6070 -4304
rect 6154 -4338 6188 -4304
rect 6272 -4338 6306 -4304
rect 6390 -4338 6424 -4304
rect 6508 -4338 6542 -4304
rect 5745 -4776 5779 -4376
rect 5190 -6030 5300 -5640
rect 5420 -6030 5530 -5640
rect 5745 -6376 5779 -5976
rect 5859 -6364 5893 -4388
rect 5977 -6364 6011 -4388
rect 6095 -6364 6129 -4388
rect 6213 -6364 6247 -4388
rect 6331 -6364 6365 -4388
rect 6449 -6364 6483 -4388
rect 6567 -6364 6601 -4388
rect 6681 -4776 6715 -4376
rect 6953 -5260 6987 -4860
rect 7067 -5248 7101 -3272
rect 7525 -5248 7559 -3272
rect 7983 -5248 8017 -3272
rect 8441 -5248 8475 -3272
rect 8899 -5248 8933 -3272
rect 9013 -3660 9047 -3260
rect 10542 -3860 10602 -2940
rect 10980 -3192 11396 -3139
rect 11396 -3192 11412 -3139
rect 10864 -3518 11340 -3484
rect 10864 -3614 11340 -3580
rect 11390 -3644 11424 -3610
rect 10864 -3710 11340 -3676
rect 10864 -3806 11340 -3772
rect 11390 -3836 11424 -3802
rect 10864 -3902 11340 -3868
rect 9013 -5260 9047 -4860
rect 7129 -5332 7497 -5298
rect 7587 -5332 7955 -5298
rect 8045 -5332 8413 -5298
rect 8503 -5332 8871 -5298
rect 9459 -4338 9493 -4304
rect 9577 -4338 9611 -4304
rect 9695 -4338 9729 -4304
rect 9813 -4338 9847 -4304
rect 9931 -4338 9965 -4304
rect 10049 -4338 10083 -4304
rect 9286 -4776 9320 -4376
rect 6681 -6376 6715 -5976
rect 7311 -5650 7345 -5616
rect 7503 -5650 7537 -5616
rect 7695 -5650 7729 -5616
rect 7887 -5650 7921 -5616
rect 8079 -5650 8113 -5616
rect 8271 -5650 8305 -5616
rect 8463 -5650 8497 -5616
rect 8655 -5650 8689 -5616
rect 6909 -6200 6943 -5700
rect 7023 -6188 7057 -5712
rect 7119 -6188 7153 -5712
rect 7215 -6188 7249 -5712
rect 7311 -6188 7345 -5712
rect 7407 -6188 7441 -5712
rect 7503 -6188 7537 -5712
rect 7599 -6188 7633 -5712
rect 7695 -6188 7729 -5712
rect 7791 -6188 7825 -5712
rect 7887 -6188 7921 -5712
rect 7983 -6188 8017 -5712
rect 8079 -6188 8113 -5712
rect 8175 -6188 8209 -5712
rect 8271 -6188 8305 -5712
rect 8367 -6188 8401 -5712
rect 8463 -6188 8497 -5712
rect 8559 -6188 8593 -5712
rect 8655 -6188 8689 -5712
rect 8751 -6188 8785 -5712
rect 8847 -6188 8881 -5712
rect 8943 -6188 8977 -5712
rect 9057 -6200 9091 -5700
rect 7119 -6276 7153 -6242
rect 8847 -6276 8881 -6242
rect 5918 -6448 5952 -6414
rect 6036 -6448 6070 -6414
rect 6154 -6448 6188 -6414
rect 6272 -6448 6306 -6414
rect 6390 -6448 6424 -6414
rect 6508 -6448 6542 -6414
rect 9286 -6376 9320 -5976
rect 9400 -6364 9434 -4388
rect 9518 -6364 9552 -4388
rect 9636 -6364 9670 -4388
rect 9754 -6364 9788 -4388
rect 9872 -6364 9906 -4388
rect 9990 -6364 10024 -4388
rect 10108 -6364 10142 -4388
rect 10222 -4776 10256 -4376
rect 10222 -6376 10256 -5976
rect 9459 -6448 9493 -6414
rect 9577 -6448 9611 -6414
rect 9695 -6448 9729 -6414
rect 9813 -6448 9847 -6414
rect 9931 -6448 9965 -6414
rect 10049 -6448 10083 -6414
rect 6154 -6838 6188 -6804
rect 6272 -6838 6306 -6804
rect 6390 -6838 6424 -6804
rect 6508 -6838 6542 -6804
rect 6626 -6838 6660 -6804
rect 6744 -6838 6778 -6804
rect 6862 -6838 6896 -6804
rect 6980 -6838 7014 -6804
rect 7098 -6838 7132 -6804
rect 7216 -6838 7250 -6804
rect 7334 -6838 7368 -6804
rect 7452 -6838 7486 -6804
rect 7570 -6838 7604 -6804
rect 7688 -6838 7722 -6804
rect 7806 -6838 7840 -6804
rect 7924 -6838 7958 -6804
rect 8042 -6838 8076 -6804
rect 8160 -6838 8194 -6804
rect 8278 -6838 8312 -6804
rect 8396 -6838 8430 -6804
rect 8514 -6838 8548 -6804
rect 8632 -6838 8666 -6804
rect 8750 -6838 8784 -6804
rect 8868 -6838 8902 -6804
rect 8986 -6838 9020 -6804
rect 9104 -6838 9138 -6804
rect 9222 -6838 9256 -6804
rect 9340 -6838 9374 -6804
rect 9458 -6838 9492 -6804
rect 9576 -6838 9610 -6804
rect 9694 -6838 9728 -6804
rect 9812 -6838 9846 -6804
rect 5981 -7285 6015 -6885
rect 5981 -8885 6015 -8485
rect 6095 -8873 6129 -6897
rect 6213 -8873 6247 -6897
rect 6331 -8873 6365 -6897
rect 6449 -8873 6483 -6897
rect 6567 -8873 6601 -6897
rect 6685 -8873 6719 -6897
rect 6803 -8873 6837 -6897
rect 6921 -8873 6955 -6897
rect 7039 -8873 7073 -6897
rect 7157 -8873 7191 -6897
rect 7275 -8873 7309 -6897
rect 7393 -8873 7427 -6897
rect 7511 -8873 7545 -6897
rect 7629 -8873 7663 -6897
rect 7747 -8873 7781 -6897
rect 7865 -8873 7899 -6897
rect 7983 -8873 8017 -6897
rect 8101 -8873 8135 -6897
rect 8219 -8873 8253 -6897
rect 8337 -8873 8371 -6897
rect 8455 -8873 8489 -6897
rect 8573 -8873 8607 -6897
rect 8691 -8873 8725 -6897
rect 8809 -8873 8843 -6897
rect 8927 -8873 8961 -6897
rect 9045 -8873 9079 -6897
rect 9163 -8873 9197 -6897
rect 9281 -8873 9315 -6897
rect 9399 -8873 9433 -6897
rect 9517 -8873 9551 -6897
rect 9635 -8873 9669 -6897
rect 9753 -8873 9787 -6897
rect 9871 -8873 9905 -6897
rect 9985 -7285 10019 -6885
rect 9985 -8885 10019 -8485
rect 6154 -8966 6188 -8932
rect 6272 -8966 6306 -8932
rect 6390 -8966 6424 -8932
rect 6508 -8966 6542 -8932
rect 6626 -8966 6660 -8932
rect 6744 -8966 6778 -8932
rect 6862 -8966 6896 -8932
rect 6980 -8966 7014 -8932
rect 7098 -8966 7132 -8932
rect 7216 -8966 7250 -8932
rect 7334 -8966 7368 -8932
rect 7452 -8966 7486 -8932
rect 8514 -8966 8548 -8932
rect 8632 -8966 8666 -8932
rect 8750 -8966 8784 -8932
rect 8868 -8966 8902 -8932
rect 8986 -8966 9020 -8932
rect 9104 -8966 9138 -8932
rect 9222 -8966 9256 -8932
rect 9340 -8966 9374 -8932
rect 9458 -8966 9492 -8932
rect 9576 -8966 9610 -8932
rect 9694 -8966 9728 -8932
rect 9812 -8966 9846 -8932
<< metal1 >>
rect 6086 12366 6204 12372
rect 6086 12332 6154 12366
rect 6188 12332 6204 12366
rect 6086 12326 6204 12332
rect 6256 12366 7502 12372
rect 6256 12332 6272 12366
rect 6306 12332 6390 12366
rect 6424 12332 6508 12366
rect 6542 12332 6626 12366
rect 6660 12332 6744 12366
rect 6778 12332 6862 12366
rect 6896 12332 6980 12366
rect 7014 12332 7098 12366
rect 7132 12332 7216 12366
rect 7250 12332 7334 12366
rect 7368 12332 7452 12366
rect 7486 12332 7502 12366
rect 6256 12326 7502 12332
rect 8498 12366 9744 12372
rect 8498 12332 8514 12366
rect 8548 12332 8632 12366
rect 8666 12332 8750 12366
rect 8784 12332 8868 12366
rect 8902 12332 8986 12366
rect 9020 12332 9104 12366
rect 9138 12332 9222 12366
rect 9256 12332 9340 12366
rect 9374 12332 9458 12366
rect 9492 12332 9576 12366
rect 9610 12332 9694 12366
rect 9728 12332 9744 12366
rect 8498 12326 9744 12332
rect 9796 12366 9914 12372
rect 9796 12332 9812 12366
rect 9846 12332 9914 12366
rect 9796 12326 9914 12332
rect 5975 12285 6021 12297
rect 6086 12285 6138 12326
rect 5975 11885 5981 12285
rect 6015 12273 6138 12285
rect 6015 11885 6086 12273
rect 5975 11873 6021 11885
rect 5975 10685 6021 10697
rect 5975 10285 5981 10685
rect 6015 10297 6086 10685
rect 6015 10285 6138 10297
rect 6204 12273 6256 12285
rect 6204 10285 6256 10297
rect 6322 12273 6374 12285
rect 6322 10285 6374 10297
rect 6440 12273 6492 12285
rect 6440 10285 6492 10297
rect 6558 12273 6610 12285
rect 6558 10285 6610 10297
rect 6676 12273 6728 12285
rect 6676 10285 6728 10297
rect 6794 12273 6846 12285
rect 6794 10285 6846 10297
rect 6912 12273 6964 12285
rect 6912 10285 6964 10297
rect 7030 12273 7082 12285
rect 7030 10285 7082 10297
rect 7148 12273 7200 12285
rect 7148 10285 7200 10297
rect 7266 12273 7318 12285
rect 7266 10285 7318 10297
rect 7384 12273 7436 12326
rect 5975 10273 6021 10285
rect 6086 10244 6138 10285
rect 7384 10244 7436 10297
rect 7502 12273 7554 12285
rect 7502 10285 7554 10297
rect 7620 12273 7672 12286
rect 7620 10285 7672 10297
rect 7738 12273 7790 12285
rect 7738 10285 7790 10297
rect 7856 12273 7908 12285
rect 7856 10285 7908 10297
rect 7974 12273 8026 12285
rect 7974 10285 8026 10297
rect 8092 12273 8144 12285
rect 8092 10285 8144 10297
rect 8210 12273 8262 12285
rect 8210 10285 8262 10297
rect 8328 12273 8380 12286
rect 8328 10285 8380 10297
rect 8446 12273 8498 12285
rect 8446 10285 8498 10297
rect 8564 12273 8616 12326
rect 9862 12285 9914 12326
rect 9979 12285 10025 12297
rect 8026 10244 8092 10250
rect 8564 10244 8616 10297
rect 8682 12273 8734 12285
rect 8682 10285 8734 10297
rect 8800 12273 8852 12285
rect 8800 10285 8852 10297
rect 8918 12273 8970 12285
rect 8918 10285 8970 10297
rect 9036 12273 9088 12285
rect 9036 10285 9088 10297
rect 9154 12273 9206 12285
rect 9154 10285 9206 10297
rect 9272 12273 9324 12285
rect 9272 10285 9324 10297
rect 9390 12273 9442 12285
rect 9390 10285 9442 10297
rect 9508 12273 9560 12285
rect 9508 10285 9560 10297
rect 9626 12273 9678 12285
rect 9626 10285 9678 10297
rect 9744 12273 9796 12285
rect 9744 10284 9796 10297
rect 9862 12273 9985 12285
rect 9914 11885 9985 12273
rect 10019 11885 10025 12285
rect 9979 11873 10025 11885
rect 9979 10685 10025 10697
rect 9914 10297 9985 10685
rect 9862 10285 9985 10297
rect 10019 10285 10025 10685
rect 9862 10244 9914 10285
rect 9979 10273 10025 10285
rect 6086 10238 6204 10244
rect 6086 10204 6154 10238
rect 6188 10204 6204 10238
rect 6086 10198 6204 10204
rect 6256 10238 7502 10244
rect 6256 10204 6272 10238
rect 6306 10204 6390 10238
rect 6424 10204 6508 10238
rect 6542 10204 6626 10238
rect 6660 10204 6744 10238
rect 6778 10204 6862 10238
rect 6896 10204 6980 10238
rect 7014 10204 7098 10238
rect 7132 10204 7216 10238
rect 7250 10204 7334 10238
rect 7368 10204 7452 10238
rect 7486 10204 7502 10238
rect 6256 10198 7502 10204
rect 7554 10238 7970 10244
rect 7554 10204 7570 10238
rect 7604 10204 7688 10238
rect 7722 10204 7806 10238
rect 7840 10204 7924 10238
rect 7958 10204 7970 10238
rect 7554 10200 7970 10204
rect 7554 10198 7917 10200
rect 7911 10148 7917 10198
rect 7969 10148 7975 10200
rect 8026 10192 8032 10244
rect 8084 10238 8446 10244
rect 8084 10204 8160 10238
rect 8194 10204 8278 10238
rect 8312 10204 8396 10238
rect 8430 10204 8446 10238
rect 8084 10198 8446 10204
rect 8498 10238 9744 10244
rect 8498 10204 8514 10238
rect 8548 10204 8632 10238
rect 8666 10204 8750 10238
rect 8784 10204 8868 10238
rect 8902 10204 8986 10238
rect 9020 10204 9104 10238
rect 9138 10204 9222 10238
rect 9256 10204 9340 10238
rect 9374 10204 9458 10238
rect 9492 10204 9576 10238
rect 9610 10204 9694 10238
rect 9728 10204 9744 10238
rect 8498 10198 9744 10204
rect 9796 10238 9914 10244
rect 9796 10204 9812 10238
rect 9846 10204 9914 10238
rect 9796 10198 9914 10204
rect 8084 10192 8092 10198
rect 8026 10181 8092 10192
rect 6204 9958 6256 9964
rect 6204 9854 6256 9906
rect 9745 9958 9797 9964
rect 9745 9854 9797 9906
rect 5850 9848 5964 9854
rect 5850 9814 5918 9848
rect 5952 9814 5964 9848
rect 5850 9808 5964 9814
rect 6020 9848 6436 9854
rect 6020 9814 6036 9848
rect 6070 9814 6154 9848
rect 6188 9814 6272 9848
rect 6306 9814 6390 9848
rect 6424 9814 6436 9848
rect 6020 9808 6436 9814
rect 6496 9848 6610 9854
rect 6496 9814 6508 9848
rect 6542 9814 6610 9848
rect 6496 9808 6610 9814
rect 5739 9776 5785 9788
rect 5850 9776 5902 9808
rect 6558 9776 6610 9808
rect 9391 9848 9505 9854
rect 9391 9814 9459 9848
rect 9493 9814 9505 9848
rect 9391 9808 9505 9814
rect 9565 9848 9981 9854
rect 9565 9814 9577 9848
rect 9611 9814 9695 9848
rect 9729 9814 9813 9848
rect 9847 9814 9931 9848
rect 9965 9814 9981 9848
rect 9565 9808 9981 9814
rect 10033 9848 10151 9854
rect 10033 9814 10049 9848
rect 10083 9814 10151 9848
rect 10033 9808 10151 9814
rect 6700 9788 6800 9800
rect 6675 9776 6800 9788
rect 5170 9430 5320 9450
rect 5170 9040 5190 9430
rect 5300 9040 5320 9430
rect 5170 9020 5320 9040
rect 5400 9430 5550 9450
rect 5400 9040 5420 9430
rect 5530 9040 5550 9430
rect 5739 9376 5745 9776
rect 5779 9764 5902 9776
rect 5779 9376 5850 9764
rect 5739 9364 5785 9376
rect 5400 9020 5550 9040
rect 5739 8176 5785 8188
rect 5739 7776 5745 8176
rect 5779 7788 5850 8176
rect 5779 7776 5902 7788
rect 5968 9764 6020 9776
rect 5968 7776 6020 7788
rect 6086 9764 6138 9776
rect 6086 7776 6138 7788
rect 6204 9764 6256 9776
rect 6204 7776 6256 7788
rect 6322 9764 6374 9776
rect 6322 7776 6374 7788
rect 6440 9764 6492 9776
rect 6440 7776 6492 7788
rect 6558 9764 6681 9776
rect 6610 9376 6681 9764
rect 6715 9700 6800 9776
rect 9200 9788 9300 9800
rect 9200 9776 9326 9788
rect 9391 9776 9443 9808
rect 10099 9776 10151 9808
rect 10216 9776 10262 9788
rect 9200 9700 9286 9776
rect 6715 9600 6960 9700
rect 7017 9676 7169 9682
rect 7017 9642 7119 9676
rect 7153 9642 7169 9676
rect 7017 9636 7169 9642
rect 8831 9676 8983 9682
rect 8831 9642 8847 9676
rect 8881 9642 8983 9676
rect 8831 9636 8983 9642
rect 7017 9600 7063 9636
rect 7113 9600 7159 9636
rect 8841 9600 8887 9636
rect 8937 9600 8983 9636
rect 9040 9600 9286 9700
rect 6715 9376 6909 9600
rect 6675 9364 6909 9376
rect 6700 9200 6909 9364
rect 6800 9100 6909 9200
rect 6943 9100 7013 9600
rect 7067 9100 7073 9600
rect 7103 9100 7109 9600
rect 7163 9100 7169 9600
rect 7199 9100 7205 9600
rect 7259 9100 7265 9600
rect 7295 9100 7301 9600
rect 7355 9100 7361 9600
rect 7391 9100 7397 9600
rect 7451 9100 7457 9600
rect 7487 9100 7493 9600
rect 7547 9100 7553 9600
rect 7583 9100 7589 9600
rect 7643 9100 7649 9600
rect 7679 9100 7685 9600
rect 7739 9100 7745 9600
rect 7775 9100 7781 9600
rect 7835 9100 7841 9600
rect 7871 9100 7877 9600
rect 7931 9100 7937 9600
rect 7967 9100 7973 9600
rect 8027 9100 8033 9600
rect 8063 9100 8069 9600
rect 8123 9100 8129 9600
rect 8159 9100 8165 9600
rect 8219 9100 8225 9600
rect 8255 9100 8261 9600
rect 8315 9100 8321 9600
rect 8351 9100 8357 9600
rect 8411 9100 8417 9600
rect 8447 9100 8453 9600
rect 8507 9100 8513 9600
rect 8543 9100 8549 9600
rect 8603 9100 8609 9600
rect 8639 9100 8645 9600
rect 8699 9100 8705 9600
rect 8735 9100 8741 9600
rect 8795 9100 8801 9600
rect 8831 9100 8837 9600
rect 8891 9100 8897 9600
rect 8927 9100 8933 9600
rect 8987 9100 9057 9600
rect 9091 9376 9286 9600
rect 9320 9764 9443 9776
rect 9320 9376 9391 9764
rect 9091 9364 9326 9376
rect 9091 9200 9300 9364
rect 9091 9100 9200 9200
rect 6800 8672 6960 9100
rect 7289 9000 7295 9056
rect 7361 9000 7367 9056
rect 7481 9000 7487 9056
rect 7553 9000 7559 9056
rect 7673 9000 7679 9056
rect 7745 9000 7751 9056
rect 7865 9000 7871 9056
rect 7937 9000 7943 9056
rect 8057 9000 8063 9056
rect 8129 9000 8135 9056
rect 8249 9000 8255 9056
rect 8321 9000 8327 9056
rect 8441 9000 8447 9056
rect 8513 9000 8519 9056
rect 8633 9000 8639 9056
rect 8705 9000 8711 9056
rect 9040 8800 9200 9100
rect 8880 8762 8944 8770
rect 7117 8732 8880 8738
rect 7117 8698 7129 8732
rect 7497 8698 7587 8732
rect 7955 8698 8045 8732
rect 8413 8698 8503 8732
rect 8871 8698 8880 8732
rect 7117 8692 8944 8698
rect 8880 8690 8944 8692
rect 6800 8660 6993 8672
rect 9000 8660 9200 8800
rect 6800 8300 6953 8660
rect 6700 8260 6953 8300
rect 6987 8648 7110 8660
rect 6987 8260 7058 8648
rect 6700 8248 6993 8260
rect 6700 8188 6960 8248
rect 6675 8176 6960 8188
rect 6610 7788 6681 8176
rect 6558 7776 6681 7788
rect 6715 7776 6960 8176
rect 5739 7764 5785 7776
rect 5850 7744 5902 7776
rect 6558 7744 6610 7776
rect 6675 7764 6960 7776
rect 5850 7738 5964 7744
rect 5850 7704 5918 7738
rect 5952 7704 5964 7738
rect 5850 7698 5964 7704
rect 6020 7738 6436 7744
rect 6020 7704 6036 7738
rect 6070 7704 6154 7738
rect 6188 7704 6272 7738
rect 6306 7704 6390 7738
rect 6424 7704 6436 7738
rect 6020 7698 6436 7704
rect 6496 7738 6610 7744
rect 6496 7704 6508 7738
rect 6542 7704 6610 7738
rect 6496 7698 6610 7704
rect 6700 7700 6960 7764
rect 6800 7640 6960 7700
rect 6800 6420 6820 7640
rect 6880 7072 6960 7640
rect 6880 7060 6993 7072
rect 6880 6660 6953 7060
rect 6987 6672 7058 7060
rect 6987 6660 7110 6672
rect 7516 8648 7568 8660
rect 7516 6660 7568 6672
rect 7974 8648 8026 8660
rect 7974 6660 8026 6672
rect 8432 8648 8484 8660
rect 8432 6660 8484 6672
rect 8890 8648 9013 8660
rect 8942 8260 9013 8648
rect 9047 8300 9200 8660
rect 9047 8260 9300 8300
rect 9000 8200 9300 8260
rect 9040 8188 9300 8200
rect 9040 8176 9326 8188
rect 9040 7776 9286 8176
rect 9320 7788 9391 8176
rect 9320 7776 9443 7788
rect 9509 9764 9561 9776
rect 9509 7776 9561 7788
rect 9627 9764 9679 9776
rect 9627 7776 9679 7788
rect 9745 9764 9797 9776
rect 9745 7776 9797 7788
rect 9863 9764 9915 9776
rect 9863 7776 9915 7788
rect 9981 9764 10033 9776
rect 9981 7776 10033 7788
rect 10099 9764 10222 9776
rect 10151 9376 10222 9764
rect 10256 9376 10262 9776
rect 10216 9364 10262 9376
rect 10216 8176 10262 8188
rect 10151 7788 10222 8176
rect 10099 7776 10222 7788
rect 10256 7776 10262 8176
rect 9040 7764 9326 7776
rect 9040 7700 9300 7764
rect 9391 7744 9443 7776
rect 10099 7744 10151 7776
rect 10216 7764 10262 7776
rect 9391 7738 9505 7744
rect 9391 7704 9459 7738
rect 9493 7704 9505 7738
rect 9040 7640 9200 7700
rect 9391 7698 9505 7704
rect 9565 7738 9981 7744
rect 9565 7704 9577 7738
rect 9611 7704 9695 7738
rect 9729 7704 9813 7738
rect 9847 7704 9931 7738
rect 9965 7704 9981 7738
rect 9565 7698 9981 7704
rect 10033 7738 10151 7744
rect 10033 7704 10049 7738
rect 10083 7704 10151 7738
rect 10033 7698 10151 7704
rect 9040 7072 9120 7640
rect 9007 7060 9120 7072
rect 8942 6672 9013 7060
rect 8890 6660 9013 6672
rect 9047 6660 9120 7060
rect 6880 6648 6993 6660
rect 9007 6648 9120 6660
rect 6880 6420 6960 6648
rect 7117 6622 8883 6628
rect 7117 6588 7129 6622
rect 7497 6588 7587 6622
rect 7955 6588 8045 6622
rect 8413 6588 8503 6622
rect 8871 6588 8883 6622
rect 7117 6582 8883 6588
rect 6800 6400 6960 6420
rect 9040 6420 9120 6648
rect 9180 6420 9200 7640
rect 10744 7302 11352 7308
rect 9040 6400 9200 6420
rect 10382 7260 10622 7280
rect 10382 6340 10402 7260
rect 10602 6340 10622 7260
rect 10744 7268 10864 7302
rect 11340 7268 11352 7302
rect 10744 7262 11352 7268
rect 10744 7116 10784 7262
rect 11384 7236 11430 7252
rect 10852 7206 10867 7215
rect 11336 7206 11353 7215
rect 10852 7172 10864 7206
rect 11340 7172 11353 7206
rect 11384 7202 11390 7236
rect 11424 7206 11430 7236
rect 11424 7202 11565 7206
rect 11384 7172 11565 7202
rect 10852 7163 10867 7172
rect 11336 7163 11353 7172
rect 10744 7110 11352 7116
rect 10744 7076 10864 7110
rect 11340 7076 11352 7110
rect 10744 7070 11352 7076
rect 10744 6924 10784 7070
rect 11384 7044 11430 7060
rect 10852 7014 11352 7020
rect 10852 6980 10864 7014
rect 11340 6980 11352 7014
rect 11384 7010 11390 7044
rect 11424 7014 11430 7044
rect 11424 7010 11503 7014
rect 11384 6980 11503 7010
rect 10852 6974 11352 6980
rect 10744 6918 11352 6924
rect 10744 6884 10864 6918
rect 11340 6884 11352 6918
rect 10744 6878 11352 6884
rect 10964 6592 10983 6600
rect 10964 6539 10980 6592
rect 10964 6530 10983 6539
rect 11412 6530 11435 6600
rect 10382 6320 10622 6340
rect 11469 6316 11503 6980
rect 11463 5180 11503 6316
rect 11050 5140 11503 5180
rect 11531 6316 11565 7172
rect 11050 4920 11090 5140
rect 11531 5100 11571 6316
rect 11210 5060 11571 5100
rect 11210 4920 11250 5060
rect 11020 4910 11120 4920
rect 11020 4830 11030 4910
rect 11110 4830 11120 4910
rect 11020 4820 11120 4830
rect 11180 4910 11280 4920
rect 11180 4830 11190 4910
rect 11270 4830 11280 4910
rect 11180 4820 11280 4830
rect 3348 4352 3468 4355
rect 4374 4352 4494 4355
rect 3348 4345 3509 4352
rect 3348 3975 3358 4345
rect 3458 4340 3509 4345
rect 3458 3975 3469 4340
rect 3348 3965 3469 3975
rect 3463 3964 3469 3965
rect 3503 3964 3509 4340
rect 3463 3952 3509 3964
rect 3551 4346 3739 4352
rect 3551 4340 3671 4346
rect 3551 3964 3557 4340
rect 3591 4332 3671 4340
rect 3641 3972 3671 4332
rect 3591 3964 3671 3972
rect 3551 3958 3671 3964
rect 3705 3958 3739 4346
rect 3551 3952 3739 3958
rect 4103 4346 4291 4352
rect 4103 3958 4137 4346
rect 4171 4340 4291 4346
rect 4171 4332 4251 4340
rect 4171 3972 4201 4332
rect 4171 3964 4251 3972
rect 4285 3964 4291 4340
rect 4171 3958 4291 3964
rect 4103 3952 4291 3958
rect 4333 4345 4494 4352
rect 4333 4340 4384 4345
rect 4333 3964 4339 4340
rect 4373 3975 4384 4340
rect 4484 3975 4494 4345
rect 4373 3965 4494 3975
rect 10308 3978 14448 3998
rect 4373 3964 4379 3965
rect 4333 3952 4379 3964
rect 3497 3914 3643 3920
rect 3497 3880 3513 3914
rect 3547 3906 3643 3914
rect 3547 3880 3577 3906
rect 3497 3864 3577 3880
rect 3563 3854 3577 3864
rect 3629 3854 3643 3906
rect 3563 3840 3643 3854
rect 4199 3914 4345 3920
rect 4199 3906 4295 3914
rect 4199 3854 4213 3906
rect 4265 3880 4295 3906
rect 4329 3880 4345 3914
rect 10308 3908 11278 3978
rect 14428 3908 14448 3978
rect 10308 3888 14448 3908
rect 4265 3864 4345 3880
rect 4265 3854 4279 3864
rect 4199 3840 4279 3854
rect 11424 3824 11464 3888
rect 11776 3824 11816 3888
rect 12692 3824 12732 3888
rect 13608 3824 13648 3888
rect 11424 3818 11816 3824
rect 11424 3784 11436 3818
rect 11804 3784 11816 3818
rect 11424 3778 11816 3784
rect 11882 3818 12274 3824
rect 11882 3784 11894 3818
rect 12262 3784 12274 3818
rect 11882 3778 12274 3784
rect 12340 3818 12732 3824
rect 12340 3784 12352 3818
rect 12720 3784 12732 3818
rect 12340 3778 12732 3784
rect 12798 3818 13190 3824
rect 12798 3784 12810 3818
rect 13178 3784 13190 3818
rect 12798 3778 13190 3784
rect 13256 3818 13648 3824
rect 13256 3784 13268 3818
rect 13636 3784 13648 3818
rect 13256 3778 13648 3784
rect 11424 3737 11464 3778
rect 11365 3725 11464 3737
rect 3463 3631 3509 3638
rect 3348 3626 3509 3631
rect 3348 3621 3469 3626
rect 3348 3251 3358 3621
rect 3458 3251 3469 3621
rect 3348 3250 3469 3251
rect 3503 3250 3509 3626
rect 3348 3241 3509 3250
rect 3463 3238 3509 3241
rect 3551 3632 3739 3638
rect 3551 3626 3671 3632
rect 3551 3250 3557 3626
rect 3591 3614 3671 3626
rect 3591 3250 3671 3264
rect 3551 3244 3671 3250
rect 3705 3244 3739 3632
rect 3551 3238 3739 3244
rect 4103 3632 4291 3638
rect 4103 3244 4137 3632
rect 4171 3626 4291 3632
rect 4171 3614 4251 3626
rect 4171 3250 4251 3264
rect 4285 3250 4291 3626
rect 4171 3244 4291 3250
rect 4103 3238 4291 3244
rect 4333 3631 4379 3638
rect 4333 3626 4494 3631
rect 4333 3250 4339 3626
rect 4373 3621 4494 3626
rect 4373 3251 4384 3621
rect 4484 3251 4494 3621
rect 4373 3250 4494 3251
rect 4333 3241 4494 3250
rect 4333 3238 4379 3241
rect 3497 3200 3643 3206
rect 3497 3166 3513 3200
rect 3547 3192 3643 3200
rect 3547 3166 3577 3192
rect 3497 3150 3577 3166
rect 3563 3140 3577 3150
rect 3629 3140 3643 3192
rect 3563 3126 3643 3140
rect 4199 3200 4345 3206
rect 4199 3192 4295 3200
rect 4199 3140 4213 3192
rect 4265 3166 4295 3192
rect 4329 3166 4345 3200
rect 4265 3150 4345 3166
rect 4265 3140 4279 3150
rect 4199 3126 4279 3140
rect 2039 2920 10199 2927
rect 2039 2895 5447 2920
rect 5867 2895 6647 2920
rect 7067 2895 7847 2920
rect 8267 2895 9047 2920
rect 9467 2895 10199 2920
rect 2039 2861 2070 2895
rect 2104 2861 2166 2895
rect 2200 2861 2262 2895
rect 2296 2861 2358 2895
rect 2392 2861 2454 2895
rect 2488 2861 2550 2895
rect 2584 2861 2646 2895
rect 2680 2861 2742 2895
rect 2776 2861 2838 2895
rect 2872 2861 2934 2895
rect 2968 2861 3030 2895
rect 3064 2861 3126 2895
rect 3160 2861 3222 2895
rect 3256 2861 3318 2895
rect 3352 2861 3414 2895
rect 3448 2861 3510 2895
rect 3544 2861 3606 2895
rect 3640 2861 3702 2895
rect 3736 2861 3798 2895
rect 3832 2861 3894 2895
rect 3928 2861 3990 2895
rect 4024 2861 4086 2895
rect 4120 2861 4182 2895
rect 4216 2861 4278 2895
rect 4312 2861 4374 2895
rect 4408 2861 4470 2895
rect 4504 2861 4566 2895
rect 4600 2861 4662 2895
rect 4696 2861 4758 2895
rect 4792 2861 4854 2895
rect 4888 2861 4950 2895
rect 4984 2861 5046 2895
rect 5080 2861 5142 2895
rect 5176 2861 5238 2895
rect 5272 2861 5334 2895
rect 5368 2861 5430 2895
rect 5867 2861 5910 2895
rect 5944 2861 6006 2895
rect 6040 2861 6102 2895
rect 6136 2861 6198 2895
rect 6232 2861 6294 2895
rect 6328 2861 6390 2895
rect 6424 2861 6486 2895
rect 6520 2861 6582 2895
rect 6616 2861 6647 2895
rect 7096 2861 7158 2895
rect 7192 2861 7254 2895
rect 7288 2861 7350 2895
rect 7384 2861 7446 2895
rect 7480 2861 7542 2895
rect 7576 2861 7638 2895
rect 7672 2861 7734 2895
rect 7768 2861 7830 2895
rect 8267 2861 8310 2895
rect 8344 2861 8406 2895
rect 8440 2861 8502 2895
rect 8536 2861 8598 2895
rect 8632 2861 8694 2895
rect 8728 2861 8790 2895
rect 8824 2861 8886 2895
rect 8920 2861 8982 2895
rect 9016 2861 9047 2895
rect 9496 2861 9558 2895
rect 9592 2861 9654 2895
rect 9688 2861 9750 2895
rect 9784 2861 9846 2895
rect 9880 2861 9942 2895
rect 9976 2861 10038 2895
rect 10072 2861 10134 2895
rect 10168 2861 10199 2895
rect 2039 2840 5447 2861
rect 5867 2840 6647 2861
rect 7067 2840 7847 2861
rect 8267 2840 9047 2861
rect 9467 2840 10199 2861
rect 2039 2829 10199 2840
rect 5319 2784 5383 2793
rect 5319 2750 5334 2784
rect 5368 2750 5383 2784
rect 5319 2741 5383 2750
rect 2530 2670 4034 2736
rect 2530 2553 2596 2670
rect 2426 2531 2596 2553
rect 2353 2479 2359 2531
rect 2411 2479 2431 2531
rect 2483 2487 2596 2531
rect 2697 2613 3118 2619
rect 2483 2479 2489 2487
rect 2697 2363 2709 2613
rect 3106 2363 3118 2613
rect 2697 2357 3118 2363
rect 3228 2613 3649 2619
rect 3228 2363 3240 2613
rect 3637 2363 3649 2613
rect 3968 2506 4034 2670
rect 3968 2472 3984 2506
rect 4018 2472 4034 2506
rect 3968 2456 4034 2472
rect 3228 2357 3649 2363
rect 3965 2347 4017 2358
rect 5223 2340 5287 2349
rect 5223 2306 5238 2340
rect 5272 2306 5287 2340
rect 5223 2297 5287 2306
rect 3965 2289 4017 2295
rect 2039 2260 10199 2261
rect 2039 2229 4747 2260
rect 5167 2240 10199 2260
rect 5167 2229 6047 2240
rect 6467 2229 7247 2240
rect 7667 2229 8447 2240
rect 8867 2229 9647 2240
rect 10067 2229 10199 2240
rect 2039 2195 2070 2229
rect 2104 2195 2166 2229
rect 2200 2195 2262 2229
rect 2296 2195 2358 2229
rect 2392 2195 2454 2229
rect 2488 2195 2550 2229
rect 2584 2195 2646 2229
rect 2680 2195 2742 2229
rect 2776 2195 2838 2229
rect 2872 2195 2934 2229
rect 2968 2195 3030 2229
rect 3064 2195 3126 2229
rect 3160 2195 3222 2229
rect 3256 2195 3318 2229
rect 3352 2195 3414 2229
rect 3448 2195 3510 2229
rect 3544 2195 3606 2229
rect 3640 2195 3702 2229
rect 3736 2195 3798 2229
rect 3832 2195 3894 2229
rect 3928 2195 3990 2229
rect 4024 2195 4086 2229
rect 4120 2195 4182 2229
rect 4216 2195 4278 2229
rect 4312 2195 4374 2229
rect 4408 2195 4470 2229
rect 4504 2195 4566 2229
rect 4600 2195 4662 2229
rect 4696 2195 4747 2229
rect 5176 2195 5238 2229
rect 5272 2195 5334 2229
rect 5368 2195 5430 2229
rect 5464 2195 5526 2229
rect 5560 2195 5622 2229
rect 5656 2195 5718 2229
rect 5752 2195 5814 2229
rect 5848 2195 5910 2229
rect 5944 2195 6006 2229
rect 6040 2195 6047 2229
rect 6467 2195 6486 2229
rect 6520 2195 6582 2229
rect 6616 2195 6678 2229
rect 6712 2195 6774 2229
rect 6808 2195 6870 2229
rect 6904 2195 6966 2229
rect 7000 2195 7062 2229
rect 7096 2195 7158 2229
rect 7192 2195 7247 2229
rect 7672 2195 7734 2229
rect 7768 2195 7830 2229
rect 7864 2195 7926 2229
rect 7960 2195 8022 2229
rect 8056 2195 8118 2229
rect 8152 2195 8214 2229
rect 8248 2195 8310 2229
rect 8344 2195 8406 2229
rect 8440 2195 8447 2229
rect 8867 2195 8886 2229
rect 8920 2195 8982 2229
rect 9016 2195 9078 2229
rect 9112 2195 9174 2229
rect 9208 2195 9270 2229
rect 9304 2195 9366 2229
rect 9400 2195 9462 2229
rect 9496 2195 9558 2229
rect 9592 2195 9647 2229
rect 10072 2195 10134 2229
rect 10168 2195 10199 2229
rect 2039 2180 4747 2195
rect 5167 2180 6047 2195
rect 6467 2180 7247 2195
rect 7667 2180 8447 2195
rect 8867 2180 9647 2195
rect 10067 2180 10199 2195
rect 2039 2163 10199 2180
rect 3965 2129 4017 2135
rect 2697 2061 3118 2067
rect 2353 1893 2359 1945
rect 2411 1893 2431 1945
rect 2483 1937 2489 1945
rect 2483 1893 2596 1937
rect 2426 1871 2596 1893
rect 2530 1754 2596 1871
rect 2697 1811 2709 2061
rect 3106 1811 3118 2061
rect 2697 1805 3118 1811
rect 3228 2061 3649 2067
rect 3965 2066 4017 2077
rect 5223 2118 5287 2127
rect 5223 2084 5238 2118
rect 5272 2084 5287 2118
rect 5223 2075 5287 2084
rect 10818 2108 10898 2118
rect 3228 1811 3240 2061
rect 3637 1811 3649 2061
rect 6570 1970 6628 1976
rect 3228 1805 3649 1811
rect 3968 1952 4034 1968
rect 3968 1918 3984 1952
rect 4018 1918 4034 1952
rect 3968 1754 4034 1918
rect 4156 1886 4162 1938
rect 4214 1886 4220 1938
rect 4433 1909 4439 1961
rect 4491 1909 4497 1961
rect 4547 1911 4553 1963
rect 4605 1911 4611 1963
rect 4940 1898 4946 1950
rect 4998 1898 5004 1950
rect 6570 1936 6582 1970
rect 6616 1967 6628 1970
rect 7434 1970 7492 1976
rect 7434 1967 7446 1970
rect 6616 1939 7446 1967
rect 6616 1936 6628 1939
rect 5704 1905 5762 1914
rect 5704 1871 5716 1905
rect 5750 1871 5762 1905
rect 6109 1883 6115 1935
rect 6167 1883 6173 1935
rect 6570 1930 6628 1936
rect 7434 1936 7446 1939
rect 7480 1936 7492 1970
rect 7434 1930 7492 1936
rect 7242 1896 7300 1902
rect 5704 1862 5762 1871
rect 7242 1862 7254 1896
rect 7288 1893 7300 1896
rect 7818 1896 7876 1902
rect 7818 1893 7830 1896
rect 7288 1865 7830 1893
rect 7288 1862 7300 1865
rect 2530 1688 4034 1754
rect 4832 1724 4838 1776
rect 4890 1724 4896 1776
rect 5040 1704 5092 1710
rect 5040 1646 5092 1652
rect 5319 1674 5383 1683
rect 5319 1640 5334 1674
rect 5368 1640 5383 1674
rect 5319 1631 5383 1640
rect 5708 1595 5754 1862
rect 7242 1856 7300 1862
rect 7818 1862 7830 1865
rect 7864 1862 7876 1896
rect 7818 1856 7876 1862
rect 7839 1595 7867 1856
rect 8188 1851 8194 1903
rect 8246 1851 8252 1903
rect 9474 1883 9480 1935
rect 9532 1883 9552 1935
rect 9604 1883 9610 1935
rect 9861 1883 9867 1935
rect 9919 1883 9939 1935
rect 9991 1883 9997 1935
rect 10180 1930 10280 1950
rect 10180 1850 10200 1930
rect 10260 1850 10280 1930
rect 8878 1832 8930 1838
rect 10180 1830 10280 1850
rect 8878 1760 8930 1780
rect 8878 1702 8930 1708
rect 10818 1678 10828 2108
rect 10888 1678 10898 2108
rect 10818 1668 10898 1678
rect 10988 2108 11068 2118
rect 10988 1678 10998 2108
rect 11058 1678 11068 2108
rect 11417 3701 11464 3725
rect 11776 3737 11816 3778
rect 12228 3748 12268 3778
rect 12228 3737 12308 3748
rect 12692 3737 12732 3778
rect 13608 3737 13648 3778
rect 14328 3737 14408 3888
rect 11776 3725 11875 3737
rect 11776 3701 11823 3725
rect 11417 1749 11464 1828
rect 11365 1737 11464 1749
rect 10988 1668 11068 1678
rect 11424 1696 11464 1737
rect 11776 1749 11823 1819
rect 12228 3725 12333 3737
rect 12228 3668 12281 3725
rect 11776 1737 11875 1749
rect 12238 1749 12281 1818
rect 12692 3725 12791 3737
rect 12692 3655 12739 3725
rect 12238 1737 12333 1749
rect 12692 1749 12739 1819
rect 13197 3725 13249 3737
rect 13188 1768 13197 1958
rect 12692 1737 12791 1749
rect 13608 3725 13704 3737
rect 13886 3728 13932 3737
rect 13608 3655 13664 3725
rect 13249 1948 13268 1958
rect 13258 1778 13268 1948
rect 13658 1819 13664 3655
rect 13249 1768 13268 1778
rect 13197 1737 13249 1749
rect 13608 1749 13664 1819
rect 13698 1749 13704 3725
rect 13608 1737 13704 1749
rect 13848 3725 13932 3728
rect 13848 2098 13892 3725
rect 13848 1888 13858 2098
rect 13848 1749 13892 1888
rect 13926 1749 13932 3725
rect 13848 1748 13932 1749
rect 13886 1737 13932 1748
rect 13974 3728 14020 3737
rect 14202 3728 14248 3737
rect 13974 3725 14058 3728
rect 13974 1749 13980 3725
rect 14014 2338 14058 3725
rect 14168 3725 14248 3728
rect 14014 2328 14068 2338
rect 14048 2118 14068 2328
rect 14014 2108 14068 2118
rect 14014 1749 14058 2108
rect 14168 1790 14208 3725
rect 13974 1748 14058 1749
rect 14116 1749 14208 1790
rect 14242 1749 14248 3725
rect 13974 1737 14020 1748
rect 14116 1746 14248 1749
rect 11776 1696 11816 1737
rect 12238 1728 12298 1737
rect 12238 1698 12278 1728
rect 11424 1690 11816 1696
rect 11424 1656 11436 1690
rect 11804 1656 11816 1690
rect 11424 1650 11816 1656
rect 11878 1690 12278 1698
rect 12692 1696 12732 1737
rect 12810 1698 13180 1700
rect 11878 1656 11894 1690
rect 12262 1656 12278 1690
rect 11878 1638 12278 1656
rect 12340 1690 12732 1696
rect 12340 1656 12352 1690
rect 12720 1656 12732 1690
rect 12340 1650 12732 1656
rect 12798 1690 13198 1698
rect 13608 1696 13648 1737
rect 12798 1656 12810 1690
rect 13178 1656 13198 1690
rect 2039 1580 10199 1595
rect 2039 1563 5447 1580
rect 5867 1563 6647 1580
rect 7067 1563 7847 1580
rect 8267 1563 9047 1580
rect 9467 1563 10199 1580
rect 11878 1578 12108 1638
rect 12208 1618 12278 1638
rect 12798 1618 12820 1656
rect 12208 1610 12820 1618
rect 13170 1610 13198 1656
rect 13256 1690 13648 1696
rect 13256 1656 13268 1690
rect 13636 1656 13648 1690
rect 13256 1650 13648 1656
rect 13908 1698 13988 1708
rect 13908 1638 13918 1698
rect 13978 1638 13988 1698
rect 13908 1628 13988 1638
rect 12208 1578 13198 1610
rect 2039 1529 2070 1563
rect 2104 1529 2166 1563
rect 2200 1529 2262 1563
rect 2296 1529 2358 1563
rect 2392 1529 2454 1563
rect 2488 1529 2550 1563
rect 2584 1529 2646 1563
rect 2680 1529 2742 1563
rect 2776 1529 2838 1563
rect 2872 1529 2934 1563
rect 2968 1529 3030 1563
rect 3064 1529 3126 1563
rect 3160 1529 3222 1563
rect 3256 1529 3318 1563
rect 3352 1529 3414 1563
rect 3448 1529 3510 1563
rect 3544 1529 3606 1563
rect 3640 1529 3702 1563
rect 3736 1529 3798 1563
rect 3832 1529 3894 1563
rect 3928 1529 3990 1563
rect 4024 1529 4086 1563
rect 4120 1529 4182 1563
rect 4216 1529 4278 1563
rect 4312 1529 4374 1563
rect 4408 1529 4470 1563
rect 4504 1529 4566 1563
rect 4600 1529 4662 1563
rect 4696 1529 4758 1563
rect 4792 1529 4854 1563
rect 4888 1529 4950 1563
rect 4984 1529 5046 1563
rect 5080 1529 5142 1563
rect 5176 1529 5238 1563
rect 5272 1529 5334 1563
rect 5368 1529 5430 1563
rect 5867 1529 5910 1563
rect 5944 1529 6006 1563
rect 6040 1529 6102 1563
rect 6136 1529 6198 1563
rect 6232 1529 6294 1563
rect 6328 1529 6390 1563
rect 6424 1529 6486 1563
rect 6520 1529 6582 1563
rect 6616 1529 6647 1563
rect 7096 1529 7158 1563
rect 7192 1529 7254 1563
rect 7288 1529 7350 1563
rect 7384 1529 7446 1563
rect 7480 1529 7542 1563
rect 7576 1529 7638 1563
rect 7672 1529 7734 1563
rect 7768 1529 7830 1563
rect 8267 1529 8310 1563
rect 8344 1529 8406 1563
rect 8440 1529 8502 1563
rect 8536 1529 8598 1563
rect 8632 1529 8694 1563
rect 8728 1529 8790 1563
rect 8824 1529 8886 1563
rect 8920 1529 8982 1563
rect 9016 1529 9047 1563
rect 9496 1529 9558 1563
rect 9592 1529 9654 1563
rect 9688 1529 9750 1563
rect 9784 1529 9846 1563
rect 9880 1529 9942 1563
rect 9976 1529 10038 1563
rect 10072 1529 10134 1563
rect 10168 1529 10199 1563
rect 14116 1548 14160 1746
rect 14202 1737 14248 1746
rect 14290 3725 14408 3737
rect 14290 1749 14296 3725
rect 14330 1749 14408 3725
rect 14290 1748 14408 1749
rect 14290 1737 14336 1748
rect 14238 1698 14318 1708
rect 14238 1638 14248 1698
rect 14308 1638 14318 1698
rect 14238 1628 14318 1638
rect 2039 1520 5447 1529
rect 5867 1520 6647 1529
rect 7067 1520 7847 1529
rect 8267 1520 9047 1529
rect 9467 1520 10199 1529
rect 2039 1498 10199 1520
rect 1767 1497 10199 1498
rect 13828 1498 14160 1548
rect 1767 1467 2871 1497
rect 1767 1433 1796 1467
rect 1830 1433 1888 1467
rect 1922 1433 1980 1467
rect 2014 1433 2072 1467
rect 2106 1433 2164 1467
rect 2198 1433 2256 1467
rect 2290 1433 2348 1467
rect 2382 1433 2440 1467
rect 2474 1433 2532 1467
rect 2566 1433 2624 1467
rect 2658 1433 2716 1467
rect 2750 1433 2808 1467
rect 2842 1433 2871 1467
rect 1767 1402 2871 1433
rect 5319 1452 5383 1461
rect 5319 1418 5334 1452
rect 5368 1418 5383 1452
rect 5319 1409 5383 1418
rect 3682 1338 5186 1404
rect 1880 1220 2020 1240
rect 1880 1167 1900 1220
rect 1876 1158 1900 1167
rect 2000 1167 2020 1220
rect 2240 1220 2380 1240
rect 2000 1158 2026 1167
rect 1876 1118 1891 1158
rect 2011 1118 2026 1158
rect 1876 1109 2026 1118
rect 2240 1158 2260 1220
rect 2360 1167 2380 1220
rect 2620 1220 2760 1240
rect 3682 1221 3748 1338
rect 2620 1167 2640 1220
rect 2360 1158 2394 1167
rect 2240 1118 2259 1158
rect 2379 1118 2394 1158
rect 2240 1109 2394 1118
rect 2612 1158 2640 1167
rect 2740 1167 2760 1220
rect 3578 1199 3748 1221
rect 2740 1158 2762 1167
rect 2612 1118 2627 1158
rect 2747 1118 2762 1158
rect 3505 1147 3511 1199
rect 3563 1147 3583 1199
rect 3635 1155 3748 1199
rect 3849 1281 4270 1287
rect 3635 1147 3641 1155
rect 2612 1109 2762 1118
rect 1880 1100 2020 1109
rect 2240 1100 2380 1109
rect 2620 1100 2760 1109
rect 3849 1031 3861 1281
rect 4258 1031 4270 1281
rect 3849 1025 4270 1031
rect 4380 1281 4801 1287
rect 4380 1031 4392 1281
rect 4789 1031 4801 1281
rect 5120 1174 5186 1338
rect 7839 1236 7867 1497
rect 10958 1440 13188 1458
rect 10958 1418 12820 1440
rect 10458 1386 10518 1388
rect 8472 1379 8524 1385
rect 8472 1307 8524 1327
rect 8472 1249 8524 1255
rect 8881 1375 8933 1381
rect 8881 1303 8933 1323
rect 10458 1380 10928 1386
rect 10458 1346 10520 1380
rect 10888 1346 10928 1380
rect 10958 1380 11358 1418
rect 10958 1378 10978 1380
rect 10458 1340 10928 1346
rect 10966 1346 10978 1378
rect 11346 1346 11358 1380
rect 10966 1340 11358 1346
rect 11424 1380 11816 1386
rect 11424 1346 11436 1380
rect 11804 1346 11816 1380
rect 11424 1340 11816 1346
rect 10458 1338 10518 1340
rect 10458 1308 10488 1338
rect 10888 1308 10928 1340
rect 11318 1308 11358 1340
rect 11776 1309 11816 1340
rect 11878 1380 12278 1418
rect 11878 1346 11894 1380
rect 12262 1346 12278 1380
rect 11878 1338 12278 1346
rect 12340 1380 12732 1386
rect 12340 1346 12352 1380
rect 12720 1346 12732 1380
rect 12340 1340 12732 1346
rect 11776 1308 11833 1309
rect 12692 1308 12732 1340
rect 12798 1380 12820 1418
rect 13170 1386 13188 1440
rect 13170 1380 13190 1386
rect 12798 1346 12810 1380
rect 13178 1346 13190 1380
rect 12798 1340 13190 1346
rect 13256 1380 13648 1386
rect 13256 1346 13268 1380
rect 13636 1346 13648 1380
rect 13256 1340 13648 1346
rect 12798 1338 13188 1340
rect 13608 1308 13648 1340
rect 13828 1308 13868 1498
rect 14130 1496 14160 1498
rect 13908 1408 13988 1418
rect 13908 1348 13918 1408
rect 13978 1348 13988 1408
rect 13908 1346 13936 1348
rect 13970 1346 13988 1348
rect 13908 1338 13988 1346
rect 14238 1408 14318 1418
rect 14238 1348 14248 1408
rect 14308 1348 14318 1408
rect 14238 1346 14252 1348
rect 14286 1346 14318 1348
rect 14238 1338 14318 1346
rect 10449 1296 10501 1308
rect 8881 1245 8933 1251
rect 5697 1179 5703 1231
rect 5755 1179 5761 1231
rect 7242 1230 7300 1236
rect 5120 1140 5136 1174
rect 5170 1140 5186 1174
rect 6113 1157 6119 1209
rect 6171 1157 6177 1209
rect 7242 1196 7254 1230
rect 7288 1227 7300 1230
rect 7818 1230 7876 1236
rect 7818 1227 7830 1230
rect 7288 1199 7830 1227
rect 7288 1196 7300 1199
rect 7242 1190 7300 1196
rect 7818 1196 7830 1199
rect 7864 1196 7876 1230
rect 7818 1190 7876 1196
rect 8190 1190 8196 1242
rect 8248 1190 8254 1242
rect 10180 1240 10280 1260
rect 9452 1230 9518 1236
rect 9452 1178 9460 1230
rect 9512 1178 9518 1230
rect 9452 1170 9518 1178
rect 9579 1171 9585 1223
rect 9637 1171 9657 1223
rect 5120 1124 5186 1140
rect 6570 1156 6628 1162
rect 6570 1122 6582 1156
rect 6616 1153 6628 1156
rect 7434 1156 7492 1162
rect 7434 1153 7446 1156
rect 6616 1125 7446 1153
rect 6616 1122 6628 1125
rect 6570 1116 6628 1122
rect 7434 1122 7446 1125
rect 7480 1122 7492 1156
rect 10180 1160 10200 1240
rect 10260 1160 10280 1240
rect 10180 1140 10280 1160
rect 7434 1116 7492 1122
rect 4380 1025 4801 1031
rect 5117 1015 5169 1026
rect 5223 1008 5287 1017
rect 5223 974 5238 1008
rect 5272 974 5287 1008
rect 5223 965 5287 974
rect 5117 957 5169 963
rect 1680 929 3287 954
rect 1680 923 10199 929
rect 1680 920 1796 923
rect 1680 858 1740 920
rect 1830 889 1888 923
rect 1922 889 1980 923
rect 2014 889 2072 923
rect 2106 920 2164 923
rect 2160 889 2164 920
rect 2198 889 2256 923
rect 2290 889 2348 923
rect 2382 889 2440 923
rect 2474 889 2532 923
rect 2566 889 2624 923
rect 2658 889 2716 923
rect 2750 889 2808 923
rect 2842 900 10199 923
rect 2842 897 6047 900
rect 6467 897 7247 900
rect 7667 897 8447 900
rect 8867 897 9647 900
rect 10067 897 10199 900
rect 2842 889 3222 897
rect 1720 800 1740 858
rect 1820 858 2080 889
rect 1820 800 1840 858
rect 1720 780 1840 800
rect 2060 800 2080 858
rect 2160 863 3222 889
rect 3256 863 3318 897
rect 3352 863 3414 897
rect 3448 863 3510 897
rect 3544 863 3606 897
rect 3640 863 3702 897
rect 3736 863 3798 897
rect 3832 863 3894 897
rect 3928 863 3990 897
rect 4024 863 4086 897
rect 4120 863 4182 897
rect 4216 863 4278 897
rect 4312 863 4374 897
rect 4408 863 4470 897
rect 4504 863 4566 897
rect 4600 863 4662 897
rect 4696 863 4758 897
rect 4792 863 4854 897
rect 4888 863 4950 897
rect 4984 863 5046 897
rect 5080 863 5142 897
rect 5176 863 5238 897
rect 5272 863 5334 897
rect 5368 863 5430 897
rect 5464 863 5526 897
rect 5560 863 5622 897
rect 5656 863 5718 897
rect 5752 863 5814 897
rect 5848 863 5910 897
rect 5944 863 6006 897
rect 6040 863 6047 897
rect 6467 863 6486 897
rect 6520 863 6582 897
rect 6616 863 6678 897
rect 6712 863 6774 897
rect 6808 863 6870 897
rect 6904 863 6966 897
rect 7000 863 7062 897
rect 7096 863 7158 897
rect 7192 863 7247 897
rect 7672 863 7734 897
rect 7768 863 7830 897
rect 7864 863 7926 897
rect 7960 863 8022 897
rect 8056 863 8118 897
rect 8152 863 8214 897
rect 8248 863 8310 897
rect 8344 863 8406 897
rect 8440 863 8447 897
rect 8867 863 8886 897
rect 8920 863 8982 897
rect 9016 863 9078 897
rect 9112 863 9174 897
rect 9208 863 9270 897
rect 9304 863 9366 897
rect 9400 863 9462 897
rect 9496 863 9558 897
rect 9592 863 9647 897
rect 10072 863 10134 897
rect 10168 863 10199 897
rect 2160 858 6047 863
rect 2160 800 2180 858
rect 3191 840 6047 858
rect 6467 840 7247 863
rect 7667 840 8447 863
rect 8867 840 9647 863
rect 10067 840 10199 863
rect 3191 831 10199 840
rect 2060 780 2180 800
rect 3941 582 4061 585
rect 3670 576 3858 582
rect 3670 188 3704 576
rect 3738 570 3858 576
rect 3738 562 3818 570
rect 3738 202 3768 562
rect 3738 194 3818 202
rect 3852 194 3858 570
rect 3738 188 3858 194
rect 3670 182 3858 188
rect 3900 575 4061 582
rect 3900 570 3951 575
rect 3900 194 3906 570
rect 3940 205 3951 570
rect 4051 205 4061 575
rect 10888 1296 10959 1308
rect 10888 1278 10907 1296
rect 10449 308 10501 320
rect 10860 320 10907 374
rect 11318 1296 11417 1308
rect 11318 1218 11365 1296
rect 10860 308 10959 320
rect 11318 320 11365 398
rect 11776 1296 11875 1308
rect 11776 1218 11823 1296
rect 11318 308 11417 320
rect 11776 320 11823 399
rect 12281 1296 12333 1308
rect 12268 1268 12281 1278
rect 12268 1168 12278 1268
rect 12268 1158 12281 1168
rect 11776 308 11875 320
rect 12692 1296 12791 1308
rect 12333 1268 12348 1278
rect 12338 1168 12348 1268
rect 12692 1217 12739 1296
rect 12333 1158 12348 1168
rect 12281 308 12333 320
rect 12692 320 12739 399
rect 13197 1296 13249 1308
rect 13188 1088 13197 1278
rect 12692 308 12791 320
rect 13608 1296 13704 1308
rect 13249 1268 13268 1278
rect 13258 1098 13268 1268
rect 13608 1242 13664 1296
rect 13249 1088 13268 1098
rect 13658 374 13664 1242
rect 13197 308 13249 320
rect 13608 320 13664 374
rect 13698 320 13704 1296
rect 13828 1296 13932 1308
rect 13828 1158 13892 1296
rect 13608 308 13704 320
rect 13848 948 13858 1158
rect 13848 320 13892 948
rect 13926 320 13932 1296
rect 13848 318 13932 320
rect 13886 308 13932 318
rect 13974 1296 14058 1308
rect 13974 320 13980 1296
rect 14014 938 14058 1296
rect 14158 1298 14248 1308
rect 14158 1238 14168 1298
rect 14228 1296 14248 1298
rect 14158 1228 14208 1238
rect 14014 928 14068 938
rect 14058 718 14068 928
rect 14014 708 14068 718
rect 14014 320 14058 708
rect 13974 318 14058 320
rect 14168 320 14208 1228
rect 14242 320 14248 1296
rect 14168 318 14248 320
rect 13974 308 14020 318
rect 14202 308 14248 318
rect 14290 1298 14336 1308
rect 14290 1296 14408 1298
rect 14290 320 14296 1296
rect 14330 320 14408 1296
rect 39370 1035 39390 1040
rect 39369 1029 39390 1035
rect 39770 1029 39790 1040
rect 37681 1012 38071 1022
rect 15547 1002 15927 1012
rect 15547 912 15557 1002
rect 15917 912 15927 1002
rect 15547 907 15927 912
rect 16261 1002 16641 1012
rect 16261 912 16271 1002
rect 16631 912 16641 1002
rect 16261 907 16641 912
rect 16975 1002 17355 1012
rect 16975 912 16985 1002
rect 17345 912 17355 1002
rect 16975 907 17355 912
rect 17689 1002 18069 1012
rect 17689 912 17699 1002
rect 18059 912 18069 1002
rect 17689 907 18069 912
rect 18403 1002 18783 1012
rect 18403 912 18413 1002
rect 18773 912 18783 1002
rect 18403 907 18783 912
rect 19117 1002 19497 1012
rect 19117 912 19127 1002
rect 19487 912 19497 1002
rect 19117 907 19497 912
rect 19831 1002 20211 1012
rect 19831 912 19841 1002
rect 20201 912 20211 1002
rect 19831 907 20211 912
rect 20545 1002 20925 1012
rect 20545 912 20555 1002
rect 20915 912 20925 1002
rect 20545 907 20925 912
rect 21259 1002 21639 1012
rect 21259 912 21269 1002
rect 21629 912 21639 1002
rect 21259 907 21639 912
rect 21973 1002 22353 1012
rect 21973 912 21983 1002
rect 22343 912 22353 1002
rect 21973 907 22353 912
rect 22687 1002 23067 1012
rect 22687 912 22697 1002
rect 23057 912 23067 1002
rect 22687 907 23067 912
rect 23401 1002 23781 1012
rect 23401 912 23411 1002
rect 23771 912 23781 1002
rect 23401 907 23781 912
rect 24115 1002 24495 1012
rect 24115 912 24125 1002
rect 24485 912 24495 1002
rect 24115 907 24495 912
rect 24829 1002 25209 1012
rect 24829 912 24839 1002
rect 25199 912 25209 1002
rect 24829 907 25209 912
rect 25543 1002 25923 1012
rect 25543 912 25553 1002
rect 25913 912 25923 1002
rect 25543 907 25923 912
rect 26257 1002 26637 1012
rect 26257 912 26267 1002
rect 26627 912 26637 1002
rect 26257 907 26637 912
rect 26971 1002 27351 1012
rect 26971 912 26981 1002
rect 27341 912 27351 1002
rect 26971 907 27351 912
rect 27685 1002 28065 1012
rect 27685 912 27695 1002
rect 28055 912 28065 1002
rect 27685 907 28065 912
rect 28399 1002 28779 1012
rect 28399 912 28409 1002
rect 28769 912 28779 1002
rect 28399 907 28779 912
rect 29113 1002 29493 1012
rect 29113 912 29123 1002
rect 29483 912 29493 1002
rect 29113 907 29493 912
rect 29827 1002 30207 1012
rect 29827 912 29837 1002
rect 30197 912 30207 1002
rect 29827 907 30207 912
rect 30541 1002 30921 1012
rect 30541 912 30551 1002
rect 30911 912 30921 1002
rect 30541 907 30921 912
rect 31255 1002 31635 1012
rect 31255 912 31265 1002
rect 31625 912 31635 1002
rect 31255 907 31635 912
rect 31969 1002 32349 1012
rect 31969 912 31979 1002
rect 32339 912 32349 1002
rect 31969 907 32349 912
rect 32683 1002 33063 1012
rect 32683 912 32693 1002
rect 33053 912 33063 1002
rect 32683 907 33063 912
rect 33397 1002 33777 1012
rect 33397 912 33407 1002
rect 33767 912 33777 1002
rect 33397 907 33777 912
rect 34111 1002 34491 1012
rect 34111 912 34121 1002
rect 34481 912 34491 1002
rect 34111 907 34491 912
rect 34825 1002 35205 1012
rect 34825 912 34835 1002
rect 35195 912 35205 1002
rect 34825 907 35205 912
rect 35539 1002 35919 1012
rect 35539 912 35549 1002
rect 35909 912 35919 1002
rect 35539 907 35919 912
rect 36253 1002 36633 1012
rect 36253 912 36263 1002
rect 36623 912 36633 1002
rect 36253 907 36633 912
rect 36967 1002 37347 1012
rect 36967 912 36977 1002
rect 37337 912 37347 1002
rect 36967 907 37347 912
rect 37681 912 37691 1012
rect 38061 912 38071 1012
rect 37681 907 38071 912
rect 38385 1012 38775 1022
rect 38385 912 38395 1012
rect 38765 912 38775 1012
rect 39369 991 39381 1029
rect 39778 991 39790 1029
rect 39369 985 39390 991
rect 39370 980 39390 985
rect 39770 980 39790 991
rect 39900 1029 39920 1040
rect 40300 1035 40320 1040
rect 40300 1029 40321 1035
rect 39900 991 39912 1029
rect 40309 991 40321 1029
rect 39900 980 39920 991
rect 40300 985 40321 991
rect 40300 980 40320 985
rect 38385 907 38775 912
rect 15540 901 15940 907
rect 15540 867 15552 901
rect 15928 867 15940 901
rect 16254 901 16654 907
rect 15540 861 15940 867
rect 15972 857 16028 873
rect 16254 867 16266 901
rect 16642 867 16654 901
rect 16968 901 17368 907
rect 16254 861 16654 867
rect 15972 823 15978 857
rect 16012 823 16028 857
rect 15540 813 15940 819
rect 15540 779 15552 813
rect 15928 779 15940 813
rect 15540 733 15558 779
rect 15918 733 15940 779
rect 15540 699 15940 733
rect 15972 807 16028 823
rect 16686 857 16742 873
rect 16968 867 16980 901
rect 17356 867 17368 901
rect 17682 901 18082 907
rect 16968 861 17368 867
rect 16686 823 16692 857
rect 16726 823 16742 857
rect 16254 813 16654 819
rect 15972 793 16052 807
rect 15972 741 15986 793
rect 16038 741 16052 793
rect 15972 727 16052 741
rect 16254 779 16266 813
rect 16642 779 16654 813
rect 16254 733 16272 779
rect 16632 733 16654 779
rect 15540 665 15546 699
rect 15934 665 15940 699
rect 15540 649 15940 665
rect 16254 699 16654 733
rect 16686 807 16742 823
rect 17400 857 17456 873
rect 17682 867 17694 901
rect 18070 867 18082 901
rect 18396 901 18796 907
rect 17682 861 18082 867
rect 17400 823 17406 857
rect 17440 823 17456 857
rect 16968 813 17368 819
rect 16686 793 16766 807
rect 16686 741 16700 793
rect 16752 741 16766 793
rect 16686 727 16766 741
rect 16968 779 16980 813
rect 17356 779 17368 813
rect 16968 733 16986 779
rect 17346 733 17368 779
rect 16254 665 16260 699
rect 16648 665 16654 699
rect 16254 649 16654 665
rect 16968 699 17368 733
rect 17400 807 17456 823
rect 18114 857 18170 873
rect 18396 867 18408 901
rect 18784 867 18796 901
rect 19110 901 19510 907
rect 18396 861 18796 867
rect 18114 823 18120 857
rect 18154 823 18170 857
rect 17682 813 18082 819
rect 17400 793 17480 807
rect 17400 741 17414 793
rect 17466 741 17480 793
rect 17400 727 17480 741
rect 17682 779 17694 813
rect 18070 779 18082 813
rect 17682 733 17700 779
rect 18060 733 18082 779
rect 16968 665 16974 699
rect 17362 665 17368 699
rect 16968 649 17368 665
rect 17682 699 18082 733
rect 18114 807 18170 823
rect 18828 857 18884 873
rect 19110 867 19122 901
rect 19498 867 19510 901
rect 19824 901 20224 907
rect 19110 861 19510 867
rect 18828 823 18834 857
rect 18868 823 18884 857
rect 18396 813 18796 819
rect 18114 793 18194 807
rect 18114 741 18128 793
rect 18180 741 18194 793
rect 18114 727 18194 741
rect 18396 779 18408 813
rect 18784 779 18796 813
rect 18396 733 18414 779
rect 18774 733 18796 779
rect 17682 665 17688 699
rect 18076 665 18082 699
rect 17682 649 18082 665
rect 18396 699 18796 733
rect 18828 807 18884 823
rect 19542 857 19598 873
rect 19824 867 19836 901
rect 20212 867 20224 901
rect 20538 901 20938 907
rect 19824 861 20224 867
rect 19542 823 19548 857
rect 19582 823 19598 857
rect 19110 813 19510 819
rect 18828 793 18908 807
rect 18828 741 18842 793
rect 18894 741 18908 793
rect 18828 727 18908 741
rect 19110 779 19122 813
rect 19498 779 19510 813
rect 19110 733 19128 779
rect 19488 733 19510 779
rect 18396 665 18402 699
rect 18790 665 18796 699
rect 18396 649 18796 665
rect 19110 699 19510 733
rect 19542 807 19598 823
rect 20256 857 20312 873
rect 20538 867 20550 901
rect 20926 867 20938 901
rect 21252 901 21652 907
rect 20538 861 20938 867
rect 20256 823 20262 857
rect 20296 823 20312 857
rect 19824 813 20224 819
rect 19542 793 19622 807
rect 19542 741 19556 793
rect 19608 741 19622 793
rect 19542 727 19622 741
rect 19824 779 19836 813
rect 20212 779 20224 813
rect 19824 733 19842 779
rect 20202 733 20224 779
rect 19110 665 19116 699
rect 19504 665 19510 699
rect 19110 649 19510 665
rect 19824 699 20224 733
rect 20256 807 20312 823
rect 20970 857 21026 873
rect 21252 867 21264 901
rect 21640 867 21652 901
rect 21966 901 22366 907
rect 21252 861 21652 867
rect 20970 823 20976 857
rect 21010 823 21026 857
rect 20538 813 20938 819
rect 20256 793 20336 807
rect 20256 741 20270 793
rect 20322 741 20336 793
rect 20256 727 20336 741
rect 20538 779 20550 813
rect 20926 779 20938 813
rect 20538 733 20556 779
rect 20916 733 20938 779
rect 19824 665 19830 699
rect 20218 665 20224 699
rect 19824 649 20224 665
rect 20538 699 20938 733
rect 20970 807 21026 823
rect 21684 857 21740 873
rect 21966 867 21978 901
rect 22354 867 22366 901
rect 22680 901 23080 907
rect 21966 861 22366 867
rect 21684 823 21690 857
rect 21724 823 21740 857
rect 21252 813 21652 819
rect 20970 793 21050 807
rect 20970 741 20984 793
rect 21036 741 21050 793
rect 20970 727 21050 741
rect 21252 779 21264 813
rect 21640 779 21652 813
rect 21252 733 21270 779
rect 21630 733 21652 779
rect 20538 665 20544 699
rect 20932 665 20938 699
rect 20538 649 20938 665
rect 21252 699 21652 733
rect 21684 807 21740 823
rect 22398 857 22454 873
rect 22680 867 22692 901
rect 23068 867 23080 901
rect 23394 901 23794 907
rect 22680 861 23080 867
rect 22398 823 22404 857
rect 22438 823 22454 857
rect 21966 813 22366 819
rect 21684 793 21764 807
rect 21684 741 21698 793
rect 21750 741 21764 793
rect 21684 727 21764 741
rect 21966 779 21978 813
rect 22354 779 22366 813
rect 21966 733 21984 779
rect 22344 733 22366 779
rect 21252 665 21258 699
rect 21646 665 21652 699
rect 21252 649 21652 665
rect 21966 699 22366 733
rect 22398 807 22454 823
rect 23112 857 23168 873
rect 23394 867 23406 901
rect 23782 867 23794 901
rect 24108 901 24508 907
rect 23394 861 23794 867
rect 23112 823 23118 857
rect 23152 823 23168 857
rect 22680 813 23080 819
rect 22398 793 22478 807
rect 22398 741 22412 793
rect 22464 741 22478 793
rect 22398 727 22478 741
rect 22680 779 22692 813
rect 23068 779 23080 813
rect 22680 733 22698 779
rect 23058 733 23080 779
rect 21966 665 21972 699
rect 22360 665 22366 699
rect 21966 649 22366 665
rect 22680 699 23080 733
rect 23112 807 23168 823
rect 23826 857 23882 873
rect 24108 867 24120 901
rect 24496 867 24508 901
rect 24822 901 25222 907
rect 24108 861 24508 867
rect 23826 823 23832 857
rect 23866 823 23882 857
rect 23394 813 23794 819
rect 23112 793 23192 807
rect 23112 741 23126 793
rect 23178 741 23192 793
rect 23112 727 23192 741
rect 23394 779 23406 813
rect 23782 779 23794 813
rect 23394 733 23412 779
rect 23772 733 23794 779
rect 22680 665 22686 699
rect 23074 665 23080 699
rect 22680 649 23080 665
rect 23394 699 23794 733
rect 23826 807 23882 823
rect 24540 857 24596 873
rect 24822 867 24834 901
rect 25210 867 25222 901
rect 25536 901 25936 907
rect 24822 861 25222 867
rect 24540 823 24546 857
rect 24580 823 24596 857
rect 24108 813 24508 819
rect 23826 793 23906 807
rect 23826 741 23840 793
rect 23892 741 23906 793
rect 23826 727 23906 741
rect 24108 779 24120 813
rect 24496 779 24508 813
rect 24108 733 24126 779
rect 24486 733 24508 779
rect 23394 665 23400 699
rect 23788 665 23794 699
rect 23394 649 23794 665
rect 24108 699 24508 733
rect 24540 807 24596 823
rect 25254 857 25310 873
rect 25536 867 25548 901
rect 25924 867 25936 901
rect 26250 901 26650 907
rect 25536 861 25936 867
rect 25254 823 25260 857
rect 25294 823 25310 857
rect 24822 813 25222 819
rect 24540 793 24620 807
rect 24540 741 24554 793
rect 24606 741 24620 793
rect 24540 727 24620 741
rect 24822 779 24834 813
rect 25210 779 25222 813
rect 24822 733 24840 779
rect 25200 733 25222 779
rect 24108 665 24114 699
rect 24502 665 24508 699
rect 24108 649 24508 665
rect 24822 699 25222 733
rect 25254 807 25310 823
rect 25968 857 26024 873
rect 26250 867 26262 901
rect 26638 867 26650 901
rect 26964 901 27364 907
rect 26250 861 26650 867
rect 25968 823 25974 857
rect 26008 823 26024 857
rect 25536 813 25936 819
rect 25254 793 25334 807
rect 25254 741 25268 793
rect 25320 741 25334 793
rect 25254 727 25334 741
rect 25536 779 25548 813
rect 25924 779 25936 813
rect 25536 733 25554 779
rect 25914 733 25936 779
rect 24822 665 24828 699
rect 25216 665 25222 699
rect 24822 649 25222 665
rect 25536 699 25936 733
rect 25968 807 26024 823
rect 26682 857 26738 873
rect 26964 867 26976 901
rect 27352 867 27364 901
rect 27678 901 28078 907
rect 26964 861 27364 867
rect 26682 823 26688 857
rect 26722 823 26738 857
rect 26250 813 26650 819
rect 25968 793 26048 807
rect 25968 741 25982 793
rect 26034 741 26048 793
rect 25968 727 26048 741
rect 26250 779 26262 813
rect 26638 779 26650 813
rect 26250 733 26268 779
rect 26628 733 26650 779
rect 25536 665 25542 699
rect 25930 665 25936 699
rect 25536 649 25936 665
rect 26250 699 26650 733
rect 26682 807 26738 823
rect 27396 857 27452 873
rect 27678 867 27690 901
rect 28066 867 28078 901
rect 28392 901 28792 907
rect 27678 861 28078 867
rect 27396 823 27402 857
rect 27436 823 27452 857
rect 26964 813 27364 819
rect 26682 793 26762 807
rect 26682 741 26696 793
rect 26748 741 26762 793
rect 26682 727 26762 741
rect 26964 779 26976 813
rect 27352 779 27364 813
rect 26964 733 26982 779
rect 27342 733 27364 779
rect 26250 665 26256 699
rect 26644 665 26650 699
rect 26250 649 26650 665
rect 26964 699 27364 733
rect 27396 807 27452 823
rect 28110 857 28166 873
rect 28392 867 28404 901
rect 28780 867 28792 901
rect 29106 901 29506 907
rect 28392 861 28792 867
rect 28110 823 28116 857
rect 28150 823 28166 857
rect 27678 813 28078 819
rect 27396 793 27476 807
rect 27396 741 27410 793
rect 27462 741 27476 793
rect 27396 727 27476 741
rect 27678 779 27690 813
rect 28066 779 28078 813
rect 27678 733 27696 779
rect 28056 733 28078 779
rect 26964 665 26970 699
rect 27358 665 27364 699
rect 26964 649 27364 665
rect 27678 699 28078 733
rect 28110 807 28166 823
rect 28824 857 28880 873
rect 29106 867 29118 901
rect 29494 867 29506 901
rect 29820 901 30220 907
rect 29106 861 29506 867
rect 28824 823 28830 857
rect 28864 823 28880 857
rect 28392 813 28792 819
rect 28110 793 28190 807
rect 28110 741 28124 793
rect 28176 741 28190 793
rect 28110 727 28190 741
rect 28392 779 28404 813
rect 28780 779 28792 813
rect 28392 733 28410 779
rect 28770 733 28792 779
rect 27678 665 27684 699
rect 28072 665 28078 699
rect 27678 649 28078 665
rect 28392 699 28792 733
rect 28824 807 28880 823
rect 29538 857 29594 873
rect 29820 867 29832 901
rect 30208 867 30220 901
rect 30534 901 30934 907
rect 29820 861 30220 867
rect 29538 823 29544 857
rect 29578 823 29594 857
rect 29106 813 29506 819
rect 28824 793 28904 807
rect 28824 741 28838 793
rect 28890 741 28904 793
rect 28824 727 28904 741
rect 29106 779 29118 813
rect 29494 779 29506 813
rect 29106 733 29124 779
rect 29484 733 29506 779
rect 28392 665 28398 699
rect 28786 665 28792 699
rect 28392 649 28792 665
rect 29106 699 29506 733
rect 29538 807 29594 823
rect 30252 857 30308 873
rect 30534 867 30546 901
rect 30922 867 30934 901
rect 31248 901 31648 907
rect 30534 861 30934 867
rect 30252 823 30258 857
rect 30292 823 30308 857
rect 29820 813 30220 819
rect 29538 793 29618 807
rect 29538 741 29552 793
rect 29604 741 29618 793
rect 29538 727 29618 741
rect 29820 779 29832 813
rect 30208 779 30220 813
rect 29820 733 29838 779
rect 30198 733 30220 779
rect 29106 665 29112 699
rect 29500 665 29506 699
rect 29106 649 29506 665
rect 29820 699 30220 733
rect 30252 807 30308 823
rect 30966 857 31022 873
rect 31248 867 31260 901
rect 31636 867 31648 901
rect 31962 901 32362 907
rect 31248 861 31648 867
rect 30966 823 30972 857
rect 31006 823 31022 857
rect 30534 813 30934 819
rect 30252 793 30332 807
rect 30252 741 30266 793
rect 30318 741 30332 793
rect 30252 727 30332 741
rect 30534 779 30546 813
rect 30922 779 30934 813
rect 30534 733 30552 779
rect 30912 733 30934 779
rect 29820 665 29826 699
rect 30214 665 30220 699
rect 29820 649 30220 665
rect 30534 699 30934 733
rect 30966 807 31022 823
rect 31680 857 31736 873
rect 31962 867 31974 901
rect 32350 867 32362 901
rect 32676 901 33076 907
rect 31962 861 32362 867
rect 31680 823 31686 857
rect 31720 823 31736 857
rect 31248 813 31648 819
rect 30966 793 31046 807
rect 30966 741 30980 793
rect 31032 741 31046 793
rect 30966 727 31046 741
rect 31248 779 31260 813
rect 31636 779 31648 813
rect 31248 733 31266 779
rect 31626 733 31648 779
rect 30534 665 30540 699
rect 30928 665 30934 699
rect 30534 649 30934 665
rect 31248 699 31648 733
rect 31680 807 31736 823
rect 32394 857 32450 873
rect 32676 867 32688 901
rect 33064 867 33076 901
rect 33390 901 33790 907
rect 32676 861 33076 867
rect 32394 823 32400 857
rect 32434 823 32450 857
rect 31962 813 32362 819
rect 31680 793 31760 807
rect 31680 741 31694 793
rect 31746 741 31760 793
rect 31680 727 31760 741
rect 31962 779 31974 813
rect 32350 779 32362 813
rect 31962 733 31980 779
rect 32340 733 32362 779
rect 31248 665 31254 699
rect 31642 665 31648 699
rect 31248 649 31648 665
rect 31962 699 32362 733
rect 32394 807 32450 823
rect 33108 857 33164 873
rect 33390 867 33402 901
rect 33778 867 33790 901
rect 34104 901 34504 907
rect 33390 861 33790 867
rect 33108 823 33114 857
rect 33148 823 33164 857
rect 32676 813 33076 819
rect 32394 793 32474 807
rect 32394 741 32408 793
rect 32460 741 32474 793
rect 32394 727 32474 741
rect 32676 779 32688 813
rect 33064 779 33076 813
rect 32676 733 32694 779
rect 33054 733 33076 779
rect 31962 665 31968 699
rect 32356 665 32362 699
rect 31962 649 32362 665
rect 32676 699 33076 733
rect 33108 807 33164 823
rect 33822 857 33878 873
rect 34104 867 34116 901
rect 34492 867 34504 901
rect 34818 901 35218 907
rect 34104 861 34504 867
rect 33822 823 33828 857
rect 33862 823 33878 857
rect 33390 813 33790 819
rect 33108 793 33188 807
rect 33108 741 33122 793
rect 33174 741 33188 793
rect 33108 727 33188 741
rect 33390 779 33402 813
rect 33778 779 33790 813
rect 33390 733 33408 779
rect 33768 733 33790 779
rect 32676 665 32682 699
rect 33070 665 33076 699
rect 32676 649 33076 665
rect 33390 699 33790 733
rect 33822 807 33878 823
rect 34536 857 34592 873
rect 34818 867 34830 901
rect 35206 867 35218 901
rect 35532 901 35932 907
rect 34818 861 35218 867
rect 34536 823 34542 857
rect 34576 823 34592 857
rect 34104 813 34504 819
rect 33822 793 33902 807
rect 33822 741 33836 793
rect 33888 741 33902 793
rect 33822 727 33902 741
rect 34104 779 34116 813
rect 34492 779 34504 813
rect 34104 733 34122 779
rect 34482 733 34504 779
rect 33390 665 33396 699
rect 33784 665 33790 699
rect 33390 649 33790 665
rect 34104 699 34504 733
rect 34536 807 34592 823
rect 35250 857 35306 873
rect 35532 867 35544 901
rect 35920 867 35932 901
rect 36246 901 36646 907
rect 35532 861 35932 867
rect 35250 823 35256 857
rect 35290 823 35306 857
rect 34818 813 35218 819
rect 34536 793 34616 807
rect 34536 741 34550 793
rect 34602 741 34616 793
rect 34536 727 34616 741
rect 34818 779 34830 813
rect 35206 779 35218 813
rect 34818 733 34836 779
rect 35196 733 35218 779
rect 34104 665 34110 699
rect 34498 665 34504 699
rect 34104 649 34504 665
rect 34818 699 35218 733
rect 35250 807 35306 823
rect 35964 857 36020 873
rect 36246 867 36258 901
rect 36634 867 36646 901
rect 36960 901 37360 907
rect 36246 861 36646 867
rect 35964 823 35970 857
rect 36004 823 36020 857
rect 35532 813 35932 819
rect 35250 793 35330 807
rect 35250 741 35264 793
rect 35316 741 35330 793
rect 35250 727 35330 741
rect 35532 779 35544 813
rect 35920 779 35932 813
rect 35532 733 35550 779
rect 35910 733 35932 779
rect 34818 665 34824 699
rect 35212 665 35218 699
rect 34818 649 35218 665
rect 35532 699 35932 733
rect 35964 807 36020 823
rect 36678 857 36734 873
rect 36960 867 36972 901
rect 37348 867 37360 901
rect 37674 901 38074 907
rect 38385 902 38788 907
rect 36960 861 37360 867
rect 36678 823 36684 857
rect 36718 823 36734 857
rect 36246 813 36646 819
rect 35964 793 36044 807
rect 35964 741 35978 793
rect 36030 741 36044 793
rect 35964 727 36044 741
rect 36246 779 36258 813
rect 36634 779 36646 813
rect 36246 733 36264 779
rect 36624 733 36646 779
rect 35532 665 35538 699
rect 35926 665 35932 699
rect 35532 649 35932 665
rect 36246 699 36646 733
rect 36678 807 36734 823
rect 37392 857 37448 873
rect 37674 867 37686 901
rect 38062 867 38074 901
rect 38388 901 38788 902
rect 37674 861 38074 867
rect 37392 823 37398 857
rect 37432 823 37448 857
rect 36960 813 37360 819
rect 36678 793 36758 807
rect 36678 741 36692 793
rect 36744 741 36758 793
rect 36678 727 36758 741
rect 36960 779 36972 813
rect 37348 779 37360 813
rect 36960 733 36978 779
rect 37338 733 37360 779
rect 36246 665 36252 699
rect 36640 665 36646 699
rect 36246 649 36646 665
rect 36960 699 37360 733
rect 37392 807 37448 823
rect 38106 857 38162 873
rect 38388 867 38400 901
rect 38776 867 38788 901
rect 38388 861 38788 867
rect 38106 823 38112 857
rect 38146 823 38162 857
rect 37674 813 38074 819
rect 37392 793 37472 807
rect 37392 741 37406 793
rect 37458 741 37472 793
rect 37392 727 37472 741
rect 37674 779 37686 813
rect 38062 779 38074 813
rect 36960 665 36966 699
rect 37354 665 37360 699
rect 36960 649 37360 665
rect 37674 699 37698 779
rect 38048 699 38074 779
rect 38106 807 38162 823
rect 38820 857 38876 873
rect 39370 869 39390 880
rect 38820 823 38826 857
rect 38860 823 38876 857
rect 38388 813 38788 819
rect 38106 793 38186 807
rect 38106 741 38120 793
rect 38172 741 38186 793
rect 38106 727 38186 741
rect 38388 779 38400 813
rect 38776 779 38788 813
rect 38388 729 38408 779
rect 38768 729 38788 779
rect 37674 665 37680 699
rect 38068 665 38074 699
rect 37674 649 38074 665
rect 38388 699 38788 729
rect 38820 807 38876 823
rect 39369 863 39390 869
rect 39770 863 39790 880
rect 39369 825 39381 863
rect 39778 825 39790 863
rect 39369 820 39390 825
rect 39770 820 39790 825
rect 39369 819 39790 820
rect 39900 863 39920 880
rect 40300 869 40320 880
rect 40300 863 40321 869
rect 39900 825 39912 863
rect 40309 825 40321 863
rect 39900 820 39920 825
rect 40300 820 40321 825
rect 39900 819 40321 820
rect 38820 793 38900 807
rect 38820 741 38834 793
rect 38886 741 38900 793
rect 38820 727 38900 741
rect 39370 703 39390 710
rect 38388 665 38394 699
rect 38782 665 38788 699
rect 38388 649 38788 665
rect 39369 697 39390 703
rect 39770 697 39790 710
rect 39369 659 39381 697
rect 39778 659 39790 697
rect 39369 653 39390 659
rect 39370 650 39390 653
rect 39770 650 39790 659
rect 39900 697 39920 710
rect 40300 703 40320 710
rect 40300 697 40321 703
rect 39900 659 39912 697
rect 40309 659 40321 697
rect 39900 650 39920 659
rect 40300 653 40321 659
rect 40300 650 40320 653
rect 14290 308 14408 320
rect 3940 195 4061 205
rect 10458 278 10488 308
rect 10458 276 10518 278
rect 10860 276 10900 308
rect 11318 276 11358 308
rect 11776 276 11816 308
rect 12692 276 12732 308
rect 13608 276 13648 308
rect 10458 270 10900 276
rect 10458 236 10520 270
rect 10888 236 10900 270
rect 10458 230 10900 236
rect 10966 270 11358 276
rect 10966 236 10978 270
rect 11346 236 11358 270
rect 10966 230 11358 236
rect 11424 270 11816 276
rect 11424 236 11436 270
rect 11804 236 11816 270
rect 11424 230 11816 236
rect 11882 270 12274 276
rect 11882 236 11894 270
rect 12262 236 12274 270
rect 11882 230 12274 236
rect 12340 270 12732 276
rect 12340 236 12352 270
rect 12720 236 12732 270
rect 12340 230 12732 236
rect 12798 270 13190 276
rect 12798 236 12810 270
rect 13178 236 13190 270
rect 12798 230 13190 236
rect 13256 270 13648 276
rect 13256 236 13268 270
rect 13636 236 13648 270
rect 13256 230 13648 236
rect 10458 228 10518 230
rect 3940 194 3946 195
rect 3900 182 3946 194
rect 10458 168 10488 228
rect 10860 168 10900 230
rect 11318 228 11358 230
rect 11776 168 11816 230
rect 12692 168 12732 230
rect 13608 168 13648 230
rect 14328 168 14408 308
rect 15318 480 38998 649
rect 39370 537 39390 550
rect 39369 531 39390 537
rect 39770 531 39790 550
rect 39369 493 39381 531
rect 39778 493 39790 531
rect 39369 490 39390 493
rect 39770 490 39790 493
rect 39150 480 39270 490
rect 39369 487 39790 490
rect 39900 531 39920 540
rect 40300 537 40320 540
rect 40300 531 40321 537
rect 39900 493 39912 531
rect 40309 493 40321 531
rect 39900 480 39920 493
rect 40300 487 40321 493
rect 40300 480 40320 487
rect 15318 470 39270 480
rect 15318 380 39170 470
rect 39250 380 39270 470
rect 15318 370 39270 380
rect 39370 371 39390 380
rect 15318 209 38998 370
rect 39150 360 39270 370
rect 39369 365 39390 371
rect 39770 365 39790 380
rect 39369 327 39381 365
rect 39778 327 39790 365
rect 39369 321 39390 327
rect 39370 320 39390 321
rect 39770 320 39790 327
rect 39900 370 40321 371
rect 39900 365 39920 370
rect 40300 365 40321 370
rect 39900 327 39912 365
rect 40309 327 40321 365
rect 39900 310 39920 327
rect 40300 321 40321 327
rect 40300 310 40320 321
rect 15540 197 15940 209
rect 10308 158 14448 168
rect 3766 144 3912 150
rect 3766 136 3862 144
rect 3766 84 3780 136
rect 3832 110 3862 136
rect 3896 110 3912 144
rect 3832 94 3912 110
rect 3832 84 3846 94
rect 3766 70 3846 84
rect 10308 78 10358 158
rect 14428 78 14448 158
rect 10308 58 14448 78
rect 15540 163 15546 197
rect 15934 163 15940 197
rect 15540 129 15940 163
rect 16254 197 16654 209
rect 16254 163 16260 197
rect 16648 163 16654 197
rect 15540 83 15558 129
rect 15918 83 15940 129
rect 15540 49 15552 83
rect 15928 49 15940 83
rect 15540 43 15940 49
rect 15972 121 16052 135
rect 15972 69 15986 121
rect 16038 69 16052 121
rect 15972 55 16052 69
rect 16254 129 16654 163
rect 16968 197 17368 209
rect 16968 163 16974 197
rect 17362 163 17368 197
rect 16254 83 16272 129
rect 16632 83 16654 129
rect 15972 39 16028 55
rect 16254 49 16266 83
rect 16642 49 16654 83
rect 16254 43 16654 49
rect 16686 121 16766 135
rect 16686 69 16700 121
rect 16752 69 16766 121
rect 16686 55 16766 69
rect 16968 129 17368 163
rect 17682 197 18082 209
rect 17682 163 17688 197
rect 18076 163 18082 197
rect 16968 83 16986 129
rect 17346 83 17368 129
rect 15972 5 15978 39
rect 16012 5 16028 39
rect 15540 -5 15940 1
rect 15540 -39 15552 -5
rect 15928 -39 15940 -5
rect 15972 -11 16028 5
rect 16686 39 16742 55
rect 16968 49 16980 83
rect 17356 49 17368 83
rect 16968 43 17368 49
rect 17400 121 17480 135
rect 17400 69 17414 121
rect 17466 69 17480 121
rect 17400 55 17480 69
rect 17682 129 18082 163
rect 18396 197 18796 209
rect 18396 163 18402 197
rect 18790 163 18796 197
rect 17682 83 17700 129
rect 18060 83 18082 129
rect 16686 5 16692 39
rect 16726 5 16742 39
rect 16254 -5 16654 1
rect 15540 -45 15940 -39
rect 16254 -39 16266 -5
rect 16642 -39 16654 -5
rect 16686 -11 16742 5
rect 17400 39 17456 55
rect 17682 49 17694 83
rect 18070 49 18082 83
rect 17682 43 18082 49
rect 18114 121 18194 135
rect 18114 69 18128 121
rect 18180 69 18194 121
rect 18114 55 18194 69
rect 18396 129 18796 163
rect 19110 197 19510 209
rect 19110 163 19116 197
rect 19504 163 19510 197
rect 18396 83 18414 129
rect 18774 83 18796 129
rect 17400 5 17406 39
rect 17440 5 17456 39
rect 16968 -5 17368 1
rect 16254 -45 16654 -39
rect 16968 -39 16980 -5
rect 17356 -39 17368 -5
rect 17400 -11 17456 5
rect 18114 39 18170 55
rect 18396 49 18408 83
rect 18784 49 18796 83
rect 18396 43 18796 49
rect 18828 121 18908 135
rect 18828 69 18842 121
rect 18894 69 18908 121
rect 18828 55 18908 69
rect 19110 129 19510 163
rect 19824 197 20224 209
rect 19824 163 19830 197
rect 20218 163 20224 197
rect 19110 83 19128 129
rect 19488 83 19510 129
rect 18114 5 18120 39
rect 18154 5 18170 39
rect 17682 -5 18082 1
rect 16968 -45 17368 -39
rect 17682 -39 17694 -5
rect 18070 -39 18082 -5
rect 18114 -11 18170 5
rect 18828 39 18884 55
rect 19110 49 19122 83
rect 19498 49 19510 83
rect 19110 43 19510 49
rect 19542 121 19622 135
rect 19542 69 19556 121
rect 19608 69 19622 121
rect 19542 55 19622 69
rect 19824 129 20224 163
rect 20538 197 20938 209
rect 20538 163 20544 197
rect 20932 163 20938 197
rect 19824 83 19842 129
rect 20202 83 20224 129
rect 18828 5 18834 39
rect 18868 5 18884 39
rect 18396 -5 18796 1
rect 17682 -45 18082 -39
rect 18396 -39 18408 -5
rect 18784 -39 18796 -5
rect 18828 -11 18884 5
rect 19542 39 19598 55
rect 19824 49 19836 83
rect 20212 49 20224 83
rect 19824 43 20224 49
rect 20256 121 20336 135
rect 20256 69 20270 121
rect 20322 69 20336 121
rect 20256 55 20336 69
rect 20538 129 20938 163
rect 21252 197 21652 209
rect 21252 163 21258 197
rect 21646 163 21652 197
rect 20538 83 20556 129
rect 20916 83 20938 129
rect 19542 5 19548 39
rect 19582 5 19598 39
rect 19110 -5 19510 1
rect 18396 -45 18796 -39
rect 19110 -39 19122 -5
rect 19498 -39 19510 -5
rect 19542 -11 19598 5
rect 20256 39 20312 55
rect 20538 49 20550 83
rect 20926 49 20938 83
rect 20538 43 20938 49
rect 20970 121 21050 135
rect 20970 69 20984 121
rect 21036 69 21050 121
rect 20970 55 21050 69
rect 21252 129 21652 163
rect 21966 197 22366 209
rect 21966 163 21972 197
rect 22360 163 22366 197
rect 21252 83 21270 129
rect 21630 83 21652 129
rect 20256 5 20262 39
rect 20296 5 20312 39
rect 19824 -5 20224 1
rect 19110 -45 19510 -39
rect 19824 -39 19836 -5
rect 20212 -39 20224 -5
rect 20256 -11 20312 5
rect 20970 39 21026 55
rect 21252 49 21264 83
rect 21640 49 21652 83
rect 21252 43 21652 49
rect 21684 121 21764 135
rect 21684 69 21698 121
rect 21750 69 21764 121
rect 21684 55 21764 69
rect 21966 129 22366 163
rect 22680 197 23080 209
rect 22680 163 22686 197
rect 23074 163 23080 197
rect 21966 83 21984 129
rect 22344 83 22366 129
rect 20970 5 20976 39
rect 21010 5 21026 39
rect 20538 -5 20938 1
rect 19824 -45 20224 -39
rect 20538 -39 20550 -5
rect 20926 -39 20938 -5
rect 20970 -11 21026 5
rect 21684 39 21740 55
rect 21966 49 21978 83
rect 22354 49 22366 83
rect 21966 43 22366 49
rect 22398 121 22478 135
rect 22398 69 22412 121
rect 22464 69 22478 121
rect 22398 55 22478 69
rect 22680 129 23080 163
rect 23394 197 23794 209
rect 23394 163 23400 197
rect 23788 163 23794 197
rect 22680 83 22698 129
rect 23058 83 23080 129
rect 21684 5 21690 39
rect 21724 5 21740 39
rect 21252 -5 21652 1
rect 20538 -45 20938 -39
rect 21252 -39 21264 -5
rect 21640 -39 21652 -5
rect 21684 -11 21740 5
rect 22398 39 22454 55
rect 22680 49 22692 83
rect 23068 49 23080 83
rect 22680 43 23080 49
rect 23112 121 23192 135
rect 23112 69 23126 121
rect 23178 69 23192 121
rect 23112 55 23192 69
rect 23394 129 23794 163
rect 24108 197 24508 209
rect 24108 163 24114 197
rect 24502 163 24508 197
rect 23394 83 23412 129
rect 23772 83 23794 129
rect 22398 5 22404 39
rect 22438 5 22454 39
rect 21966 -5 22366 1
rect 21252 -45 21652 -39
rect 21966 -39 21978 -5
rect 22354 -39 22366 -5
rect 22398 -11 22454 5
rect 23112 39 23168 55
rect 23394 49 23406 83
rect 23782 49 23794 83
rect 23394 43 23794 49
rect 23826 121 23906 135
rect 23826 69 23840 121
rect 23892 69 23906 121
rect 23826 55 23906 69
rect 24108 129 24508 163
rect 24822 197 25222 209
rect 24822 163 24828 197
rect 25216 163 25222 197
rect 24108 83 24126 129
rect 24486 83 24508 129
rect 23112 5 23118 39
rect 23152 5 23168 39
rect 22680 -5 23080 1
rect 21966 -45 22366 -39
rect 22680 -39 22692 -5
rect 23068 -39 23080 -5
rect 23112 -11 23168 5
rect 23826 39 23882 55
rect 24108 49 24120 83
rect 24496 49 24508 83
rect 24108 43 24508 49
rect 24540 121 24620 135
rect 24540 69 24554 121
rect 24606 69 24620 121
rect 24540 55 24620 69
rect 24822 129 25222 163
rect 25536 197 25936 209
rect 25536 163 25542 197
rect 25930 163 25936 197
rect 24822 83 24840 129
rect 25200 83 25222 129
rect 23826 5 23832 39
rect 23866 5 23882 39
rect 23394 -5 23794 1
rect 22680 -45 23080 -39
rect 23394 -39 23406 -5
rect 23782 -39 23794 -5
rect 23826 -11 23882 5
rect 24540 39 24596 55
rect 24822 49 24834 83
rect 25210 49 25222 83
rect 24822 43 25222 49
rect 25254 121 25334 135
rect 25254 69 25268 121
rect 25320 69 25334 121
rect 25254 55 25334 69
rect 25536 129 25936 163
rect 26250 197 26650 209
rect 26250 163 26256 197
rect 26644 163 26650 197
rect 25536 83 25554 129
rect 25914 83 25936 129
rect 24540 5 24546 39
rect 24580 5 24596 39
rect 24108 -5 24508 1
rect 23394 -45 23794 -39
rect 24108 -39 24120 -5
rect 24496 -39 24508 -5
rect 24540 -11 24596 5
rect 25254 39 25310 55
rect 25536 49 25548 83
rect 25924 49 25936 83
rect 25536 43 25936 49
rect 25968 121 26048 135
rect 25968 69 25982 121
rect 26034 69 26048 121
rect 25968 55 26048 69
rect 26250 129 26650 163
rect 26964 197 27364 209
rect 26964 163 26970 197
rect 27358 163 27364 197
rect 26250 83 26268 129
rect 26628 83 26650 129
rect 25254 5 25260 39
rect 25294 5 25310 39
rect 24822 -5 25222 1
rect 24108 -45 24508 -39
rect 24822 -39 24834 -5
rect 25210 -39 25222 -5
rect 25254 -11 25310 5
rect 25968 39 26024 55
rect 26250 49 26262 83
rect 26638 49 26650 83
rect 26250 43 26650 49
rect 26682 121 26762 135
rect 26682 69 26696 121
rect 26748 69 26762 121
rect 26682 55 26762 69
rect 26964 129 27364 163
rect 27678 197 28078 209
rect 27678 163 27684 197
rect 28072 163 28078 197
rect 26964 83 26982 129
rect 27342 83 27364 129
rect 25968 5 25974 39
rect 26008 5 26024 39
rect 25536 -5 25936 1
rect 24822 -45 25222 -39
rect 25536 -39 25548 -5
rect 25924 -39 25936 -5
rect 25968 -11 26024 5
rect 26682 39 26738 55
rect 26964 49 26976 83
rect 27352 49 27364 83
rect 26964 43 27364 49
rect 27396 121 27476 135
rect 27396 69 27410 121
rect 27462 69 27476 121
rect 27396 55 27476 69
rect 27678 129 28078 163
rect 28392 197 28792 209
rect 28392 163 28398 197
rect 28786 163 28792 197
rect 27678 83 27696 129
rect 28056 83 28078 129
rect 26682 5 26688 39
rect 26722 5 26738 39
rect 26250 -5 26650 1
rect 25536 -45 25936 -39
rect 26250 -39 26262 -5
rect 26638 -39 26650 -5
rect 26682 -11 26738 5
rect 27396 39 27452 55
rect 27678 49 27690 83
rect 28066 49 28078 83
rect 27678 43 28078 49
rect 28110 121 28190 135
rect 28110 69 28124 121
rect 28176 69 28190 121
rect 28110 55 28190 69
rect 28392 129 28792 163
rect 29106 197 29506 209
rect 29106 163 29112 197
rect 29500 163 29506 197
rect 28392 83 28410 129
rect 28770 83 28792 129
rect 27396 5 27402 39
rect 27436 5 27452 39
rect 26964 -5 27364 1
rect 26250 -45 26650 -39
rect 26964 -39 26976 -5
rect 27352 -39 27364 -5
rect 27396 -11 27452 5
rect 28110 39 28166 55
rect 28392 49 28404 83
rect 28780 49 28792 83
rect 28392 43 28792 49
rect 28824 121 28904 135
rect 28824 69 28838 121
rect 28890 69 28904 121
rect 28824 55 28904 69
rect 29106 129 29506 163
rect 29820 197 30220 209
rect 29820 163 29826 197
rect 30214 163 30220 197
rect 29106 83 29124 129
rect 29484 83 29506 129
rect 28110 5 28116 39
rect 28150 5 28166 39
rect 27678 -5 28078 1
rect 26964 -45 27364 -39
rect 27678 -39 27690 -5
rect 28066 -39 28078 -5
rect 28110 -11 28166 5
rect 28824 39 28880 55
rect 29106 49 29118 83
rect 29494 49 29506 83
rect 29106 43 29506 49
rect 29538 121 29618 135
rect 29538 69 29552 121
rect 29604 69 29618 121
rect 29538 55 29618 69
rect 29820 129 30220 163
rect 30534 197 30934 209
rect 30534 163 30540 197
rect 30928 163 30934 197
rect 29820 83 29838 129
rect 30198 83 30220 129
rect 28824 5 28830 39
rect 28864 5 28880 39
rect 28392 -5 28792 1
rect 27678 -45 28078 -39
rect 28392 -39 28404 -5
rect 28780 -39 28792 -5
rect 28824 -11 28880 5
rect 29538 39 29594 55
rect 29820 49 29832 83
rect 30208 49 30220 83
rect 29820 43 30220 49
rect 30252 121 30332 135
rect 30252 69 30266 121
rect 30318 69 30332 121
rect 30252 55 30332 69
rect 30534 129 30934 163
rect 31248 197 31648 209
rect 31248 163 31254 197
rect 31642 163 31648 197
rect 30534 83 30552 129
rect 30912 83 30934 129
rect 29538 5 29544 39
rect 29578 5 29594 39
rect 29106 -5 29506 1
rect 28392 -45 28792 -39
rect 29106 -39 29118 -5
rect 29494 -39 29506 -5
rect 29538 -11 29594 5
rect 30252 39 30308 55
rect 30534 49 30546 83
rect 30922 49 30934 83
rect 30534 43 30934 49
rect 30966 121 31046 135
rect 30966 69 30980 121
rect 31032 69 31046 121
rect 30966 55 31046 69
rect 31248 129 31648 163
rect 31962 197 32362 209
rect 31962 163 31968 197
rect 32356 163 32362 197
rect 31248 83 31266 129
rect 31626 83 31648 129
rect 30252 5 30258 39
rect 30292 5 30308 39
rect 29820 -5 30220 1
rect 29106 -45 29506 -39
rect 29820 -39 29832 -5
rect 30208 -39 30220 -5
rect 30252 -11 30308 5
rect 30966 39 31022 55
rect 31248 49 31260 83
rect 31636 49 31648 83
rect 31248 43 31648 49
rect 31680 121 31760 135
rect 31680 69 31694 121
rect 31746 69 31760 121
rect 31680 55 31760 69
rect 31962 129 32362 163
rect 32676 197 33076 209
rect 32676 163 32682 197
rect 33070 163 33076 197
rect 31962 83 31980 129
rect 32340 83 32362 129
rect 30966 5 30972 39
rect 31006 5 31022 39
rect 30534 -5 30934 1
rect 29820 -45 30220 -39
rect 30534 -39 30546 -5
rect 30922 -39 30934 -5
rect 30966 -11 31022 5
rect 31680 39 31736 55
rect 31962 49 31974 83
rect 32350 49 32362 83
rect 31962 43 32362 49
rect 32394 121 32474 135
rect 32394 69 32408 121
rect 32460 69 32474 121
rect 32394 55 32474 69
rect 32676 129 33076 163
rect 33390 197 33790 209
rect 33390 163 33396 197
rect 33784 163 33790 197
rect 32676 83 32694 129
rect 33054 83 33076 129
rect 31680 5 31686 39
rect 31720 5 31736 39
rect 31248 -5 31648 1
rect 30534 -45 30934 -39
rect 31248 -39 31260 -5
rect 31636 -39 31648 -5
rect 31680 -11 31736 5
rect 32394 39 32450 55
rect 32676 49 32688 83
rect 33064 49 33076 83
rect 32676 43 33076 49
rect 33108 121 33188 135
rect 33108 69 33122 121
rect 33174 69 33188 121
rect 33108 55 33188 69
rect 33390 129 33790 163
rect 34104 197 34504 209
rect 34104 163 34110 197
rect 34498 163 34504 197
rect 33390 83 33408 129
rect 33768 83 33790 129
rect 32394 5 32400 39
rect 32434 5 32450 39
rect 31962 -5 32362 1
rect 31248 -45 31648 -39
rect 31962 -39 31974 -5
rect 32350 -39 32362 -5
rect 32394 -11 32450 5
rect 33108 39 33164 55
rect 33390 49 33402 83
rect 33778 49 33790 83
rect 33390 43 33790 49
rect 33822 121 33902 135
rect 33822 69 33836 121
rect 33888 69 33902 121
rect 33822 55 33902 69
rect 34104 129 34504 163
rect 34818 197 35218 209
rect 34818 163 34824 197
rect 35212 163 35218 197
rect 34104 83 34122 129
rect 34482 83 34504 129
rect 33108 5 33114 39
rect 33148 5 33164 39
rect 32676 -5 33076 1
rect 31962 -45 32362 -39
rect 32676 -39 32688 -5
rect 33064 -39 33076 -5
rect 33108 -11 33164 5
rect 33822 39 33878 55
rect 34104 49 34116 83
rect 34492 49 34504 83
rect 34104 43 34504 49
rect 34536 121 34616 135
rect 34536 69 34550 121
rect 34602 69 34616 121
rect 34536 55 34616 69
rect 34818 129 35218 163
rect 35532 197 35932 209
rect 35532 163 35538 197
rect 35926 163 35932 197
rect 34818 83 34836 129
rect 35196 83 35218 129
rect 33822 5 33828 39
rect 33862 5 33878 39
rect 33390 -5 33790 1
rect 32676 -45 33076 -39
rect 33390 -39 33402 -5
rect 33778 -39 33790 -5
rect 33822 -11 33878 5
rect 34536 39 34592 55
rect 34818 49 34830 83
rect 35206 49 35218 83
rect 34818 43 35218 49
rect 35250 121 35330 135
rect 35250 69 35264 121
rect 35316 69 35330 121
rect 35250 55 35330 69
rect 35532 129 35932 163
rect 36246 197 36646 209
rect 36246 163 36252 197
rect 36640 163 36646 197
rect 35532 83 35550 129
rect 35910 83 35932 129
rect 34536 5 34542 39
rect 34576 5 34592 39
rect 34104 -5 34504 1
rect 33390 -45 33790 -39
rect 34104 -39 34116 -5
rect 34492 -39 34504 -5
rect 34536 -11 34592 5
rect 35250 39 35306 55
rect 35532 49 35544 83
rect 35920 49 35932 83
rect 35532 43 35932 49
rect 35964 121 36044 135
rect 35964 69 35978 121
rect 36030 69 36044 121
rect 35964 55 36044 69
rect 36246 129 36646 163
rect 36960 197 37360 209
rect 36960 163 36966 197
rect 37354 163 37360 197
rect 36246 83 36264 129
rect 36624 83 36646 129
rect 35250 5 35256 39
rect 35290 5 35306 39
rect 34818 -5 35218 1
rect 34104 -45 34504 -39
rect 34818 -39 34830 -5
rect 35206 -39 35218 -5
rect 35250 -11 35306 5
rect 35964 39 36020 55
rect 36246 49 36258 83
rect 36634 49 36646 83
rect 36246 43 36646 49
rect 36678 121 36758 135
rect 36678 69 36692 121
rect 36744 69 36758 121
rect 36678 55 36758 69
rect 36960 129 37360 163
rect 37674 197 38074 209
rect 37674 163 37680 197
rect 38068 163 38074 197
rect 36960 83 36978 129
rect 37338 83 37360 129
rect 35964 5 35970 39
rect 36004 5 36020 39
rect 35532 -5 35932 1
rect 34818 -45 35218 -39
rect 35532 -39 35544 -5
rect 35920 -39 35932 -5
rect 35964 -11 36020 5
rect 36678 39 36734 55
rect 36960 49 36972 83
rect 37348 49 37360 83
rect 36960 43 37360 49
rect 37392 121 37472 135
rect 37392 69 37406 121
rect 37458 69 37472 121
rect 37392 55 37472 69
rect 37674 129 38074 163
rect 38388 197 38788 209
rect 39370 205 39390 220
rect 38388 163 38394 197
rect 38782 163 38788 197
rect 37674 83 37692 129
rect 38052 83 38074 129
rect 36678 5 36684 39
rect 36718 5 36734 39
rect 36246 -5 36646 1
rect 35532 -45 35932 -39
rect 36246 -39 36258 -5
rect 36634 -39 36646 -5
rect 36678 -11 36734 5
rect 37392 39 37448 55
rect 37674 49 37686 83
rect 38062 49 38074 83
rect 37674 43 38074 49
rect 38106 121 38186 135
rect 38106 69 38120 121
rect 38172 69 38186 121
rect 38106 55 38186 69
rect 38388 129 38788 163
rect 39369 199 39390 205
rect 39770 199 39790 220
rect 39369 161 39381 199
rect 39778 161 39790 199
rect 39369 160 39390 161
rect 39770 160 39790 161
rect 39369 155 39790 160
rect 39900 210 40320 211
rect 39900 199 39920 210
rect 40300 205 40320 210
rect 40300 199 40321 205
rect 39900 161 39912 199
rect 40309 161 40321 199
rect 39900 150 39920 161
rect 40300 155 40321 161
rect 40300 150 40320 155
rect 38388 83 38406 129
rect 38766 83 38788 129
rect 37392 5 37398 39
rect 37432 5 37448 39
rect 36960 -5 37360 1
rect 36246 -45 36646 -39
rect 36960 -39 36972 -5
rect 37348 -39 37360 -5
rect 37392 -11 37448 5
rect 38106 39 38162 55
rect 38388 49 38400 83
rect 38776 49 38788 83
rect 38388 43 38788 49
rect 38820 121 38900 135
rect 38820 69 38834 121
rect 38886 69 38900 121
rect 38820 55 38900 69
rect 38106 5 38112 39
rect 38146 5 38162 39
rect 37674 -5 38074 1
rect 36960 -45 37360 -39
rect 37674 -39 37686 -5
rect 38062 -39 38074 -5
rect 38106 -11 38162 5
rect 38820 39 38876 55
rect 39900 50 40320 51
rect 39370 39 39390 50
rect 38820 5 38826 39
rect 38860 5 38876 39
rect 38388 -5 38788 1
rect 37674 -45 38074 -39
rect 38388 -39 38400 -5
rect 38776 -39 38788 -5
rect 38820 -11 38876 5
rect 39369 33 39390 39
rect 39770 33 39790 50
rect 39369 -5 39381 33
rect 39778 -5 39790 33
rect 39369 -10 39390 -5
rect 39770 -10 39790 -5
rect 39369 -11 39790 -10
rect 39900 33 39920 50
rect 40300 39 40320 50
rect 40300 33 40321 39
rect 39900 -5 39912 33
rect 40309 -5 40321 33
rect 39900 -10 39920 -5
rect 40300 -10 40321 -5
rect 39900 -11 40321 -10
rect 38388 -45 38788 -39
rect 15547 -50 15927 -45
rect 3670 -138 3858 -132
rect 3670 -526 3704 -138
rect 3738 -144 3858 -138
rect 3738 -156 3818 -144
rect 3738 -520 3818 -506
rect 3852 -520 3858 -144
rect 3738 -526 3858 -520
rect 3670 -532 3858 -526
rect 3900 -139 3946 -132
rect 3900 -144 4061 -139
rect 3900 -520 3906 -144
rect 3940 -149 4061 -144
rect 3940 -519 3951 -149
rect 4051 -519 4061 -149
rect 15547 -140 15557 -50
rect 15917 -140 15927 -50
rect 15547 -150 15927 -140
rect 16261 -50 16641 -45
rect 16261 -140 16271 -50
rect 16631 -140 16641 -50
rect 16261 -150 16641 -140
rect 16975 -50 17355 -45
rect 16975 -140 16985 -50
rect 17345 -140 17355 -50
rect 16975 -150 17355 -140
rect 17689 -50 18069 -45
rect 17689 -140 17699 -50
rect 18059 -140 18069 -50
rect 17689 -150 18069 -140
rect 18403 -50 18783 -45
rect 18403 -140 18413 -50
rect 18773 -140 18783 -50
rect 18403 -150 18783 -140
rect 19117 -50 19497 -45
rect 19117 -140 19127 -50
rect 19487 -140 19497 -50
rect 19117 -150 19497 -140
rect 19831 -50 20211 -45
rect 19831 -140 19841 -50
rect 20201 -140 20211 -50
rect 19831 -150 20211 -140
rect 20545 -50 20925 -45
rect 20545 -140 20555 -50
rect 20915 -140 20925 -50
rect 20545 -150 20925 -140
rect 21259 -50 21639 -45
rect 21259 -140 21269 -50
rect 21629 -140 21639 -50
rect 21259 -150 21639 -140
rect 21973 -50 22353 -45
rect 21973 -140 21983 -50
rect 22343 -140 22353 -50
rect 21973 -150 22353 -140
rect 22687 -50 23067 -45
rect 22687 -140 22697 -50
rect 23057 -140 23067 -50
rect 22687 -150 23067 -140
rect 23401 -50 23781 -45
rect 23401 -140 23411 -50
rect 23771 -140 23781 -50
rect 23401 -150 23781 -140
rect 24115 -50 24495 -45
rect 24115 -140 24125 -50
rect 24485 -140 24495 -50
rect 24115 -150 24495 -140
rect 24829 -50 25209 -45
rect 24829 -140 24839 -50
rect 25199 -140 25209 -50
rect 24829 -150 25209 -140
rect 25543 -50 25923 -45
rect 25543 -140 25553 -50
rect 25913 -140 25923 -50
rect 25543 -150 25923 -140
rect 26257 -50 26637 -45
rect 26257 -140 26267 -50
rect 26627 -140 26637 -50
rect 26257 -150 26637 -140
rect 26971 -50 27351 -45
rect 26971 -140 26981 -50
rect 27341 -140 27351 -50
rect 26971 -150 27351 -140
rect 27685 -50 28065 -45
rect 27685 -140 27695 -50
rect 28055 -140 28065 -50
rect 27685 -150 28065 -140
rect 28399 -50 28779 -45
rect 28399 -140 28409 -50
rect 28769 -140 28779 -50
rect 28399 -150 28779 -140
rect 29113 -50 29493 -45
rect 29113 -140 29123 -50
rect 29483 -140 29493 -50
rect 29113 -150 29493 -140
rect 29827 -50 30207 -45
rect 29827 -140 29837 -50
rect 30197 -140 30207 -50
rect 29827 -150 30207 -140
rect 30541 -50 30921 -45
rect 30541 -140 30551 -50
rect 30911 -140 30921 -50
rect 30541 -150 30921 -140
rect 31255 -50 31635 -45
rect 31255 -140 31265 -50
rect 31625 -140 31635 -50
rect 31255 -150 31635 -140
rect 31969 -50 32349 -45
rect 31969 -140 31979 -50
rect 32339 -140 32349 -50
rect 31969 -150 32349 -140
rect 32683 -50 33063 -45
rect 32683 -140 32693 -50
rect 33053 -140 33063 -50
rect 32683 -150 33063 -140
rect 33397 -50 33777 -45
rect 33397 -140 33407 -50
rect 33767 -140 33777 -50
rect 33397 -150 33777 -140
rect 34111 -50 34491 -45
rect 34111 -140 34121 -50
rect 34481 -140 34491 -50
rect 34111 -150 34491 -140
rect 34825 -50 35205 -45
rect 34825 -140 34835 -50
rect 35195 -140 35205 -50
rect 34825 -150 35205 -140
rect 35539 -50 35919 -45
rect 35539 -140 35549 -50
rect 35909 -140 35919 -50
rect 35539 -150 35919 -140
rect 36253 -50 36633 -45
rect 36253 -140 36263 -50
rect 36623 -140 36633 -50
rect 36253 -150 36633 -140
rect 36967 -50 37347 -45
rect 36967 -140 36977 -50
rect 37337 -140 37347 -50
rect 36967 -150 37347 -140
rect 37681 -50 38061 -45
rect 37681 -140 37691 -50
rect 38051 -140 38061 -50
rect 37681 -150 38061 -140
rect 38395 -50 38775 -45
rect 38395 -140 38405 -50
rect 38765 -140 38775 -50
rect 39900 -120 40320 -119
rect 39370 -127 39390 -120
rect 38395 -150 38775 -140
rect 39369 -133 39390 -127
rect 39770 -133 39790 -120
rect 39369 -171 39381 -133
rect 39778 -171 39790 -133
rect 39369 -177 39390 -171
rect 39370 -180 39390 -177
rect 39770 -180 39790 -171
rect 39900 -133 39920 -120
rect 40300 -127 40320 -120
rect 40300 -133 40321 -127
rect 39900 -171 39912 -133
rect 40309 -171 40321 -133
rect 39900 -180 39920 -171
rect 40300 -177 40321 -171
rect 40300 -180 40320 -177
rect 10200 -383 10296 -354
rect 10200 -400 10231 -383
rect 3940 -520 4061 -519
rect 3900 -529 4061 -520
rect 10020 -417 10231 -400
rect 10265 -417 10296 -383
rect 10020 -420 10296 -417
rect 10744 -383 10840 -354
rect 10744 -417 10775 -383
rect 10809 -400 10840 -383
rect 10809 -417 10980 -400
rect 10744 -420 10980 -417
rect 3900 -532 3946 -529
rect 3766 -570 3912 -564
rect 3766 -578 3862 -570
rect 3766 -630 3780 -578
rect 3832 -604 3862 -578
rect 3896 -604 3912 -570
rect 3832 -620 3912 -604
rect 3832 -630 3846 -620
rect 3766 -644 3846 -630
rect 10020 -740 10040 -420
rect 10160 -475 10296 -420
rect 10160 -509 10231 -475
rect 10265 -509 10296 -475
rect 10160 -567 10296 -509
rect 10160 -601 10231 -567
rect 10265 -601 10296 -567
rect 10160 -659 10296 -601
rect 10160 -693 10231 -659
rect 10265 -693 10296 -659
rect 10160 -740 10296 -693
rect 10480 -440 10640 -420
rect 10480 -700 10500 -440
rect 10620 -700 10640 -440
rect 10480 -720 10640 -700
rect 10744 -475 10800 -420
rect 10744 -509 10775 -475
rect 10744 -567 10800 -509
rect 10744 -601 10775 -567
rect 10744 -659 10800 -601
rect 10744 -693 10775 -659
rect 10020 -751 10296 -740
rect 10020 -760 10231 -751
rect 10200 -785 10231 -760
rect 10265 -785 10296 -751
rect 10744 -740 10800 -693
rect 10960 -740 10980 -420
rect 10744 -751 10980 -740
rect 10200 -843 10296 -785
rect 10546 -786 10552 -775
rect 10514 -827 10552 -786
rect 10604 -786 10610 -775
rect 10744 -785 10775 -751
rect 10809 -760 10980 -751
rect 10809 -785 10840 -760
rect 10604 -827 10616 -786
rect 10514 -834 10616 -827
rect 10200 -877 10231 -843
rect 10265 -877 10296 -843
rect 10200 -935 10296 -877
rect 10200 -969 10231 -935
rect 10265 -969 10296 -935
rect 10200 -1027 10296 -969
rect 10200 -1061 10231 -1027
rect 10265 -1061 10296 -1027
rect 10200 -1119 10296 -1061
rect 10744 -843 10840 -785
rect 10744 -877 10775 -843
rect 10809 -877 10840 -843
rect 10744 -935 10840 -877
rect 11200 -790 11300 -780
rect 11200 -870 11210 -790
rect 11290 -870 11300 -790
rect 11200 -880 11300 -870
rect 10744 -969 10775 -935
rect 10809 -969 10840 -935
rect 10744 -1027 10840 -969
rect 10744 -1061 10775 -1027
rect 10809 -1061 10840 -1027
rect 10200 -1153 10231 -1119
rect 10265 -1153 10296 -1119
rect 10531 -1120 10589 -1107
rect 10744 -1119 10840 -1061
rect 10200 -1211 10296 -1153
rect 10200 -1245 10231 -1211
rect 10265 -1245 10296 -1211
rect 10200 -1303 10296 -1245
rect 10480 -1122 10640 -1120
rect 10480 -1130 10540 -1122
rect 10580 -1130 10640 -1122
rect 10480 -1240 10490 -1130
rect 10630 -1240 10640 -1130
rect 10480 -1242 10540 -1240
rect 10580 -1242 10640 -1240
rect 10480 -1250 10640 -1242
rect 10744 -1153 10775 -1119
rect 10809 -1153 10840 -1119
rect 10744 -1211 10840 -1153
rect 10744 -1245 10775 -1211
rect 10809 -1245 10840 -1211
rect 10531 -1257 10589 -1250
rect 10200 -1337 10231 -1303
rect 10265 -1337 10296 -1303
rect 10200 -1366 10296 -1337
rect 10744 -1303 10840 -1245
rect 11230 -1210 11270 -880
rect 11380 -1090 11480 -1080
rect 11380 -1170 11390 -1090
rect 11470 -1110 11480 -1090
rect 11470 -1150 11571 -1110
rect 11470 -1170 11480 -1150
rect 11380 -1180 11480 -1170
rect 11230 -1250 11503 -1210
rect 10744 -1337 10775 -1303
rect 10809 -1337 10840 -1303
rect 10744 -1366 10840 -1337
rect 11463 -2916 11503 -1250
rect 10382 -2940 10622 -2920
rect 6800 -3020 6960 -3000
rect 6800 -4240 6820 -3020
rect 6880 -3248 6960 -3020
rect 9040 -3020 9200 -3000
rect 7117 -3188 8883 -3182
rect 7117 -3222 7129 -3188
rect 7497 -3222 7587 -3188
rect 7955 -3222 8045 -3188
rect 8413 -3222 8503 -3188
rect 8871 -3222 8883 -3188
rect 7117 -3228 8883 -3222
rect 9040 -3248 9120 -3020
rect 6880 -3260 6993 -3248
rect 9007 -3260 9120 -3248
rect 6880 -3660 6953 -3260
rect 6987 -3272 7110 -3260
rect 6987 -3660 7058 -3272
rect 6880 -3672 6993 -3660
rect 6880 -4240 6960 -3672
rect 5850 -4304 5964 -4298
rect 5850 -4338 5918 -4304
rect 5952 -4338 5964 -4304
rect 5850 -4344 5964 -4338
rect 6020 -4304 6436 -4298
rect 6020 -4338 6036 -4304
rect 6070 -4338 6154 -4304
rect 6188 -4338 6272 -4304
rect 6306 -4338 6390 -4304
rect 6424 -4338 6436 -4304
rect 6020 -4344 6436 -4338
rect 6496 -4304 6610 -4298
rect 6800 -4300 6960 -4240
rect 6496 -4338 6508 -4304
rect 6542 -4338 6610 -4304
rect 6496 -4344 6610 -4338
rect 5739 -4376 5785 -4364
rect 5850 -4376 5902 -4344
rect 6558 -4376 6610 -4344
rect 6700 -4364 6960 -4300
rect 6675 -4376 6960 -4364
rect 5739 -4776 5745 -4376
rect 5779 -4388 5902 -4376
rect 5779 -4776 5850 -4388
rect 5739 -4788 5785 -4776
rect 5170 -5640 5320 -5620
rect 5170 -6030 5190 -5640
rect 5300 -6030 5320 -5640
rect 5170 -6050 5320 -6030
rect 5400 -5640 5550 -5620
rect 5400 -6030 5420 -5640
rect 5530 -6030 5550 -5640
rect 5400 -6050 5550 -6030
rect 5739 -5976 5785 -5964
rect 5739 -6376 5745 -5976
rect 5779 -6364 5850 -5976
rect 5779 -6376 5902 -6364
rect 5968 -4388 6020 -4376
rect 5968 -6376 6020 -6364
rect 6086 -4388 6138 -4376
rect 6086 -6376 6138 -6364
rect 6204 -4388 6256 -4376
rect 6204 -6376 6256 -6364
rect 6322 -4388 6374 -4376
rect 6322 -6376 6374 -6364
rect 6440 -4388 6492 -4376
rect 6440 -6376 6492 -6364
rect 6558 -4388 6681 -4376
rect 6610 -4776 6681 -4388
rect 6715 -4776 6960 -4376
rect 6675 -4788 6960 -4776
rect 6700 -4848 6960 -4788
rect 6700 -4860 6993 -4848
rect 6700 -4900 6953 -4860
rect 6800 -5260 6953 -4900
rect 6987 -5248 7058 -4860
rect 6987 -5260 7110 -5248
rect 7516 -3272 7568 -3260
rect 7516 -5260 7568 -5248
rect 7974 -3272 8026 -3260
rect 7974 -5260 8026 -5248
rect 8432 -3272 8484 -3260
rect 8432 -5260 8484 -5248
rect 8890 -3272 9013 -3260
rect 8942 -3660 9013 -3272
rect 9047 -3660 9120 -3260
rect 9007 -3672 9120 -3660
rect 9040 -4240 9120 -3672
rect 9180 -4240 9200 -3020
rect 10382 -3860 10402 -2940
rect 10602 -3860 10622 -2940
rect 10964 -3139 10983 -3130
rect 10964 -3192 10980 -3139
rect 10964 -3200 10983 -3192
rect 11412 -3200 11435 -3130
rect 10382 -3880 10622 -3860
rect 10744 -3484 11352 -3478
rect 10744 -3518 10864 -3484
rect 11340 -3518 11352 -3484
rect 10744 -3524 11352 -3518
rect 10744 -3670 10784 -3524
rect 10852 -3580 11352 -3574
rect 11469 -3580 11503 -2916
rect 10852 -3614 10864 -3580
rect 11340 -3614 11352 -3580
rect 10852 -3620 11352 -3614
rect 11384 -3610 11503 -3580
rect 11384 -3644 11390 -3610
rect 11424 -3614 11503 -3610
rect 11531 -2916 11571 -1150
rect 11424 -3644 11430 -3614
rect 11384 -3660 11430 -3644
rect 10744 -3676 11352 -3670
rect 10744 -3710 10864 -3676
rect 11340 -3710 11352 -3676
rect 10744 -3716 11352 -3710
rect 10744 -3862 10784 -3716
rect 10852 -3772 10867 -3763
rect 11336 -3772 11353 -3763
rect 11531 -3772 11565 -2916
rect 10852 -3806 10864 -3772
rect 11340 -3806 11353 -3772
rect 10852 -3815 10867 -3806
rect 11336 -3815 11353 -3806
rect 11384 -3802 11565 -3772
rect 11384 -3836 11390 -3802
rect 11424 -3806 11565 -3802
rect 11424 -3836 11430 -3806
rect 11384 -3852 11430 -3836
rect 10744 -3868 11352 -3862
rect 10744 -3902 10864 -3868
rect 11340 -3902 11352 -3868
rect 10744 -3908 11352 -3902
rect 9040 -4300 9200 -4240
rect 9040 -4364 9300 -4300
rect 9391 -4304 9505 -4298
rect 9391 -4338 9459 -4304
rect 9493 -4338 9505 -4304
rect 9391 -4344 9505 -4338
rect 9565 -4304 9981 -4298
rect 9565 -4338 9577 -4304
rect 9611 -4338 9695 -4304
rect 9729 -4338 9813 -4304
rect 9847 -4338 9931 -4304
rect 9965 -4338 9981 -4304
rect 9565 -4344 9981 -4338
rect 10033 -4304 10151 -4298
rect 10033 -4338 10049 -4304
rect 10083 -4338 10151 -4304
rect 10033 -4344 10151 -4338
rect 9040 -4376 9326 -4364
rect 9391 -4376 9443 -4344
rect 10099 -4376 10151 -4344
rect 10216 -4376 10262 -4364
rect 9040 -4776 9286 -4376
rect 9320 -4388 9443 -4376
rect 9320 -4776 9391 -4388
rect 9040 -4788 9326 -4776
rect 9040 -4800 9300 -4788
rect 9000 -4860 9300 -4800
rect 8942 -5248 9013 -4860
rect 8890 -5260 9013 -5248
rect 9047 -4900 9300 -4860
rect 9047 -5260 9200 -4900
rect 6800 -5272 6993 -5260
rect 6800 -5700 6960 -5272
rect 8880 -5292 8944 -5290
rect 7117 -5298 8944 -5292
rect 7117 -5332 7129 -5298
rect 7497 -5332 7587 -5298
rect 7955 -5332 8045 -5298
rect 8413 -5332 8503 -5298
rect 8871 -5332 8880 -5298
rect 7117 -5338 8880 -5332
rect 8880 -5370 8944 -5362
rect 9000 -5400 9200 -5260
rect 7289 -5656 7295 -5600
rect 7361 -5656 7367 -5600
rect 7481 -5656 7487 -5600
rect 7553 -5656 7559 -5600
rect 7673 -5656 7679 -5600
rect 7745 -5656 7751 -5600
rect 7865 -5656 7871 -5600
rect 7937 -5656 7943 -5600
rect 8057 -5656 8063 -5600
rect 8129 -5656 8135 -5600
rect 8249 -5656 8255 -5600
rect 8321 -5656 8327 -5600
rect 8441 -5656 8447 -5600
rect 8513 -5656 8519 -5600
rect 8633 -5656 8639 -5600
rect 8705 -5656 8711 -5600
rect 9040 -5700 9200 -5400
rect 6800 -5800 6909 -5700
rect 6700 -5964 6909 -5800
rect 6675 -5976 6909 -5964
rect 6610 -6364 6681 -5976
rect 6558 -6376 6681 -6364
rect 6715 -6200 6909 -5976
rect 6943 -6200 7013 -5700
rect 7067 -6200 7073 -5700
rect 7103 -6200 7109 -5700
rect 7163 -6200 7169 -5700
rect 7199 -6200 7205 -5700
rect 7259 -6200 7265 -5700
rect 7295 -6200 7301 -5700
rect 7355 -6200 7361 -5700
rect 7391 -6200 7397 -5700
rect 7451 -6200 7457 -5700
rect 7487 -6200 7493 -5700
rect 7547 -6200 7553 -5700
rect 7583 -6200 7589 -5700
rect 7643 -6200 7649 -5700
rect 7679 -6200 7685 -5700
rect 7739 -6200 7745 -5700
rect 7775 -6200 7781 -5700
rect 7835 -6200 7841 -5700
rect 7871 -6200 7877 -5700
rect 7931 -6200 7937 -5700
rect 7967 -6200 7973 -5700
rect 8027 -6200 8033 -5700
rect 8063 -6200 8069 -5700
rect 8123 -6200 8129 -5700
rect 8159 -6200 8165 -5700
rect 8219 -6200 8225 -5700
rect 8255 -6200 8261 -5700
rect 8315 -6200 8321 -5700
rect 8351 -6200 8357 -5700
rect 8411 -6200 8417 -5700
rect 8447 -6200 8453 -5700
rect 8507 -6200 8513 -5700
rect 8543 -6200 8549 -5700
rect 8603 -6200 8609 -5700
rect 8639 -6200 8645 -5700
rect 8699 -6200 8705 -5700
rect 8735 -6200 8741 -5700
rect 8795 -6200 8801 -5700
rect 8831 -6200 8837 -5700
rect 8891 -6200 8897 -5700
rect 8927 -6200 8933 -5700
rect 8987 -6200 9057 -5700
rect 9091 -5800 9200 -5700
rect 9091 -5964 9300 -5800
rect 9091 -5976 9326 -5964
rect 9091 -6200 9286 -5976
rect 6715 -6300 6960 -6200
rect 7017 -6236 7063 -6200
rect 7113 -6236 7159 -6200
rect 8841 -6236 8887 -6200
rect 8937 -6236 8983 -6200
rect 7017 -6242 7169 -6236
rect 7017 -6276 7119 -6242
rect 7153 -6276 7169 -6242
rect 7017 -6282 7169 -6276
rect 8831 -6242 8983 -6236
rect 8831 -6276 8847 -6242
rect 8881 -6276 8983 -6242
rect 8831 -6282 8983 -6276
rect 9040 -6300 9286 -6200
rect 6715 -6376 6800 -6300
rect 5739 -6388 5785 -6376
rect 5850 -6408 5902 -6376
rect 6558 -6408 6610 -6376
rect 6675 -6388 6800 -6376
rect 6700 -6400 6800 -6388
rect 9200 -6376 9286 -6300
rect 9320 -6364 9391 -5976
rect 9320 -6376 9443 -6364
rect 9509 -4388 9561 -4376
rect 9509 -6376 9561 -6364
rect 9627 -4388 9679 -4376
rect 9627 -6376 9679 -6364
rect 9745 -4388 9797 -4376
rect 9745 -6376 9797 -6364
rect 9863 -4388 9915 -4376
rect 9863 -6376 9915 -6364
rect 9981 -4388 10033 -4376
rect 9981 -6376 10033 -6364
rect 10099 -4388 10222 -4376
rect 10151 -4776 10222 -4388
rect 10256 -4776 10262 -4376
rect 10216 -4788 10262 -4776
rect 10216 -5976 10262 -5964
rect 10151 -6364 10222 -5976
rect 10099 -6376 10222 -6364
rect 10256 -6376 10262 -5976
rect 9200 -6388 9326 -6376
rect 9200 -6400 9300 -6388
rect 5850 -6414 5964 -6408
rect 5850 -6448 5918 -6414
rect 5952 -6448 5964 -6414
rect 5850 -6454 5964 -6448
rect 6020 -6414 6436 -6408
rect 6020 -6448 6036 -6414
rect 6070 -6448 6154 -6414
rect 6188 -6448 6272 -6414
rect 6306 -6448 6390 -6414
rect 6424 -6448 6436 -6414
rect 6020 -6454 6436 -6448
rect 6496 -6414 6610 -6408
rect 6496 -6448 6508 -6414
rect 6542 -6448 6610 -6414
rect 6496 -6454 6610 -6448
rect 9391 -6408 9443 -6376
rect 10099 -6408 10151 -6376
rect 10216 -6388 10262 -6376
rect 9391 -6414 9505 -6408
rect 9391 -6448 9459 -6414
rect 9493 -6448 9505 -6414
rect 9391 -6454 9505 -6448
rect 9565 -6414 9981 -6408
rect 9565 -6448 9577 -6414
rect 9611 -6448 9695 -6414
rect 9729 -6448 9813 -6414
rect 9847 -6448 9931 -6414
rect 9965 -6448 9981 -6414
rect 9565 -6454 9981 -6448
rect 10033 -6414 10151 -6408
rect 10033 -6448 10049 -6414
rect 10083 -6448 10151 -6414
rect 10033 -6454 10151 -6448
rect 6204 -6506 6256 -6454
rect 6204 -6564 6256 -6558
rect 9745 -6506 9797 -6454
rect 9745 -6564 9797 -6558
rect 7911 -6798 7917 -6748
rect 6086 -6804 6204 -6798
rect 6086 -6838 6154 -6804
rect 6188 -6838 6204 -6804
rect 6086 -6844 6204 -6838
rect 6256 -6804 7502 -6798
rect 6256 -6838 6272 -6804
rect 6306 -6838 6390 -6804
rect 6424 -6838 6508 -6804
rect 6542 -6838 6626 -6804
rect 6660 -6838 6744 -6804
rect 6778 -6838 6862 -6804
rect 6896 -6838 6980 -6804
rect 7014 -6838 7098 -6804
rect 7132 -6838 7216 -6804
rect 7250 -6838 7334 -6804
rect 7368 -6838 7452 -6804
rect 7486 -6838 7502 -6804
rect 6256 -6844 7502 -6838
rect 7554 -6800 7917 -6798
rect 7969 -6800 7975 -6748
rect 8026 -6792 8092 -6781
rect 7554 -6804 7970 -6800
rect 7554 -6838 7570 -6804
rect 7604 -6838 7688 -6804
rect 7722 -6838 7806 -6804
rect 7840 -6838 7924 -6804
rect 7958 -6838 7970 -6804
rect 7554 -6844 7970 -6838
rect 8026 -6844 8032 -6792
rect 8084 -6798 8092 -6792
rect 8084 -6804 8446 -6798
rect 8084 -6838 8160 -6804
rect 8194 -6838 8278 -6804
rect 8312 -6838 8396 -6804
rect 8430 -6838 8446 -6804
rect 8084 -6844 8446 -6838
rect 8498 -6804 9744 -6798
rect 8498 -6838 8514 -6804
rect 8548 -6838 8632 -6804
rect 8666 -6838 8750 -6804
rect 8784 -6838 8868 -6804
rect 8902 -6838 8986 -6804
rect 9020 -6838 9104 -6804
rect 9138 -6838 9222 -6804
rect 9256 -6838 9340 -6804
rect 9374 -6838 9458 -6804
rect 9492 -6838 9576 -6804
rect 9610 -6838 9694 -6804
rect 9728 -6838 9744 -6804
rect 8498 -6844 9744 -6838
rect 9796 -6804 9914 -6798
rect 9796 -6838 9812 -6804
rect 9846 -6838 9914 -6804
rect 9796 -6844 9914 -6838
rect 5975 -6885 6021 -6873
rect 6086 -6885 6138 -6844
rect 5975 -7285 5981 -6885
rect 6015 -6897 6138 -6885
rect 6015 -7285 6086 -6897
rect 5975 -7297 6021 -7285
rect 5975 -8485 6021 -8473
rect 5975 -8885 5981 -8485
rect 6015 -8873 6086 -8485
rect 6015 -8885 6138 -8873
rect 6204 -6897 6256 -6885
rect 6204 -8885 6256 -8873
rect 6322 -6897 6374 -6885
rect 6322 -8885 6374 -8873
rect 6440 -6897 6492 -6885
rect 6440 -8885 6492 -8873
rect 6558 -6897 6610 -6885
rect 6558 -8885 6610 -8873
rect 6676 -6897 6728 -6885
rect 6676 -8885 6728 -8873
rect 6794 -6897 6846 -6885
rect 6794 -8885 6846 -8873
rect 6912 -6897 6964 -6885
rect 6912 -8885 6964 -8873
rect 7030 -6897 7082 -6885
rect 7030 -8885 7082 -8873
rect 7148 -6897 7200 -6885
rect 7148 -8885 7200 -8873
rect 7266 -6897 7318 -6885
rect 7266 -8885 7318 -8873
rect 7384 -6897 7436 -6844
rect 8026 -6850 8092 -6844
rect 5975 -8897 6021 -8885
rect 6086 -8926 6138 -8885
rect 7384 -8926 7436 -8873
rect 7502 -6897 7554 -6885
rect 7502 -8885 7554 -8873
rect 7620 -6897 7672 -6885
rect 7620 -8886 7672 -8873
rect 7738 -6897 7790 -6885
rect 7738 -8885 7790 -8873
rect 7856 -6897 7908 -6885
rect 7856 -8885 7908 -8873
rect 7974 -6897 8026 -6885
rect 7974 -8885 8026 -8873
rect 8092 -6897 8144 -6885
rect 8092 -8885 8144 -8873
rect 8210 -6897 8262 -6885
rect 8210 -8885 8262 -8873
rect 8328 -6897 8380 -6885
rect 8328 -8886 8380 -8873
rect 8446 -6897 8498 -6885
rect 8446 -8885 8498 -8873
rect 8564 -6897 8616 -6844
rect 8564 -8926 8616 -8873
rect 8682 -6897 8734 -6885
rect 8682 -8885 8734 -8873
rect 8800 -6897 8852 -6885
rect 8800 -8885 8852 -8873
rect 8918 -6897 8970 -6885
rect 8918 -8885 8970 -8873
rect 9036 -6897 9088 -6885
rect 9036 -8885 9088 -8873
rect 9154 -6897 9206 -6885
rect 9154 -8885 9206 -8873
rect 9272 -6897 9324 -6885
rect 9272 -8885 9324 -8873
rect 9390 -6897 9442 -6885
rect 9390 -8885 9442 -8873
rect 9508 -6897 9560 -6885
rect 9508 -8885 9560 -8873
rect 9626 -6897 9678 -6885
rect 9626 -8885 9678 -8873
rect 9744 -6897 9796 -6884
rect 9744 -8885 9796 -8873
rect 9862 -6885 9914 -6844
rect 9979 -6885 10025 -6873
rect 9862 -6897 9985 -6885
rect 9914 -7285 9985 -6897
rect 10019 -7285 10025 -6885
rect 9979 -7297 10025 -7285
rect 9979 -8485 10025 -8473
rect 9914 -8873 9985 -8485
rect 9862 -8885 9985 -8873
rect 10019 -8885 10025 -8485
rect 9862 -8926 9914 -8885
rect 9979 -8897 10025 -8885
rect 6086 -8932 6204 -8926
rect 6086 -8966 6154 -8932
rect 6188 -8966 6204 -8932
rect 6086 -8972 6204 -8966
rect 6256 -8932 7502 -8926
rect 6256 -8966 6272 -8932
rect 6306 -8966 6390 -8932
rect 6424 -8966 6508 -8932
rect 6542 -8966 6626 -8932
rect 6660 -8966 6744 -8932
rect 6778 -8966 6862 -8932
rect 6896 -8966 6980 -8932
rect 7014 -8966 7098 -8932
rect 7132 -8966 7216 -8932
rect 7250 -8966 7334 -8932
rect 7368 -8966 7452 -8932
rect 7486 -8966 7502 -8932
rect 6256 -8972 7502 -8966
rect 8498 -8932 9744 -8926
rect 8498 -8966 8514 -8932
rect 8548 -8966 8632 -8932
rect 8666 -8966 8750 -8932
rect 8784 -8966 8868 -8932
rect 8902 -8966 8986 -8932
rect 9020 -8966 9104 -8932
rect 9138 -8966 9222 -8932
rect 9256 -8966 9340 -8932
rect 9374 -8966 9458 -8932
rect 9492 -8966 9576 -8932
rect 9610 -8966 9694 -8932
rect 9728 -8966 9744 -8932
rect 8498 -8972 9744 -8966
rect 9796 -8932 9914 -8926
rect 9796 -8966 9812 -8932
rect 9846 -8966 9914 -8932
rect 9796 -8972 9914 -8966
<< via1 >>
rect 6086 10297 6095 12273
rect 6095 10297 6129 12273
rect 6129 10297 6138 12273
rect 6204 10297 6213 12273
rect 6213 10297 6247 12273
rect 6247 10297 6256 12273
rect 6322 10297 6331 12273
rect 6331 10297 6365 12273
rect 6365 10297 6374 12273
rect 6440 10297 6449 12273
rect 6449 10297 6483 12273
rect 6483 10297 6492 12273
rect 6558 10297 6567 12273
rect 6567 10297 6601 12273
rect 6601 10297 6610 12273
rect 6676 10297 6685 12273
rect 6685 10297 6719 12273
rect 6719 10297 6728 12273
rect 6794 10297 6803 12273
rect 6803 10297 6837 12273
rect 6837 10297 6846 12273
rect 6912 10297 6921 12273
rect 6921 10297 6955 12273
rect 6955 10297 6964 12273
rect 7030 10297 7039 12273
rect 7039 10297 7073 12273
rect 7073 10297 7082 12273
rect 7148 10297 7157 12273
rect 7157 10297 7191 12273
rect 7191 10297 7200 12273
rect 7266 10297 7275 12273
rect 7275 10297 7309 12273
rect 7309 10297 7318 12273
rect 7384 10297 7393 12273
rect 7393 10297 7427 12273
rect 7427 10297 7436 12273
rect 7502 10297 7511 12273
rect 7511 10297 7545 12273
rect 7545 10297 7554 12273
rect 7620 10297 7629 12273
rect 7629 10297 7663 12273
rect 7663 10297 7672 12273
rect 7738 10297 7747 12273
rect 7747 10297 7781 12273
rect 7781 10297 7790 12273
rect 7856 10297 7865 12273
rect 7865 10297 7899 12273
rect 7899 10297 7908 12273
rect 7974 10297 7983 12273
rect 7983 10297 8017 12273
rect 8017 10297 8026 12273
rect 8092 10297 8101 12273
rect 8101 10297 8135 12273
rect 8135 10297 8144 12273
rect 8210 10297 8219 12273
rect 8219 10297 8253 12273
rect 8253 10297 8262 12273
rect 8328 10297 8337 12273
rect 8337 10297 8371 12273
rect 8371 10297 8380 12273
rect 8446 10297 8455 12273
rect 8455 10297 8489 12273
rect 8489 10297 8498 12273
rect 8564 10297 8573 12273
rect 8573 10297 8607 12273
rect 8607 10297 8616 12273
rect 8682 10297 8691 12273
rect 8691 10297 8725 12273
rect 8725 10297 8734 12273
rect 8800 10297 8809 12273
rect 8809 10297 8843 12273
rect 8843 10297 8852 12273
rect 8918 10297 8927 12273
rect 8927 10297 8961 12273
rect 8961 10297 8970 12273
rect 9036 10297 9045 12273
rect 9045 10297 9079 12273
rect 9079 10297 9088 12273
rect 9154 10297 9163 12273
rect 9163 10297 9197 12273
rect 9197 10297 9206 12273
rect 9272 10297 9281 12273
rect 9281 10297 9315 12273
rect 9315 10297 9324 12273
rect 9390 10297 9399 12273
rect 9399 10297 9433 12273
rect 9433 10297 9442 12273
rect 9508 10297 9517 12273
rect 9517 10297 9551 12273
rect 9551 10297 9560 12273
rect 9626 10297 9635 12273
rect 9635 10297 9669 12273
rect 9669 10297 9678 12273
rect 9744 10297 9753 12273
rect 9753 10297 9787 12273
rect 9787 10297 9796 12273
rect 9862 10297 9871 12273
rect 9871 10297 9905 12273
rect 9905 10297 9914 12273
rect 7917 10148 7969 10200
rect 8032 10238 8084 10244
rect 8032 10204 8042 10238
rect 8042 10204 8076 10238
rect 8076 10204 8084 10238
rect 8032 10192 8084 10204
rect 6204 9906 6256 9958
rect 9745 9906 9797 9958
rect 5190 9040 5300 9430
rect 5420 9040 5530 9430
rect 5850 7788 5859 9764
rect 5859 7788 5893 9764
rect 5893 7788 5902 9764
rect 5968 7788 5977 9764
rect 5977 7788 6011 9764
rect 6011 7788 6020 9764
rect 6086 7788 6095 9764
rect 6095 7788 6129 9764
rect 6129 7788 6138 9764
rect 6204 7788 6213 9764
rect 6213 7788 6247 9764
rect 6247 7788 6256 9764
rect 6322 7788 6331 9764
rect 6331 7788 6365 9764
rect 6365 7788 6374 9764
rect 6440 7788 6449 9764
rect 6449 7788 6483 9764
rect 6483 7788 6492 9764
rect 6558 7788 6567 9764
rect 6567 7788 6601 9764
rect 6601 7788 6610 9764
rect 7013 9588 7067 9600
rect 7013 9112 7023 9588
rect 7023 9112 7057 9588
rect 7057 9112 7067 9588
rect 7013 9100 7067 9112
rect 7109 9588 7163 9600
rect 7109 9112 7119 9588
rect 7119 9112 7153 9588
rect 7153 9112 7163 9588
rect 7109 9100 7163 9112
rect 7205 9588 7259 9600
rect 7205 9112 7215 9588
rect 7215 9112 7249 9588
rect 7249 9112 7259 9588
rect 7205 9100 7259 9112
rect 7301 9588 7355 9600
rect 7301 9112 7311 9588
rect 7311 9112 7345 9588
rect 7345 9112 7355 9588
rect 7301 9100 7355 9112
rect 7397 9588 7451 9600
rect 7397 9112 7407 9588
rect 7407 9112 7441 9588
rect 7441 9112 7451 9588
rect 7397 9100 7451 9112
rect 7493 9588 7547 9600
rect 7493 9112 7503 9588
rect 7503 9112 7537 9588
rect 7537 9112 7547 9588
rect 7493 9100 7547 9112
rect 7589 9588 7643 9600
rect 7589 9112 7599 9588
rect 7599 9112 7633 9588
rect 7633 9112 7643 9588
rect 7589 9100 7643 9112
rect 7685 9588 7739 9600
rect 7685 9112 7695 9588
rect 7695 9112 7729 9588
rect 7729 9112 7739 9588
rect 7685 9100 7739 9112
rect 7781 9588 7835 9600
rect 7781 9112 7791 9588
rect 7791 9112 7825 9588
rect 7825 9112 7835 9588
rect 7781 9100 7835 9112
rect 7877 9588 7931 9600
rect 7877 9112 7887 9588
rect 7887 9112 7921 9588
rect 7921 9112 7931 9588
rect 7877 9100 7931 9112
rect 7973 9588 8027 9600
rect 7973 9112 7983 9588
rect 7983 9112 8017 9588
rect 8017 9112 8027 9588
rect 7973 9100 8027 9112
rect 8069 9588 8123 9600
rect 8069 9112 8079 9588
rect 8079 9112 8113 9588
rect 8113 9112 8123 9588
rect 8069 9100 8123 9112
rect 8165 9588 8219 9600
rect 8165 9112 8175 9588
rect 8175 9112 8209 9588
rect 8209 9112 8219 9588
rect 8165 9100 8219 9112
rect 8261 9588 8315 9600
rect 8261 9112 8271 9588
rect 8271 9112 8305 9588
rect 8305 9112 8315 9588
rect 8261 9100 8315 9112
rect 8357 9588 8411 9600
rect 8357 9112 8367 9588
rect 8367 9112 8401 9588
rect 8401 9112 8411 9588
rect 8357 9100 8411 9112
rect 8453 9588 8507 9600
rect 8453 9112 8463 9588
rect 8463 9112 8497 9588
rect 8497 9112 8507 9588
rect 8453 9100 8507 9112
rect 8549 9588 8603 9600
rect 8549 9112 8559 9588
rect 8559 9112 8593 9588
rect 8593 9112 8603 9588
rect 8549 9100 8603 9112
rect 8645 9588 8699 9600
rect 8645 9112 8655 9588
rect 8655 9112 8689 9588
rect 8689 9112 8699 9588
rect 8645 9100 8699 9112
rect 8741 9588 8795 9600
rect 8741 9112 8751 9588
rect 8751 9112 8785 9588
rect 8785 9112 8795 9588
rect 8741 9100 8795 9112
rect 8837 9588 8891 9600
rect 8837 9112 8847 9588
rect 8847 9112 8881 9588
rect 8881 9112 8891 9588
rect 8837 9100 8891 9112
rect 8933 9588 8987 9600
rect 8933 9112 8943 9588
rect 8943 9112 8977 9588
rect 8977 9112 8987 9588
rect 8933 9100 8987 9112
rect 7295 9050 7361 9056
rect 7295 9016 7311 9050
rect 7311 9016 7345 9050
rect 7345 9016 7361 9050
rect 7295 9000 7361 9016
rect 7487 9050 7553 9056
rect 7487 9016 7503 9050
rect 7503 9016 7537 9050
rect 7537 9016 7553 9050
rect 7487 9000 7553 9016
rect 7679 9050 7745 9056
rect 7679 9016 7695 9050
rect 7695 9016 7729 9050
rect 7729 9016 7745 9050
rect 7679 9000 7745 9016
rect 7871 9050 7937 9056
rect 7871 9016 7887 9050
rect 7887 9016 7921 9050
rect 7921 9016 7937 9050
rect 7871 9000 7937 9016
rect 8063 9050 8129 9056
rect 8063 9016 8079 9050
rect 8079 9016 8113 9050
rect 8113 9016 8129 9050
rect 8063 9000 8129 9016
rect 8255 9050 8321 9056
rect 8255 9016 8271 9050
rect 8271 9016 8305 9050
rect 8305 9016 8321 9050
rect 8255 9000 8321 9016
rect 8447 9050 8513 9056
rect 8447 9016 8463 9050
rect 8463 9016 8497 9050
rect 8497 9016 8513 9050
rect 8447 9000 8513 9016
rect 8639 9050 8705 9056
rect 8639 9016 8655 9050
rect 8655 9016 8689 9050
rect 8689 9016 8705 9050
rect 8639 9000 8705 9016
rect 8880 8698 8944 8762
rect 6820 6420 6880 7640
rect 7058 6672 7067 8648
rect 7067 6672 7101 8648
rect 7101 6672 7110 8648
rect 7516 6672 7525 8648
rect 7525 6672 7559 8648
rect 7559 6672 7568 8648
rect 7974 6672 7983 8648
rect 7983 6672 8017 8648
rect 8017 6672 8026 8648
rect 8432 6672 8441 8648
rect 8441 6672 8475 8648
rect 8475 6672 8484 8648
rect 8890 6672 8899 8648
rect 8899 6672 8933 8648
rect 8933 6672 8942 8648
rect 9391 7788 9400 9764
rect 9400 7788 9434 9764
rect 9434 7788 9443 9764
rect 9509 7788 9518 9764
rect 9518 7788 9552 9764
rect 9552 7788 9561 9764
rect 9627 7788 9636 9764
rect 9636 7788 9670 9764
rect 9670 7788 9679 9764
rect 9745 7788 9754 9764
rect 9754 7788 9788 9764
rect 9788 7788 9797 9764
rect 9863 7788 9872 9764
rect 9872 7788 9906 9764
rect 9906 7788 9915 9764
rect 9981 7788 9990 9764
rect 9990 7788 10024 9764
rect 10024 7788 10033 9764
rect 10099 7788 10108 9764
rect 10108 7788 10142 9764
rect 10142 7788 10151 9764
rect 9120 6420 9180 7640
rect 10402 6340 10542 7260
rect 10542 6340 10602 7260
rect 10867 7206 11336 7215
rect 10867 7172 11336 7206
rect 10867 7163 11336 7172
rect 10983 6592 11412 6600
rect 10983 6539 11412 6592
rect 10983 6530 11412 6539
rect 11030 4830 11110 4910
rect 11190 4830 11270 4910
rect 3358 3975 3458 4345
rect 3571 3972 3591 4332
rect 3591 3972 3641 4332
rect 4201 3972 4251 4332
rect 4251 3972 4271 4332
rect 4384 3975 4484 4345
rect 3577 3854 3629 3906
rect 4213 3854 4265 3906
rect 11278 3908 14428 3978
rect 3358 3251 3458 3621
rect 3571 3264 3591 3614
rect 3591 3264 3671 3614
rect 3671 3264 3681 3614
rect 4161 3264 4171 3614
rect 4171 3264 4251 3614
rect 4251 3264 4271 3614
rect 4384 3251 4484 3621
rect 3577 3140 3629 3192
rect 4213 3140 4265 3192
rect 5447 2895 5867 2920
rect 6647 2895 7067 2920
rect 7847 2895 8267 2920
rect 9047 2895 9467 2920
rect 5447 2861 5464 2895
rect 5464 2861 5526 2895
rect 5526 2861 5560 2895
rect 5560 2861 5622 2895
rect 5622 2861 5656 2895
rect 5656 2861 5718 2895
rect 5718 2861 5752 2895
rect 5752 2861 5814 2895
rect 5814 2861 5848 2895
rect 5848 2861 5867 2895
rect 6647 2861 6678 2895
rect 6678 2861 6712 2895
rect 6712 2861 6774 2895
rect 6774 2861 6808 2895
rect 6808 2861 6870 2895
rect 6870 2861 6904 2895
rect 6904 2861 6966 2895
rect 6966 2861 7000 2895
rect 7000 2861 7062 2895
rect 7062 2861 7067 2895
rect 7847 2861 7864 2895
rect 7864 2861 7926 2895
rect 7926 2861 7960 2895
rect 7960 2861 8022 2895
rect 8022 2861 8056 2895
rect 8056 2861 8118 2895
rect 8118 2861 8152 2895
rect 8152 2861 8214 2895
rect 8214 2861 8248 2895
rect 8248 2861 8267 2895
rect 9047 2861 9078 2895
rect 9078 2861 9112 2895
rect 9112 2861 9174 2895
rect 9174 2861 9208 2895
rect 9208 2861 9270 2895
rect 9270 2861 9304 2895
rect 9304 2861 9366 2895
rect 9366 2861 9400 2895
rect 9400 2861 9462 2895
rect 9462 2861 9467 2895
rect 5447 2840 5867 2861
rect 6647 2840 7067 2861
rect 7847 2840 8267 2861
rect 9047 2840 9467 2861
rect 2359 2522 2411 2531
rect 2359 2488 2368 2522
rect 2368 2488 2402 2522
rect 2402 2488 2411 2522
rect 2359 2479 2411 2488
rect 2431 2522 2483 2531
rect 2431 2488 2440 2522
rect 2440 2488 2474 2522
rect 2474 2488 2483 2522
rect 2431 2479 2483 2488
rect 3250 2368 3630 2608
rect 3965 2338 4017 2347
rect 3965 2304 3974 2338
rect 3974 2304 4008 2338
rect 4008 2304 4017 2338
rect 3965 2295 4017 2304
rect 4747 2229 5167 2260
rect 6047 2229 6467 2240
rect 7247 2229 7667 2240
rect 8447 2229 8867 2240
rect 9647 2229 10067 2240
rect 4747 2195 4758 2229
rect 4758 2195 4792 2229
rect 4792 2195 4854 2229
rect 4854 2195 4888 2229
rect 4888 2195 4950 2229
rect 4950 2195 4984 2229
rect 4984 2195 5046 2229
rect 5046 2195 5080 2229
rect 5080 2195 5142 2229
rect 5142 2195 5167 2229
rect 6047 2195 6102 2229
rect 6102 2195 6136 2229
rect 6136 2195 6198 2229
rect 6198 2195 6232 2229
rect 6232 2195 6294 2229
rect 6294 2195 6328 2229
rect 6328 2195 6390 2229
rect 6390 2195 6424 2229
rect 6424 2195 6467 2229
rect 7247 2195 7254 2229
rect 7254 2195 7288 2229
rect 7288 2195 7350 2229
rect 7350 2195 7384 2229
rect 7384 2195 7446 2229
rect 7446 2195 7480 2229
rect 7480 2195 7542 2229
rect 7542 2195 7576 2229
rect 7576 2195 7638 2229
rect 7638 2195 7667 2229
rect 8447 2195 8502 2229
rect 8502 2195 8536 2229
rect 8536 2195 8598 2229
rect 8598 2195 8632 2229
rect 8632 2195 8694 2229
rect 8694 2195 8728 2229
rect 8728 2195 8790 2229
rect 8790 2195 8824 2229
rect 8824 2195 8867 2229
rect 9647 2195 9654 2229
rect 9654 2195 9688 2229
rect 9688 2195 9750 2229
rect 9750 2195 9784 2229
rect 9784 2195 9846 2229
rect 9846 2195 9880 2229
rect 9880 2195 9942 2229
rect 9942 2195 9976 2229
rect 9976 2195 10038 2229
rect 10038 2195 10067 2229
rect 4747 2180 5167 2195
rect 6047 2180 6467 2195
rect 7247 2180 7667 2195
rect 8447 2180 8867 2195
rect 9647 2180 10067 2195
rect 3965 2120 4017 2129
rect 3965 2086 3974 2120
rect 3974 2086 4008 2120
rect 4008 2086 4017 2120
rect 3965 2077 4017 2086
rect 2359 1936 2411 1945
rect 2359 1902 2368 1936
rect 2368 1902 2402 1936
rect 2402 1902 2411 1936
rect 2359 1893 2411 1902
rect 2431 1936 2483 1945
rect 2431 1902 2440 1936
rect 2440 1902 2474 1936
rect 2474 1902 2483 1936
rect 2431 1893 2483 1902
rect 3250 1816 3630 2056
rect 4162 1929 4214 1938
rect 4162 1895 4171 1929
rect 4171 1895 4205 1929
rect 4205 1895 4214 1929
rect 4162 1886 4214 1895
rect 4439 1952 4491 1961
rect 4439 1918 4448 1952
rect 4448 1918 4482 1952
rect 4482 1918 4491 1952
rect 4439 1909 4491 1918
rect 4553 1954 4605 1963
rect 4553 1920 4562 1954
rect 4562 1920 4596 1954
rect 4596 1920 4605 1954
rect 4553 1911 4605 1920
rect 4946 1941 4998 1950
rect 4946 1907 4955 1941
rect 4955 1907 4989 1941
rect 4989 1907 4998 1941
rect 4946 1898 4998 1907
rect 6115 1926 6167 1935
rect 6115 1892 6124 1926
rect 6124 1892 6158 1926
rect 6158 1892 6167 1926
rect 6115 1883 6167 1892
rect 4838 1767 4890 1776
rect 4838 1733 4847 1767
rect 4847 1733 4881 1767
rect 4881 1733 4890 1767
rect 4838 1724 4890 1733
rect 5040 1695 5092 1704
rect 5040 1661 5049 1695
rect 5049 1661 5083 1695
rect 5083 1661 5092 1695
rect 5040 1652 5092 1661
rect 8194 1894 8246 1903
rect 8194 1860 8203 1894
rect 8203 1860 8237 1894
rect 8237 1860 8246 1894
rect 8194 1851 8246 1860
rect 9480 1926 9532 1935
rect 9480 1892 9489 1926
rect 9489 1892 9523 1926
rect 9523 1892 9532 1926
rect 9480 1883 9532 1892
rect 9552 1926 9604 1935
rect 9552 1892 9561 1926
rect 9561 1892 9595 1926
rect 9595 1892 9604 1926
rect 9552 1883 9604 1892
rect 9867 1926 9919 1935
rect 9867 1892 9876 1926
rect 9876 1892 9910 1926
rect 9910 1892 9919 1926
rect 9867 1883 9919 1892
rect 9939 1926 9991 1935
rect 9939 1892 9948 1926
rect 9948 1892 9982 1926
rect 9982 1892 9991 1926
rect 9939 1883 9991 1892
rect 10200 1850 10260 1930
rect 8878 1823 8930 1832
rect 8878 1789 8887 1823
rect 8887 1789 8921 1823
rect 8921 1789 8930 1823
rect 8878 1780 8930 1789
rect 8878 1751 8930 1760
rect 8878 1717 8887 1751
rect 8887 1717 8921 1751
rect 8921 1717 8930 1751
rect 8878 1708 8930 1717
rect 10828 2098 10888 2108
rect 10828 1688 10888 2098
rect 10828 1678 10888 1688
rect 10998 2098 11058 2108
rect 10998 1688 11058 2098
rect 10998 1678 11058 1688
rect 11365 1749 11374 3725
rect 11374 1749 11408 3725
rect 11408 1749 11417 3725
rect 11823 1749 11832 3725
rect 11832 1749 11866 3725
rect 11866 1749 11875 3725
rect 12281 1749 12290 3725
rect 12290 1749 12324 3725
rect 12324 1749 12333 3725
rect 12739 1749 12748 3725
rect 12748 1749 12782 3725
rect 12782 1749 12791 3725
rect 13197 1749 13206 3725
rect 13206 1749 13240 3725
rect 13240 1948 13249 3725
rect 13240 1778 13258 1948
rect 13240 1749 13249 1778
rect 13858 1888 13892 2098
rect 13892 1888 13918 2098
rect 13988 2118 14014 2328
rect 14014 2118 14048 2328
rect 12820 1656 13170 1690
rect 5447 1563 5867 1580
rect 6647 1563 7067 1580
rect 7847 1563 8267 1580
rect 9047 1563 9467 1580
rect 12108 1578 12208 1638
rect 12820 1610 13170 1656
rect 13918 1690 13978 1698
rect 13918 1656 13936 1690
rect 13936 1656 13970 1690
rect 13970 1656 13978 1690
rect 13918 1638 13978 1656
rect 5447 1529 5464 1563
rect 5464 1529 5526 1563
rect 5526 1529 5560 1563
rect 5560 1529 5622 1563
rect 5622 1529 5656 1563
rect 5656 1529 5718 1563
rect 5718 1529 5752 1563
rect 5752 1529 5814 1563
rect 5814 1529 5848 1563
rect 5848 1529 5867 1563
rect 6647 1529 6678 1563
rect 6678 1529 6712 1563
rect 6712 1529 6774 1563
rect 6774 1529 6808 1563
rect 6808 1529 6870 1563
rect 6870 1529 6904 1563
rect 6904 1529 6966 1563
rect 6966 1529 7000 1563
rect 7000 1529 7062 1563
rect 7062 1529 7067 1563
rect 7847 1529 7864 1563
rect 7864 1529 7926 1563
rect 7926 1529 7960 1563
rect 7960 1529 8022 1563
rect 8022 1529 8056 1563
rect 8056 1529 8118 1563
rect 8118 1529 8152 1563
rect 8152 1529 8214 1563
rect 8214 1529 8248 1563
rect 8248 1529 8267 1563
rect 9047 1529 9078 1563
rect 9078 1529 9112 1563
rect 9112 1529 9174 1563
rect 9174 1529 9208 1563
rect 9208 1529 9270 1563
rect 9270 1529 9304 1563
rect 9304 1529 9366 1563
rect 9366 1529 9400 1563
rect 9400 1529 9462 1563
rect 9462 1529 9467 1563
rect 14248 1690 14308 1698
rect 14248 1656 14252 1690
rect 14252 1656 14286 1690
rect 14286 1656 14308 1690
rect 14248 1638 14308 1656
rect 5447 1520 5867 1529
rect 6647 1520 7067 1529
rect 7847 1520 8267 1529
rect 9047 1520 9467 1529
rect 1900 1158 2000 1220
rect 1900 1120 2000 1158
rect 2260 1158 2360 1220
rect 2260 1120 2360 1158
rect 2640 1158 2740 1220
rect 2640 1120 2740 1158
rect 3511 1190 3563 1199
rect 3511 1156 3520 1190
rect 3520 1156 3554 1190
rect 3554 1156 3563 1190
rect 3511 1147 3563 1156
rect 3583 1190 3635 1199
rect 3583 1156 3592 1190
rect 3592 1156 3626 1190
rect 3626 1156 3635 1190
rect 3583 1147 3635 1156
rect 4402 1036 4782 1276
rect 8472 1370 8524 1379
rect 8472 1336 8481 1370
rect 8481 1336 8515 1370
rect 8515 1336 8524 1370
rect 8472 1327 8524 1336
rect 8472 1298 8524 1307
rect 8472 1264 8481 1298
rect 8481 1264 8515 1298
rect 8515 1264 8524 1298
rect 8472 1255 8524 1264
rect 8881 1366 8933 1375
rect 8881 1332 8890 1366
rect 8890 1332 8924 1366
rect 8924 1332 8933 1366
rect 8881 1323 8933 1332
rect 12820 1380 13170 1440
rect 12820 1360 13170 1380
rect 13918 1380 13978 1408
rect 13918 1348 13936 1380
rect 13936 1348 13970 1380
rect 13970 1348 13978 1380
rect 14248 1380 14308 1408
rect 14248 1348 14252 1380
rect 14252 1348 14286 1380
rect 14286 1348 14308 1380
rect 8881 1294 8933 1303
rect 8881 1260 8890 1294
rect 8890 1260 8924 1294
rect 8924 1260 8933 1294
rect 8881 1251 8933 1260
rect 5703 1222 5755 1231
rect 5703 1188 5712 1222
rect 5712 1188 5746 1222
rect 5746 1188 5755 1222
rect 5703 1179 5755 1188
rect 6119 1200 6171 1209
rect 6119 1166 6128 1200
rect 6128 1166 6162 1200
rect 6162 1166 6171 1200
rect 6119 1157 6171 1166
rect 8196 1233 8248 1242
rect 8196 1199 8205 1233
rect 8205 1199 8239 1233
rect 8239 1199 8248 1233
rect 8196 1190 8248 1199
rect 9460 1221 9512 1230
rect 9460 1187 9469 1221
rect 9469 1187 9503 1221
rect 9503 1187 9512 1221
rect 9460 1178 9512 1187
rect 9585 1214 9637 1223
rect 9585 1180 9594 1214
rect 9594 1180 9628 1214
rect 9628 1180 9637 1214
rect 9585 1171 9637 1180
rect 10200 1160 10260 1240
rect 5117 1006 5169 1015
rect 5117 972 5126 1006
rect 5126 972 5160 1006
rect 5160 972 5169 1006
rect 5117 963 5169 972
rect 1740 889 1796 920
rect 1796 889 1820 920
rect 2080 889 2106 920
rect 2106 889 2160 920
rect 6047 897 6467 900
rect 7247 897 7667 900
rect 8447 897 8867 900
rect 9647 897 10067 900
rect 1740 800 1820 889
rect 2080 800 2160 889
rect 6047 863 6102 897
rect 6102 863 6136 897
rect 6136 863 6198 897
rect 6198 863 6232 897
rect 6232 863 6294 897
rect 6294 863 6328 897
rect 6328 863 6390 897
rect 6390 863 6424 897
rect 6424 863 6467 897
rect 7247 863 7254 897
rect 7254 863 7288 897
rect 7288 863 7350 897
rect 7350 863 7384 897
rect 7384 863 7446 897
rect 7446 863 7480 897
rect 7480 863 7542 897
rect 7542 863 7576 897
rect 7576 863 7638 897
rect 7638 863 7667 897
rect 8447 863 8502 897
rect 8502 863 8536 897
rect 8536 863 8598 897
rect 8598 863 8632 897
rect 8632 863 8694 897
rect 8694 863 8728 897
rect 8728 863 8790 897
rect 8790 863 8824 897
rect 8824 863 8867 897
rect 9647 863 9654 897
rect 9654 863 9688 897
rect 9688 863 9750 897
rect 9750 863 9784 897
rect 9784 863 9846 897
rect 9846 863 9880 897
rect 9880 863 9942 897
rect 9942 863 9976 897
rect 9976 863 10038 897
rect 10038 863 10067 897
rect 6047 840 6467 863
rect 7247 840 7667 863
rect 8447 840 8867 863
rect 9647 840 10067 863
rect 3768 202 3818 562
rect 3818 202 3838 562
rect 3951 205 4051 575
rect 10449 320 10458 1296
rect 10458 320 10492 1296
rect 10492 320 10501 1296
rect 10907 320 10916 1296
rect 10916 320 10950 1296
rect 10950 320 10959 1296
rect 11365 320 11374 1296
rect 11374 320 11408 1296
rect 11408 320 11417 1296
rect 11823 320 11832 1296
rect 11832 320 11866 1296
rect 11866 320 11875 1296
rect 12281 1268 12290 1296
rect 12278 1168 12290 1268
rect 12281 320 12290 1168
rect 12290 320 12324 1296
rect 12324 1268 12333 1296
rect 12324 1168 12338 1268
rect 12324 320 12333 1168
rect 12739 320 12748 1296
rect 12748 320 12782 1296
rect 12782 320 12791 1296
rect 13197 320 13206 1296
rect 13206 320 13240 1296
rect 13240 1268 13249 1296
rect 13240 1098 13258 1268
rect 13240 320 13249 1098
rect 13858 948 13892 1158
rect 13892 948 13918 1158
rect 14168 1296 14228 1298
rect 14168 1238 14208 1296
rect 14208 1238 14228 1296
rect 13988 718 14014 928
rect 14014 718 14058 928
rect 39390 1029 39770 1040
rect 15557 912 15917 1002
rect 16271 912 16631 1002
rect 16985 912 17345 1002
rect 17699 912 18059 1002
rect 18413 912 18773 1002
rect 19127 912 19487 1002
rect 19841 912 20201 1002
rect 20555 912 20915 1002
rect 21269 912 21629 1002
rect 21983 912 22343 1002
rect 22697 912 23057 1002
rect 23411 912 23771 1002
rect 24125 912 24485 1002
rect 24839 912 25199 1002
rect 25553 912 25913 1002
rect 26267 912 26627 1002
rect 26981 912 27341 1002
rect 27695 912 28055 1002
rect 28409 912 28769 1002
rect 29123 912 29483 1002
rect 29837 912 30197 1002
rect 30551 912 30911 1002
rect 31265 912 31625 1002
rect 31979 912 32339 1002
rect 32693 912 33053 1002
rect 33407 912 33767 1002
rect 34121 912 34481 1002
rect 34835 912 35195 1002
rect 35549 912 35909 1002
rect 36263 912 36623 1002
rect 36977 912 37337 1002
rect 37691 912 38061 1012
rect 38395 912 38765 1012
rect 39390 991 39770 1029
rect 39390 980 39770 991
rect 39920 1029 40300 1040
rect 39920 991 40300 1029
rect 39920 980 40300 991
rect 15558 779 15918 803
rect 15558 733 15918 779
rect 15986 741 16038 793
rect 16272 779 16632 803
rect 16272 733 16632 779
rect 16700 741 16752 793
rect 16986 779 17346 803
rect 16986 733 17346 779
rect 17414 741 17466 793
rect 17700 779 18060 803
rect 17700 733 18060 779
rect 18128 741 18180 793
rect 18414 779 18774 803
rect 18414 733 18774 779
rect 18842 741 18894 793
rect 19128 779 19488 803
rect 19128 733 19488 779
rect 19556 741 19608 793
rect 19842 779 20202 803
rect 19842 733 20202 779
rect 20270 741 20322 793
rect 20556 779 20916 803
rect 20556 733 20916 779
rect 20984 741 21036 793
rect 21270 779 21630 803
rect 21270 733 21630 779
rect 21698 741 21750 793
rect 21984 779 22344 803
rect 21984 733 22344 779
rect 22412 741 22464 793
rect 22698 779 23058 803
rect 22698 733 23058 779
rect 23126 741 23178 793
rect 23412 779 23772 803
rect 23412 733 23772 779
rect 23840 741 23892 793
rect 24126 779 24486 803
rect 24126 733 24486 779
rect 24554 741 24606 793
rect 24840 779 25200 803
rect 24840 733 25200 779
rect 25268 741 25320 793
rect 25554 779 25914 803
rect 25554 733 25914 779
rect 25982 741 26034 793
rect 26268 779 26628 803
rect 26268 733 26628 779
rect 26696 741 26748 793
rect 26982 779 27342 803
rect 26982 733 27342 779
rect 27410 741 27462 793
rect 27696 779 28056 803
rect 27696 733 28056 779
rect 28124 741 28176 793
rect 28410 779 28770 803
rect 28410 733 28770 779
rect 28838 741 28890 793
rect 29124 779 29484 803
rect 29124 733 29484 779
rect 29552 741 29604 793
rect 29838 779 30198 803
rect 29838 733 30198 779
rect 30266 741 30318 793
rect 30552 779 30912 803
rect 30552 733 30912 779
rect 30980 741 31032 793
rect 31266 779 31626 803
rect 31266 733 31626 779
rect 31694 741 31746 793
rect 31980 779 32340 803
rect 31980 733 32340 779
rect 32408 741 32460 793
rect 32694 779 33054 803
rect 32694 733 33054 779
rect 33122 741 33174 793
rect 33408 779 33768 803
rect 33408 733 33768 779
rect 33836 741 33888 793
rect 34122 779 34482 803
rect 34122 733 34482 779
rect 34550 741 34602 793
rect 34836 779 35196 803
rect 34836 733 35196 779
rect 35264 741 35316 793
rect 35550 779 35910 803
rect 35550 733 35910 779
rect 35978 741 36030 793
rect 36264 779 36624 803
rect 36264 733 36624 779
rect 36692 741 36744 793
rect 36978 779 37338 803
rect 36978 733 37338 779
rect 37406 741 37458 793
rect 37698 779 38048 799
rect 37698 699 38048 779
rect 38120 741 38172 793
rect 38408 779 38768 799
rect 38408 729 38768 779
rect 37698 689 38048 699
rect 39390 863 39770 880
rect 39390 825 39770 863
rect 39390 820 39770 825
rect 39920 863 40300 880
rect 39920 825 40300 863
rect 39920 820 40300 825
rect 38834 741 38886 793
rect 39390 697 39770 710
rect 39390 659 39770 697
rect 39390 650 39770 659
rect 39920 697 40300 710
rect 39920 659 40300 697
rect 39920 650 40300 659
rect 39390 531 39770 550
rect 39390 493 39770 531
rect 39390 490 39770 493
rect 39920 531 40300 540
rect 39920 493 40300 531
rect 39920 480 40300 493
rect 39390 365 39770 380
rect 39390 327 39770 365
rect 39390 320 39770 327
rect 39920 365 40300 370
rect 39920 327 40300 365
rect 39920 310 40300 327
rect 3780 84 3832 136
rect 10358 78 14428 158
rect 15558 83 15918 129
rect 15558 59 15918 83
rect 15986 69 16038 121
rect 16272 83 16632 129
rect 16272 59 16632 83
rect 16700 69 16752 121
rect 16986 83 17346 129
rect 16986 59 17346 83
rect 17414 69 17466 121
rect 17700 83 18060 129
rect 17700 59 18060 83
rect 18128 69 18180 121
rect 18414 83 18774 129
rect 18414 59 18774 83
rect 18842 69 18894 121
rect 19128 83 19488 129
rect 19128 59 19488 83
rect 19556 69 19608 121
rect 19842 83 20202 129
rect 19842 59 20202 83
rect 20270 69 20322 121
rect 20556 83 20916 129
rect 20556 59 20916 83
rect 20984 69 21036 121
rect 21270 83 21630 129
rect 21270 59 21630 83
rect 21698 69 21750 121
rect 21984 83 22344 129
rect 21984 59 22344 83
rect 22412 69 22464 121
rect 22698 83 23058 129
rect 22698 59 23058 83
rect 23126 69 23178 121
rect 23412 83 23772 129
rect 23412 59 23772 83
rect 23840 69 23892 121
rect 24126 83 24486 129
rect 24126 59 24486 83
rect 24554 69 24606 121
rect 24840 83 25200 129
rect 24840 59 25200 83
rect 25268 69 25320 121
rect 25554 83 25914 129
rect 25554 59 25914 83
rect 25982 69 26034 121
rect 26268 83 26628 129
rect 26268 59 26628 83
rect 26696 69 26748 121
rect 26982 83 27342 129
rect 26982 59 27342 83
rect 27410 69 27462 121
rect 27696 83 28056 129
rect 27696 59 28056 83
rect 28124 69 28176 121
rect 28410 83 28770 129
rect 28410 59 28770 83
rect 28838 69 28890 121
rect 29124 83 29484 129
rect 29124 59 29484 83
rect 29552 69 29604 121
rect 29838 83 30198 129
rect 29838 59 30198 83
rect 30266 69 30318 121
rect 30552 83 30912 129
rect 30552 59 30912 83
rect 30980 69 31032 121
rect 31266 83 31626 129
rect 31266 59 31626 83
rect 31694 69 31746 121
rect 31980 83 32340 129
rect 31980 59 32340 83
rect 32408 69 32460 121
rect 32694 83 33054 129
rect 32694 59 33054 83
rect 33122 69 33174 121
rect 33408 83 33768 129
rect 33408 59 33768 83
rect 33836 69 33888 121
rect 34122 83 34482 129
rect 34122 59 34482 83
rect 34550 69 34602 121
rect 34836 83 35196 129
rect 34836 59 35196 83
rect 35264 69 35316 121
rect 35550 83 35910 129
rect 35550 59 35910 83
rect 35978 69 36030 121
rect 36264 83 36624 129
rect 36264 59 36624 83
rect 36692 69 36744 121
rect 36978 83 37338 129
rect 36978 59 37338 83
rect 37406 69 37458 121
rect 37692 83 38052 129
rect 37692 59 38052 83
rect 38120 69 38172 121
rect 39390 199 39770 220
rect 39390 161 39770 199
rect 39390 160 39770 161
rect 39920 199 40300 210
rect 39920 161 40300 199
rect 39920 150 40300 161
rect 38406 83 38766 129
rect 38406 59 38766 83
rect 38834 69 38886 121
rect 39390 33 39770 50
rect 39390 -5 39770 33
rect 39390 -10 39770 -5
rect 39920 33 40300 50
rect 39920 -5 40300 33
rect 39920 -10 40300 -5
rect 3728 -506 3738 -156
rect 3738 -506 3818 -156
rect 3818 -506 3838 -156
rect 3951 -519 4051 -149
rect 15557 -140 15917 -50
rect 16271 -140 16631 -50
rect 16985 -140 17345 -50
rect 17699 -140 18059 -50
rect 18413 -140 18773 -50
rect 19127 -140 19487 -50
rect 19841 -140 20201 -50
rect 20555 -140 20915 -50
rect 21269 -140 21629 -50
rect 21983 -140 22343 -50
rect 22697 -140 23057 -50
rect 23411 -140 23771 -50
rect 24125 -140 24485 -50
rect 24839 -140 25199 -50
rect 25553 -140 25913 -50
rect 26267 -140 26627 -50
rect 26981 -140 27341 -50
rect 27695 -140 28055 -50
rect 28409 -140 28769 -50
rect 29123 -140 29483 -50
rect 29837 -140 30197 -50
rect 30551 -140 30911 -50
rect 31265 -140 31625 -50
rect 31979 -140 32339 -50
rect 32693 -140 33053 -50
rect 33407 -140 33767 -50
rect 34121 -140 34481 -50
rect 34835 -140 35195 -50
rect 35549 -140 35909 -50
rect 36263 -140 36623 -50
rect 36977 -140 37337 -50
rect 37691 -140 38051 -50
rect 38405 -140 38765 -50
rect 39390 -133 39770 -120
rect 39390 -171 39770 -133
rect 39390 -180 39770 -171
rect 39920 -133 40300 -120
rect 39920 -171 40300 -133
rect 39920 -180 40300 -171
rect 3780 -630 3832 -578
rect 10040 -740 10160 -420
rect 10500 -478 10620 -440
rect 10500 -598 10540 -478
rect 10540 -598 10580 -478
rect 10580 -598 10620 -478
rect 10500 -700 10620 -598
rect 10800 -475 10960 -420
rect 10800 -509 10809 -475
rect 10809 -509 10960 -475
rect 10800 -567 10960 -509
rect 10800 -601 10809 -567
rect 10809 -601 10960 -567
rect 10800 -659 10960 -601
rect 10800 -693 10809 -659
rect 10809 -693 10960 -659
rect 10800 -740 10960 -693
rect 10552 -793 10604 -775
rect 10552 -827 10570 -793
rect 10570 -827 10604 -793
rect 11210 -870 11290 -790
rect 10490 -1240 10540 -1130
rect 10540 -1240 10580 -1130
rect 10580 -1240 10630 -1130
rect 11390 -1170 11470 -1090
rect 6820 -4240 6880 -3020
rect 5190 -6030 5300 -5640
rect 5420 -6030 5530 -5640
rect 5850 -6364 5859 -4388
rect 5859 -6364 5893 -4388
rect 5893 -6364 5902 -4388
rect 5968 -6364 5977 -4388
rect 5977 -6364 6011 -4388
rect 6011 -6364 6020 -4388
rect 6086 -6364 6095 -4388
rect 6095 -6364 6129 -4388
rect 6129 -6364 6138 -4388
rect 6204 -6364 6213 -4388
rect 6213 -6364 6247 -4388
rect 6247 -6364 6256 -4388
rect 6322 -6364 6331 -4388
rect 6331 -6364 6365 -4388
rect 6365 -6364 6374 -4388
rect 6440 -6364 6449 -4388
rect 6449 -6364 6483 -4388
rect 6483 -6364 6492 -4388
rect 6558 -6364 6567 -4388
rect 6567 -6364 6601 -4388
rect 6601 -6364 6610 -4388
rect 7058 -5248 7067 -3272
rect 7067 -5248 7101 -3272
rect 7101 -5248 7110 -3272
rect 7516 -5248 7525 -3272
rect 7525 -5248 7559 -3272
rect 7559 -5248 7568 -3272
rect 7974 -5248 7983 -3272
rect 7983 -5248 8017 -3272
rect 8017 -5248 8026 -3272
rect 8432 -5248 8441 -3272
rect 8441 -5248 8475 -3272
rect 8475 -5248 8484 -3272
rect 8890 -5248 8899 -3272
rect 8899 -5248 8933 -3272
rect 8933 -5248 8942 -3272
rect 9120 -4240 9180 -3020
rect 10402 -3860 10542 -2940
rect 10542 -3860 10602 -2940
rect 10983 -3139 11412 -3130
rect 10983 -3192 11412 -3139
rect 10983 -3200 11412 -3192
rect 10867 -3772 11336 -3763
rect 10867 -3806 11336 -3772
rect 10867 -3815 11336 -3806
rect 8880 -5362 8944 -5298
rect 7295 -5616 7361 -5600
rect 7295 -5650 7311 -5616
rect 7311 -5650 7345 -5616
rect 7345 -5650 7361 -5616
rect 7295 -5656 7361 -5650
rect 7487 -5616 7553 -5600
rect 7487 -5650 7503 -5616
rect 7503 -5650 7537 -5616
rect 7537 -5650 7553 -5616
rect 7487 -5656 7553 -5650
rect 7679 -5616 7745 -5600
rect 7679 -5650 7695 -5616
rect 7695 -5650 7729 -5616
rect 7729 -5650 7745 -5616
rect 7679 -5656 7745 -5650
rect 7871 -5616 7937 -5600
rect 7871 -5650 7887 -5616
rect 7887 -5650 7921 -5616
rect 7921 -5650 7937 -5616
rect 7871 -5656 7937 -5650
rect 8063 -5616 8129 -5600
rect 8063 -5650 8079 -5616
rect 8079 -5650 8113 -5616
rect 8113 -5650 8129 -5616
rect 8063 -5656 8129 -5650
rect 8255 -5616 8321 -5600
rect 8255 -5650 8271 -5616
rect 8271 -5650 8305 -5616
rect 8305 -5650 8321 -5616
rect 8255 -5656 8321 -5650
rect 8447 -5616 8513 -5600
rect 8447 -5650 8463 -5616
rect 8463 -5650 8497 -5616
rect 8497 -5650 8513 -5616
rect 8447 -5656 8513 -5650
rect 8639 -5616 8705 -5600
rect 8639 -5650 8655 -5616
rect 8655 -5650 8689 -5616
rect 8689 -5650 8705 -5616
rect 8639 -5656 8705 -5650
rect 7013 -5712 7067 -5700
rect 7013 -6188 7023 -5712
rect 7023 -6188 7057 -5712
rect 7057 -6188 7067 -5712
rect 7013 -6200 7067 -6188
rect 7109 -5712 7163 -5700
rect 7109 -6188 7119 -5712
rect 7119 -6188 7153 -5712
rect 7153 -6188 7163 -5712
rect 7109 -6200 7163 -6188
rect 7205 -5712 7259 -5700
rect 7205 -6188 7215 -5712
rect 7215 -6188 7249 -5712
rect 7249 -6188 7259 -5712
rect 7205 -6200 7259 -6188
rect 7301 -5712 7355 -5700
rect 7301 -6188 7311 -5712
rect 7311 -6188 7345 -5712
rect 7345 -6188 7355 -5712
rect 7301 -6200 7355 -6188
rect 7397 -5712 7451 -5700
rect 7397 -6188 7407 -5712
rect 7407 -6188 7441 -5712
rect 7441 -6188 7451 -5712
rect 7397 -6200 7451 -6188
rect 7493 -5712 7547 -5700
rect 7493 -6188 7503 -5712
rect 7503 -6188 7537 -5712
rect 7537 -6188 7547 -5712
rect 7493 -6200 7547 -6188
rect 7589 -5712 7643 -5700
rect 7589 -6188 7599 -5712
rect 7599 -6188 7633 -5712
rect 7633 -6188 7643 -5712
rect 7589 -6200 7643 -6188
rect 7685 -5712 7739 -5700
rect 7685 -6188 7695 -5712
rect 7695 -6188 7729 -5712
rect 7729 -6188 7739 -5712
rect 7685 -6200 7739 -6188
rect 7781 -5712 7835 -5700
rect 7781 -6188 7791 -5712
rect 7791 -6188 7825 -5712
rect 7825 -6188 7835 -5712
rect 7781 -6200 7835 -6188
rect 7877 -5712 7931 -5700
rect 7877 -6188 7887 -5712
rect 7887 -6188 7921 -5712
rect 7921 -6188 7931 -5712
rect 7877 -6200 7931 -6188
rect 7973 -5712 8027 -5700
rect 7973 -6188 7983 -5712
rect 7983 -6188 8017 -5712
rect 8017 -6188 8027 -5712
rect 7973 -6200 8027 -6188
rect 8069 -5712 8123 -5700
rect 8069 -6188 8079 -5712
rect 8079 -6188 8113 -5712
rect 8113 -6188 8123 -5712
rect 8069 -6200 8123 -6188
rect 8165 -5712 8219 -5700
rect 8165 -6188 8175 -5712
rect 8175 -6188 8209 -5712
rect 8209 -6188 8219 -5712
rect 8165 -6200 8219 -6188
rect 8261 -5712 8315 -5700
rect 8261 -6188 8271 -5712
rect 8271 -6188 8305 -5712
rect 8305 -6188 8315 -5712
rect 8261 -6200 8315 -6188
rect 8357 -5712 8411 -5700
rect 8357 -6188 8367 -5712
rect 8367 -6188 8401 -5712
rect 8401 -6188 8411 -5712
rect 8357 -6200 8411 -6188
rect 8453 -5712 8507 -5700
rect 8453 -6188 8463 -5712
rect 8463 -6188 8497 -5712
rect 8497 -6188 8507 -5712
rect 8453 -6200 8507 -6188
rect 8549 -5712 8603 -5700
rect 8549 -6188 8559 -5712
rect 8559 -6188 8593 -5712
rect 8593 -6188 8603 -5712
rect 8549 -6200 8603 -6188
rect 8645 -5712 8699 -5700
rect 8645 -6188 8655 -5712
rect 8655 -6188 8689 -5712
rect 8689 -6188 8699 -5712
rect 8645 -6200 8699 -6188
rect 8741 -5712 8795 -5700
rect 8741 -6188 8751 -5712
rect 8751 -6188 8785 -5712
rect 8785 -6188 8795 -5712
rect 8741 -6200 8795 -6188
rect 8837 -5712 8891 -5700
rect 8837 -6188 8847 -5712
rect 8847 -6188 8881 -5712
rect 8881 -6188 8891 -5712
rect 8837 -6200 8891 -6188
rect 8933 -5712 8987 -5700
rect 8933 -6188 8943 -5712
rect 8943 -6188 8977 -5712
rect 8977 -6188 8987 -5712
rect 8933 -6200 8987 -6188
rect 9391 -6364 9400 -4388
rect 9400 -6364 9434 -4388
rect 9434 -6364 9443 -4388
rect 9509 -6364 9518 -4388
rect 9518 -6364 9552 -4388
rect 9552 -6364 9561 -4388
rect 9627 -6364 9636 -4388
rect 9636 -6364 9670 -4388
rect 9670 -6364 9679 -4388
rect 9745 -6364 9754 -4388
rect 9754 -6364 9788 -4388
rect 9788 -6364 9797 -4388
rect 9863 -6364 9872 -4388
rect 9872 -6364 9906 -4388
rect 9906 -6364 9915 -4388
rect 9981 -6364 9990 -4388
rect 9990 -6364 10024 -4388
rect 10024 -6364 10033 -4388
rect 10099 -6364 10108 -4388
rect 10108 -6364 10142 -4388
rect 10142 -6364 10151 -4388
rect 6204 -6558 6256 -6506
rect 9745 -6558 9797 -6506
rect 7917 -6800 7969 -6748
rect 8032 -6804 8084 -6792
rect 8032 -6838 8042 -6804
rect 8042 -6838 8076 -6804
rect 8076 -6838 8084 -6804
rect 8032 -6844 8084 -6838
rect 6086 -8873 6095 -6897
rect 6095 -8873 6129 -6897
rect 6129 -8873 6138 -6897
rect 6204 -8873 6213 -6897
rect 6213 -8873 6247 -6897
rect 6247 -8873 6256 -6897
rect 6322 -8873 6331 -6897
rect 6331 -8873 6365 -6897
rect 6365 -8873 6374 -6897
rect 6440 -8873 6449 -6897
rect 6449 -8873 6483 -6897
rect 6483 -8873 6492 -6897
rect 6558 -8873 6567 -6897
rect 6567 -8873 6601 -6897
rect 6601 -8873 6610 -6897
rect 6676 -8873 6685 -6897
rect 6685 -8873 6719 -6897
rect 6719 -8873 6728 -6897
rect 6794 -8873 6803 -6897
rect 6803 -8873 6837 -6897
rect 6837 -8873 6846 -6897
rect 6912 -8873 6921 -6897
rect 6921 -8873 6955 -6897
rect 6955 -8873 6964 -6897
rect 7030 -8873 7039 -6897
rect 7039 -8873 7073 -6897
rect 7073 -8873 7082 -6897
rect 7148 -8873 7157 -6897
rect 7157 -8873 7191 -6897
rect 7191 -8873 7200 -6897
rect 7266 -8873 7275 -6897
rect 7275 -8873 7309 -6897
rect 7309 -8873 7318 -6897
rect 7384 -8873 7393 -6897
rect 7393 -8873 7427 -6897
rect 7427 -8873 7436 -6897
rect 7502 -8873 7511 -6897
rect 7511 -8873 7545 -6897
rect 7545 -8873 7554 -6897
rect 7620 -8873 7629 -6897
rect 7629 -8873 7663 -6897
rect 7663 -8873 7672 -6897
rect 7738 -8873 7747 -6897
rect 7747 -8873 7781 -6897
rect 7781 -8873 7790 -6897
rect 7856 -8873 7865 -6897
rect 7865 -8873 7899 -6897
rect 7899 -8873 7908 -6897
rect 7974 -8873 7983 -6897
rect 7983 -8873 8017 -6897
rect 8017 -8873 8026 -6897
rect 8092 -8873 8101 -6897
rect 8101 -8873 8135 -6897
rect 8135 -8873 8144 -6897
rect 8210 -8873 8219 -6897
rect 8219 -8873 8253 -6897
rect 8253 -8873 8262 -6897
rect 8328 -8873 8337 -6897
rect 8337 -8873 8371 -6897
rect 8371 -8873 8380 -6897
rect 8446 -8873 8455 -6897
rect 8455 -8873 8489 -6897
rect 8489 -8873 8498 -6897
rect 8564 -8873 8573 -6897
rect 8573 -8873 8607 -6897
rect 8607 -8873 8616 -6897
rect 8682 -8873 8691 -6897
rect 8691 -8873 8725 -6897
rect 8725 -8873 8734 -6897
rect 8800 -8873 8809 -6897
rect 8809 -8873 8843 -6897
rect 8843 -8873 8852 -6897
rect 8918 -8873 8927 -6897
rect 8927 -8873 8961 -6897
rect 8961 -8873 8970 -6897
rect 9036 -8873 9045 -6897
rect 9045 -8873 9079 -6897
rect 9079 -8873 9088 -6897
rect 9154 -8873 9163 -6897
rect 9163 -8873 9197 -6897
rect 9197 -8873 9206 -6897
rect 9272 -8873 9281 -6897
rect 9281 -8873 9315 -6897
rect 9315 -8873 9324 -6897
rect 9390 -8873 9399 -6897
rect 9399 -8873 9433 -6897
rect 9433 -8873 9442 -6897
rect 9508 -8873 9517 -6897
rect 9517 -8873 9551 -6897
rect 9551 -8873 9560 -6897
rect 9626 -8873 9635 -6897
rect 9635 -8873 9669 -6897
rect 9669 -8873 9678 -6897
rect 9744 -8873 9753 -6897
rect 9753 -8873 9787 -6897
rect 9787 -8873 9796 -6897
rect 9862 -8873 9871 -6897
rect 9871 -8873 9905 -6897
rect 9905 -8873 9914 -6897
<< metal2 >>
rect 6402 13200 9802 13300
rect 6402 12800 6502 13200
rect 6108 12700 6502 12800
rect 9702 12800 9802 13200
rect 9702 12700 9892 12800
rect 6108 12600 9892 12700
rect 6108 12536 6208 12600
rect 6600 12536 6700 12600
rect 7000 12536 7100 12600
rect 7400 12536 7500 12600
rect 7800 12536 7900 12600
rect 8100 12536 8200 12600
rect 8500 12536 8600 12600
rect 8900 12536 9000 12600
rect 9300 12536 9400 12600
rect 9792 12536 9892 12600
rect 6086 12434 9914 12536
rect 6086 12273 6138 12434
rect 6086 10285 6138 10297
rect 6204 12273 6256 12285
rect 6322 12273 6374 12434
rect 6256 10297 6257 10365
rect 6204 10188 6257 10297
rect 6322 10285 6374 10297
rect 6440 12273 6492 12285
rect 6558 12273 6610 12434
rect 6492 10297 6493 10365
rect 6440 10285 6493 10297
rect 6558 10285 6610 10297
rect 6676 12273 6728 12285
rect 6794 12273 6846 12434
rect 6728 10297 6729 10365
rect 6676 10285 6729 10297
rect 6794 10285 6846 10297
rect 6912 12273 6964 12285
rect 7030 12273 7082 12434
rect 6964 10297 6965 10365
rect 6912 10285 6965 10297
rect 7030 10285 7082 10297
rect 7148 12273 7200 12285
rect 7266 12273 7318 12434
rect 7200 10297 7201 10365
rect 7148 10285 7201 10297
rect 7266 10285 7318 10297
rect 7384 12273 7436 12285
rect 6441 10188 6493 10285
rect 6677 10188 6729 10285
rect 6913 10188 6965 10285
rect 6000 10140 6130 10150
rect 6000 10050 6010 10140
rect 6120 10066 6130 10140
rect 6204 10136 6965 10188
rect 7149 10189 7201 10285
rect 7384 10190 7436 10297
rect 7502 12273 7554 12434
rect 7502 10285 7554 10297
rect 7620 12273 7672 12285
rect 7620 10285 7672 10297
rect 7738 12273 7790 12434
rect 7738 10285 7790 10297
rect 7856 12273 7908 12285
rect 7856 10256 7908 10297
rect 7974 12273 8026 12434
rect 7974 10284 8026 10297
rect 8092 12273 8144 12285
rect 8092 10278 8144 10297
rect 8210 12273 8262 12434
rect 8210 10285 8262 10297
rect 8328 12273 8380 12285
rect 8328 10285 8380 10297
rect 8446 12273 8498 12434
rect 8446 10285 8498 10297
rect 8564 12273 8616 12285
rect 7854 10250 8060 10256
rect 7854 10244 8084 10250
rect 7854 10228 8032 10244
rect 7384 10189 7620 10190
rect 7149 10188 7620 10189
rect 7854 10188 7883 10228
rect 7149 10138 7883 10188
rect 7149 10137 7436 10138
rect 6441 10066 6493 10136
rect 6120 10050 6493 10066
rect 6000 10014 6493 10050
rect 5850 9764 5902 9776
rect 5170 9430 5320 9450
rect 5170 9040 5190 9430
rect 5300 9040 5320 9430
rect 5170 9020 5320 9040
rect 5400 9430 5550 9450
rect 5400 9040 5420 9430
rect 5530 9040 5550 9430
rect 5400 9020 5550 9040
rect 5850 7636 5902 7788
rect 5968 9764 6020 9776
rect 5968 7636 6020 7788
rect 6086 9764 6138 10014
rect 6200 9960 6261 9969
rect 6200 9904 6202 9960
rect 6258 9904 6261 9960
rect 6200 9895 6261 9904
rect 6086 7776 6138 7788
rect 6204 9764 6256 9776
rect 6204 7636 6256 7788
rect 6322 9764 6374 10014
rect 7384 9810 7436 10137
rect 7620 10136 7883 10138
rect 7911 10148 7917 10200
rect 7969 10158 7975 10200
rect 8032 10186 8084 10192
rect 8112 10188 8144 10278
rect 8564 10188 8616 10297
rect 8682 12273 8734 12434
rect 8682 10285 8734 10297
rect 8800 12273 8852 12285
rect 8800 10188 8852 10297
rect 8918 12273 8970 12434
rect 8918 10285 8970 10297
rect 9036 12273 9088 12285
rect 8112 10158 8852 10188
rect 7969 10148 8852 10158
rect 7911 10136 8852 10148
rect 9036 10188 9088 10297
rect 9154 12273 9206 12434
rect 9154 10285 9206 10297
rect 9272 12273 9324 12285
rect 9272 10188 9324 10297
rect 9390 12273 9442 12434
rect 9390 10285 9442 10297
rect 9508 12273 9560 12285
rect 9508 10188 9560 10297
rect 9626 12273 9678 12434
rect 9626 10285 9678 10297
rect 9744 12273 9796 12285
rect 9744 10188 9796 10297
rect 9862 12273 9914 12434
rect 9862 10285 9914 10297
rect 9036 10136 9796 10188
rect 7911 10130 8144 10136
rect 8564 9810 8616 10136
rect 9508 10066 9560 10136
rect 9508 10014 9915 10066
rect 9627 9969 9679 10014
rect 9863 9969 9915 10014
rect 9627 9960 9915 9969
rect 9627 9904 9743 9960
rect 9799 9904 9915 9960
rect 9627 9895 9915 9904
rect 6322 7776 6374 7788
rect 6440 9764 6492 9776
rect 6440 7660 6492 7788
rect 6558 9764 6610 9776
rect 7295 9670 7937 9810
rect 7295 9600 7361 9670
rect 7487 9600 7553 9670
rect 7679 9600 7745 9670
rect 7871 9600 7937 9670
rect 8063 9670 8705 9810
rect 8063 9600 8129 9670
rect 8255 9600 8321 9670
rect 8447 9600 8513 9670
rect 8639 9600 8705 9670
rect 9391 9764 9443 9776
rect 7007 9100 7013 9600
rect 7067 9100 7073 9600
rect 7103 9100 7109 9600
rect 7163 9100 7169 9600
rect 7199 9100 7205 9600
rect 7259 9100 7265 9600
rect 7295 9100 7301 9600
rect 7355 9100 7361 9600
rect 7391 9100 7397 9600
rect 7451 9100 7457 9600
rect 7487 9100 7493 9600
rect 7547 9100 7553 9600
rect 7583 9100 7589 9600
rect 7643 9100 7649 9600
rect 7679 9100 7685 9600
rect 7739 9100 7745 9600
rect 7775 9100 7781 9600
rect 7835 9100 7841 9600
rect 7871 9100 7877 9600
rect 7931 9100 7937 9600
rect 7967 9100 7973 9600
rect 8027 9100 8033 9600
rect 8063 9100 8069 9600
rect 8123 9100 8129 9600
rect 8159 9100 8165 9600
rect 8219 9100 8225 9600
rect 8255 9100 8261 9600
rect 8315 9100 8321 9600
rect 8351 9100 8357 9600
rect 8411 9100 8417 9600
rect 8447 9100 8453 9600
rect 8507 9100 8513 9600
rect 8543 9100 8549 9600
rect 8603 9100 8609 9600
rect 8639 9100 8645 9600
rect 8699 9100 8705 9600
rect 8735 9100 8741 9600
rect 8795 9100 8801 9600
rect 8831 9100 8837 9600
rect 8891 9100 8897 9600
rect 8927 9100 8933 9600
rect 8987 9100 8993 9600
rect 7205 8940 7259 9100
rect 7295 9056 7361 9062
rect 7295 8980 7361 8994
rect 7397 8940 7451 9100
rect 7487 9056 7553 9062
rect 7487 8980 7553 8994
rect 7589 8940 7643 9100
rect 7679 9056 7745 9062
rect 7679 8980 7745 8994
rect 7781 8940 7835 9100
rect 7871 9056 7937 9062
rect 7871 8980 7937 8994
rect 7973 8940 8027 9100
rect 8063 9056 8129 9062
rect 8063 8980 8129 8994
rect 8165 8940 8219 9100
rect 8255 9056 8321 9062
rect 8255 8980 8321 8994
rect 8357 8940 8411 9100
rect 8447 9056 8513 9062
rect 8447 8980 8513 8994
rect 8549 8940 8603 9100
rect 8639 9056 8705 9062
rect 8639 8980 8705 8994
rect 8741 8940 8795 9100
rect 7205 8870 8795 8940
rect 7205 8784 7259 8870
rect 7397 8784 7451 8870
rect 7589 8784 7643 8870
rect 7781 8784 7835 8870
rect 7973 8784 8027 8870
rect 8165 8784 8219 8870
rect 8357 8784 8411 8870
rect 8549 8784 8603 8870
rect 8741 8784 8795 8870
rect 7205 8692 8795 8784
rect 8880 8762 9202 8770
rect 8944 8760 9202 8762
rect 8944 8700 9032 8760
rect 9192 8700 9202 8760
rect 8944 8698 9202 8700
rect 6558 7660 6610 7788
rect 7058 8648 7110 8660
rect 6440 7640 6900 7660
rect 6440 7636 6820 7640
rect 5850 7566 6820 7636
rect 6000 7400 6100 7566
rect 6200 7400 6300 7566
rect 6400 7560 6820 7566
rect 6400 7400 6500 7560
rect 6600 7400 6700 7560
rect 5802 7300 6700 7400
rect 6800 7300 6820 7560
rect 5802 7200 6820 7300
rect 5802 6900 6700 7200
rect 6800 6900 6820 7200
rect 5802 6800 6820 6900
rect 5802 6500 6700 6800
rect 6800 6500 6820 6800
rect 5802 6420 6820 6500
rect 6880 6500 6900 7640
rect 7058 6520 7110 6672
rect 7516 8648 7568 8692
rect 7516 6660 7568 6672
rect 7974 8648 8026 8660
rect 7974 6520 8026 6672
rect 8432 8648 8484 8692
rect 8880 8690 9202 8698
rect 8432 6660 8484 6672
rect 8890 8648 8942 8660
rect 9391 7660 9443 7788
rect 9509 9764 9561 9776
rect 9509 7660 9561 7788
rect 9627 9764 9679 9895
rect 9627 7776 9679 7788
rect 9745 9764 9797 9776
rect 8890 6520 8942 6672
rect 7058 6500 8942 6520
rect 9100 7640 9561 7660
rect 9100 6500 9120 7640
rect 6880 6420 9120 6500
rect 9180 7636 9561 7640
rect 9745 7636 9797 7788
rect 9863 9764 9915 9895
rect 9863 7776 9915 7788
rect 9981 9764 10033 9776
rect 9981 7636 10033 7788
rect 10099 9764 10151 9776
rect 10099 7636 10151 7788
rect 9180 7566 10200 7636
rect 9180 7560 9600 7566
rect 9180 7400 9200 7560
rect 9300 7400 9400 7560
rect 9500 7400 9600 7560
rect 9700 7400 9800 7566
rect 9900 7400 10000 7566
rect 10100 7400 10200 7566
rect 10852 7432 11102 7451
rect 9180 7200 10242 7400
rect 9180 6900 9200 7200
rect 9300 6900 10242 7200
rect 9180 6800 10242 6900
rect 9180 6500 9200 6800
rect 9300 6500 10242 6800
rect 10382 7260 10622 7280
rect 10382 6500 10402 7260
rect 9180 6420 10402 6500
rect 5802 6340 10402 6420
rect 10602 6340 10622 7260
rect 10852 7215 10872 7432
rect 11082 7215 11102 7432
rect 10852 7163 10867 7215
rect 11336 7163 11353 7215
rect 10964 6530 10983 6600
rect 11412 6530 11435 6600
rect 11202 6352 11402 6530
rect 5802 6200 10622 6340
rect 5802 6100 7202 6200
rect 5802 5500 5902 6100
rect 7102 5500 7202 6100
rect 5802 5400 7202 5500
rect 9002 6100 10402 6200
rect 9002 5500 9102 6100
rect 10302 5500 10402 6100
rect 9002 5400 10402 5500
rect 11020 4910 11120 4920
rect 11020 4830 11030 4910
rect 11110 4830 11120 4910
rect 11020 4820 11120 4830
rect 11180 4910 11280 4920
rect 11180 4830 11190 4910
rect 11270 4830 11280 4910
rect 11180 4820 11280 4830
rect 11322 4770 11402 6352
rect 11320 4760 11420 4770
rect 11320 4680 11330 4760
rect 11410 4680 11420 4760
rect 11320 4670 11420 4680
rect 3348 4345 3468 4355
rect 3348 3975 3358 4345
rect 3458 3975 3468 4345
rect 4374 4345 4494 4355
rect 3348 3965 3468 3975
rect 3561 4332 3651 4342
rect 3561 3972 3571 4332
rect 3641 3972 3651 4332
rect 3561 3962 3651 3972
rect 4191 4332 4281 4342
rect 4191 3972 4201 4332
rect 4271 3972 4281 4332
rect 4191 3962 4281 3972
rect 4374 3975 4384 4345
rect 4484 3975 4494 4345
rect 4374 3965 4494 3975
rect 9240 4260 14440 4280
rect 2927 3906 4279 3920
rect 2927 3854 3577 3906
rect 3629 3854 4213 3906
rect 4265 3854 4279 3906
rect 2927 3840 4279 3854
rect 1920 2540 2040 2560
rect 1920 2460 1940 2540
rect 2020 2531 2387 2540
rect 2020 2479 2359 2531
rect 2411 2479 2431 2531
rect 2483 2479 2489 2531
rect 2020 2460 2387 2479
rect 1920 2440 2040 2460
rect 1920 1960 2040 1980
rect 1920 1880 1940 1960
rect 2020 1945 2367 1960
rect 2020 1893 2359 1945
rect 2411 1893 2431 1945
rect 2483 1893 2489 1945
rect 2020 1880 2367 1893
rect 1920 1860 2040 1880
rect 1880 1220 2020 1240
rect 1880 1120 1900 1220
rect 2000 1120 2020 1220
rect 1880 1100 2020 1120
rect 2240 1220 2380 1240
rect 2240 1120 2260 1220
rect 2360 1120 2380 1220
rect 2240 1040 2380 1120
rect 2240 960 2260 1040
rect 2360 960 2380 1040
rect 2240 940 2380 960
rect 2620 1220 2760 1240
rect 2620 1120 2640 1220
rect 2740 1120 2760 1220
rect 1720 920 1840 940
rect 1720 800 1740 920
rect 1820 800 1840 920
rect 1720 780 1840 800
rect 2060 920 2180 940
rect 2060 800 2080 920
rect 2160 800 2180 920
rect 2060 780 2180 800
rect 2620 860 2760 1120
rect 2927 1060 3007 3840
rect 3348 3621 3468 3631
rect 3348 3251 3358 3621
rect 3458 3251 3468 3621
rect 3561 3614 3691 3624
rect 3561 3264 3571 3614
rect 3681 3264 3691 3614
rect 3561 3254 3691 3264
rect 4151 3614 4281 3624
rect 4151 3264 4161 3614
rect 4271 3264 4281 3614
rect 4151 3254 4281 3264
rect 4374 3621 4494 3631
rect 3348 3241 3468 3251
rect 4374 3251 4384 3621
rect 4484 3251 4494 3621
rect 4374 3241 4494 3251
rect 2887 1040 3007 1060
rect 2887 960 2907 1040
rect 2987 960 3007 1040
rect 2887 940 3007 960
rect 2620 780 2640 860
rect 2740 780 2760 860
rect 2620 760 2760 780
rect 2927 -580 3007 940
rect 3067 3192 4279 3206
rect 3067 3140 3577 3192
rect 3629 3140 4213 3192
rect 4265 3140 4279 3192
rect 3067 3126 4279 3140
rect 3067 880 3147 3126
rect 9240 2960 9260 4260
rect 14420 3998 14440 4260
rect 14420 3978 14448 3998
rect 9460 3908 11278 3960
rect 14428 3908 14448 3978
rect 9460 3888 14448 3908
rect 9460 3880 10460 3888
rect 9460 2960 9480 3880
rect 9240 2940 9480 2960
rect 11365 3725 11417 3737
rect 5427 2920 5887 2940
rect 5427 2840 5447 2920
rect 5867 2840 5887 2920
rect 5427 2820 5887 2840
rect 6627 2920 7087 2940
rect 6627 2840 6647 2920
rect 7067 2840 7087 2920
rect 6627 2820 7087 2840
rect 7827 2920 8287 2940
rect 7827 2840 7847 2920
rect 8267 2840 8287 2920
rect 7827 2820 8287 2840
rect 9027 2920 9487 2940
rect 9027 2840 9047 2920
rect 9467 2840 9487 2920
rect 9027 2820 9487 2840
rect 3240 2608 3640 2618
rect 3240 2600 3250 2608
rect 3240 2380 3247 2600
rect 3240 2368 3250 2380
rect 3630 2368 3640 2608
rect 3240 2358 3640 2368
rect 3965 2347 4017 2358
rect 4017 2319 4066 2341
rect 4017 2295 4594 2319
rect 3965 2289 4594 2295
rect 3965 2129 4017 2135
rect 4017 2118 4066 2129
rect 4017 2088 4481 2118
rect 4017 2077 4066 2088
rect 3965 2066 4017 2077
rect 3240 2056 3640 2066
rect 3240 2040 3250 2056
rect 3240 1820 3247 2040
rect 3240 1816 3250 1820
rect 3630 1816 3640 2056
rect 3240 1806 3640 1816
rect 4063 2008 4297 2045
rect 3714 1430 3766 1432
rect 4063 1430 4100 2008
rect 4156 1886 4162 1938
rect 4214 1886 4220 1938
rect 4162 1850 4214 1886
rect 4260 1857 4297 2008
rect 4451 1961 4481 2088
rect 4564 1963 4594 2289
rect 4727 2260 5187 2280
rect 4727 2180 4747 2260
rect 5167 2180 5187 2260
rect 4727 2160 5187 2180
rect 6027 2240 6487 2260
rect 6027 2160 6047 2240
rect 6467 2160 6487 2240
rect 6027 2140 6487 2160
rect 7227 2240 7687 2260
rect 7227 2160 7247 2240
rect 7667 2160 7687 2240
rect 7227 2140 7687 2160
rect 8427 2240 8887 2260
rect 8427 2160 8447 2240
rect 8867 2160 8887 2240
rect 8427 2140 8887 2160
rect 9627 2240 10087 2260
rect 9627 2160 9647 2240
rect 10067 2160 10087 2240
rect 9627 2140 10087 2160
rect 10818 2108 10898 2118
rect 5974 1981 8240 2021
rect 4433 1909 4439 1961
rect 4491 1909 4497 1961
rect 4547 1911 4553 1963
rect 4605 1911 4611 1963
rect 4940 1898 4946 1950
rect 4998 1898 5004 1950
rect 4948 1857 4985 1898
rect 4169 1461 4210 1850
rect 4260 1820 4985 1857
rect 5974 1788 6014 1981
rect 6109 1921 6115 1935
rect 4832 1776 6014 1788
rect 4832 1724 4838 1776
rect 4890 1748 6014 1776
rect 6063 1883 6115 1921
rect 6167 1883 6173 1935
rect 8200 1903 8240 1981
rect 9256 1987 9921 2024
rect 4890 1724 4897 1748
rect 6063 1710 6101 1883
rect 8188 1851 8194 1903
rect 8246 1851 8252 1903
rect 5040 1704 6101 1710
rect 5092 1672 6101 1704
rect 8878 1832 8930 1838
rect 8930 1823 8947 1832
rect 9256 1823 9293 1987
rect 9884 1935 9921 1987
rect 9474 1883 9480 1935
rect 9532 1883 9552 1935
rect 9604 1883 9610 1935
rect 9861 1883 9867 1935
rect 9919 1883 9939 1935
rect 9991 1883 9997 1935
rect 10180 1930 10280 1950
rect 8930 1786 9293 1823
rect 8930 1780 8947 1786
rect 8878 1760 8930 1780
rect 8878 1702 8930 1708
rect 5040 1646 5092 1652
rect 5427 1600 5887 1620
rect 5427 1520 5447 1600
rect 5867 1520 5887 1600
rect 5427 1500 5887 1520
rect 6627 1600 7087 1620
rect 6627 1520 6647 1600
rect 7067 1520 7087 1600
rect 6627 1500 7087 1520
rect 7827 1600 8287 1620
rect 7827 1520 7847 1600
rect 8267 1520 8287 1600
rect 7827 1500 8287 1520
rect 9027 1600 9487 1620
rect 9027 1520 9047 1600
rect 9467 1520 9487 1600
rect 9027 1500 9487 1520
rect 3714 1378 4107 1430
rect 4169 1420 8577 1461
rect 3227 1220 3347 1240
rect 3227 1140 3247 1220
rect 3327 1199 3567 1220
rect 3714 1199 3766 1378
rect 3327 1147 3511 1199
rect 3563 1147 3583 1199
rect 3635 1147 3766 1199
rect 4387 1280 4807 1300
rect 4387 1276 4407 1280
rect 3327 1140 3567 1147
rect 3227 1120 3347 1140
rect 4387 1036 4402 1276
rect 4787 1040 4807 1280
rect 5709 1231 5750 1420
rect 8472 1379 8577 1420
rect 8524 1327 8577 1379
rect 8472 1307 8577 1327
rect 8524 1296 8577 1307
rect 8881 1375 8933 1381
rect 8881 1303 8933 1323
rect 9537 1303 9570 1883
rect 8524 1255 8801 1296
rect 8472 1249 8524 1255
rect 5697 1179 5703 1231
rect 5755 1179 5761 1231
rect 6113 1205 6119 1209
rect 4782 1036 4807 1040
rect 4387 1020 4807 1036
rect 5991 1157 6119 1205
rect 6171 1157 6177 1209
rect 8190 1190 8196 1242
rect 8248 1190 8254 1242
rect 5117 1015 5169 1026
rect 5991 1011 6039 1157
rect 8190 1154 8254 1190
rect 8756 1207 8797 1255
rect 8933 1270 9570 1303
rect 8933 1251 8966 1270
rect 8881 1245 8933 1251
rect 9412 1230 9518 1236
rect 9412 1207 9460 1230
rect 8756 1178 9460 1207
rect 9512 1178 9518 1230
rect 9907 1223 9940 1883
rect 10180 1850 10200 1930
rect 10260 1850 10280 1930
rect 10180 1830 10280 1850
rect 10818 1678 10828 2108
rect 10888 1678 10898 2108
rect 10818 1668 10898 1678
rect 10988 2108 11068 2118
rect 10988 1678 10998 2108
rect 11058 1678 11068 2108
rect 11365 1737 11417 1749
rect 11823 3725 11875 3737
rect 11823 1737 11875 1749
rect 12281 3725 12333 3737
rect 12281 1737 12333 1749
rect 12739 3725 12791 3737
rect 13197 3725 13249 3737
rect 13188 1768 13197 1958
rect 13978 2328 14068 2338
rect 13978 2118 13988 2328
rect 14048 2118 14068 2328
rect 13978 2108 14068 2118
rect 13848 2098 13928 2108
rect 13848 1958 13858 2098
rect 13249 1948 13858 1958
rect 13258 1888 13858 1948
rect 13918 1888 13928 2098
rect 13258 1878 13928 1888
rect 13258 1778 13268 1878
rect 12739 1737 12791 1749
rect 13249 1768 13268 1778
rect 13197 1737 13249 1749
rect 10988 1668 11068 1678
rect 12810 1690 13180 1700
rect 10838 1438 10878 1668
rect 11008 1538 11048 1668
rect 12098 1638 12218 1648
rect 12098 1578 12108 1638
rect 12208 1608 12218 1638
rect 12810 1610 12820 1690
rect 13170 1610 13180 1690
rect 12208 1578 12288 1608
rect 12810 1600 13180 1610
rect 12098 1568 12288 1578
rect 12248 1538 12288 1568
rect 13828 1598 13878 1878
rect 13908 1698 13988 1708
rect 13908 1638 13918 1698
rect 13978 1638 13988 1698
rect 13908 1628 13988 1638
rect 14238 1698 14318 1708
rect 14238 1638 14248 1698
rect 14308 1638 14318 1698
rect 14238 1628 14318 1638
rect 13828 1548 14128 1598
rect 11008 1498 12288 1538
rect 12810 1440 13180 1450
rect 10838 1398 12328 1438
rect 12288 1308 12328 1398
rect 12810 1360 12820 1440
rect 13170 1360 13180 1440
rect 12810 1350 13180 1360
rect 13908 1408 13988 1418
rect 13908 1348 13918 1408
rect 13978 1348 13988 1408
rect 13908 1338 13988 1348
rect 14088 1308 14128 1548
rect 14238 1408 14318 1418
rect 14238 1348 14248 1408
rect 14308 1348 14318 1408
rect 14238 1338 14318 1348
rect 10449 1296 10501 1308
rect 8756 1170 9518 1178
rect 9579 1171 9585 1223
rect 9637 1171 9940 1223
rect 10180 1240 10280 1260
rect 8756 1166 9412 1170
rect 10180 1160 10200 1240
rect 10260 1160 10280 1240
rect 10180 1140 10280 1160
rect 5169 963 6039 1011
rect 5117 957 5169 963
rect 6027 900 6487 920
rect 3067 860 3187 880
rect 3067 780 3087 860
rect 3167 780 3187 860
rect 6027 820 6047 900
rect 6467 820 6487 900
rect 6027 800 6487 820
rect 7227 900 7687 920
rect 7227 820 7247 900
rect 7667 820 7687 900
rect 7227 800 7687 820
rect 8427 900 8887 920
rect 8427 820 8447 900
rect 8867 820 8887 900
rect 8427 800 8887 820
rect 9627 900 10087 920
rect 9627 820 9647 900
rect 10067 820 10087 900
rect 9627 800 10087 820
rect 3067 760 3187 780
rect 3067 140 3147 760
rect 3941 575 4061 585
rect 3758 562 3848 572
rect 3758 202 3768 562
rect 3838 202 3848 562
rect 3758 192 3848 202
rect 3941 205 3951 575
rect 4051 205 4061 575
rect 3941 195 4061 205
rect 3766 145 3846 150
rect 3761 140 3846 145
rect 3067 136 3846 140
rect 3067 84 3780 136
rect 3832 84 3846 136
rect 3067 70 3846 84
rect 9880 120 10080 800
rect 10449 308 10501 320
rect 10907 1296 10959 1308
rect 11365 1296 11417 1308
rect 11070 920 11365 940
rect 11070 840 11090 920
rect 11190 840 11365 920
rect 11070 820 11365 840
rect 10907 308 10959 320
rect 11365 308 11417 320
rect 11823 1296 11875 1308
rect 12281 1296 12333 1308
rect 12268 1268 12281 1278
rect 12739 1296 12791 1308
rect 12333 1268 12348 1278
rect 12268 1168 12278 1268
rect 12338 1168 12348 1268
rect 12268 1158 12281 1168
rect 11823 308 11875 320
rect 12333 1158 12348 1168
rect 12281 308 12333 320
rect 13197 1296 13249 1308
rect 13188 1088 13197 1278
rect 14088 1298 14238 1308
rect 13249 1268 13268 1278
rect 14088 1268 14168 1298
rect 13258 1168 13268 1268
rect 14158 1238 14168 1268
rect 14228 1238 14238 1298
rect 14158 1228 14238 1238
rect 13258 1158 13928 1168
rect 13258 1098 13858 1158
rect 12739 308 12791 320
rect 13249 1088 13858 1098
rect 13848 948 13858 1088
rect 13918 948 13928 1158
rect 39900 1040 40320 1050
rect 39370 1030 39390 1040
rect 37681 1012 38071 1022
rect 13848 938 13928 948
rect 15547 1002 15927 1012
rect 13978 928 14068 938
rect 13978 718 13988 928
rect 14058 718 14068 928
rect 15547 912 15557 1002
rect 15917 912 15927 1002
rect 15547 902 15927 912
rect 16261 1002 16641 1012
rect 16261 912 16271 1002
rect 16631 912 16641 1002
rect 16261 902 16641 912
rect 16975 1002 17355 1012
rect 16975 912 16985 1002
rect 17345 912 17355 1002
rect 16975 902 17355 912
rect 17689 1002 18069 1012
rect 17689 912 17699 1002
rect 18059 912 18069 1002
rect 17689 902 18069 912
rect 18403 1002 18783 1012
rect 18403 912 18413 1002
rect 18773 912 18783 1002
rect 18403 902 18783 912
rect 19117 1002 19497 1012
rect 19117 912 19127 1002
rect 19487 912 19497 1002
rect 19117 902 19497 912
rect 19831 1002 20211 1012
rect 19831 912 19841 1002
rect 20201 912 20211 1002
rect 19831 902 20211 912
rect 20545 1002 20925 1012
rect 20545 912 20555 1002
rect 20915 912 20925 1002
rect 20545 902 20925 912
rect 21259 1002 21639 1012
rect 21259 912 21269 1002
rect 21629 912 21639 1002
rect 21259 902 21639 912
rect 21973 1002 22353 1012
rect 21973 912 21983 1002
rect 22343 912 22353 1002
rect 21973 902 22353 912
rect 22687 1002 23067 1012
rect 22687 912 22697 1002
rect 23057 912 23067 1002
rect 22687 902 23067 912
rect 23401 1002 23781 1012
rect 23401 912 23411 1002
rect 23771 912 23781 1002
rect 23401 902 23781 912
rect 24115 1002 24495 1012
rect 24115 912 24125 1002
rect 24485 912 24495 1002
rect 24115 902 24495 912
rect 24829 1002 25209 1012
rect 24829 912 24839 1002
rect 25199 912 25209 1002
rect 24829 902 25209 912
rect 25543 1002 25923 1012
rect 25543 912 25553 1002
rect 25913 912 25923 1002
rect 25543 902 25923 912
rect 26257 1002 26637 1012
rect 26257 912 26267 1002
rect 26627 912 26637 1002
rect 26257 902 26637 912
rect 26971 1002 27351 1012
rect 26971 912 26981 1002
rect 27341 912 27351 1002
rect 26971 902 27351 912
rect 27685 1002 28065 1012
rect 27685 912 27695 1002
rect 28055 912 28065 1002
rect 27685 902 28065 912
rect 28399 1002 28779 1012
rect 28399 912 28409 1002
rect 28769 912 28779 1002
rect 28399 902 28779 912
rect 29113 1002 29493 1012
rect 29113 912 29123 1002
rect 29483 912 29493 1002
rect 29113 902 29493 912
rect 29827 1002 30207 1012
rect 29827 912 29837 1002
rect 30197 912 30207 1002
rect 29827 902 30207 912
rect 30541 1002 30921 1012
rect 30541 912 30551 1002
rect 30911 912 30921 1002
rect 30541 902 30921 912
rect 31255 1002 31635 1012
rect 31255 912 31265 1002
rect 31625 912 31635 1002
rect 31255 902 31635 912
rect 31969 1002 32349 1012
rect 31969 912 31979 1002
rect 32339 912 32349 1002
rect 31969 902 32349 912
rect 32683 1002 33063 1012
rect 32683 912 32693 1002
rect 33053 912 33063 1002
rect 32683 902 33063 912
rect 33397 1002 33777 1012
rect 33397 912 33407 1002
rect 33767 912 33777 1002
rect 33397 902 33777 912
rect 34111 1002 34491 1012
rect 34111 912 34121 1002
rect 34481 912 34491 1002
rect 34111 902 34491 912
rect 34825 1002 35205 1012
rect 34825 912 34835 1002
rect 35195 912 35205 1002
rect 34825 902 35205 912
rect 35539 1002 35919 1012
rect 35539 912 35549 1002
rect 35909 912 35919 1002
rect 35539 902 35919 912
rect 36253 1002 36633 1012
rect 36253 912 36263 1002
rect 36623 912 36633 1002
rect 36253 902 36633 912
rect 36967 1002 37347 1012
rect 36967 912 36977 1002
rect 37337 912 37347 1002
rect 36967 902 37347 912
rect 37681 912 37691 1012
rect 38061 912 38071 1012
rect 37681 902 38071 912
rect 38385 1012 38775 1022
rect 38385 912 38395 1012
rect 38765 912 38775 1012
rect 38385 902 38775 912
rect 39140 990 39390 1030
rect 15548 803 15928 813
rect 15548 733 15558 803
rect 15918 733 15928 803
rect 15548 723 15928 733
rect 15972 793 16052 807
rect 15972 741 15986 793
rect 16038 741 16052 793
rect 15972 727 16052 741
rect 16262 803 16642 813
rect 16262 733 16272 803
rect 16632 733 16642 803
rect 15977 722 16047 727
rect 16262 723 16642 733
rect 16686 793 16766 807
rect 16686 741 16700 793
rect 16752 741 16766 793
rect 16686 727 16766 741
rect 16976 803 17356 813
rect 16976 733 16986 803
rect 17346 733 17356 803
rect 16691 722 16761 727
rect 16976 723 17356 733
rect 17400 793 17480 807
rect 17400 741 17414 793
rect 17466 741 17480 793
rect 17400 727 17480 741
rect 17690 803 18070 813
rect 17690 733 17700 803
rect 18060 733 18070 803
rect 17405 722 17475 727
rect 17690 723 18070 733
rect 18114 793 18194 807
rect 18114 741 18128 793
rect 18180 741 18194 793
rect 18114 727 18194 741
rect 18404 803 18784 813
rect 18404 733 18414 803
rect 18774 733 18784 803
rect 18119 722 18189 727
rect 18404 723 18784 733
rect 18828 793 18908 807
rect 18828 741 18842 793
rect 18894 741 18908 793
rect 18828 727 18908 741
rect 19118 803 19498 813
rect 19118 733 19128 803
rect 19488 733 19498 803
rect 18833 722 18903 727
rect 19118 723 19498 733
rect 19542 793 19622 807
rect 19542 741 19556 793
rect 19608 741 19622 793
rect 19542 727 19622 741
rect 19832 803 20212 813
rect 19832 733 19842 803
rect 20202 733 20212 803
rect 19547 722 19617 727
rect 19832 723 20212 733
rect 20256 793 20336 807
rect 20256 741 20270 793
rect 20322 741 20336 793
rect 20256 727 20336 741
rect 20546 803 20926 813
rect 20546 733 20556 803
rect 20916 733 20926 803
rect 20261 722 20331 727
rect 20546 723 20926 733
rect 20970 793 21050 807
rect 20970 741 20984 793
rect 21036 741 21050 793
rect 20970 727 21050 741
rect 21260 803 21640 813
rect 21260 733 21270 803
rect 21630 733 21640 803
rect 20975 722 21045 727
rect 21260 723 21640 733
rect 21684 793 21764 807
rect 21684 741 21698 793
rect 21750 741 21764 793
rect 21684 727 21764 741
rect 21974 803 22354 813
rect 21974 733 21984 803
rect 22344 733 22354 803
rect 21689 722 21759 727
rect 21974 723 22354 733
rect 22398 793 22478 807
rect 22398 741 22412 793
rect 22464 741 22478 793
rect 22398 727 22478 741
rect 22688 803 23068 813
rect 22688 733 22698 803
rect 23058 733 23068 803
rect 22403 722 22473 727
rect 22688 723 23068 733
rect 23112 793 23192 807
rect 23112 741 23126 793
rect 23178 741 23192 793
rect 23112 727 23192 741
rect 23402 803 23782 813
rect 23402 733 23412 803
rect 23772 733 23782 803
rect 23117 722 23187 727
rect 23402 723 23782 733
rect 23826 793 23906 807
rect 23826 741 23840 793
rect 23892 741 23906 793
rect 23826 727 23906 741
rect 24116 803 24496 813
rect 24116 733 24126 803
rect 24486 733 24496 803
rect 23831 722 23901 727
rect 24116 723 24496 733
rect 24540 793 24620 807
rect 24540 741 24554 793
rect 24606 741 24620 793
rect 24540 727 24620 741
rect 24830 803 25210 813
rect 24830 733 24840 803
rect 25200 733 25210 803
rect 24545 722 24615 727
rect 24830 723 25210 733
rect 25254 793 25334 807
rect 25254 741 25268 793
rect 25320 741 25334 793
rect 25254 727 25334 741
rect 25544 803 25924 813
rect 25544 733 25554 803
rect 25914 733 25924 803
rect 25259 722 25329 727
rect 25544 723 25924 733
rect 25968 793 26048 807
rect 25968 741 25982 793
rect 26034 741 26048 793
rect 25968 727 26048 741
rect 26258 803 26638 813
rect 26258 733 26268 803
rect 26628 733 26638 803
rect 25973 722 26043 727
rect 26258 723 26638 733
rect 26682 793 26762 807
rect 26682 741 26696 793
rect 26748 741 26762 793
rect 26682 727 26762 741
rect 26972 803 27352 813
rect 26972 733 26982 803
rect 27342 733 27352 803
rect 26687 722 26757 727
rect 26972 723 27352 733
rect 27396 793 27476 807
rect 27396 741 27410 793
rect 27462 741 27476 793
rect 27396 727 27476 741
rect 27686 803 28066 813
rect 27686 733 27696 803
rect 28056 733 28066 803
rect 27401 722 27471 727
rect 27686 723 28066 733
rect 28110 793 28190 807
rect 28110 741 28124 793
rect 28176 741 28190 793
rect 28110 727 28190 741
rect 28400 803 28780 813
rect 28400 733 28410 803
rect 28770 733 28780 803
rect 28115 722 28185 727
rect 28400 723 28780 733
rect 28824 793 28904 807
rect 28824 741 28838 793
rect 28890 741 28904 793
rect 28824 727 28904 741
rect 29114 803 29494 813
rect 29114 733 29124 803
rect 29484 733 29494 803
rect 28829 722 28899 727
rect 29114 723 29494 733
rect 29538 793 29618 807
rect 29538 741 29552 793
rect 29604 741 29618 793
rect 29538 727 29618 741
rect 29828 803 30208 813
rect 29828 733 29838 803
rect 30198 733 30208 803
rect 29543 722 29613 727
rect 29828 723 30208 733
rect 30252 793 30332 807
rect 30252 741 30266 793
rect 30318 741 30332 793
rect 30252 727 30332 741
rect 30542 803 30922 813
rect 30542 733 30552 803
rect 30912 733 30922 803
rect 30257 722 30327 727
rect 30542 723 30922 733
rect 30966 793 31046 807
rect 30966 741 30980 793
rect 31032 741 31046 793
rect 30966 727 31046 741
rect 31256 803 31636 813
rect 31256 733 31266 803
rect 31626 733 31636 803
rect 30971 722 31041 727
rect 31256 723 31636 733
rect 31680 793 31760 807
rect 31680 741 31694 793
rect 31746 741 31760 793
rect 31680 727 31760 741
rect 31970 803 32350 813
rect 31970 733 31980 803
rect 32340 733 32350 803
rect 31685 722 31755 727
rect 31970 723 32350 733
rect 32394 793 32474 807
rect 32394 741 32408 793
rect 32460 741 32474 793
rect 32394 727 32474 741
rect 32684 803 33064 813
rect 32684 733 32694 803
rect 33054 733 33064 803
rect 32399 722 32469 727
rect 32684 723 33064 733
rect 33108 793 33188 807
rect 33108 741 33122 793
rect 33174 741 33188 793
rect 33108 727 33188 741
rect 33398 803 33778 813
rect 33398 733 33408 803
rect 33768 733 33778 803
rect 33113 722 33183 727
rect 33398 723 33778 733
rect 33822 793 33902 807
rect 33822 741 33836 793
rect 33888 741 33902 793
rect 33822 727 33902 741
rect 34112 803 34492 813
rect 34112 733 34122 803
rect 34482 733 34492 803
rect 33827 722 33897 727
rect 34112 723 34492 733
rect 34536 793 34616 807
rect 34536 741 34550 793
rect 34602 741 34616 793
rect 34536 727 34616 741
rect 34826 803 35206 813
rect 34826 733 34836 803
rect 35196 733 35206 803
rect 34541 722 34611 727
rect 34826 723 35206 733
rect 35250 793 35330 807
rect 35250 741 35264 793
rect 35316 741 35330 793
rect 35250 727 35330 741
rect 35540 803 35920 813
rect 35540 733 35550 803
rect 35910 733 35920 803
rect 35255 722 35325 727
rect 35540 723 35920 733
rect 35964 793 36044 807
rect 35964 741 35978 793
rect 36030 741 36044 793
rect 35964 727 36044 741
rect 36254 803 36634 813
rect 36254 733 36264 803
rect 36624 733 36634 803
rect 35969 722 36039 727
rect 36254 723 36634 733
rect 36678 793 36758 807
rect 36678 741 36692 793
rect 36744 741 36758 793
rect 36678 727 36758 741
rect 36968 803 37348 813
rect 39140 809 39180 990
rect 39370 980 39390 990
rect 39770 980 39790 1040
rect 39900 980 39920 1040
rect 40300 980 40320 1040
rect 39900 970 40320 980
rect 39900 880 40320 890
rect 39370 870 39390 880
rect 36968 733 36978 803
rect 37338 733 37348 803
rect 36683 722 36753 727
rect 36968 723 37348 733
rect 37392 793 37472 807
rect 37392 741 37406 793
rect 37458 741 37472 793
rect 37392 727 37472 741
rect 37688 799 38058 809
rect 37397 722 37467 727
rect 13978 708 14068 718
rect 13197 308 13249 320
rect 15988 339 16028 722
rect 16702 339 16742 722
rect 17416 339 17456 722
rect 18130 339 18170 722
rect 18844 339 18884 722
rect 19558 339 19598 722
rect 20272 339 20312 722
rect 20986 339 21026 722
rect 21700 339 21740 722
rect 22414 339 22454 722
rect 23128 339 23168 722
rect 23842 339 23882 722
rect 24556 339 24596 722
rect 25270 339 25310 722
rect 25984 339 26024 722
rect 26698 339 26738 722
rect 27418 409 27458 722
rect 28128 409 28168 722
rect 28848 409 28888 722
rect 29558 409 29598 722
rect 30268 409 30308 722
rect 30988 409 31028 722
rect 31708 409 31748 722
rect 32418 409 32458 722
rect 33128 479 33168 722
rect 33848 479 33888 722
rect 34558 479 34598 722
rect 35268 479 35308 722
rect 35988 549 36028 722
rect 36698 549 36738 722
rect 37418 619 37458 722
rect 37688 689 37698 799
rect 38048 689 38058 799
rect 38106 793 38186 807
rect 38106 741 38120 793
rect 38172 741 38186 793
rect 38106 727 38186 741
rect 38398 799 38778 809
rect 38838 807 39180 809
rect 38398 729 38408 799
rect 38768 729 38778 799
rect 38111 722 38181 727
rect 37688 679 38058 689
rect 38118 689 38158 722
rect 38398 719 38778 729
rect 38820 793 39180 807
rect 38820 741 38834 793
rect 38886 769 39180 793
rect 39210 830 39390 870
rect 38886 741 38900 769
rect 38820 727 38900 741
rect 38825 722 38895 727
rect 39210 689 39250 830
rect 39370 820 39390 830
rect 39770 820 39790 880
rect 39900 820 39920 880
rect 40300 820 40320 880
rect 39900 810 40320 820
rect 39900 710 40320 720
rect 39370 700 39390 710
rect 38118 649 39250 689
rect 39280 660 39390 700
rect 39280 619 39320 660
rect 39370 650 39390 660
rect 39770 650 39790 710
rect 39900 650 39920 710
rect 40300 650 40320 710
rect 39900 640 40320 650
rect 37418 579 39320 619
rect 39370 549 39390 550
rect 35988 509 39390 549
rect 39370 490 39390 509
rect 39770 490 39790 550
rect 39900 540 40320 550
rect 39900 480 39920 540
rect 40300 480 40320 540
rect 33128 439 39330 479
rect 39900 470 40320 480
rect 27418 369 39260 409
rect 15988 299 39190 339
rect 15994 229 39120 269
rect 10308 158 14448 168
rect 10308 120 10358 158
rect 9880 100 10358 120
rect 3067 60 3767 70
rect 3718 -156 3848 -146
rect 3718 -506 3728 -156
rect 3838 -506 3848 -156
rect 3718 -516 3848 -506
rect 3941 -149 4061 -139
rect 3941 -519 3951 -149
rect 4051 -519 4061 -149
rect 9880 -180 9900 100
rect 14428 78 14448 158
rect 15994 140 16034 229
rect 16708 140 16748 229
rect 17422 140 17462 229
rect 18136 140 18176 229
rect 18850 140 18890 229
rect 19564 140 19604 229
rect 20278 140 20318 229
rect 20992 140 21032 229
rect 21706 140 21746 229
rect 22420 140 22460 229
rect 23134 140 23174 229
rect 23848 140 23888 229
rect 24562 140 24602 229
rect 25276 140 25316 229
rect 25990 140 26030 229
rect 26704 140 26744 229
rect 27418 140 27458 229
rect 28132 140 28172 229
rect 28846 140 28886 229
rect 29560 140 29600 229
rect 30274 140 30314 229
rect 30988 140 31028 229
rect 31702 140 31742 229
rect 32416 140 32456 229
rect 33130 140 33170 229
rect 33844 140 33884 229
rect 34558 140 34598 229
rect 35272 140 35312 229
rect 35986 140 36026 229
rect 36700 140 36740 229
rect 37414 140 37454 229
rect 38128 140 38168 229
rect 38838 140 38878 229
rect 14380 58 14448 78
rect 15548 129 15928 139
rect 15977 135 16047 140
rect 15548 59 15558 129
rect 15918 59 15928 129
rect 14380 -180 14400 58
rect 15548 49 15928 59
rect 15972 121 16052 135
rect 15972 69 15986 121
rect 16038 69 16052 121
rect 15972 55 16052 69
rect 16262 129 16642 139
rect 16691 135 16761 140
rect 16262 59 16272 129
rect 16632 59 16642 129
rect 16262 49 16642 59
rect 16686 121 16766 135
rect 16686 69 16700 121
rect 16752 69 16766 121
rect 16686 55 16766 69
rect 16976 129 17356 139
rect 17405 135 17475 140
rect 16976 59 16986 129
rect 17346 59 17356 129
rect 16976 49 17356 59
rect 17400 121 17480 135
rect 17400 69 17414 121
rect 17466 69 17480 121
rect 17400 55 17480 69
rect 17690 129 18070 139
rect 18119 135 18189 140
rect 17690 59 17700 129
rect 18060 59 18070 129
rect 17690 49 18070 59
rect 18114 121 18194 135
rect 18114 69 18128 121
rect 18180 69 18194 121
rect 18114 55 18194 69
rect 18404 129 18784 139
rect 18833 135 18903 140
rect 18404 59 18414 129
rect 18774 59 18784 129
rect 18404 49 18784 59
rect 18828 121 18908 135
rect 18828 69 18842 121
rect 18894 69 18908 121
rect 18828 55 18908 69
rect 19118 129 19498 139
rect 19547 135 19617 140
rect 19118 59 19128 129
rect 19488 59 19498 129
rect 19118 49 19498 59
rect 19542 121 19622 135
rect 19542 69 19556 121
rect 19608 69 19622 121
rect 19542 55 19622 69
rect 19832 129 20212 139
rect 20261 135 20331 140
rect 19832 59 19842 129
rect 20202 59 20212 129
rect 19832 49 20212 59
rect 20256 121 20336 135
rect 20256 69 20270 121
rect 20322 69 20336 121
rect 20256 55 20336 69
rect 20546 129 20926 139
rect 20975 135 21045 140
rect 20546 59 20556 129
rect 20916 59 20926 129
rect 20546 49 20926 59
rect 20970 121 21050 135
rect 20970 69 20984 121
rect 21036 69 21050 121
rect 20970 55 21050 69
rect 21260 129 21640 139
rect 21689 135 21759 140
rect 21260 59 21270 129
rect 21630 59 21640 129
rect 21260 49 21640 59
rect 21684 121 21764 135
rect 21684 69 21698 121
rect 21750 69 21764 121
rect 21684 55 21764 69
rect 21974 129 22354 139
rect 22403 135 22473 140
rect 21974 59 21984 129
rect 22344 59 22354 129
rect 21974 49 22354 59
rect 22398 121 22478 135
rect 22398 69 22412 121
rect 22464 69 22478 121
rect 22398 55 22478 69
rect 22688 129 23068 139
rect 23117 135 23187 140
rect 22688 59 22698 129
rect 23058 59 23068 129
rect 22688 49 23068 59
rect 23112 121 23192 135
rect 23112 69 23126 121
rect 23178 69 23192 121
rect 23112 55 23192 69
rect 23402 129 23782 139
rect 23831 135 23901 140
rect 23402 59 23412 129
rect 23772 59 23782 129
rect 23402 49 23782 59
rect 23826 121 23906 135
rect 23826 69 23840 121
rect 23892 69 23906 121
rect 23826 55 23906 69
rect 24116 129 24496 139
rect 24545 135 24615 140
rect 24116 59 24126 129
rect 24486 59 24496 129
rect 24116 49 24496 59
rect 24540 121 24620 135
rect 24540 69 24554 121
rect 24606 69 24620 121
rect 24540 55 24620 69
rect 24830 129 25210 139
rect 25259 135 25329 140
rect 24830 59 24840 129
rect 25200 59 25210 129
rect 24830 49 25210 59
rect 25254 121 25334 135
rect 25254 69 25268 121
rect 25320 69 25334 121
rect 25254 55 25334 69
rect 25544 129 25924 139
rect 25973 135 26043 140
rect 25544 59 25554 129
rect 25914 59 25924 129
rect 25544 49 25924 59
rect 25968 121 26048 135
rect 25968 69 25982 121
rect 26034 69 26048 121
rect 25968 55 26048 69
rect 26258 129 26638 139
rect 26687 135 26757 140
rect 26258 59 26268 129
rect 26628 59 26638 129
rect 26258 49 26638 59
rect 26682 121 26762 135
rect 26682 69 26696 121
rect 26748 69 26762 121
rect 26682 55 26762 69
rect 26972 129 27352 139
rect 27401 135 27471 140
rect 26972 59 26982 129
rect 27342 59 27352 129
rect 26972 49 27352 59
rect 27396 121 27476 135
rect 27396 69 27410 121
rect 27462 69 27476 121
rect 27396 55 27476 69
rect 27686 129 28066 139
rect 28115 135 28185 140
rect 27686 59 27696 129
rect 28056 59 28066 129
rect 27686 49 28066 59
rect 28110 121 28190 135
rect 28110 69 28124 121
rect 28176 69 28190 121
rect 28110 55 28190 69
rect 28400 129 28780 139
rect 28829 135 28899 140
rect 28400 59 28410 129
rect 28770 59 28780 129
rect 28400 49 28780 59
rect 28824 121 28904 135
rect 28824 69 28838 121
rect 28890 69 28904 121
rect 28824 55 28904 69
rect 29114 129 29494 139
rect 29543 135 29613 140
rect 29114 59 29124 129
rect 29484 59 29494 129
rect 29114 49 29494 59
rect 29538 121 29618 135
rect 29538 69 29552 121
rect 29604 69 29618 121
rect 29538 55 29618 69
rect 29828 129 30208 139
rect 30257 135 30327 140
rect 29828 59 29838 129
rect 30198 59 30208 129
rect 29828 49 30208 59
rect 30252 121 30332 135
rect 30252 69 30266 121
rect 30318 69 30332 121
rect 30252 55 30332 69
rect 30542 129 30922 139
rect 30971 135 31041 140
rect 30542 59 30552 129
rect 30912 59 30922 129
rect 30542 49 30922 59
rect 30966 121 31046 135
rect 30966 69 30980 121
rect 31032 69 31046 121
rect 30966 55 31046 69
rect 31256 129 31636 139
rect 31685 135 31755 140
rect 31256 59 31266 129
rect 31626 59 31636 129
rect 31256 49 31636 59
rect 31680 121 31760 135
rect 31680 69 31694 121
rect 31746 69 31760 121
rect 31680 55 31760 69
rect 31970 129 32350 139
rect 32399 135 32469 140
rect 31970 59 31980 129
rect 32340 59 32350 129
rect 31970 49 32350 59
rect 32394 121 32474 135
rect 32394 69 32408 121
rect 32460 69 32474 121
rect 32394 55 32474 69
rect 32684 129 33064 139
rect 33113 135 33183 140
rect 32684 59 32694 129
rect 33054 59 33064 129
rect 32684 49 33064 59
rect 33108 121 33188 135
rect 33108 69 33122 121
rect 33174 69 33188 121
rect 33108 55 33188 69
rect 33398 129 33778 139
rect 33827 135 33897 140
rect 33398 59 33408 129
rect 33768 59 33778 129
rect 33398 49 33778 59
rect 33822 121 33902 135
rect 33822 69 33836 121
rect 33888 69 33902 121
rect 33822 55 33902 69
rect 34112 129 34492 139
rect 34541 135 34611 140
rect 34112 59 34122 129
rect 34482 59 34492 129
rect 34112 49 34492 59
rect 34536 121 34616 135
rect 34536 69 34550 121
rect 34602 69 34616 121
rect 34536 55 34616 69
rect 34826 129 35206 139
rect 35255 135 35325 140
rect 34826 59 34836 129
rect 35196 59 35206 129
rect 34826 49 35206 59
rect 35250 121 35330 135
rect 35250 69 35264 121
rect 35316 69 35330 121
rect 35250 55 35330 69
rect 35540 129 35920 139
rect 35969 135 36039 140
rect 35540 59 35550 129
rect 35910 59 35920 129
rect 35540 49 35920 59
rect 35964 121 36044 135
rect 35964 69 35978 121
rect 36030 69 36044 121
rect 35964 55 36044 69
rect 36254 129 36634 139
rect 36683 135 36753 140
rect 36254 59 36264 129
rect 36624 59 36634 129
rect 36254 49 36634 59
rect 36678 121 36758 135
rect 36678 69 36692 121
rect 36744 69 36758 121
rect 36678 55 36758 69
rect 36968 129 37348 139
rect 37397 135 37467 140
rect 36968 59 36978 129
rect 37338 59 37348 129
rect 36968 49 37348 59
rect 37392 121 37472 135
rect 37392 69 37406 121
rect 37458 69 37472 121
rect 37392 55 37472 69
rect 37682 129 38062 139
rect 38111 135 38181 140
rect 37682 59 37692 129
rect 38052 59 38062 129
rect 37682 49 38062 59
rect 38106 121 38186 135
rect 38106 69 38120 121
rect 38172 69 38186 121
rect 38106 55 38186 69
rect 38396 129 38776 139
rect 38825 135 38895 140
rect 38396 59 38406 129
rect 38766 59 38776 129
rect 38396 49 38776 59
rect 38820 121 38900 135
rect 38820 69 38834 121
rect 38886 69 38900 121
rect 38820 55 38900 69
rect 15547 -50 15927 -40
rect 15547 -140 15557 -50
rect 15917 -140 15927 -50
rect 15547 -150 15927 -140
rect 16261 -50 16641 -40
rect 16261 -140 16271 -50
rect 16631 -140 16641 -50
rect 16261 -150 16641 -140
rect 16975 -50 17355 -40
rect 16975 -140 16985 -50
rect 17345 -140 17355 -50
rect 16975 -150 17355 -140
rect 17689 -50 18069 -40
rect 17689 -140 17699 -50
rect 18059 -140 18069 -50
rect 17689 -150 18069 -140
rect 18403 -50 18783 -40
rect 18403 -140 18413 -50
rect 18773 -140 18783 -50
rect 18403 -150 18783 -140
rect 19117 -50 19497 -40
rect 19117 -140 19127 -50
rect 19487 -140 19497 -50
rect 19117 -150 19497 -140
rect 19831 -50 20211 -40
rect 19831 -140 19841 -50
rect 20201 -140 20211 -50
rect 19831 -150 20211 -140
rect 20545 -50 20925 -40
rect 20545 -140 20555 -50
rect 20915 -140 20925 -50
rect 20545 -150 20925 -140
rect 21259 -50 21639 -40
rect 21259 -140 21269 -50
rect 21629 -140 21639 -50
rect 21259 -150 21639 -140
rect 21973 -50 22353 -40
rect 21973 -140 21983 -50
rect 22343 -140 22353 -50
rect 21973 -150 22353 -140
rect 22687 -50 23067 -40
rect 22687 -140 22697 -50
rect 23057 -140 23067 -50
rect 22687 -150 23067 -140
rect 23401 -50 23781 -40
rect 23401 -140 23411 -50
rect 23771 -140 23781 -50
rect 23401 -150 23781 -140
rect 24115 -50 24495 -40
rect 24115 -140 24125 -50
rect 24485 -140 24495 -50
rect 24115 -150 24495 -140
rect 24829 -50 25209 -40
rect 24829 -140 24839 -50
rect 25199 -140 25209 -50
rect 24829 -150 25209 -140
rect 25543 -50 25923 -40
rect 25543 -140 25553 -50
rect 25913 -140 25923 -50
rect 25543 -150 25923 -140
rect 26257 -50 26637 -40
rect 26257 -140 26267 -50
rect 26627 -140 26637 -50
rect 26257 -150 26637 -140
rect 26971 -50 27351 -40
rect 26971 -140 26981 -50
rect 27341 -140 27351 -50
rect 26971 -150 27351 -140
rect 27685 -50 28065 -40
rect 27685 -140 27695 -50
rect 28055 -140 28065 -50
rect 27685 -150 28065 -140
rect 28399 -50 28779 -40
rect 28399 -140 28409 -50
rect 28769 -140 28779 -50
rect 28399 -150 28779 -140
rect 29113 -50 29493 -40
rect 29113 -140 29123 -50
rect 29483 -140 29493 -50
rect 29113 -150 29493 -140
rect 29827 -50 30207 -40
rect 29827 -140 29837 -50
rect 30197 -140 30207 -50
rect 29827 -150 30207 -140
rect 30541 -50 30921 -40
rect 30541 -140 30551 -50
rect 30911 -140 30921 -50
rect 30541 -150 30921 -140
rect 31255 -50 31635 -40
rect 31255 -140 31265 -50
rect 31625 -140 31635 -50
rect 31255 -150 31635 -140
rect 31969 -50 32349 -40
rect 31969 -140 31979 -50
rect 32339 -140 32349 -50
rect 31969 -150 32349 -140
rect 32683 -50 33063 -40
rect 32683 -140 32693 -50
rect 33053 -140 33063 -50
rect 32683 -150 33063 -140
rect 33397 -50 33777 -40
rect 33397 -140 33407 -50
rect 33767 -140 33777 -50
rect 33397 -150 33777 -140
rect 34111 -50 34491 -40
rect 34111 -140 34121 -50
rect 34481 -140 34491 -50
rect 34111 -150 34491 -140
rect 34825 -50 35205 -40
rect 34825 -140 34835 -50
rect 35195 -140 35205 -50
rect 34825 -150 35205 -140
rect 35539 -50 35919 -40
rect 35539 -140 35549 -50
rect 35909 -140 35919 -50
rect 35539 -150 35919 -140
rect 36253 -50 36633 -40
rect 36253 -140 36263 -50
rect 36623 -140 36633 -50
rect 36253 -150 36633 -140
rect 36967 -50 37347 -40
rect 36967 -140 36977 -50
rect 37337 -140 37347 -50
rect 36967 -150 37347 -140
rect 37681 -50 38061 -40
rect 37681 -140 37691 -50
rect 38051 -140 38061 -50
rect 37681 -150 38061 -140
rect 38395 -50 38775 -40
rect 38395 -140 38405 -50
rect 38765 -140 38775 -50
rect 38395 -150 38775 -140
rect 39080 -130 39120 229
rect 39150 40 39190 299
rect 39220 210 39260 369
rect 39290 370 39330 439
rect 39370 370 39390 380
rect 39290 330 39390 370
rect 39370 320 39390 330
rect 39770 320 39790 380
rect 39900 370 40320 380
rect 39900 310 39920 370
rect 40300 310 40320 370
rect 39900 300 40320 310
rect 39370 210 39390 220
rect 39220 170 39390 210
rect 39370 160 39390 170
rect 39770 160 39790 220
rect 39900 210 40320 220
rect 39900 150 39920 210
rect 40300 150 40320 210
rect 39900 140 40320 150
rect 39900 50 40320 60
rect 39370 40 39390 50
rect 39150 0 39390 40
rect 39370 -10 39390 0
rect 39770 -10 39790 50
rect 39900 -10 39920 50
rect 40300 -10 40320 50
rect 39900 -20 40320 -10
rect 39900 -120 40320 -110
rect 39370 -130 39390 -120
rect 39080 -170 39390 -130
rect 39370 -180 39390 -170
rect 39770 -180 39790 -120
rect 39900 -180 39920 -120
rect 40300 -180 40320 -120
rect 9880 -200 14400 -180
rect 39900 -190 40320 -180
rect 3941 -529 4061 -519
rect 10020 -420 10280 -400
rect 10780 -420 10980 -400
rect 3766 -569 3846 -564
rect 3761 -578 3846 -569
rect 3761 -580 3780 -578
rect 2927 -630 3780 -580
rect 3832 -630 3846 -578
rect 2927 -644 3846 -630
rect 2927 -660 3827 -644
rect 10020 -740 10040 -420
rect 10160 -740 10280 -420
rect 10480 -440 10640 -420
rect 10480 -700 10500 -440
rect 10620 -700 10640 -440
rect 10480 -720 10640 -700
rect 10020 -760 10280 -740
rect 10780 -740 10800 -420
rect 10960 -740 10980 -420
rect 10780 -760 10980 -740
rect 10546 -786 10552 -775
rect 10514 -827 10552 -786
rect 10604 -786 10610 -775
rect 10604 -800 10616 -786
rect 11200 -790 11300 -780
rect 10604 -827 10960 -800
rect 10514 -830 10960 -827
rect 10514 -834 10880 -830
rect 10550 -840 10880 -834
rect 10870 -890 10880 -840
rect 10950 -890 10960 -830
rect 11200 -870 11210 -790
rect 11290 -870 11300 -790
rect 11200 -880 11300 -870
rect 10870 -900 10960 -890
rect 11380 -1090 11480 -1080
rect 10480 -1130 10640 -1120
rect 10480 -1240 10490 -1130
rect 10630 -1240 10640 -1130
rect 11380 -1170 11390 -1090
rect 11470 -1170 11480 -1090
rect 11380 -1180 11480 -1170
rect 10480 -1250 10640 -1240
rect 11310 -1490 11410 -1480
rect 11310 -1570 11320 -1490
rect 11400 -1570 11410 -1490
rect 11310 -1580 11410 -1570
rect 5802 -2100 7202 -2000
rect 5802 -2580 5902 -2100
rect 1720 -2600 5902 -2580
rect 1720 -2780 1760 -2600
rect 1820 -2780 2080 -2600
rect 2140 -2700 5902 -2600
rect 7102 -2700 7202 -2100
rect 2140 -2780 7202 -2700
rect 1720 -2800 7202 -2780
rect 9002 -2100 10402 -2000
rect 9002 -2700 9102 -2100
rect 10302 -2700 10402 -2100
rect 9002 -2800 10402 -2700
rect 5802 -2940 10622 -2800
rect 11321 -2831 11404 -1580
rect 5802 -3020 10402 -2940
rect 5802 -3100 6820 -3020
rect 5802 -3400 6700 -3100
rect 6800 -3400 6820 -3100
rect 5802 -3500 6820 -3400
rect 5802 -3800 6700 -3500
rect 6800 -3800 6820 -3500
rect 5802 -3900 6820 -3800
rect 5802 -4000 6700 -3900
rect 6000 -4166 6100 -4000
rect 6200 -4166 6300 -4000
rect 6400 -4160 6500 -4000
rect 6600 -4160 6700 -4000
rect 6800 -4160 6820 -3900
rect 6400 -4166 6820 -4160
rect 5850 -4236 6820 -4166
rect 5850 -4388 5902 -4236
rect 5170 -5640 5320 -5620
rect 5170 -6030 5190 -5640
rect 5300 -6030 5320 -5640
rect 5170 -6050 5320 -6030
rect 5400 -5640 5550 -5620
rect 5400 -6030 5420 -5640
rect 5530 -6030 5550 -5640
rect 5400 -6050 5550 -6030
rect 5850 -6376 5902 -6364
rect 5968 -4388 6020 -4236
rect 5968 -6376 6020 -6364
rect 6086 -4388 6138 -4376
rect 6086 -6614 6138 -6364
rect 6204 -4388 6256 -4236
rect 6440 -4240 6820 -4236
rect 6880 -3100 9120 -3020
rect 6880 -4240 6900 -3100
rect 6440 -4260 6900 -4240
rect 7058 -3120 8942 -3100
rect 7058 -3272 7110 -3120
rect 6204 -6376 6256 -6364
rect 6322 -4388 6374 -4376
rect 6200 -6504 6261 -6495
rect 6200 -6560 6202 -6504
rect 6258 -6560 6261 -6504
rect 6200 -6569 6261 -6560
rect 6322 -6614 6374 -6364
rect 6440 -4388 6492 -4260
rect 6440 -6376 6492 -6364
rect 6558 -4388 6610 -4260
rect 7058 -5260 7110 -5248
rect 7516 -3272 7568 -3260
rect 7516 -5292 7568 -5248
rect 7974 -3272 8026 -3120
rect 7974 -5260 8026 -5248
rect 8432 -3272 8484 -3260
rect 8432 -5292 8484 -5248
rect 8890 -3272 8942 -3120
rect 9100 -4240 9120 -3100
rect 9180 -3100 10402 -3020
rect 9180 -3400 9200 -3100
rect 9300 -3400 10242 -3100
rect 9180 -3500 10242 -3400
rect 9180 -3800 9200 -3500
rect 9300 -3800 10242 -3500
rect 9180 -4000 10242 -3800
rect 10382 -3860 10402 -3100
rect 10602 -3860 10622 -2940
rect 11322 -2952 11402 -2831
rect 11202 -3130 11402 -2952
rect 10964 -3200 10983 -3130
rect 11412 -3200 11435 -3130
rect 10382 -3880 10622 -3860
rect 10852 -3815 10867 -3763
rect 11336 -3815 11353 -3763
rect 9180 -4160 9200 -4000
rect 9300 -4160 9400 -4000
rect 9500 -4160 9600 -4000
rect 9180 -4166 9600 -4160
rect 9700 -4166 9800 -4000
rect 9900 -4166 10000 -4000
rect 10100 -4166 10200 -4000
rect 10852 -4032 10872 -3815
rect 11082 -4032 11102 -3815
rect 10852 -4051 11102 -4032
rect 9180 -4236 10200 -4166
rect 9180 -4240 9561 -4236
rect 9100 -4260 9561 -4240
rect 8890 -5260 8942 -5248
rect 9391 -4388 9443 -4260
rect 7205 -5384 8795 -5292
rect 8880 -5298 9202 -5290
rect 8944 -5300 9202 -5298
rect 8944 -5360 9032 -5300
rect 9192 -5360 9202 -5300
rect 8944 -5362 9202 -5360
rect 8880 -5370 9202 -5362
rect 7205 -5470 7259 -5384
rect 7397 -5470 7451 -5384
rect 7589 -5470 7643 -5384
rect 7781 -5470 7835 -5384
rect 7973 -5470 8027 -5384
rect 8165 -5470 8219 -5384
rect 8357 -5470 8411 -5384
rect 8549 -5470 8603 -5384
rect 8741 -5470 8795 -5384
rect 7205 -5540 8795 -5470
rect 7205 -5700 7259 -5540
rect 7295 -5594 7361 -5580
rect 7295 -5662 7361 -5656
rect 7397 -5700 7451 -5540
rect 7487 -5594 7553 -5580
rect 7487 -5662 7553 -5656
rect 7589 -5700 7643 -5540
rect 7679 -5594 7745 -5580
rect 7679 -5662 7745 -5656
rect 7781 -5700 7835 -5540
rect 7871 -5594 7937 -5580
rect 7871 -5662 7937 -5656
rect 7973 -5700 8027 -5540
rect 8063 -5594 8129 -5580
rect 8063 -5662 8129 -5656
rect 8165 -5700 8219 -5540
rect 8255 -5594 8321 -5580
rect 8255 -5662 8321 -5656
rect 8357 -5700 8411 -5540
rect 8447 -5594 8513 -5580
rect 8447 -5662 8513 -5656
rect 8549 -5700 8603 -5540
rect 8639 -5594 8705 -5580
rect 8639 -5662 8705 -5656
rect 8741 -5700 8795 -5540
rect 7007 -6200 7013 -5700
rect 7067 -6200 7073 -5700
rect 7103 -6200 7109 -5700
rect 7163 -6200 7169 -5700
rect 7199 -6200 7205 -5700
rect 7259 -6200 7265 -5700
rect 7295 -6200 7301 -5700
rect 7355 -6200 7361 -5700
rect 7391 -6200 7397 -5700
rect 7451 -6200 7457 -5700
rect 7487 -6200 7493 -5700
rect 7547 -6200 7553 -5700
rect 7583 -6200 7589 -5700
rect 7643 -6200 7649 -5700
rect 7679 -6200 7685 -5700
rect 7739 -6200 7745 -5700
rect 7775 -6200 7781 -5700
rect 7835 -6200 7841 -5700
rect 7871 -6200 7877 -5700
rect 7931 -6200 7937 -5700
rect 7967 -6200 7973 -5700
rect 8027 -6200 8033 -5700
rect 8063 -6200 8069 -5700
rect 8123 -6200 8129 -5700
rect 8159 -6200 8165 -5700
rect 8219 -6200 8225 -5700
rect 8255 -6200 8261 -5700
rect 8315 -6200 8321 -5700
rect 8351 -6200 8357 -5700
rect 8411 -6200 8417 -5700
rect 8447 -6200 8453 -5700
rect 8507 -6200 8513 -5700
rect 8543 -6200 8549 -5700
rect 8603 -6200 8609 -5700
rect 8639 -6200 8645 -5700
rect 8699 -6200 8705 -5700
rect 8735 -6200 8741 -5700
rect 8795 -6200 8801 -5700
rect 8831 -6200 8837 -5700
rect 8891 -6200 8897 -5700
rect 8927 -6200 8933 -5700
rect 8987 -6200 8993 -5700
rect 6558 -6376 6610 -6364
rect 7295 -6270 7361 -6200
rect 7487 -6270 7553 -6200
rect 7679 -6270 7745 -6200
rect 7871 -6270 7937 -6200
rect 7295 -6410 7937 -6270
rect 8063 -6270 8129 -6200
rect 8255 -6270 8321 -6200
rect 8447 -6270 8513 -6200
rect 8639 -6270 8705 -6200
rect 8063 -6410 8705 -6270
rect 9391 -6376 9443 -6364
rect 9509 -4388 9561 -4260
rect 9509 -6376 9561 -6364
rect 9627 -4388 9679 -4376
rect 6000 -6650 6493 -6614
rect 6000 -6740 6010 -6650
rect 6120 -6666 6493 -6650
rect 6120 -6740 6130 -6666
rect 6441 -6736 6493 -6666
rect 6000 -6750 6130 -6740
rect 6204 -6788 6965 -6736
rect 7384 -6737 7436 -6410
rect 7911 -6736 8144 -6730
rect 8564 -6736 8616 -6410
rect 9627 -6495 9679 -6364
rect 9745 -4388 9797 -4236
rect 9745 -6376 9797 -6364
rect 9863 -4388 9915 -4376
rect 9863 -6495 9915 -6364
rect 9981 -4388 10033 -4236
rect 9981 -6376 10033 -6364
rect 10099 -4388 10151 -4236
rect 10099 -6376 10151 -6364
rect 9627 -6504 9915 -6495
rect 9627 -6560 9743 -6504
rect 9799 -6560 9915 -6504
rect 9627 -6569 9915 -6560
rect 9627 -6614 9679 -6569
rect 9863 -6614 9915 -6569
rect 9508 -6666 9915 -6614
rect 9508 -6736 9560 -6666
rect 6086 -6897 6138 -6885
rect 6086 -9034 6138 -8873
rect 6204 -6897 6257 -6788
rect 6441 -6885 6493 -6788
rect 6677 -6885 6729 -6788
rect 6913 -6885 6965 -6788
rect 7149 -6738 7436 -6737
rect 7620 -6738 7883 -6736
rect 7149 -6788 7883 -6738
rect 7149 -6789 7620 -6788
rect 7149 -6885 7201 -6789
rect 7384 -6790 7620 -6789
rect 6256 -6965 6257 -6897
rect 6322 -6897 6374 -6885
rect 6204 -8885 6256 -8873
rect 6322 -9034 6374 -8873
rect 6440 -6897 6493 -6885
rect 6492 -6965 6493 -6897
rect 6558 -6897 6610 -6885
rect 6440 -8885 6492 -8873
rect 6558 -9034 6610 -8873
rect 6676 -6897 6729 -6885
rect 6728 -6965 6729 -6897
rect 6794 -6897 6846 -6885
rect 6676 -8885 6728 -8873
rect 6794 -9034 6846 -8873
rect 6912 -6897 6965 -6885
rect 6964 -6965 6965 -6897
rect 7030 -6897 7082 -6885
rect 6912 -8885 6964 -8873
rect 7030 -9034 7082 -8873
rect 7148 -6897 7201 -6885
rect 7200 -6965 7201 -6897
rect 7266 -6897 7318 -6885
rect 7148 -8885 7200 -8873
rect 7266 -9034 7318 -8873
rect 7384 -6897 7436 -6790
rect 7854 -6828 7883 -6788
rect 7911 -6748 8852 -6736
rect 7911 -6800 7917 -6748
rect 7969 -6758 8852 -6748
rect 7969 -6800 7975 -6758
rect 8032 -6792 8084 -6786
rect 7854 -6844 8032 -6828
rect 7854 -6850 8084 -6844
rect 8112 -6788 8852 -6758
rect 7854 -6856 8060 -6850
rect 7384 -8885 7436 -8873
rect 7502 -6897 7554 -6885
rect 7502 -9034 7554 -8873
rect 7620 -6897 7672 -6885
rect 7620 -8885 7672 -8873
rect 7738 -6897 7790 -6885
rect 7738 -9034 7790 -8873
rect 7856 -6897 7908 -6856
rect 8112 -6878 8144 -6788
rect 7856 -8885 7908 -8873
rect 7974 -6897 8026 -6884
rect 7974 -9034 8026 -8873
rect 8092 -6897 8144 -6878
rect 8092 -8885 8144 -8873
rect 8210 -6897 8262 -6885
rect 8210 -9034 8262 -8873
rect 8328 -6897 8380 -6885
rect 8328 -8885 8380 -8873
rect 8446 -6897 8498 -6885
rect 8446 -9034 8498 -8873
rect 8564 -6897 8616 -6788
rect 8564 -8885 8616 -8873
rect 8682 -6897 8734 -6885
rect 8682 -9034 8734 -8873
rect 8800 -6897 8852 -6788
rect 9036 -6788 9796 -6736
rect 8800 -8885 8852 -8873
rect 8918 -6897 8970 -6885
rect 8918 -9034 8970 -8873
rect 9036 -6897 9088 -6788
rect 9036 -8885 9088 -8873
rect 9154 -6897 9206 -6885
rect 9154 -9034 9206 -8873
rect 9272 -6897 9324 -6788
rect 9272 -8885 9324 -8873
rect 9390 -6897 9442 -6885
rect 9390 -9034 9442 -8873
rect 9508 -6897 9560 -6788
rect 9508 -8885 9560 -8873
rect 9626 -6897 9678 -6885
rect 9626 -9034 9678 -8873
rect 9744 -6897 9796 -6788
rect 9744 -8885 9796 -8873
rect 9862 -6897 9914 -6885
rect 9862 -9034 9914 -8873
rect 6086 -9136 9914 -9034
rect 6108 -9200 6208 -9136
rect 6600 -9200 6700 -9136
rect 7000 -9200 7100 -9136
rect 7400 -9200 7500 -9136
rect 7800 -9200 7900 -9136
rect 8100 -9200 8200 -9136
rect 8500 -9200 8600 -9136
rect 8900 -9200 9000 -9136
rect 9300 -9200 9400 -9136
rect 9792 -9200 9892 -9136
rect 6108 -9300 9892 -9200
rect 6108 -9400 6502 -9300
rect 6402 -9800 6502 -9400
rect 9702 -9400 9892 -9300
rect 9702 -9800 9802 -9400
rect 6402 -9900 9802 -9800
<< via2 >>
rect 6502 12700 9702 13200
rect 6010 10050 6120 10140
rect 5190 9040 5300 9430
rect 5420 9040 5530 9430
rect 6202 9958 6258 9960
rect 6202 9906 6204 9958
rect 6204 9906 6256 9958
rect 6256 9906 6258 9958
rect 6202 9904 6258 9906
rect 9743 9958 9799 9960
rect 9743 9906 9745 9958
rect 9745 9906 9797 9958
rect 9797 9906 9799 9958
rect 9743 9904 9799 9906
rect 7295 9000 7361 9050
rect 7295 8994 7361 9000
rect 7487 9000 7553 9050
rect 7487 8994 7553 9000
rect 7679 9000 7745 9050
rect 7679 8994 7745 9000
rect 7871 9000 7937 9050
rect 7871 8994 7937 9000
rect 8063 9000 8129 9050
rect 8063 8994 8129 9000
rect 8255 9000 8321 9050
rect 8255 8994 8321 9000
rect 8447 9000 8513 9050
rect 8447 8994 8513 9000
rect 8639 9000 8705 9050
rect 8639 8994 8705 9000
rect 9032 8700 9192 8760
rect 10402 6340 10602 7260
rect 10872 7215 11082 7432
rect 10872 7212 11082 7215
rect 5902 5500 7102 6100
rect 9102 5500 10302 6100
rect 11030 4830 11110 4910
rect 11190 4830 11270 4910
rect 11330 4680 11410 4760
rect 3358 3975 3458 4345
rect 3581 3972 3641 4332
rect 4201 3972 4261 4332
rect 4384 3975 4484 4345
rect 1940 2460 2020 2540
rect 1940 1880 2020 1960
rect 1900 1120 2000 1220
rect 2260 960 2360 1040
rect 1740 800 1820 920
rect 2080 800 2160 920
rect 3358 3251 3458 3621
rect 3581 3264 3681 3614
rect 4161 3264 4261 3614
rect 4384 3251 4484 3621
rect 2907 960 2987 1040
rect 2640 780 2740 860
rect 9260 3978 14420 4260
rect 9260 3960 11278 3978
rect 11278 3960 14420 3978
rect 9260 2960 9460 3960
rect 5447 2840 5867 2920
rect 6647 2840 7067 2920
rect 7847 2840 8267 2920
rect 9047 2840 9467 2920
rect 3247 2380 3250 2600
rect 3250 2380 3627 2600
rect 3247 1820 3250 2040
rect 3250 1820 3627 2040
rect 4747 2180 5167 2260
rect 6047 2180 6467 2240
rect 6047 2160 6467 2180
rect 7247 2180 7667 2240
rect 7247 2160 7667 2180
rect 8447 2180 8867 2240
rect 8447 2160 8867 2180
rect 9647 2180 10067 2240
rect 9647 2160 10067 2180
rect 5447 1580 5867 1600
rect 5447 1520 5867 1580
rect 6647 1580 7067 1600
rect 6647 1520 7067 1580
rect 7847 1580 8267 1600
rect 7847 1520 8267 1580
rect 9047 1580 9467 1600
rect 9047 1520 9467 1580
rect 3247 1140 3327 1220
rect 4407 1276 4787 1280
rect 4407 1040 4782 1276
rect 4782 1040 4787 1276
rect 10200 1850 10260 1930
rect 13988 2118 14048 2328
rect 12820 1610 13170 1690
rect 13918 1638 13978 1698
rect 14248 1638 14308 1698
rect 12820 1360 13170 1440
rect 13918 1348 13978 1408
rect 14248 1348 14308 1408
rect 10200 1160 10260 1240
rect 3087 780 3167 860
rect 6047 840 6467 900
rect 6047 820 6467 840
rect 7247 840 7667 900
rect 7247 820 7667 840
rect 8447 840 8867 900
rect 8447 820 8867 840
rect 9647 840 10067 900
rect 9647 820 10067 840
rect 3768 202 3828 562
rect 3951 205 4051 575
rect 11090 840 11190 920
rect 13988 718 14058 928
rect 15557 912 15917 1002
rect 16271 912 16631 1002
rect 16985 912 17345 1002
rect 17699 912 18059 1002
rect 18413 912 18773 1002
rect 19127 912 19487 1002
rect 19841 912 20201 1002
rect 20555 912 20915 1002
rect 21269 912 21629 1002
rect 21983 912 22343 1002
rect 22697 912 23057 1002
rect 23411 912 23771 1002
rect 24125 912 24485 1002
rect 24839 912 25199 1002
rect 25553 912 25913 1002
rect 26267 912 26627 1002
rect 26981 912 27341 1002
rect 27695 912 28055 1002
rect 28409 912 28769 1002
rect 29123 912 29483 1002
rect 29837 912 30197 1002
rect 30551 912 30911 1002
rect 31265 912 31625 1002
rect 31979 912 32339 1002
rect 32693 912 33053 1002
rect 33407 912 33767 1002
rect 34121 912 34481 1002
rect 34835 912 35195 1002
rect 35549 912 35909 1002
rect 36263 912 36623 1002
rect 36977 912 37337 1002
rect 37691 912 38061 1012
rect 38395 912 38765 1012
rect 15558 733 15918 793
rect 16272 733 16632 793
rect 16986 733 17346 793
rect 17700 733 18060 793
rect 18414 733 18774 793
rect 19128 733 19488 793
rect 19842 733 20202 793
rect 20556 733 20916 793
rect 21270 733 21630 793
rect 21984 733 22344 793
rect 22698 733 23058 793
rect 23412 733 23772 793
rect 24126 733 24486 793
rect 24840 733 25200 793
rect 25554 733 25914 793
rect 26268 733 26628 793
rect 26982 733 27342 793
rect 27696 733 28056 793
rect 28410 733 28770 793
rect 29124 733 29484 793
rect 29838 733 30198 793
rect 30552 733 30912 793
rect 31266 733 31626 793
rect 31980 733 32340 793
rect 32694 733 33054 793
rect 33408 733 33768 793
rect 34122 733 34482 793
rect 34836 733 35196 793
rect 35550 733 35910 793
rect 36264 733 36624 793
rect 39920 980 40300 1040
rect 36978 733 37338 793
rect 37698 689 38048 789
rect 38408 729 38768 789
rect 39920 820 40300 880
rect 39920 650 40300 710
rect 39920 480 40300 540
rect 3728 -506 3828 -156
rect 3951 -519 4051 -149
rect 9900 78 10358 100
rect 10358 78 14380 100
rect 9900 -180 14380 78
rect 15558 69 15918 129
rect 16272 69 16632 129
rect 16986 69 17346 129
rect 17700 69 18060 129
rect 18414 69 18774 129
rect 19128 69 19488 129
rect 19842 69 20202 129
rect 20556 69 20916 129
rect 21270 69 21630 129
rect 21984 69 22344 129
rect 22698 69 23058 129
rect 23412 69 23772 129
rect 24126 69 24486 129
rect 24840 69 25200 129
rect 25554 69 25914 129
rect 26268 69 26628 129
rect 26982 69 27342 129
rect 27696 69 28056 129
rect 28410 69 28770 129
rect 29124 69 29484 129
rect 29838 69 30198 129
rect 30552 69 30912 129
rect 31266 69 31626 129
rect 31980 69 32340 129
rect 32694 69 33054 129
rect 33408 69 33768 129
rect 34122 69 34482 129
rect 34836 69 35196 129
rect 35550 69 35910 129
rect 36264 69 36624 129
rect 36978 69 37338 129
rect 37692 69 38052 129
rect 38406 69 38766 129
rect 15557 -140 15917 -50
rect 16271 -140 16631 -50
rect 16985 -140 17345 -50
rect 17699 -140 18059 -50
rect 18413 -140 18773 -50
rect 19127 -140 19487 -50
rect 19841 -140 20201 -50
rect 20555 -140 20915 -50
rect 21269 -140 21629 -50
rect 21983 -140 22343 -50
rect 22697 -140 23057 -50
rect 23411 -140 23771 -50
rect 24125 -140 24485 -50
rect 24839 -140 25199 -50
rect 25553 -140 25913 -50
rect 26267 -140 26627 -50
rect 26981 -140 27341 -50
rect 27695 -140 28055 -50
rect 28409 -140 28769 -50
rect 29123 -140 29483 -50
rect 29837 -140 30197 -50
rect 30551 -140 30911 -50
rect 31265 -140 31625 -50
rect 31979 -140 32339 -50
rect 32693 -140 33053 -50
rect 33407 -140 33767 -50
rect 34121 -140 34481 -50
rect 34835 -140 35195 -50
rect 35549 -140 35909 -50
rect 36263 -140 36623 -50
rect 36977 -140 37337 -50
rect 37691 -140 38051 -50
rect 38405 -140 38765 -50
rect 39920 310 40300 370
rect 39920 150 40300 210
rect 39920 -10 40300 50
rect 39920 -180 40300 -120
rect 10040 -740 10160 -420
rect 10500 -700 10620 -440
rect 10880 -740 10960 -420
rect 10880 -890 10950 -830
rect 11210 -870 11290 -790
rect 10490 -1240 10630 -1130
rect 11390 -1170 11470 -1090
rect 11320 -1570 11400 -1490
rect 1760 -2780 1820 -2600
rect 2080 -2780 2140 -2600
rect 5902 -2700 7102 -2100
rect 9102 -2700 10302 -2100
rect 5190 -6030 5300 -5640
rect 5420 -6030 5530 -5640
rect 6202 -6506 6258 -6504
rect 6202 -6558 6204 -6506
rect 6204 -6558 6256 -6506
rect 6256 -6558 6258 -6506
rect 6202 -6560 6258 -6558
rect 10402 -3860 10602 -2940
rect 10872 -3815 11082 -3812
rect 10872 -4032 11082 -3815
rect 9032 -5360 9192 -5300
rect 7295 -5600 7361 -5594
rect 7295 -5650 7361 -5600
rect 7487 -5600 7553 -5594
rect 7487 -5650 7553 -5600
rect 7679 -5600 7745 -5594
rect 7679 -5650 7745 -5600
rect 7871 -5600 7937 -5594
rect 7871 -5650 7937 -5600
rect 8063 -5600 8129 -5594
rect 8063 -5650 8129 -5600
rect 8255 -5600 8321 -5594
rect 8255 -5650 8321 -5600
rect 8447 -5600 8513 -5594
rect 8447 -5650 8513 -5600
rect 8639 -5600 8705 -5594
rect 8639 -5650 8705 -5600
rect 6010 -6740 6120 -6650
rect 9743 -6506 9799 -6504
rect 9743 -6558 9745 -6506
rect 9745 -6558 9797 -6506
rect 9797 -6558 9799 -6506
rect 9743 -6560 9799 -6558
rect 6502 -9800 9702 -9300
<< metal3 >>
rect 6402 13200 9802 13300
rect 5000 10100 5800 12800
rect 6402 12700 6502 13200
rect 9702 12700 9802 13200
rect 6402 12600 9802 12700
rect 6000 10140 6130 10150
rect 5000 9980 5600 10100
rect 6000 10050 6010 10140
rect 6120 10050 6130 10140
rect 6000 10040 6130 10050
rect 5000 9820 5020 9980
rect 5580 9820 5600 9980
rect 5000 9740 5030 9820
rect 5570 9740 5600 9820
rect 5000 9710 5600 9740
rect 5660 9960 9807 9969
rect 5660 9904 6202 9960
rect 6258 9904 9743 9960
rect 9799 9904 9807 9960
rect 5660 9895 9807 9904
rect 5220 9450 5290 9710
rect 5170 9430 5320 9450
rect 5170 9040 5190 9430
rect 5300 9040 5320 9430
rect 5170 9020 5320 9040
rect 5400 9449 5550 9450
rect 5660 9449 5734 9895
rect 6261 9864 9740 9895
rect 5400 9430 5734 9449
rect 5400 9040 5420 9430
rect 5530 9375 5734 9430
rect 5530 9040 5550 9375
rect 5400 9020 5550 9040
rect 7289 9050 7943 9062
rect 7289 8994 7295 9050
rect 7361 8994 7487 9050
rect 7553 8994 7679 9050
rect 7745 8994 7871 9050
rect 7937 8994 7943 9050
rect 7289 8980 7943 8994
rect 8057 9050 8711 9062
rect 8057 8994 8063 9050
rect 8129 8994 8255 9050
rect 8321 8994 8447 9050
rect 8513 8994 8639 9050
rect 8705 8994 8711 9050
rect 8057 8980 8711 8994
rect 7300 7240 7500 8980
rect -1020 7180 -520 7240
rect -40 7180 7500 7240
rect -1020 7100 7500 7180
rect -1020 7040 -520 7100
rect -40 7040 7500 7100
rect -1020 -7320 -820 7040
rect 5802 6100 7202 6200
rect 5802 5500 5902 6100
rect 7102 5500 7202 6100
rect 5802 5400 7202 5500
rect 8480 5180 8680 8980
rect 9022 8760 9202 8770
rect 9022 8700 9032 8760
rect 9192 8700 9202 8760
rect 9022 7500 9202 8700
rect 10302 7700 11602 13052
rect 9902 7500 11602 7700
rect 9022 7200 10202 7500
rect 10302 7452 11602 7500
rect 10702 7432 11602 7452
rect 10302 7260 10622 7280
rect 10302 6340 10322 7260
rect 10602 6340 10622 7260
rect 10702 7212 10872 7432
rect 11082 7212 11602 7432
rect 10702 6952 11602 7212
rect 10702 6552 10802 6952
rect 11502 6552 11602 6952
rect 10702 6452 11602 6552
rect 10302 6320 10622 6340
rect 9002 6100 10402 6200
rect 9002 5500 9102 6100
rect 10302 5500 10402 6100
rect 9002 5400 10402 5500
rect 12002 6100 14802 13000
rect 12002 5500 12102 6100
rect 14702 5500 14802 6100
rect 12002 5400 14802 5500
rect 8480 4980 14900 5180
rect 11020 4910 11120 4920
rect 11020 4830 11030 4910
rect 11110 4830 11120 4910
rect 11020 4820 11120 4830
rect 11180 4910 11280 4920
rect 11180 4830 11190 4910
rect 11270 4830 11280 4910
rect 11180 4820 11280 4830
rect 11320 4760 11420 4770
rect 11320 4680 11330 4760
rect 11410 4680 11420 4760
rect 11320 4670 11420 4680
rect -380 4440 -180 4460
rect -380 4280 -360 4440
rect -200 4280 -180 4440
rect -380 4260 -180 4280
rect 1478 4345 3508 4355
rect 1478 4315 3358 4345
rect 3458 4315 3508 4345
rect -340 2560 -220 4260
rect 1478 3995 3228 4315
rect 3468 3995 3508 4315
rect 1478 3975 3358 3995
rect 3458 3975 3508 3995
rect 1478 3961 3508 3975
rect 3571 4332 4271 4352
rect 3571 3972 3581 4332
rect 3641 4212 4201 4332
rect 3641 4112 3651 4212
rect 3787 4112 3947 4212
rect 4191 4112 4201 4212
rect 3641 3972 4201 4112
rect 4261 3972 4271 4332
rect 3571 3962 3651 3972
rect -92 3621 3508 3641
rect 3787 3634 3947 3972
rect 4191 3962 4271 3972
rect 4334 4345 6364 4355
rect 4334 4315 4384 4345
rect 4484 4315 6364 4345
rect 4334 3995 4374 4315
rect 4614 3995 6364 4315
rect 4334 3975 4384 3995
rect 4484 3975 6364 3995
rect 4334 3961 6364 3975
rect 8600 4260 14440 4280
rect 8600 3960 8620 4260
rect 14420 3960 14440 4260
rect 8600 3940 9260 3960
rect -92 3601 3358 3621
rect 3458 3601 3508 3621
rect -92 3281 3228 3601
rect 3468 3281 3508 3601
rect -92 3251 3358 3281
rect 3458 3251 3508 3281
rect 3571 3614 4271 3634
rect 3571 3264 3581 3614
rect 3681 3494 4161 3614
rect 3681 3394 3691 3494
rect 3787 3394 3947 3494
rect 4151 3394 4161 3494
rect 3681 3264 4161 3394
rect 4261 3264 4271 3614
rect 3571 3254 4271 3264
rect 4334 3621 7934 3641
rect 4334 3601 4384 3621
rect 4484 3601 7934 3621
rect 4334 3281 4374 3601
rect 4614 3281 7934 3601
rect -92 3247 3508 3251
rect 3348 3241 3468 3247
rect 3227 2600 3647 2620
rect -340 2540 2040 2560
rect -340 2460 1940 2540
rect 2020 2460 2040 2540
rect -340 2440 2040 2460
rect 3227 2380 3247 2600
rect 3627 2380 3647 2600
rect 3227 2360 3647 2380
rect 3787 2300 3947 3254
rect 4334 3251 4384 3281
rect 4484 3251 7934 3281
rect 4334 3247 7934 3251
rect 4374 3241 4494 3247
rect 9240 2960 9260 3940
rect 9460 3940 14440 3960
rect 9460 2960 9480 3940
rect 9240 2940 9480 2960
rect 5427 2920 9487 2940
rect 5427 2840 5447 2920
rect 5867 2840 6647 2920
rect 7067 2840 7847 2920
rect 8267 2840 9047 2920
rect 9467 2840 9487 2920
rect 5427 2820 9487 2840
rect 3787 2260 5247 2300
rect 3787 2180 4747 2260
rect 5167 2180 5247 2260
rect 3787 2140 5247 2180
rect 3227 2040 3647 2060
rect -340 1960 2040 1980
rect -340 1880 1940 1960
rect 2020 1880 2040 1960
rect -340 1860 2040 1880
rect -340 0 -220 1860
rect 3227 1820 3247 2040
rect 3627 1820 3647 2040
rect 3227 1800 3647 1820
rect 3787 1700 3947 2140
rect 3427 1540 3947 1700
rect 5427 1620 5547 2820
rect 5767 1620 5887 2820
rect 5427 1600 5887 1620
rect 1880 1220 3347 1240
rect 1880 1120 1900 1220
rect 2000 1140 3247 1220
rect 3327 1140 3347 1220
rect 2000 1120 3347 1140
rect 1880 1100 2020 1120
rect 1720 920 1840 940
rect 1720 800 1740 920
rect 1820 800 1840 920
rect 1720 780 1840 800
rect -380 -20 -180 0
rect -380 -180 -360 -20
rect -200 -180 -180 -20
rect -380 -200 -180 -180
rect 1740 -2600 1840 780
rect 1740 -2780 1760 -2600
rect 1820 -2780 1840 -2600
rect 1740 -6680 1840 -2780
rect 1900 -6680 2000 1100
rect 2240 1040 3007 1060
rect 2240 960 2260 1040
rect 2360 960 2907 1040
rect 2987 960 3007 1040
rect 2240 940 3007 960
rect 2060 920 2180 940
rect 2060 800 2080 920
rect 2160 800 2180 920
rect 2060 780 2180 800
rect 2060 -2600 2160 780
rect 2060 -2780 2080 -2600
rect 2140 -2780 2160 -2600
rect 2060 -6680 2160 -2780
rect 2240 -6680 2360 940
rect 3427 920 3587 1540
rect 5427 1520 5447 1600
rect 5867 1520 5887 1600
rect 5427 1500 5887 1520
rect 6027 2240 6487 2260
rect 6027 2160 6047 2240
rect 6467 2160 6487 2240
rect 6027 2140 6487 2160
rect 4387 1280 4807 1300
rect 4387 1040 4407 1280
rect 4787 1040 4807 1280
rect 4387 1020 4807 1040
rect 6027 920 6147 2140
rect 6367 920 6487 2140
rect 6627 1620 6747 2820
rect 6967 1620 7087 2820
rect 6627 1600 7087 1620
rect 6627 1520 6647 1600
rect 7067 1520 7087 1600
rect 6627 1500 7087 1520
rect 7227 2240 7687 2260
rect 7227 2160 7247 2240
rect 7667 2160 7687 2240
rect 7227 2140 7687 2160
rect 7227 920 7347 2140
rect 7567 920 7687 2140
rect 7827 1620 7947 2820
rect 8167 1620 8287 2820
rect 7827 1600 8287 1620
rect 7827 1520 7847 1600
rect 8267 1520 8287 1600
rect 7827 1500 8287 1520
rect 8427 2240 8887 2260
rect 8427 2160 8447 2240
rect 8867 2160 8887 2240
rect 8427 2140 8887 2160
rect 8427 920 8547 2140
rect 8767 920 8887 2140
rect 9027 1620 9147 2820
rect 9367 1620 9487 2820
rect 14700 2660 14900 4980
rect 14600 2620 15000 2660
rect 13978 2328 14068 2338
rect 9027 1600 9487 1620
rect 9027 1520 9047 1600
rect 9467 1520 9487 1600
rect 9027 1500 9487 1520
rect 9627 2240 10087 2260
rect 9627 2160 9647 2240
rect 10067 2160 10087 2240
rect 9627 2140 10087 2160
rect 9627 920 9747 2140
rect 9967 920 10087 2140
rect 13978 2118 13988 2328
rect 14058 2118 14068 2328
rect 14600 2300 14640 2620
rect 14960 2300 15000 2620
rect 14600 2260 15000 2300
rect 13978 2108 14068 2118
rect 13520 1980 14460 2040
rect 10280 1950 14460 1980
rect 10180 1930 13620 1950
rect 10180 1850 10200 1930
rect 10260 1880 13620 1930
rect 10260 1850 10280 1880
rect 10180 1830 10280 1850
rect 13748 1788 14308 1848
rect 12810 1690 13180 1700
rect 12810 1610 12820 1690
rect 13170 1610 13180 1690
rect 12810 1600 13180 1610
rect 10970 1410 11730 1510
rect 10180 1240 10280 1260
rect 10180 1160 10200 1240
rect 10260 1230 10280 1240
rect 10970 1230 11070 1410
rect 10260 1160 11070 1230
rect 10180 1140 11070 1160
rect 10280 1130 11070 1140
rect 11630 1160 11730 1410
rect 12810 1440 13180 1450
rect 12810 1360 12820 1440
rect 13170 1360 13180 1440
rect 12810 1350 13180 1360
rect 13748 1408 13808 1788
rect 14248 1708 14308 1788
rect 13908 1698 14038 1708
rect 14238 1698 14318 1708
rect 13908 1638 13918 1698
rect 13978 1638 14158 1698
rect 13908 1628 14038 1638
rect 13908 1408 13988 1418
rect 13748 1348 13918 1408
rect 13978 1348 13988 1408
rect 14098 1408 14158 1638
rect 14238 1638 14248 1698
rect 14308 1638 14318 1698
rect 14238 1628 14318 1638
rect 14238 1410 14318 1418
rect 14400 1410 14460 1950
rect 14238 1408 14460 1410
rect 14098 1348 14248 1408
rect 14308 1350 14460 1408
rect 14308 1348 14318 1350
rect 13748 1160 13808 1348
rect 13908 1338 13988 1348
rect 14238 1338 14318 1348
rect 11630 1060 13830 1160
rect 15537 1142 15931 7602
rect 15537 1002 15577 1142
rect 15897 1002 15931 1142
rect 3427 900 10087 920
rect 2620 860 3187 880
rect 2620 840 2640 860
rect 1760 -7320 1820 -6680
rect 1920 -7320 1980 -6680
rect 2080 -7320 2140 -6680
rect 2300 -7320 2360 -6680
rect -1020 -7520 1520 -7320
rect 1400 -9060 1520 -7520
rect 1740 -9060 1840 -7320
rect 1900 -9060 2000 -7320
rect 2060 -9060 2160 -7320
rect 2240 -9060 2360 -7320
rect 2420 780 2640 840
rect 2740 780 3087 860
rect 3167 780 3187 860
rect 2420 760 3187 780
rect 3427 820 6047 900
rect 6467 820 7247 900
rect 7667 820 8447 900
rect 8867 820 9647 900
rect 10067 820 10087 900
rect 11070 920 11210 940
rect 11070 840 11090 920
rect 11190 840 11210 920
rect 11070 820 11210 840
rect 13978 928 14068 938
rect 3427 800 10087 820
rect 2420 -6680 2540 760
rect 3427 582 3587 800
rect 13978 718 13988 928
rect 14058 718 14068 928
rect 15537 912 15557 1002
rect 15917 912 15931 1002
rect 15537 902 15577 912
rect 15897 902 15931 912
rect 15537 863 15931 902
rect 16251 1142 16645 7602
rect 16251 1002 16291 1142
rect 16611 1002 16645 1142
rect 16251 912 16271 1002
rect 16631 912 16645 1002
rect 16251 902 16291 912
rect 16611 902 16645 912
rect 16251 863 16645 902
rect 16965 1142 17359 7602
rect 16965 1002 17005 1142
rect 17325 1002 17359 1142
rect 16965 912 16985 1002
rect 17345 912 17359 1002
rect 16965 902 17005 912
rect 17325 902 17359 912
rect 16965 863 17359 902
rect 17679 1142 18073 7602
rect 17679 1002 17719 1142
rect 18039 1002 18073 1142
rect 17679 912 17699 1002
rect 18059 912 18073 1002
rect 17679 902 17719 912
rect 18039 902 18073 912
rect 17679 863 18073 902
rect 18393 1142 18787 7602
rect 18393 1002 18433 1142
rect 18753 1002 18787 1142
rect 18393 912 18413 1002
rect 18773 912 18787 1002
rect 18393 902 18433 912
rect 18753 902 18787 912
rect 18393 863 18787 902
rect 19107 1142 19501 7602
rect 19107 1002 19147 1142
rect 19467 1002 19501 1142
rect 19107 912 19127 1002
rect 19487 912 19501 1002
rect 19107 902 19147 912
rect 19467 902 19501 912
rect 19107 863 19501 902
rect 19821 1142 20215 7602
rect 19821 1002 19861 1142
rect 20181 1002 20215 1142
rect 19821 912 19841 1002
rect 20201 912 20215 1002
rect 19821 902 19861 912
rect 20181 902 20215 912
rect 19821 863 20215 902
rect 20535 1142 20929 7602
rect 20535 1002 20575 1142
rect 20895 1002 20929 1142
rect 20535 912 20555 1002
rect 20915 912 20929 1002
rect 20535 902 20575 912
rect 20895 902 20929 912
rect 20535 863 20929 902
rect 21249 1142 21643 7602
rect 21249 1002 21289 1142
rect 21609 1002 21643 1142
rect 21249 912 21269 1002
rect 21629 912 21643 1002
rect 21249 902 21289 912
rect 21609 902 21643 912
rect 21249 863 21643 902
rect 21963 1142 22357 7602
rect 21963 1002 22003 1142
rect 22323 1002 22357 1142
rect 21963 912 21983 1002
rect 22343 912 22357 1002
rect 21963 902 22003 912
rect 22323 902 22357 912
rect 21963 863 22357 902
rect 22677 1142 23071 7602
rect 22677 1002 22717 1142
rect 23037 1002 23071 1142
rect 22677 912 22697 1002
rect 23057 912 23071 1002
rect 22677 902 22717 912
rect 23037 902 23071 912
rect 22677 863 23071 902
rect 23391 1142 23785 7602
rect 23391 1002 23431 1142
rect 23751 1002 23785 1142
rect 23391 912 23411 1002
rect 23771 912 23785 1002
rect 23391 902 23431 912
rect 23751 902 23785 912
rect 23391 863 23785 902
rect 24105 1142 24499 7602
rect 24105 1002 24145 1142
rect 24465 1002 24499 1142
rect 24105 912 24125 1002
rect 24485 912 24499 1002
rect 24105 902 24145 912
rect 24465 902 24499 912
rect 24105 863 24499 902
rect 24819 1142 25213 7602
rect 24819 1002 24859 1142
rect 25179 1002 25213 1142
rect 24819 912 24839 1002
rect 25199 912 25213 1002
rect 24819 902 24859 912
rect 25179 902 25213 912
rect 24819 863 25213 902
rect 25533 1142 25927 7602
rect 25533 1002 25573 1142
rect 25893 1002 25927 1142
rect 25533 912 25553 1002
rect 25913 912 25927 1002
rect 25533 902 25573 912
rect 25893 902 25927 912
rect 25533 863 25927 902
rect 26247 1142 26641 7602
rect 26247 1002 26287 1142
rect 26607 1002 26641 1142
rect 26247 912 26267 1002
rect 26627 912 26641 1002
rect 26247 902 26287 912
rect 26607 902 26641 912
rect 26247 863 26641 902
rect 26961 1142 27355 7602
rect 26961 1002 27001 1142
rect 27321 1002 27355 1142
rect 26961 912 26981 1002
rect 27341 912 27355 1002
rect 26961 902 27001 912
rect 27321 902 27355 912
rect 26961 863 27355 902
rect 27675 1142 28069 7602
rect 27675 1002 27715 1142
rect 28035 1002 28069 1142
rect 27675 912 27695 1002
rect 28055 912 28069 1002
rect 27675 902 27715 912
rect 28035 902 28069 912
rect 27675 863 28069 902
rect 28389 1142 28783 7602
rect 28389 1002 28429 1142
rect 28749 1002 28783 1142
rect 28389 912 28409 1002
rect 28769 912 28783 1002
rect 28389 902 28429 912
rect 28749 902 28783 912
rect 28389 863 28783 902
rect 29103 1142 29497 7602
rect 29103 1002 29143 1142
rect 29463 1002 29497 1142
rect 29103 912 29123 1002
rect 29483 912 29497 1002
rect 29103 902 29143 912
rect 29463 902 29497 912
rect 29103 863 29497 902
rect 29817 1142 30211 7602
rect 29817 1002 29857 1142
rect 30177 1002 30211 1142
rect 29817 912 29837 1002
rect 30197 912 30211 1002
rect 29817 902 29857 912
rect 30177 902 30211 912
rect 29817 863 30211 902
rect 30531 1142 30925 7602
rect 30531 1002 30571 1142
rect 30891 1002 30925 1142
rect 30531 912 30551 1002
rect 30911 912 30925 1002
rect 30531 902 30571 912
rect 30891 902 30925 912
rect 30531 863 30925 902
rect 31245 1142 31639 7602
rect 31245 1002 31285 1142
rect 31605 1002 31639 1142
rect 31245 912 31265 1002
rect 31625 912 31639 1002
rect 31245 902 31285 912
rect 31605 902 31639 912
rect 31245 863 31639 902
rect 31959 1142 32353 7602
rect 31959 1002 31999 1142
rect 32319 1002 32353 1142
rect 31959 912 31979 1002
rect 32339 912 32353 1002
rect 31959 902 31999 912
rect 32319 902 32353 912
rect 31959 863 32353 902
rect 32673 1142 33067 7602
rect 32673 1002 32713 1142
rect 33033 1002 33067 1142
rect 32673 912 32693 1002
rect 33053 912 33067 1002
rect 32673 902 32713 912
rect 33033 902 33067 912
rect 32673 863 33067 902
rect 33387 1142 33781 7602
rect 33387 1002 33427 1142
rect 33747 1002 33781 1142
rect 33387 912 33407 1002
rect 33767 912 33781 1002
rect 33387 902 33427 912
rect 33747 902 33781 912
rect 33387 863 33781 902
rect 34101 1142 34495 7602
rect 34101 1002 34141 1142
rect 34461 1002 34495 1142
rect 34101 912 34121 1002
rect 34481 912 34495 1002
rect 34101 902 34141 912
rect 34461 902 34495 912
rect 34101 863 34495 902
rect 34815 1142 35209 7602
rect 34815 1002 34855 1142
rect 35175 1002 35209 1142
rect 34815 912 34835 1002
rect 35195 912 35209 1002
rect 34815 902 34855 912
rect 35175 902 35209 912
rect 34815 863 35209 902
rect 35529 1142 35923 7602
rect 35529 1002 35569 1142
rect 35889 1002 35923 1142
rect 35529 912 35549 1002
rect 35909 912 35923 1002
rect 35529 902 35569 912
rect 35889 902 35923 912
rect 35529 863 35923 902
rect 36243 1142 36637 7602
rect 36243 1002 36283 1142
rect 36603 1002 36637 1142
rect 36243 912 36263 1002
rect 36623 912 36637 1002
rect 36243 902 36283 912
rect 36603 902 36637 912
rect 36243 863 36637 902
rect 36957 1142 37351 7602
rect 36957 1002 36997 1142
rect 37317 1002 37351 1142
rect 36957 912 36977 1002
rect 37337 912 37351 1002
rect 36957 902 36997 912
rect 37317 902 37351 912
rect 36957 863 37351 902
rect 37671 1142 38065 4462
rect 37671 1012 37711 1142
rect 38031 1022 38065 1142
rect 38385 1142 38779 2892
rect 40000 1950 40600 2000
rect 38031 1012 38071 1022
rect 37671 912 37691 1012
rect 38061 912 38071 1012
rect 37671 902 37711 912
rect 38031 902 38071 912
rect 38385 1012 38425 1142
rect 38745 1012 38779 1142
rect 38385 912 38395 1012
rect 38765 912 38779 1012
rect 38385 902 38425 912
rect 38745 902 38779 912
rect 37671 862 38065 902
rect 38385 862 38779 902
rect 39150 1900 40600 1950
rect 39150 1700 40100 1900
rect 40500 1700 40600 1900
rect 39150 1650 40600 1700
rect 13978 708 14068 718
rect 15548 793 15928 803
rect 15548 733 15558 793
rect 15918 733 15928 793
rect 15548 723 15928 733
rect 15548 589 15688 723
rect 15788 589 15928 723
rect 16262 793 16642 803
rect 16262 733 16272 793
rect 16632 733 16642 793
rect 16262 723 16642 733
rect 16262 589 16402 723
rect 16502 589 16642 723
rect 16976 793 17356 803
rect 16976 733 16986 793
rect 17346 733 17356 793
rect 16976 723 17356 733
rect 16976 589 17116 723
rect 17216 589 17356 723
rect 17690 793 18070 803
rect 17690 733 17700 793
rect 18060 733 18070 793
rect 17690 723 18070 733
rect 17690 589 17830 723
rect 17930 589 18070 723
rect 18404 793 18784 803
rect 18404 733 18414 793
rect 18774 733 18784 793
rect 18404 723 18784 733
rect 18404 589 18544 723
rect 18644 589 18784 723
rect 19118 793 19498 803
rect 19118 733 19128 793
rect 19488 733 19498 793
rect 19118 723 19498 733
rect 19118 589 19258 723
rect 19358 589 19498 723
rect 19832 793 20212 803
rect 19832 733 19842 793
rect 20202 733 20212 793
rect 19832 723 20212 733
rect 19832 589 19972 723
rect 20072 589 20212 723
rect 20546 793 20926 803
rect 20546 733 20556 793
rect 20916 733 20926 793
rect 20546 723 20926 733
rect 20546 589 20686 723
rect 20786 589 20926 723
rect 21260 793 21640 803
rect 21260 733 21270 793
rect 21630 733 21640 793
rect 21260 723 21640 733
rect 21260 589 21400 723
rect 21500 589 21640 723
rect 21974 793 22354 803
rect 21974 733 21984 793
rect 22344 733 22354 793
rect 21974 723 22354 733
rect 21974 589 22114 723
rect 22214 589 22354 723
rect 22688 793 23068 803
rect 22688 733 22698 793
rect 23058 733 23068 793
rect 22688 723 23068 733
rect 22688 589 22828 723
rect 22928 589 23068 723
rect 23402 793 23782 803
rect 23402 733 23412 793
rect 23772 733 23782 793
rect 23402 723 23782 733
rect 23402 589 23542 723
rect 23642 589 23782 723
rect 24116 793 24496 803
rect 24116 733 24126 793
rect 24486 733 24496 793
rect 24116 723 24496 733
rect 24116 589 24256 723
rect 24356 589 24496 723
rect 24830 793 25210 803
rect 24830 733 24840 793
rect 25200 733 25210 793
rect 24830 723 25210 733
rect 24830 589 24970 723
rect 25070 589 25210 723
rect 25544 793 25924 803
rect 25544 733 25554 793
rect 25914 733 25924 793
rect 25544 723 25924 733
rect 25544 589 25684 723
rect 25784 589 25924 723
rect 26258 793 26638 803
rect 26258 733 26268 793
rect 26628 733 26638 793
rect 26258 723 26638 733
rect 26258 589 26398 723
rect 26498 589 26638 723
rect 26972 793 27352 803
rect 26972 733 26982 793
rect 27342 733 27352 793
rect 26972 723 27352 733
rect 26972 589 27112 723
rect 27212 589 27352 723
rect 27686 793 28066 803
rect 27686 733 27696 793
rect 28056 733 28066 793
rect 27686 723 28066 733
rect 27686 589 27826 723
rect 27926 589 28066 723
rect 28400 793 28780 803
rect 28400 733 28410 793
rect 28770 733 28780 793
rect 28400 723 28780 733
rect 28400 589 28540 723
rect 28640 589 28780 723
rect 29114 793 29494 803
rect 29114 733 29124 793
rect 29484 733 29494 793
rect 29114 723 29494 733
rect 29114 589 29254 723
rect 29354 589 29494 723
rect 29828 793 30208 803
rect 29828 733 29838 793
rect 30198 733 30208 793
rect 29828 723 30208 733
rect 29828 589 29968 723
rect 30068 589 30208 723
rect 30542 793 30922 803
rect 30542 733 30552 793
rect 30912 733 30922 793
rect 30542 723 30922 733
rect 30542 589 30682 723
rect 30782 589 30922 723
rect 31256 793 31636 803
rect 31256 733 31266 793
rect 31626 733 31636 793
rect 31256 723 31636 733
rect 31256 589 31396 723
rect 31496 589 31636 723
rect 31970 793 32350 803
rect 31970 733 31980 793
rect 32340 733 32350 793
rect 31970 723 32350 733
rect 31970 589 32110 723
rect 32210 589 32350 723
rect 32684 793 33064 803
rect 32684 733 32694 793
rect 33054 733 33064 793
rect 32684 723 33064 733
rect 32684 589 32824 723
rect 32924 589 33064 723
rect 33398 793 33778 803
rect 33398 733 33408 793
rect 33768 733 33778 793
rect 33398 723 33778 733
rect 33398 589 33538 723
rect 33638 589 33778 723
rect 34112 793 34492 803
rect 34112 733 34122 793
rect 34482 733 34492 793
rect 34112 723 34492 733
rect 34112 589 34252 723
rect 34352 589 34492 723
rect 34826 793 35206 803
rect 34826 733 34836 793
rect 35196 733 35206 793
rect 34826 723 35206 733
rect 34826 589 34966 723
rect 35066 589 35206 723
rect 35540 793 35920 803
rect 35540 733 35550 793
rect 35910 733 35920 793
rect 35540 723 35920 733
rect 35540 589 35680 723
rect 35780 589 35920 723
rect 36254 793 36634 803
rect 36254 733 36264 793
rect 36624 733 36634 793
rect 36254 723 36634 733
rect 36254 589 36394 723
rect 36494 589 36634 723
rect 36968 793 37348 803
rect 36968 733 36978 793
rect 37338 733 37348 793
rect 36968 723 37348 733
rect 36968 589 37108 723
rect 37208 589 37348 723
rect 37678 789 38058 799
rect 37678 689 37698 789
rect 38048 689 38058 789
rect 37678 679 38058 689
rect 37678 589 37818 679
rect 37918 589 38058 679
rect 38388 789 38778 799
rect 38388 729 38408 789
rect 38768 729 38778 789
rect 38388 719 38778 729
rect 38388 589 38528 719
rect 38628 589 38768 719
rect 39150 589 39450 1650
rect 40000 1600 40600 1650
rect 39900 1040 40320 1050
rect 39900 980 39920 1040
rect 40300 980 40530 1040
rect 39900 970 40320 980
rect 39900 880 40320 890
rect 39900 820 39920 880
rect 40300 820 40530 880
rect 39900 810 40320 820
rect 39900 710 40320 720
rect 39900 650 39920 710
rect 40300 650 40530 710
rect 39900 640 40320 650
rect 3427 562 3838 582
rect 3427 442 3768 562
rect 3427 342 3587 442
rect 3758 342 3768 442
rect 3427 202 3768 342
rect 3828 202 3838 562
rect 3427 -136 3587 202
rect 3758 192 3838 202
rect 3901 575 5931 585
rect 14428 580 39450 589
rect 3901 545 3951 575
rect 4051 545 5931 575
rect 3901 225 3941 545
rect 4181 225 5931 545
rect 3901 205 3951 225
rect 4051 205 5931 225
rect 3901 191 5931 205
rect 14380 289 39450 580
rect 39900 540 40320 550
rect 39900 480 39920 540
rect 40300 480 40530 540
rect 39900 470 40320 480
rect 39900 370 40320 380
rect 39900 310 39920 370
rect 40300 310 40530 370
rect 39900 300 40320 310
rect 14380 120 14700 289
rect 9880 100 14700 120
rect 3427 -156 3838 -136
rect 3427 -276 3728 -156
rect 3427 -376 3587 -276
rect 3718 -376 3728 -276
rect 3427 -506 3728 -376
rect 3828 -506 3838 -156
rect 3427 -516 3838 -506
rect 3901 -149 7501 -129
rect 3901 -169 3951 -149
rect 4051 -169 7501 -149
rect 3901 -489 3941 -169
rect 4181 -489 7501 -169
rect 9880 -180 9900 100
rect 14380 -180 14700 100
rect 15548 139 15688 289
rect 15788 139 15928 289
rect 15548 129 15928 139
rect 15548 69 15558 129
rect 15918 69 15928 129
rect 15548 59 15928 69
rect 16262 139 16402 289
rect 16502 139 16642 289
rect 16262 129 16642 139
rect 16262 69 16272 129
rect 16632 69 16642 129
rect 16262 59 16642 69
rect 16976 139 17116 289
rect 17216 139 17356 289
rect 16976 129 17356 139
rect 16976 69 16986 129
rect 17346 69 17356 129
rect 16976 59 17356 69
rect 17690 139 17830 289
rect 17930 139 18070 289
rect 17690 129 18070 139
rect 17690 69 17700 129
rect 18060 69 18070 129
rect 17690 59 18070 69
rect 18404 139 18544 289
rect 18644 139 18784 289
rect 18404 129 18784 139
rect 18404 69 18414 129
rect 18774 69 18784 129
rect 18404 59 18784 69
rect 19118 139 19258 289
rect 19358 139 19498 289
rect 19118 129 19498 139
rect 19118 69 19128 129
rect 19488 69 19498 129
rect 19118 59 19498 69
rect 19832 139 19972 289
rect 20072 139 20212 289
rect 19832 129 20212 139
rect 19832 69 19842 129
rect 20202 69 20212 129
rect 19832 59 20212 69
rect 20546 139 20686 289
rect 20786 139 20926 289
rect 20546 129 20926 139
rect 20546 69 20556 129
rect 20916 69 20926 129
rect 20546 59 20926 69
rect 21260 139 21400 289
rect 21500 139 21640 289
rect 21260 129 21640 139
rect 21260 69 21270 129
rect 21630 69 21640 129
rect 21260 59 21640 69
rect 21974 139 22114 289
rect 22214 139 22354 289
rect 21974 129 22354 139
rect 21974 69 21984 129
rect 22344 69 22354 129
rect 21974 59 22354 69
rect 22688 139 22828 289
rect 22928 139 23068 289
rect 22688 129 23068 139
rect 22688 69 22698 129
rect 23058 69 23068 129
rect 22688 59 23068 69
rect 23402 139 23542 289
rect 23642 139 23782 289
rect 23402 129 23782 139
rect 23402 69 23412 129
rect 23772 69 23782 129
rect 23402 59 23782 69
rect 24116 139 24256 289
rect 24356 139 24496 289
rect 24116 129 24496 139
rect 24116 69 24126 129
rect 24486 69 24496 129
rect 24116 59 24496 69
rect 24830 139 24970 289
rect 25070 139 25210 289
rect 24830 129 25210 139
rect 24830 69 24840 129
rect 25200 69 25210 129
rect 24830 59 25210 69
rect 25544 139 25684 289
rect 25784 139 25924 289
rect 25544 129 25924 139
rect 25544 69 25554 129
rect 25914 69 25924 129
rect 25544 59 25924 69
rect 26258 139 26398 289
rect 26498 139 26638 289
rect 26258 129 26638 139
rect 26258 69 26268 129
rect 26628 69 26638 129
rect 26258 59 26638 69
rect 26972 139 27112 289
rect 27212 139 27352 289
rect 26972 129 27352 139
rect 26972 69 26982 129
rect 27342 69 27352 129
rect 26972 59 27352 69
rect 27686 139 27826 289
rect 27926 139 28066 289
rect 27686 129 28066 139
rect 27686 69 27696 129
rect 28056 69 28066 129
rect 27686 59 28066 69
rect 28400 139 28540 289
rect 28640 139 28780 289
rect 28400 129 28780 139
rect 28400 69 28410 129
rect 28770 69 28780 129
rect 28400 59 28780 69
rect 29114 139 29254 289
rect 29354 139 29494 289
rect 29114 129 29494 139
rect 29114 69 29124 129
rect 29484 69 29494 129
rect 29114 59 29494 69
rect 29828 139 29968 289
rect 30068 139 30208 289
rect 29828 129 30208 139
rect 29828 69 29838 129
rect 30198 69 30208 129
rect 29828 59 30208 69
rect 30542 139 30682 289
rect 30782 139 30922 289
rect 30542 129 30922 139
rect 30542 69 30552 129
rect 30912 69 30922 129
rect 30542 59 30922 69
rect 31256 139 31396 289
rect 31496 139 31636 289
rect 31256 129 31636 139
rect 31256 69 31266 129
rect 31626 69 31636 129
rect 31256 59 31636 69
rect 31970 139 32110 289
rect 32210 139 32350 289
rect 31970 129 32350 139
rect 31970 69 31980 129
rect 32340 69 32350 129
rect 31970 59 32350 69
rect 32684 139 32824 289
rect 32924 139 33064 289
rect 32684 129 33064 139
rect 32684 69 32694 129
rect 33054 69 33064 129
rect 32684 59 33064 69
rect 33398 139 33538 289
rect 33638 139 33778 289
rect 33398 129 33778 139
rect 33398 69 33408 129
rect 33768 69 33778 129
rect 33398 59 33778 69
rect 34112 139 34252 289
rect 34352 139 34492 289
rect 34112 129 34492 139
rect 34112 69 34122 129
rect 34482 69 34492 129
rect 34112 59 34492 69
rect 34826 139 34966 289
rect 35066 139 35206 289
rect 34826 129 35206 139
rect 34826 69 34836 129
rect 35196 69 35206 129
rect 34826 59 35206 69
rect 35540 139 35680 289
rect 35780 139 35920 289
rect 35540 129 35920 139
rect 35540 69 35550 129
rect 35910 69 35920 129
rect 35540 59 35920 69
rect 36254 139 36394 289
rect 36494 139 36634 289
rect 36254 129 36634 139
rect 36254 69 36264 129
rect 36624 69 36634 129
rect 36254 59 36634 69
rect 36968 139 37108 289
rect 37208 139 37348 289
rect 36968 129 37348 139
rect 36968 69 36978 129
rect 37338 69 37348 129
rect 36968 59 37348 69
rect 37682 139 37822 289
rect 37922 139 38062 289
rect 37682 129 38062 139
rect 37682 69 37692 129
rect 38052 69 38062 129
rect 37682 59 38062 69
rect 38396 139 38536 289
rect 38636 139 38776 289
rect 38396 129 38776 139
rect 38396 69 38406 129
rect 38766 69 38776 129
rect 38396 59 38776 69
rect 9880 -200 14700 -180
rect 15537 -40 15931 -1
rect 15537 -50 15577 -40
rect 15897 -50 15931 -40
rect 15537 -140 15557 -50
rect 15917 -140 15931 -50
rect 3427 -700 3587 -516
rect 3901 -519 3951 -489
rect 4051 -519 7501 -489
rect 3901 -523 7501 -519
rect 10020 -420 10180 -400
rect 10860 -420 10980 -200
rect 3941 -529 4061 -523
rect 10020 -740 10040 -420
rect 10160 -740 10180 -420
rect 10480 -440 10640 -420
rect 10480 -540 10500 -440
rect 10020 -760 10180 -740
rect 10240 -650 10500 -540
rect 10240 -980 10300 -650
rect 10480 -700 10500 -650
rect 10620 -700 10640 -440
rect 10480 -720 10640 -700
rect 10860 -740 10880 -420
rect 10960 -740 10980 -420
rect 10860 -760 10980 -740
rect 15537 -280 15577 -140
rect 15897 -280 15931 -140
rect 11200 -790 11300 -780
rect 10870 -830 11060 -820
rect 10870 -900 10880 -830
rect 11050 -900 11060 -830
rect 11200 -870 11210 -790
rect 11290 -870 11300 -790
rect 11200 -880 11300 -870
rect 10870 -910 11060 -900
rect 2780 -1100 10300 -980
rect 14600 -1040 15000 -1000
rect 11380 -1090 11480 -1080
rect 2600 -4120 2720 -4100
rect 2600 -4280 2620 -4120
rect 2700 -4280 2720 -4120
rect 2600 -6680 2720 -4280
rect 2780 -6680 2900 -1100
rect 10480 -1130 10640 -1120
rect 10480 -1240 10490 -1130
rect 10630 -1240 10640 -1130
rect 11380 -1170 11390 -1090
rect 11470 -1170 11480 -1090
rect 11380 -1180 11480 -1170
rect 10480 -1250 10640 -1240
rect 3000 -1251 10640 -1250
rect 2960 -1370 10640 -1251
rect 14600 -1360 14640 -1040
rect 14960 -1360 15000 -1040
rect 2960 -6680 3080 -1370
rect 14600 -1400 15000 -1360
rect 11310 -1490 11410 -1480
rect 11310 -1570 11320 -1490
rect 11400 -1570 11410 -1490
rect 11310 -1580 11410 -1570
rect 14700 -1700 14900 -1400
rect 7700 -1900 14900 -1700
rect 5802 -2100 7202 -2000
rect 5802 -2700 5902 -2100
rect 7102 -2700 7202 -2100
rect 5802 -2800 7202 -2700
rect 7700 -5580 7900 -1900
rect 9002 -2100 10402 -2000
rect 9002 -2700 9102 -2100
rect 10302 -2700 10402 -2100
rect 9002 -2800 10402 -2700
rect 12002 -2100 14802 -2000
rect 12002 -2700 12102 -2100
rect 14702 -2700 14802 -2100
rect 10302 -2940 10622 -2920
rect 9022 -4100 10202 -3800
rect 10302 -3860 10322 -2940
rect 10602 -3860 10622 -2940
rect 10302 -3880 10622 -3860
rect 10702 -3152 11602 -3052
rect 10702 -3552 10802 -3152
rect 11502 -3552 11602 -3152
rect 10702 -3812 11602 -3552
rect 10702 -4032 10872 -3812
rect 11082 -4032 11602 -3812
rect 10702 -4052 11602 -4032
rect 10302 -4100 11602 -4052
rect 9022 -5300 9202 -4100
rect 9902 -4300 11602 -4100
rect 9022 -5360 9032 -5300
rect 9192 -5360 9202 -5300
rect 9022 -5370 9202 -5360
rect 8100 -5420 8300 -5400
rect 8100 -5580 8120 -5420
rect 8280 -5580 8300 -5420
rect 7289 -5594 7943 -5580
rect 5170 -5640 5320 -5620
rect 5170 -6030 5190 -5640
rect 5300 -6030 5320 -5640
rect 5170 -6050 5320 -6030
rect 5400 -5640 5550 -5620
rect 5400 -6030 5420 -5640
rect 5530 -5975 5550 -5640
rect 7289 -5650 7295 -5594
rect 7361 -5650 7487 -5594
rect 7553 -5650 7679 -5594
rect 7745 -5650 7871 -5594
rect 7937 -5650 7943 -5594
rect 7289 -5662 7943 -5650
rect 8057 -5594 8711 -5580
rect 8057 -5650 8063 -5594
rect 8129 -5650 8255 -5594
rect 8321 -5650 8447 -5594
rect 8513 -5650 8639 -5594
rect 8705 -5650 8711 -5594
rect 8057 -5662 8711 -5650
rect 5530 -6030 5734 -5975
rect 5400 -6049 5734 -6030
rect 5400 -6050 5550 -6049
rect 5220 -6310 5290 -6050
rect 5000 -6340 5600 -6310
rect 5000 -6420 5030 -6340
rect 5570 -6420 5600 -6340
rect 5000 -6580 5020 -6420
rect 5580 -6580 5600 -6420
rect 5660 -6495 5734 -6049
rect 6261 -6495 9740 -6464
rect 5660 -6504 9807 -6495
rect 5660 -6560 6202 -6504
rect 6258 -6560 9743 -6504
rect 9799 -6560 9807 -6504
rect 5660 -6569 9807 -6560
rect 2420 -7320 2480 -6680
rect 2620 -7320 2700 -6680
rect 2800 -7320 2880 -6680
rect 2980 -7320 3060 -6680
rect 5000 -6700 5600 -6580
rect 6000 -6650 6130 -6640
rect 2420 -9060 2540 -7320
rect 2600 -9060 2720 -7320
rect 2780 -9060 2900 -7320
rect 2960 -9060 3080 -7320
rect 5000 -9400 5800 -6700
rect 6000 -6740 6010 -6650
rect 6120 -6740 6130 -6650
rect 6000 -6750 6130 -6740
rect 6402 -9300 9802 -9200
rect 6402 -9800 6502 -9300
rect 9702 -9800 9802 -9300
rect 10302 -9652 11602 -4300
rect 12002 -9600 14802 -2700
rect 15537 -6740 15931 -280
rect 16251 -40 16645 -1
rect 16251 -50 16291 -40
rect 16611 -50 16645 -40
rect 16251 -140 16271 -50
rect 16631 -140 16645 -50
rect 16251 -280 16291 -140
rect 16611 -280 16645 -140
rect 16251 -6740 16645 -280
rect 16965 -40 17359 -1
rect 16965 -50 17005 -40
rect 17325 -50 17359 -40
rect 16965 -140 16985 -50
rect 17345 -140 17359 -50
rect 16965 -280 17005 -140
rect 17325 -280 17359 -140
rect 16965 -6740 17359 -280
rect 17679 -40 18073 -1
rect 17679 -50 17719 -40
rect 18039 -50 18073 -40
rect 17679 -140 17699 -50
rect 18059 -140 18073 -50
rect 17679 -280 17719 -140
rect 18039 -280 18073 -140
rect 17679 -6740 18073 -280
rect 18393 -40 18787 -1
rect 18393 -50 18433 -40
rect 18753 -50 18787 -40
rect 18393 -140 18413 -50
rect 18773 -140 18787 -50
rect 18393 -280 18433 -140
rect 18753 -280 18787 -140
rect 18393 -6740 18787 -280
rect 19107 -40 19501 -1
rect 19107 -50 19147 -40
rect 19467 -50 19501 -40
rect 19107 -140 19127 -50
rect 19487 -140 19501 -50
rect 19107 -280 19147 -140
rect 19467 -280 19501 -140
rect 19107 -6740 19501 -280
rect 19821 -40 20215 -1
rect 19821 -50 19861 -40
rect 20181 -50 20215 -40
rect 19821 -140 19841 -50
rect 20201 -140 20215 -50
rect 19821 -280 19861 -140
rect 20181 -280 20215 -140
rect 19821 -6740 20215 -280
rect 20535 -40 20929 -1
rect 20535 -50 20575 -40
rect 20895 -50 20929 -40
rect 20535 -140 20555 -50
rect 20915 -140 20929 -50
rect 20535 -280 20575 -140
rect 20895 -280 20929 -140
rect 20535 -6740 20929 -280
rect 21249 -40 21643 -1
rect 21249 -50 21289 -40
rect 21609 -50 21643 -40
rect 21249 -140 21269 -50
rect 21629 -140 21643 -50
rect 21249 -280 21289 -140
rect 21609 -280 21643 -140
rect 21249 -6740 21643 -280
rect 21963 -40 22357 -1
rect 21963 -50 22003 -40
rect 22323 -50 22357 -40
rect 21963 -140 21983 -50
rect 22343 -140 22357 -50
rect 21963 -280 22003 -140
rect 22323 -280 22357 -140
rect 21963 -6740 22357 -280
rect 22677 -40 23071 -1
rect 22677 -50 22717 -40
rect 23037 -50 23071 -40
rect 22677 -140 22697 -50
rect 23057 -140 23071 -50
rect 22677 -280 22717 -140
rect 23037 -280 23071 -140
rect 22677 -6740 23071 -280
rect 23391 -40 23785 -1
rect 23391 -50 23431 -40
rect 23751 -50 23785 -40
rect 23391 -140 23411 -50
rect 23771 -140 23785 -50
rect 23391 -280 23431 -140
rect 23751 -280 23785 -140
rect 23391 -6740 23785 -280
rect 24105 -40 24499 -1
rect 24105 -50 24145 -40
rect 24465 -50 24499 -40
rect 24105 -140 24125 -50
rect 24485 -140 24499 -50
rect 24105 -280 24145 -140
rect 24465 -280 24499 -140
rect 24105 -6740 24499 -280
rect 24819 -40 25213 -1
rect 24819 -50 24859 -40
rect 25179 -50 25213 -40
rect 24819 -140 24839 -50
rect 25199 -140 25213 -50
rect 24819 -280 24859 -140
rect 25179 -280 25213 -140
rect 24819 -6740 25213 -280
rect 25533 -40 25927 -1
rect 25533 -50 25573 -40
rect 25893 -50 25927 -40
rect 25533 -140 25553 -50
rect 25913 -140 25927 -50
rect 25533 -280 25573 -140
rect 25893 -280 25927 -140
rect 25533 -6740 25927 -280
rect 26247 -40 26641 -1
rect 26247 -50 26287 -40
rect 26607 -50 26641 -40
rect 26247 -140 26267 -50
rect 26627 -140 26641 -50
rect 26247 -280 26287 -140
rect 26607 -280 26641 -140
rect 26247 -6740 26641 -280
rect 26961 -40 27355 -1
rect 26961 -50 27001 -40
rect 27321 -50 27355 -40
rect 26961 -140 26981 -50
rect 27341 -140 27355 -50
rect 26961 -280 27001 -140
rect 27321 -280 27355 -140
rect 26961 -6740 27355 -280
rect 27675 -40 28069 -1
rect 27675 -50 27715 -40
rect 28035 -50 28069 -40
rect 27675 -140 27695 -50
rect 28055 -140 28069 -50
rect 27675 -280 27715 -140
rect 28035 -280 28069 -140
rect 27675 -6740 28069 -280
rect 28389 -40 28783 -1
rect 28389 -50 28429 -40
rect 28749 -50 28783 -40
rect 28389 -140 28409 -50
rect 28769 -140 28783 -50
rect 28389 -280 28429 -140
rect 28749 -280 28783 -140
rect 28389 -6740 28783 -280
rect 29103 -40 29497 -1
rect 29103 -50 29143 -40
rect 29463 -50 29497 -40
rect 29103 -140 29123 -50
rect 29483 -140 29497 -50
rect 29103 -280 29143 -140
rect 29463 -280 29497 -140
rect 29103 -6740 29497 -280
rect 29817 -40 30211 -1
rect 29817 -50 29857 -40
rect 30177 -50 30211 -40
rect 29817 -140 29837 -50
rect 30197 -140 30211 -50
rect 29817 -280 29857 -140
rect 30177 -280 30211 -140
rect 29817 -6740 30211 -280
rect 30531 -40 30925 -1
rect 30531 -50 30571 -40
rect 30891 -50 30925 -40
rect 30531 -140 30551 -50
rect 30911 -140 30925 -50
rect 30531 -280 30571 -140
rect 30891 -280 30925 -140
rect 30531 -6740 30925 -280
rect 31245 -40 31639 -1
rect 31245 -50 31285 -40
rect 31605 -50 31639 -40
rect 31245 -140 31265 -50
rect 31625 -140 31639 -50
rect 31245 -280 31285 -140
rect 31605 -280 31639 -140
rect 31245 -6740 31639 -280
rect 31959 -40 32353 -1
rect 31959 -50 31999 -40
rect 32319 -50 32353 -40
rect 31959 -140 31979 -50
rect 32339 -140 32353 -50
rect 31959 -280 31999 -140
rect 32319 -280 32353 -140
rect 31959 -6740 32353 -280
rect 32673 -40 33067 -1
rect 32673 -50 32713 -40
rect 33033 -50 33067 -40
rect 32673 -140 32693 -50
rect 33053 -140 33067 -50
rect 32673 -280 32713 -140
rect 33033 -280 33067 -140
rect 32673 -6740 33067 -280
rect 33387 -40 33781 -1
rect 33387 -50 33427 -40
rect 33747 -50 33781 -40
rect 33387 -140 33407 -50
rect 33767 -140 33781 -50
rect 33387 -280 33427 -140
rect 33747 -280 33781 -140
rect 33387 -6740 33781 -280
rect 34101 -40 34495 -1
rect 34101 -50 34141 -40
rect 34461 -50 34495 -40
rect 34101 -140 34121 -50
rect 34481 -140 34495 -50
rect 34101 -280 34141 -140
rect 34461 -280 34495 -140
rect 34101 -6740 34495 -280
rect 34815 -40 35209 -1
rect 34815 -50 34855 -40
rect 35175 -50 35209 -40
rect 34815 -140 34835 -50
rect 35195 -140 35209 -50
rect 34815 -280 34855 -140
rect 35175 -280 35209 -140
rect 34815 -6740 35209 -280
rect 35529 -40 35923 -1
rect 35529 -50 35569 -40
rect 35889 -50 35923 -40
rect 35529 -140 35549 -50
rect 35909 -140 35923 -50
rect 35529 -280 35569 -140
rect 35889 -280 35923 -140
rect 35529 -6740 35923 -280
rect 36243 -40 36637 -1
rect 36243 -50 36283 -40
rect 36603 -50 36637 -40
rect 36243 -140 36263 -50
rect 36623 -140 36637 -50
rect 36243 -280 36283 -140
rect 36603 -280 36637 -140
rect 36243 -6740 36637 -280
rect 36957 -40 37351 -1
rect 36957 -50 36997 -40
rect 37317 -50 37351 -40
rect 36957 -140 36977 -50
rect 37337 -140 37351 -50
rect 36957 -280 36997 -140
rect 37317 -280 37351 -140
rect 36957 -6740 37351 -280
rect 37671 -40 38065 -1
rect 37671 -50 37711 -40
rect 38031 -50 38065 -40
rect 37671 -140 37691 -50
rect 38051 -140 38065 -50
rect 37671 -280 37711 -140
rect 38031 -280 38065 -140
rect 37671 -6740 38065 -280
rect 38385 -40 38779 -1
rect 38385 -50 38425 -40
rect 38745 -50 38779 -40
rect 38385 -140 38405 -50
rect 38765 -140 38779 -50
rect 38385 -280 38425 -140
rect 38745 -280 38779 -140
rect 38385 -6740 38779 -280
rect 39150 -850 39450 289
rect 39900 210 40320 220
rect 39900 150 39920 210
rect 40300 150 40530 210
rect 39900 140 40320 150
rect 39900 50 40320 60
rect 39900 -10 39920 50
rect 40300 -10 40530 50
rect 39900 -20 40320 -10
rect 39900 -120 40320 -110
rect 39900 -180 39920 -120
rect 40300 -180 40530 -120
rect 39900 -190 40320 -180
rect 40000 -850 40600 -800
rect 39150 -900 40600 -850
rect 39150 -1100 40100 -900
rect 40500 -1100 40600 -900
rect 39150 -1150 40600 -1100
rect 40000 -1200 40600 -1150
rect 6402 -9900 9802 -9800
<< via3 >>
rect 6502 12700 9702 13200
rect 6010 10050 6120 10140
rect 5020 9820 5580 9980
rect 5030 9740 5570 9820
rect 5902 5500 7102 6100
rect 10322 6340 10402 7260
rect 10402 6340 10522 7260
rect 10802 6552 11502 6952
rect 9102 5500 10302 6100
rect 12102 5500 14702 6100
rect 11030 4830 11110 4910
rect 11190 4830 11270 4910
rect 11330 4680 11410 4760
rect -360 4280 -200 4440
rect 3228 3995 3358 4315
rect 3358 3995 3458 4315
rect 3458 3995 3468 4315
rect 4374 3995 4384 4315
rect 4384 3995 4484 4315
rect 4484 3995 4614 4315
rect 8620 3960 9260 4260
rect 9260 3960 9580 4260
rect 3228 3281 3358 3601
rect 3358 3281 3458 3601
rect 3458 3281 3468 3601
rect 4374 3281 4384 3601
rect 4384 3281 4484 3601
rect 4484 3281 4614 3601
rect 3247 2380 3627 2600
rect 3247 1820 3627 2040
rect -360 -180 -200 -20
rect 4407 1040 4787 1280
rect 13988 2118 14048 2328
rect 14048 2118 14058 2328
rect 14640 2300 14960 2620
rect 12820 1360 13170 1440
rect 15577 1002 15897 1142
rect 11090 840 11190 920
rect 13988 718 14058 928
rect 15577 912 15897 1002
rect 15577 902 15897 912
rect 16291 1002 16611 1142
rect 16291 912 16611 1002
rect 16291 902 16611 912
rect 17005 1002 17325 1142
rect 17005 912 17325 1002
rect 17005 902 17325 912
rect 17719 1002 18039 1142
rect 17719 912 18039 1002
rect 17719 902 18039 912
rect 18433 1002 18753 1142
rect 18433 912 18753 1002
rect 18433 902 18753 912
rect 19147 1002 19467 1142
rect 19147 912 19467 1002
rect 19147 902 19467 912
rect 19861 1002 20181 1142
rect 19861 912 20181 1002
rect 19861 902 20181 912
rect 20575 1002 20895 1142
rect 20575 912 20895 1002
rect 20575 902 20895 912
rect 21289 1002 21609 1142
rect 21289 912 21609 1002
rect 21289 902 21609 912
rect 22003 1002 22323 1142
rect 22003 912 22323 1002
rect 22003 902 22323 912
rect 22717 1002 23037 1142
rect 22717 912 23037 1002
rect 22717 902 23037 912
rect 23431 1002 23751 1142
rect 23431 912 23751 1002
rect 23431 902 23751 912
rect 24145 1002 24465 1142
rect 24145 912 24465 1002
rect 24145 902 24465 912
rect 24859 1002 25179 1142
rect 24859 912 25179 1002
rect 24859 902 25179 912
rect 25573 1002 25893 1142
rect 25573 912 25893 1002
rect 25573 902 25893 912
rect 26287 1002 26607 1142
rect 26287 912 26607 1002
rect 26287 902 26607 912
rect 27001 1002 27321 1142
rect 27001 912 27321 1002
rect 27001 902 27321 912
rect 27715 1002 28035 1142
rect 27715 912 28035 1002
rect 27715 902 28035 912
rect 28429 1002 28749 1142
rect 28429 912 28749 1002
rect 28429 902 28749 912
rect 29143 1002 29463 1142
rect 29143 912 29463 1002
rect 29143 902 29463 912
rect 29857 1002 30177 1142
rect 29857 912 30177 1002
rect 29857 902 30177 912
rect 30571 1002 30891 1142
rect 30571 912 30891 1002
rect 30571 902 30891 912
rect 31285 1002 31605 1142
rect 31285 912 31605 1002
rect 31285 902 31605 912
rect 31999 1002 32319 1142
rect 31999 912 32319 1002
rect 31999 902 32319 912
rect 32713 1002 33033 1142
rect 32713 912 33033 1002
rect 32713 902 33033 912
rect 33427 1002 33747 1142
rect 33427 912 33747 1002
rect 33427 902 33747 912
rect 34141 1002 34461 1142
rect 34141 912 34461 1002
rect 34141 902 34461 912
rect 34855 1002 35175 1142
rect 34855 912 35175 1002
rect 34855 902 35175 912
rect 35569 1002 35889 1142
rect 35569 912 35889 1002
rect 35569 902 35889 912
rect 36283 1002 36603 1142
rect 36283 912 36603 1002
rect 36283 902 36603 912
rect 36997 1002 37317 1142
rect 36997 912 37317 1002
rect 36997 902 37317 912
rect 37711 1012 38031 1142
rect 37711 912 38031 1012
rect 37711 902 38031 912
rect 38425 1012 38745 1142
rect 38425 912 38745 1012
rect 38425 902 38745 912
rect 40100 1700 40500 1900
rect 3941 225 3951 545
rect 3951 225 4051 545
rect 4051 225 4181 545
rect 3941 -489 3951 -169
rect 3951 -489 4051 -169
rect 4051 -489 4181 -169
rect 12020 -180 12780 100
rect 15577 -50 15897 -40
rect 15577 -140 15897 -50
rect 10040 -740 10160 -420
rect 10500 -700 10620 -440
rect 15577 -280 15897 -140
rect 10880 -890 10950 -830
rect 10950 -890 11050 -830
rect 10880 -900 11050 -890
rect 11210 -870 11290 -790
rect 2620 -4280 2700 -4120
rect 10490 -1240 10630 -1130
rect 11390 -1170 11470 -1090
rect 14640 -1360 14960 -1040
rect 11320 -1570 11400 -1490
rect 5902 -2700 7102 -2100
rect 9102 -2700 10302 -2100
rect 12102 -2700 14702 -2100
rect 10322 -3860 10402 -2940
rect 10402 -3860 10522 -2940
rect 10802 -3552 11502 -3152
rect 8120 -5580 8280 -5420
rect 5030 -6420 5570 -6340
rect 5020 -6580 5580 -6420
rect 6010 -6740 6120 -6650
rect 6502 -9800 9702 -9300
rect 16291 -50 16611 -40
rect 16291 -140 16611 -50
rect 16291 -280 16611 -140
rect 17005 -50 17325 -40
rect 17005 -140 17325 -50
rect 17005 -280 17325 -140
rect 17719 -50 18039 -40
rect 17719 -140 18039 -50
rect 17719 -280 18039 -140
rect 18433 -50 18753 -40
rect 18433 -140 18753 -50
rect 18433 -280 18753 -140
rect 19147 -50 19467 -40
rect 19147 -140 19467 -50
rect 19147 -280 19467 -140
rect 19861 -50 20181 -40
rect 19861 -140 20181 -50
rect 19861 -280 20181 -140
rect 20575 -50 20895 -40
rect 20575 -140 20895 -50
rect 20575 -280 20895 -140
rect 21289 -50 21609 -40
rect 21289 -140 21609 -50
rect 21289 -280 21609 -140
rect 22003 -50 22323 -40
rect 22003 -140 22323 -50
rect 22003 -280 22323 -140
rect 22717 -50 23037 -40
rect 22717 -140 23037 -50
rect 22717 -280 23037 -140
rect 23431 -50 23751 -40
rect 23431 -140 23751 -50
rect 23431 -280 23751 -140
rect 24145 -50 24465 -40
rect 24145 -140 24465 -50
rect 24145 -280 24465 -140
rect 24859 -50 25179 -40
rect 24859 -140 25179 -50
rect 24859 -280 25179 -140
rect 25573 -50 25893 -40
rect 25573 -140 25893 -50
rect 25573 -280 25893 -140
rect 26287 -50 26607 -40
rect 26287 -140 26607 -50
rect 26287 -280 26607 -140
rect 27001 -50 27321 -40
rect 27001 -140 27321 -50
rect 27001 -280 27321 -140
rect 27715 -50 28035 -40
rect 27715 -140 28035 -50
rect 27715 -280 28035 -140
rect 28429 -50 28749 -40
rect 28429 -140 28749 -50
rect 28429 -280 28749 -140
rect 29143 -50 29463 -40
rect 29143 -140 29463 -50
rect 29143 -280 29463 -140
rect 29857 -50 30177 -40
rect 29857 -140 30177 -50
rect 29857 -280 30177 -140
rect 30571 -50 30891 -40
rect 30571 -140 30891 -50
rect 30571 -280 30891 -140
rect 31285 -50 31605 -40
rect 31285 -140 31605 -50
rect 31285 -280 31605 -140
rect 31999 -50 32319 -40
rect 31999 -140 32319 -50
rect 31999 -280 32319 -140
rect 32713 -50 33033 -40
rect 32713 -140 33033 -50
rect 32713 -280 33033 -140
rect 33427 -50 33747 -40
rect 33427 -140 33747 -50
rect 33427 -280 33747 -140
rect 34141 -50 34461 -40
rect 34141 -140 34461 -50
rect 34141 -280 34461 -140
rect 34855 -50 35175 -40
rect 34855 -140 35175 -50
rect 34855 -280 35175 -140
rect 35569 -50 35889 -40
rect 35569 -140 35889 -50
rect 35569 -280 35889 -140
rect 36283 -50 36603 -40
rect 36283 -140 36603 -50
rect 36283 -280 36603 -140
rect 36997 -50 37317 -40
rect 36997 -140 37317 -50
rect 36997 -280 37317 -140
rect 37711 -50 38031 -40
rect 37711 -140 38031 -50
rect 37711 -280 38031 -140
rect 38425 -50 38745 -40
rect 38425 -140 38745 -50
rect 38425 -280 38745 -140
rect 40100 -1100 40500 -900
<< mimcap >>
rect 10402 12912 11502 12952
rect 5030 12750 5770 12770
rect 5030 10150 5050 12750
rect 5750 10150 5770 12750
rect 5030 10130 5770 10150
rect 10402 7592 10442 12912
rect 11462 7592 11502 12912
rect 10402 7552 11502 7592
rect 12102 12860 14702 12900
rect 12102 6740 12142 12860
rect 14662 6740 14702 12860
rect 12102 6700 14702 6740
rect 15577 7542 15897 7562
rect 1518 4295 3088 4315
rect 1518 4015 1538 4295
rect 3068 4015 3088 4295
rect 1518 3995 3088 4015
rect 4754 4295 6324 4315
rect 4754 4015 4774 4295
rect 6304 4015 6324 4295
rect 4754 3995 6324 4015
rect -52 3581 3088 3601
rect -52 3301 -32 3581
rect 3068 3301 3088 3581
rect -52 3281 3088 3301
rect 4754 3581 7894 3601
rect 4754 3301 4774 3581
rect 7874 3301 7894 3581
rect 4754 3281 7894 3301
rect 15577 1302 15597 7542
rect 15877 1302 15897 7542
rect 15577 1282 15897 1302
rect 16291 7542 16611 7562
rect 16291 1302 16311 7542
rect 16591 1302 16611 7542
rect 16291 1282 16611 1302
rect 17005 7542 17325 7562
rect 17005 1302 17025 7542
rect 17305 1302 17325 7542
rect 17005 1282 17325 1302
rect 17719 7542 18039 7562
rect 17719 1302 17739 7542
rect 18019 1302 18039 7542
rect 17719 1282 18039 1302
rect 18433 7542 18753 7562
rect 18433 1302 18453 7542
rect 18733 1302 18753 7542
rect 18433 1282 18753 1302
rect 19147 7542 19467 7562
rect 19147 1302 19167 7542
rect 19447 1302 19467 7542
rect 19147 1282 19467 1302
rect 19861 7542 20181 7562
rect 19861 1302 19881 7542
rect 20161 1302 20181 7542
rect 19861 1282 20181 1302
rect 20575 7542 20895 7562
rect 20575 1302 20595 7542
rect 20875 1302 20895 7542
rect 20575 1282 20895 1302
rect 21289 7542 21609 7562
rect 21289 1302 21309 7542
rect 21589 1302 21609 7542
rect 21289 1282 21609 1302
rect 22003 7542 22323 7562
rect 22003 1302 22023 7542
rect 22303 1302 22323 7542
rect 22003 1282 22323 1302
rect 22717 7542 23037 7562
rect 22717 1302 22737 7542
rect 23017 1302 23037 7542
rect 22717 1282 23037 1302
rect 23431 7542 23751 7562
rect 23431 1302 23451 7542
rect 23731 1302 23751 7542
rect 23431 1282 23751 1302
rect 24145 7542 24465 7562
rect 24145 1302 24165 7542
rect 24445 1302 24465 7542
rect 24145 1282 24465 1302
rect 24859 7542 25179 7562
rect 24859 1302 24879 7542
rect 25159 1302 25179 7542
rect 24859 1282 25179 1302
rect 25573 7542 25893 7562
rect 25573 1302 25593 7542
rect 25873 1302 25893 7542
rect 25573 1282 25893 1302
rect 26287 7542 26607 7562
rect 26287 1302 26307 7542
rect 26587 1302 26607 7542
rect 26287 1282 26607 1302
rect 27001 7542 27321 7562
rect 27001 1302 27021 7542
rect 27301 1302 27321 7542
rect 27001 1282 27321 1302
rect 27715 7542 28035 7562
rect 27715 1302 27735 7542
rect 28015 1302 28035 7542
rect 27715 1282 28035 1302
rect 28429 7542 28749 7562
rect 28429 1302 28449 7542
rect 28729 1302 28749 7542
rect 28429 1282 28749 1302
rect 29143 7542 29463 7562
rect 29143 1302 29163 7542
rect 29443 1302 29463 7542
rect 29143 1282 29463 1302
rect 29857 7542 30177 7562
rect 29857 1302 29877 7542
rect 30157 1302 30177 7542
rect 29857 1282 30177 1302
rect 30571 7542 30891 7562
rect 30571 1302 30591 7542
rect 30871 1302 30891 7542
rect 30571 1282 30891 1302
rect 31285 7542 31605 7562
rect 31285 1302 31305 7542
rect 31585 1302 31605 7542
rect 31285 1282 31605 1302
rect 31999 7542 32319 7562
rect 31999 1302 32019 7542
rect 32299 1302 32319 7542
rect 31999 1282 32319 1302
rect 32713 7542 33033 7562
rect 32713 1302 32733 7542
rect 33013 1302 33033 7542
rect 32713 1282 33033 1302
rect 33427 7542 33747 7562
rect 33427 1302 33447 7542
rect 33727 1302 33747 7542
rect 33427 1282 33747 1302
rect 34141 7542 34461 7562
rect 34141 1302 34161 7542
rect 34441 1302 34461 7542
rect 34141 1282 34461 1302
rect 34855 7542 35175 7562
rect 34855 1302 34875 7542
rect 35155 1302 35175 7542
rect 34855 1282 35175 1302
rect 35569 7542 35889 7562
rect 35569 1302 35589 7542
rect 35869 1302 35889 7542
rect 35569 1282 35889 1302
rect 36283 7542 36603 7562
rect 36283 1302 36303 7542
rect 36583 1302 36603 7542
rect 36283 1282 36603 1302
rect 36997 7542 37317 7562
rect 36997 1302 37017 7542
rect 37297 1302 37317 7542
rect 36997 1282 37317 1302
rect 37711 4402 38031 4422
rect 37711 1302 37731 4402
rect 38011 1302 38031 4402
rect 37711 1282 38031 1302
rect 38425 2832 38745 2852
rect 38425 1302 38445 2832
rect 38725 1302 38745 2832
rect 38425 1282 38745 1302
rect 4321 525 5891 545
rect 4321 245 4341 525
rect 5871 245 5891 525
rect 4321 225 5891 245
rect 4321 -189 7461 -169
rect 4321 -469 4341 -189
rect 7441 -469 7461 -189
rect 4321 -489 7461 -469
rect 15577 -440 15897 -420
rect 12102 -3340 14702 -3300
rect 10402 -4192 11502 -4152
rect 5030 -6750 5770 -6730
rect 5030 -9350 5050 -6750
rect 5750 -9350 5770 -6750
rect 5030 -9370 5770 -9350
rect 10402 -9512 10442 -4192
rect 11462 -9512 11502 -4192
rect 12102 -9460 12142 -3340
rect 14662 -9460 14702 -3340
rect 15577 -6680 15597 -440
rect 15877 -6680 15897 -440
rect 15577 -6700 15897 -6680
rect 16291 -440 16611 -420
rect 16291 -6680 16311 -440
rect 16591 -6680 16611 -440
rect 16291 -6700 16611 -6680
rect 17005 -440 17325 -420
rect 17005 -6680 17025 -440
rect 17305 -6680 17325 -440
rect 17005 -6700 17325 -6680
rect 17719 -440 18039 -420
rect 17719 -6680 17739 -440
rect 18019 -6680 18039 -440
rect 17719 -6700 18039 -6680
rect 18433 -440 18753 -420
rect 18433 -6680 18453 -440
rect 18733 -6680 18753 -440
rect 18433 -6700 18753 -6680
rect 19147 -440 19467 -420
rect 19147 -6680 19167 -440
rect 19447 -6680 19467 -440
rect 19147 -6700 19467 -6680
rect 19861 -440 20181 -420
rect 19861 -6680 19881 -440
rect 20161 -6680 20181 -440
rect 19861 -6700 20181 -6680
rect 20575 -440 20895 -420
rect 20575 -6680 20595 -440
rect 20875 -6680 20895 -440
rect 20575 -6700 20895 -6680
rect 21289 -440 21609 -420
rect 21289 -6680 21309 -440
rect 21589 -6680 21609 -440
rect 21289 -6700 21609 -6680
rect 22003 -440 22323 -420
rect 22003 -6680 22023 -440
rect 22303 -6680 22323 -440
rect 22003 -6700 22323 -6680
rect 22717 -440 23037 -420
rect 22717 -6680 22737 -440
rect 23017 -6680 23037 -440
rect 22717 -6700 23037 -6680
rect 23431 -440 23751 -420
rect 23431 -6680 23451 -440
rect 23731 -6680 23751 -440
rect 23431 -6700 23751 -6680
rect 24145 -440 24465 -420
rect 24145 -6680 24165 -440
rect 24445 -6680 24465 -440
rect 24145 -6700 24465 -6680
rect 24859 -440 25179 -420
rect 24859 -6680 24879 -440
rect 25159 -6680 25179 -440
rect 24859 -6700 25179 -6680
rect 25573 -440 25893 -420
rect 25573 -6680 25593 -440
rect 25873 -6680 25893 -440
rect 25573 -6700 25893 -6680
rect 26287 -440 26607 -420
rect 26287 -6680 26307 -440
rect 26587 -6680 26607 -440
rect 26287 -6700 26607 -6680
rect 27001 -440 27321 -420
rect 27001 -6680 27021 -440
rect 27301 -6680 27321 -440
rect 27001 -6700 27321 -6680
rect 27715 -440 28035 -420
rect 27715 -6680 27735 -440
rect 28015 -6680 28035 -440
rect 27715 -6700 28035 -6680
rect 28429 -440 28749 -420
rect 28429 -6680 28449 -440
rect 28729 -6680 28749 -440
rect 28429 -6700 28749 -6680
rect 29143 -440 29463 -420
rect 29143 -6680 29163 -440
rect 29443 -6680 29463 -440
rect 29143 -6700 29463 -6680
rect 29857 -440 30177 -420
rect 29857 -6680 29877 -440
rect 30157 -6680 30177 -440
rect 29857 -6700 30177 -6680
rect 30571 -440 30891 -420
rect 30571 -6680 30591 -440
rect 30871 -6680 30891 -440
rect 30571 -6700 30891 -6680
rect 31285 -440 31605 -420
rect 31285 -6680 31305 -440
rect 31585 -6680 31605 -440
rect 31285 -6700 31605 -6680
rect 31999 -440 32319 -420
rect 31999 -6680 32019 -440
rect 32299 -6680 32319 -440
rect 31999 -6700 32319 -6680
rect 32713 -440 33033 -420
rect 32713 -6680 32733 -440
rect 33013 -6680 33033 -440
rect 32713 -6700 33033 -6680
rect 33427 -440 33747 -420
rect 33427 -6680 33447 -440
rect 33727 -6680 33747 -440
rect 33427 -6700 33747 -6680
rect 34141 -440 34461 -420
rect 34141 -6680 34161 -440
rect 34441 -6680 34461 -440
rect 34141 -6700 34461 -6680
rect 34855 -440 35175 -420
rect 34855 -6680 34875 -440
rect 35155 -6680 35175 -440
rect 34855 -6700 35175 -6680
rect 35569 -440 35889 -420
rect 35569 -6680 35589 -440
rect 35869 -6680 35889 -440
rect 35569 -6700 35889 -6680
rect 36283 -440 36603 -420
rect 36283 -6680 36303 -440
rect 36583 -6680 36603 -440
rect 36283 -6700 36603 -6680
rect 36997 -440 37317 -420
rect 36997 -6680 37017 -440
rect 37297 -6680 37317 -440
rect 36997 -6700 37317 -6680
rect 37711 -440 38031 -420
rect 37711 -6680 37731 -440
rect 38011 -6680 38031 -440
rect 37711 -6700 38031 -6680
rect 38425 -440 38745 -420
rect 38425 -6680 38445 -440
rect 38725 -6680 38745 -440
rect 38425 -6700 38745 -6680
rect 12102 -9500 14702 -9460
rect 10402 -9552 11502 -9512
<< mimcapcontact >>
rect 5050 10150 5750 12750
rect 10442 7592 11462 12912
rect 12142 6740 14662 12860
rect 1538 4015 3068 4295
rect 4774 4015 6304 4295
rect -32 3301 3068 3581
rect 4774 3301 7874 3581
rect 15597 1302 15877 7542
rect 16311 1302 16591 7542
rect 17025 1302 17305 7542
rect 17739 1302 18019 7542
rect 18453 1302 18733 7542
rect 19167 1302 19447 7542
rect 19881 1302 20161 7542
rect 20595 1302 20875 7542
rect 21309 1302 21589 7542
rect 22023 1302 22303 7542
rect 22737 1302 23017 7542
rect 23451 1302 23731 7542
rect 24165 1302 24445 7542
rect 24879 1302 25159 7542
rect 25593 1302 25873 7542
rect 26307 1302 26587 7542
rect 27021 1302 27301 7542
rect 27735 1302 28015 7542
rect 28449 1302 28729 7542
rect 29163 1302 29443 7542
rect 29877 1302 30157 7542
rect 30591 1302 30871 7542
rect 31305 1302 31585 7542
rect 32019 1302 32299 7542
rect 32733 1302 33013 7542
rect 33447 1302 33727 7542
rect 34161 1302 34441 7542
rect 34875 1302 35155 7542
rect 35589 1302 35869 7542
rect 36303 1302 36583 7542
rect 37017 1302 37297 7542
rect 37731 1302 38011 4402
rect 38445 1302 38725 2832
rect 4341 245 5871 525
rect 4341 -469 7441 -189
rect 5050 -9350 5750 -6750
rect 10442 -9512 11462 -4192
rect 12142 -9460 14662 -3340
rect 15597 -6680 15877 -440
rect 16311 -6680 16591 -440
rect 17025 -6680 17305 -440
rect 17739 -6680 18019 -440
rect 18453 -6680 18733 -440
rect 19167 -6680 19447 -440
rect 19881 -6680 20161 -440
rect 20595 -6680 20875 -440
rect 21309 -6680 21589 -440
rect 22023 -6680 22303 -440
rect 22737 -6680 23017 -440
rect 23451 -6680 23731 -440
rect 24165 -6680 24445 -440
rect 24879 -6680 25159 -440
rect 25593 -6680 25873 -440
rect 26307 -6680 26587 -440
rect 27021 -6680 27301 -440
rect 27735 -6680 28015 -440
rect 28449 -6680 28729 -440
rect 29163 -6680 29443 -440
rect 29877 -6680 30157 -440
rect 30591 -6680 30871 -440
rect 31305 -6680 31585 -440
rect 32019 -6680 32299 -440
rect 32733 -6680 33013 -440
rect 33447 -6680 33727 -440
rect 34161 -6680 34441 -440
rect 34875 -6680 35155 -440
rect 35589 -6680 35869 -440
rect 36303 -6680 36583 -440
rect 37017 -6680 37297 -440
rect 37731 -6680 38011 -440
rect 38445 -6680 38725 -440
<< metal4 >>
rect 3400 13800 4600 14000
rect 3400 13200 3600 13800
rect 4400 13700 44200 13800
rect 4400 13300 43100 13700
rect 4400 13200 9802 13300
rect 3400 13000 4600 13200
rect 5000 12750 5800 12800
rect 5000 10460 5050 12750
rect -360 10300 5050 10460
rect -360 4460 -200 10300
rect 5000 10150 5050 10300
rect 5750 10160 5800 12750
rect 6402 12700 6502 13200
rect 9702 12700 9802 13200
rect 6402 12600 9802 12700
rect 10302 12912 11602 13052
rect 12202 13000 43100 13300
rect 5750 10150 6130 10160
rect 5000 10140 6130 10150
rect 5000 10100 6010 10140
rect 0 9800 100 10100
rect 200 9800 300 10100
rect 400 9800 500 10100
rect 600 9900 900 10100
rect 6000 10050 6010 10100
rect 6120 10050 6130 10140
rect 6000 10040 6130 10050
rect 600 9800 700 9900
rect 800 9800 900 9900
rect 5000 9980 5600 10000
rect 5000 9820 5020 9980
rect 5000 9740 5030 9820
rect 5580 9820 5600 9980
rect 5570 9740 5600 9820
rect 5000 9710 5600 9740
rect 10302 7592 10442 12912
rect 11462 7592 11602 12912
rect 10302 7452 11602 7592
rect 12002 12860 43100 13000
rect 10302 7260 10542 7452
rect 10302 6340 10322 7260
rect 10522 6340 10542 7260
rect 10702 6952 11602 7052
rect 10702 6552 10802 6952
rect 11502 6552 11602 6952
rect 12002 6740 12142 12860
rect 14662 12600 43100 12860
rect 44100 12600 44200 13700
rect 14662 12500 44200 12600
rect 14662 6740 14802 12500
rect 12002 6600 14802 6740
rect 15537 7542 15931 7602
rect 10702 6452 11602 6552
rect 10302 6320 10542 6340
rect 10303 6200 10542 6320
rect 5802 6100 10542 6200
rect 5802 5500 5902 6100
rect 7102 5500 9102 6100
rect 10302 5900 10542 6100
rect 12002 6100 14802 6200
rect 12002 5900 12102 6100
rect 10302 5500 12102 5900
rect 14702 5500 14802 6100
rect 5802 5400 14802 5500
rect 11020 4910 11120 4920
rect 11020 4830 11030 4910
rect 11110 4830 11120 4910
rect 11020 4820 11120 4830
rect 11060 4460 11120 4820
rect 11180 4910 11280 4920
rect 11180 4830 11190 4910
rect 11270 4830 11280 4910
rect 11180 4820 11280 4830
rect 11180 4580 11240 4820
rect 11320 4760 11990 4770
rect 11320 4680 11330 4760
rect 11410 4680 11990 4760
rect 11320 4670 11990 4680
rect 11180 4520 11620 4580
rect -380 4440 -180 4460
rect -380 4280 -360 4440
rect -200 4280 -180 4440
rect 11060 4400 11490 4460
rect 1478 4345 3128 4355
rect -380 4260 -180 4280
rect 1468 4295 3128 4345
rect 1468 4015 1538 4295
rect 3068 4015 3128 4295
rect 1468 3965 3128 4015
rect 1478 3961 3128 3965
rect 3188 4315 3508 4355
rect 3188 3995 3228 4315
rect 3468 3995 3508 4315
rect 3188 3961 3508 3995
rect 4334 4315 4654 4355
rect 4334 3995 4374 4315
rect 4614 3995 4654 4315
rect 4334 3961 4654 3995
rect 4714 4345 6364 4355
rect 4714 4295 6374 4345
rect 4714 4015 4774 4295
rect 6304 4015 6374 4295
rect 4714 3965 6374 4015
rect 8600 4260 9600 4280
rect 4714 3961 6364 3965
rect 2707 3641 2907 3961
rect 4847 3641 5047 3961
rect 8600 3960 8620 4260
rect 9580 3960 9600 4260
rect 8600 3940 9600 3960
rect -92 3631 3128 3641
rect -102 3581 3128 3631
rect -102 3301 -32 3581
rect 3068 3301 3128 3581
rect -102 3251 3128 3301
rect -92 3247 3128 3251
rect 3188 3601 3508 3641
rect 3188 3281 3228 3601
rect 3468 3281 3508 3601
rect 3188 3247 3508 3281
rect 4334 3601 4654 3641
rect 4334 3281 4374 3601
rect 4614 3281 4654 3601
rect 4334 3247 4654 3281
rect 4714 3631 7934 3641
rect 4714 3581 7944 3631
rect 4714 3301 4774 3581
rect 7874 3301 7944 3581
rect 4714 3251 7944 3301
rect 4714 3247 7934 3251
rect 2707 2080 2907 3247
rect 4847 2640 5047 3247
rect 3207 2600 5047 2640
rect 3207 2380 3247 2600
rect 3627 2440 5047 2600
rect 3627 2380 3707 2440
rect 3207 2340 3707 2380
rect 2707 2040 3707 2080
rect 2707 1880 3247 2040
rect 3207 1820 3247 1880
rect 3627 1820 3707 2040
rect 3207 1780 3707 1820
rect 4387 1280 4807 1300
rect 4387 1040 4407 1280
rect 4787 1040 4807 1280
rect 4387 1020 4807 1040
rect 4527 585 4727 1020
rect 10500 920 11210 940
rect 10500 840 11090 920
rect 11190 840 11210 920
rect 10500 820 11210 840
rect 3901 545 4221 585
rect 3901 225 3941 545
rect 4181 225 4221 545
rect 3901 191 4221 225
rect 4281 575 5931 585
rect 4281 525 5941 575
rect 4281 245 4341 525
rect 5871 245 5941 525
rect 4281 195 5941 245
rect 4281 191 5931 195
rect -380 -20 -180 0
rect -380 -180 -360 -20
rect -200 -180 -180 -20
rect 4527 -129 4727 191
rect -380 -200 -180 -180
rect 3901 -169 4221 -129
rect -360 -6920 -200 -200
rect 3901 -489 3941 -169
rect 4181 -489 4221 -169
rect 3901 -523 4221 -489
rect 4281 -139 7501 -129
rect 4281 -189 7511 -139
rect 4281 -469 4341 -189
rect 7441 -469 7511 -189
rect 4281 -519 7511 -469
rect 9900 -420 10180 -400
rect 10500 -420 10620 820
rect 11430 680 11490 4400
rect 11240 620 11490 680
rect 4281 -523 7501 -519
rect 9900 -740 9920 -420
rect 10160 -740 10180 -420
rect 10480 -440 10640 -420
rect 10480 -700 10500 -440
rect 10620 -700 10640 -440
rect 10480 -720 10640 -700
rect 9900 -760 10180 -740
rect 11240 -780 11300 620
rect 11560 560 11620 4520
rect 11200 -790 11300 -780
rect 11200 -820 11210 -790
rect 10870 -830 11210 -820
rect 10870 -900 10880 -830
rect 11050 -870 11210 -830
rect 11290 -870 11300 -790
rect 11050 -880 11300 -870
rect 11420 500 11620 560
rect 11890 1450 11990 4670
rect 14600 2620 15000 2660
rect 13978 2328 14068 2338
rect 13978 2118 13988 2328
rect 14058 2228 14068 2328
rect 14600 2300 14640 2620
rect 14960 2300 15000 2620
rect 14600 2229 15000 2300
rect 15537 2229 15597 7542
rect 14598 2228 15597 2229
rect 14058 2118 15597 2228
rect 13978 2108 15597 2118
rect 14458 1629 15597 2108
rect 11890 1440 13180 1450
rect 11890 1360 12820 1440
rect 13170 1360 13180 1440
rect 11890 1350 13180 1360
rect 11050 -900 11060 -880
rect 10870 -910 11060 -900
rect 11420 -1080 11480 500
rect 11890 370 11990 1350
rect 14458 938 15198 1629
rect 15537 1302 15597 1629
rect 15877 2229 15931 7542
rect 16251 7542 16645 7602
rect 16251 2229 16311 7542
rect 15877 1629 16311 2229
rect 15877 1302 15931 1629
rect 15537 1242 15931 1302
rect 16251 1302 16311 1629
rect 16591 2229 16645 7542
rect 16965 7542 17359 7602
rect 16965 2229 17025 7542
rect 16591 1629 17025 2229
rect 16591 1302 16645 1629
rect 16251 1242 16645 1302
rect 16965 1302 17025 1629
rect 17305 2229 17359 7542
rect 17679 7542 18073 7602
rect 17679 2229 17739 7542
rect 17305 1629 17739 2229
rect 17305 1302 17359 1629
rect 16965 1242 17359 1302
rect 17679 1302 17739 1629
rect 18019 2229 18073 7542
rect 18393 7542 18787 7602
rect 18393 2229 18453 7542
rect 18019 1629 18453 2229
rect 18019 1302 18073 1629
rect 17679 1242 18073 1302
rect 18393 1302 18453 1629
rect 18733 2229 18787 7542
rect 19107 7542 19501 7602
rect 19107 2229 19167 7542
rect 18733 1629 19167 2229
rect 18733 1302 18787 1629
rect 18393 1242 18787 1302
rect 19107 1302 19167 1629
rect 19447 2229 19501 7542
rect 19821 7542 20215 7602
rect 19821 2229 19881 7542
rect 19447 1629 19881 2229
rect 19447 1302 19501 1629
rect 19107 1242 19501 1302
rect 19821 1302 19881 1629
rect 20161 2229 20215 7542
rect 20535 7542 20929 7602
rect 20535 2229 20595 7542
rect 20161 1629 20595 2229
rect 20161 1302 20215 1629
rect 19821 1242 20215 1302
rect 20535 1302 20595 1629
rect 20875 2229 20929 7542
rect 21249 7542 21643 7602
rect 21249 2229 21309 7542
rect 20875 1629 21309 2229
rect 20875 1302 20929 1629
rect 20535 1242 20929 1302
rect 21249 1302 21309 1629
rect 21589 2229 21643 7542
rect 21963 7542 22357 7602
rect 21963 2229 22023 7542
rect 21589 1629 22023 2229
rect 21589 1302 21643 1629
rect 21249 1242 21643 1302
rect 21963 1302 22023 1629
rect 22303 2229 22357 7542
rect 22677 7542 23071 7602
rect 22677 2229 22737 7542
rect 22303 1629 22737 2229
rect 22303 1302 22357 1629
rect 21963 1242 22357 1302
rect 22677 1302 22737 1629
rect 23017 2229 23071 7542
rect 23391 7542 23785 7602
rect 23391 2229 23451 7542
rect 23017 1629 23451 2229
rect 23017 1302 23071 1629
rect 22677 1242 23071 1302
rect 23391 1302 23451 1629
rect 23731 2229 23785 7542
rect 24105 7542 24499 7602
rect 24105 2229 24165 7542
rect 23731 1629 24165 2229
rect 23731 1302 23785 1629
rect 23391 1242 23785 1302
rect 24105 1302 24165 1629
rect 24445 2229 24499 7542
rect 24819 7542 25213 7602
rect 24819 2229 24879 7542
rect 24445 1629 24879 2229
rect 24445 1302 24499 1629
rect 24105 1242 24499 1302
rect 24819 1302 24879 1629
rect 25159 2229 25213 7542
rect 25533 7542 25927 7602
rect 25533 2229 25593 7542
rect 25159 1629 25593 2229
rect 25159 1302 25213 1629
rect 24819 1242 25213 1302
rect 25533 1302 25593 1629
rect 25873 2229 25927 7542
rect 26247 7542 26641 7602
rect 26247 2229 26307 7542
rect 25873 1629 26307 2229
rect 25873 1302 25927 1629
rect 25533 1242 25927 1302
rect 26247 1302 26307 1629
rect 26587 2229 26641 7542
rect 26961 7542 27355 7602
rect 26961 2229 27021 7542
rect 26587 1629 27021 2229
rect 26587 1302 26641 1629
rect 26247 1242 26641 1302
rect 26961 1302 27021 1629
rect 27301 2229 27355 7542
rect 27675 7542 28069 7602
rect 27675 2229 27735 7542
rect 27301 1629 27735 2229
rect 27301 1302 27355 1629
rect 26961 1242 27355 1302
rect 27675 1302 27735 1629
rect 28015 2229 28069 7542
rect 28389 7542 28783 7602
rect 28389 2229 28449 7542
rect 28015 1629 28449 2229
rect 28015 1302 28069 1629
rect 27675 1242 28069 1302
rect 28389 1302 28449 1629
rect 28729 2229 28783 7542
rect 29103 7542 29497 7602
rect 29103 2229 29163 7542
rect 28729 1629 29163 2229
rect 28729 1302 28783 1629
rect 28389 1242 28783 1302
rect 29103 1302 29163 1629
rect 29443 2229 29497 7542
rect 29817 7542 30211 7602
rect 29817 2229 29877 7542
rect 29443 1629 29877 2229
rect 29443 1302 29497 1629
rect 29103 1242 29497 1302
rect 29817 1302 29877 1629
rect 30157 2229 30211 7542
rect 30531 7542 30925 7602
rect 30531 2229 30591 7542
rect 30157 1629 30591 2229
rect 30157 1302 30211 1629
rect 29817 1242 30211 1302
rect 30531 1302 30591 1629
rect 30871 2229 30925 7542
rect 31245 7542 31639 7602
rect 31245 2229 31305 7542
rect 30871 1629 31305 2229
rect 30871 1302 30925 1629
rect 30531 1242 30925 1302
rect 31245 1302 31305 1629
rect 31585 2229 31639 7542
rect 31959 7542 32353 7602
rect 31959 2229 32019 7542
rect 31585 1629 32019 2229
rect 31585 1302 31639 1629
rect 31245 1242 31639 1302
rect 31959 1302 32019 1629
rect 32299 2229 32353 7542
rect 32673 7542 33067 7602
rect 32673 2229 32733 7542
rect 32299 1629 32733 2229
rect 32299 1302 32353 1629
rect 31959 1242 32353 1302
rect 32673 1302 32733 1629
rect 33013 2229 33067 7542
rect 33387 7542 33781 7602
rect 33387 2229 33447 7542
rect 33013 1629 33447 2229
rect 33013 1302 33067 1629
rect 32673 1242 33067 1302
rect 33387 1302 33447 1629
rect 33727 2229 33781 7542
rect 34101 7542 34495 7602
rect 34101 2229 34161 7542
rect 33727 1629 34161 2229
rect 33727 1302 33781 1629
rect 33387 1242 33781 1302
rect 34101 1302 34161 1629
rect 34441 2229 34495 7542
rect 34815 7542 35209 7602
rect 34815 2229 34875 7542
rect 34441 1629 34875 2229
rect 34441 1302 34495 1629
rect 34101 1242 34495 1302
rect 34815 1302 34875 1629
rect 35155 2229 35209 7542
rect 35529 7542 35923 7602
rect 35529 2229 35589 7542
rect 35155 1629 35589 2229
rect 35155 1302 35209 1629
rect 34815 1242 35209 1302
rect 35529 1302 35589 1629
rect 35869 2229 35923 7542
rect 36243 7542 36637 7602
rect 36243 2229 36303 7542
rect 35869 1629 36303 2229
rect 35869 1302 35923 1629
rect 35529 1242 35923 1302
rect 36243 1302 36303 1629
rect 36583 2229 36637 7542
rect 36957 7542 37351 7602
rect 36957 2229 37017 7542
rect 36583 1629 37017 2229
rect 36583 1302 36637 1629
rect 36243 1242 36637 1302
rect 36957 1302 37017 1629
rect 37297 2229 37351 7542
rect 37681 4462 38061 4472
rect 37671 4402 38065 4462
rect 37671 2229 37731 4402
rect 37297 1629 37731 2229
rect 37297 1302 37351 1629
rect 36957 1242 37351 1302
rect 37671 1302 37731 1629
rect 38011 2229 38065 4402
rect 38395 2892 38775 2902
rect 38385 2832 38779 2892
rect 38385 2229 38445 2832
rect 38011 1629 38445 2229
rect 38011 1302 38065 1629
rect 37671 1242 38065 1302
rect 38385 1302 38445 1629
rect 38725 1302 38779 2832
rect 40000 2100 40600 2200
rect 40000 1700 40100 2100
rect 40500 1700 40600 2100
rect 40000 1600 40600 1700
rect 38385 1242 38779 1302
rect 13978 928 15198 938
rect 13978 718 13988 928
rect 14058 818 15198 928
rect 15537 1142 15931 1182
rect 15537 902 15577 1142
rect 15897 902 15931 1142
rect 15537 863 15931 902
rect 16251 1142 16645 1182
rect 16251 902 16291 1142
rect 16611 902 16645 1142
rect 16251 863 16645 902
rect 16965 1142 17359 1182
rect 16965 902 17005 1142
rect 17325 902 17359 1142
rect 16965 863 17359 902
rect 17679 1142 18073 1182
rect 17679 902 17719 1142
rect 18039 902 18073 1142
rect 17679 863 18073 902
rect 18393 1142 18787 1182
rect 18393 902 18433 1142
rect 18753 902 18787 1142
rect 18393 863 18787 902
rect 19107 1142 19501 1182
rect 19107 902 19147 1142
rect 19467 902 19501 1142
rect 19107 863 19501 902
rect 19821 1142 20215 1182
rect 19821 902 19861 1142
rect 20181 902 20215 1142
rect 19821 863 20215 902
rect 20535 1142 20929 1182
rect 20535 902 20575 1142
rect 20895 902 20929 1142
rect 20535 863 20929 902
rect 21249 1142 21643 1182
rect 21249 902 21289 1142
rect 21609 902 21643 1142
rect 21249 863 21643 902
rect 21963 1142 22357 1182
rect 21963 902 22003 1142
rect 22323 902 22357 1142
rect 21963 863 22357 902
rect 22677 1142 23071 1182
rect 22677 902 22717 1142
rect 23037 902 23071 1142
rect 22677 863 23071 902
rect 23391 1142 23785 1182
rect 23391 902 23431 1142
rect 23751 902 23785 1142
rect 23391 863 23785 902
rect 24105 1142 24499 1182
rect 24105 902 24145 1142
rect 24465 902 24499 1142
rect 24105 863 24499 902
rect 24819 1142 25213 1182
rect 24819 902 24859 1142
rect 25179 902 25213 1142
rect 24819 863 25213 902
rect 25533 1142 25927 1182
rect 25533 902 25573 1142
rect 25893 902 25927 1142
rect 25533 863 25927 902
rect 26247 1142 26641 1182
rect 26247 902 26287 1142
rect 26607 902 26641 1142
rect 26247 863 26641 902
rect 26961 1142 27355 1182
rect 26961 902 27001 1142
rect 27321 902 27355 1142
rect 26961 863 27355 902
rect 27675 1142 28069 1182
rect 27675 902 27715 1142
rect 28035 902 28069 1142
rect 27675 863 28069 902
rect 28389 1142 28783 1182
rect 28389 902 28429 1142
rect 28749 902 28783 1142
rect 28389 863 28783 902
rect 29103 1142 29497 1182
rect 29103 902 29143 1142
rect 29463 902 29497 1142
rect 29103 863 29497 902
rect 29817 1142 30211 1182
rect 29817 902 29857 1142
rect 30177 902 30211 1142
rect 29817 863 30211 902
rect 30531 1142 30925 1182
rect 30531 902 30571 1142
rect 30891 902 30925 1142
rect 30531 863 30925 902
rect 31245 1142 31639 1182
rect 31245 902 31285 1142
rect 31605 902 31639 1142
rect 31245 863 31639 902
rect 31959 1142 32353 1182
rect 31959 902 31999 1142
rect 32319 902 32353 1142
rect 31959 863 32353 902
rect 32673 1142 33067 1182
rect 32673 902 32713 1142
rect 33033 902 33067 1142
rect 32673 863 33067 902
rect 33387 1142 33781 1182
rect 33387 902 33427 1142
rect 33747 902 33781 1142
rect 33387 863 33781 902
rect 34101 1142 34495 1182
rect 34101 902 34141 1142
rect 34461 902 34495 1142
rect 34101 863 34495 902
rect 34815 1142 35209 1182
rect 34815 902 34855 1142
rect 35175 902 35209 1142
rect 34815 863 35209 902
rect 35529 1142 35923 1182
rect 35529 902 35569 1142
rect 35889 902 35923 1142
rect 35529 863 35923 902
rect 36243 1142 36637 1182
rect 36243 902 36283 1142
rect 36603 902 36637 1142
rect 36243 863 36637 902
rect 36957 1142 37351 1182
rect 36957 902 36997 1142
rect 37317 902 37351 1142
rect 36957 863 37351 902
rect 37671 1142 38065 1182
rect 37671 902 37711 1142
rect 38031 902 38065 1142
rect 37671 862 38065 902
rect 38385 1142 38779 1182
rect 38385 902 38425 1142
rect 38745 902 38779 1142
rect 38385 862 38779 902
rect 14058 718 14068 818
rect 13978 708 14068 718
rect 11380 -1090 11480 -1080
rect 11380 -1120 11390 -1090
rect 10480 -1130 11390 -1120
rect 10480 -1240 10490 -1130
rect 10630 -1170 11390 -1130
rect 11470 -1170 11480 -1090
rect 10630 -1180 11480 -1170
rect 11790 270 11990 370
rect 10630 -1240 10640 -1180
rect 10480 -1250 10640 -1240
rect 11790 -1480 11890 270
rect 11980 100 12820 120
rect 11980 -180 12020 100
rect 12780 -180 12820 100
rect 11980 -200 12820 -180
rect 14598 -771 15198 818
rect 15537 -40 15931 -1
rect 15537 -280 15577 -40
rect 15897 -280 15931 -40
rect 15537 -320 15931 -280
rect 16251 -40 16645 -1
rect 16251 -280 16291 -40
rect 16611 -280 16645 -40
rect 16251 -320 16645 -280
rect 16965 -40 17359 -1
rect 16965 -280 17005 -40
rect 17325 -280 17359 -40
rect 16965 -320 17359 -280
rect 17679 -40 18073 -1
rect 17679 -280 17719 -40
rect 18039 -280 18073 -40
rect 17679 -320 18073 -280
rect 18393 -40 18787 -1
rect 18393 -280 18433 -40
rect 18753 -280 18787 -40
rect 18393 -320 18787 -280
rect 19107 -40 19501 -1
rect 19107 -280 19147 -40
rect 19467 -280 19501 -40
rect 19107 -320 19501 -280
rect 19821 -40 20215 -1
rect 19821 -280 19861 -40
rect 20181 -280 20215 -40
rect 19821 -320 20215 -280
rect 20535 -40 20929 -1
rect 20535 -280 20575 -40
rect 20895 -280 20929 -40
rect 20535 -320 20929 -280
rect 21249 -40 21643 -1
rect 21249 -280 21289 -40
rect 21609 -280 21643 -40
rect 21249 -320 21643 -280
rect 21963 -40 22357 -1
rect 21963 -280 22003 -40
rect 22323 -280 22357 -40
rect 21963 -320 22357 -280
rect 22677 -40 23071 -1
rect 22677 -280 22717 -40
rect 23037 -280 23071 -40
rect 22677 -320 23071 -280
rect 23391 -40 23785 -1
rect 23391 -280 23431 -40
rect 23751 -280 23785 -40
rect 23391 -320 23785 -280
rect 24105 -40 24499 -1
rect 24105 -280 24145 -40
rect 24465 -280 24499 -40
rect 24105 -320 24499 -280
rect 24819 -40 25213 -1
rect 24819 -280 24859 -40
rect 25179 -280 25213 -40
rect 24819 -320 25213 -280
rect 25533 -40 25927 -1
rect 25533 -280 25573 -40
rect 25893 -280 25927 -40
rect 25533 -320 25927 -280
rect 26247 -40 26641 -1
rect 26247 -280 26287 -40
rect 26607 -280 26641 -40
rect 26247 -320 26641 -280
rect 26961 -40 27355 -1
rect 26961 -280 27001 -40
rect 27321 -280 27355 -40
rect 26961 -320 27355 -280
rect 27675 -40 28069 -1
rect 27675 -280 27715 -40
rect 28035 -280 28069 -40
rect 27675 -320 28069 -280
rect 28389 -40 28783 -1
rect 28389 -280 28429 -40
rect 28749 -280 28783 -40
rect 28389 -320 28783 -280
rect 29103 -40 29497 -1
rect 29103 -280 29143 -40
rect 29463 -280 29497 -40
rect 29103 -320 29497 -280
rect 29817 -40 30211 -1
rect 29817 -280 29857 -40
rect 30177 -280 30211 -40
rect 29817 -320 30211 -280
rect 30531 -40 30925 -1
rect 30531 -280 30571 -40
rect 30891 -280 30925 -40
rect 30531 -320 30925 -280
rect 31245 -40 31639 -1
rect 31245 -280 31285 -40
rect 31605 -280 31639 -40
rect 31245 -320 31639 -280
rect 31959 -40 32353 -1
rect 31959 -280 31999 -40
rect 32319 -280 32353 -40
rect 31959 -320 32353 -280
rect 32673 -40 33067 -1
rect 32673 -280 32713 -40
rect 33033 -280 33067 -40
rect 32673 -320 33067 -280
rect 33387 -40 33781 -1
rect 33387 -280 33427 -40
rect 33747 -280 33781 -40
rect 33387 -320 33781 -280
rect 34101 -40 34495 -1
rect 34101 -280 34141 -40
rect 34461 -280 34495 -40
rect 34101 -320 34495 -280
rect 34815 -40 35209 -1
rect 34815 -280 34855 -40
rect 35175 -280 35209 -40
rect 34815 -320 35209 -280
rect 35529 -40 35923 -1
rect 35529 -280 35569 -40
rect 35889 -280 35923 -40
rect 35529 -320 35923 -280
rect 36243 -40 36637 -1
rect 36243 -280 36283 -40
rect 36603 -280 36637 -40
rect 36243 -320 36637 -280
rect 36957 -40 37351 -1
rect 36957 -280 36997 -40
rect 37317 -280 37351 -40
rect 36957 -320 37351 -280
rect 37671 -40 38065 -1
rect 37671 -280 37711 -40
rect 38031 -280 38065 -40
rect 37671 -320 38065 -280
rect 38385 -40 38779 -1
rect 38385 -280 38425 -40
rect 38745 -280 38779 -40
rect 38385 -320 38779 -280
rect 15537 -440 15931 -380
rect 15537 -771 15597 -440
rect 14598 -1040 15597 -771
rect 14598 -1360 14640 -1040
rect 14960 -1360 15597 -1040
rect 14598 -1371 15597 -1360
rect 14600 -1400 15000 -1371
rect 11310 -1490 11890 -1480
rect 11310 -1570 11320 -1490
rect 11400 -1570 11890 -1490
rect 11310 -1580 11890 -1570
rect 5802 -2100 14802 -2000
rect 5802 -2700 5902 -2100
rect 7102 -2700 9102 -2100
rect 10302 -2500 12102 -2100
rect 10302 -2700 10542 -2500
rect 5802 -2800 10542 -2700
rect 12002 -2700 12102 -2500
rect 14702 -2700 14802 -2100
rect 12002 -2800 14802 -2700
rect 10303 -2920 10542 -2800
rect 10302 -2940 10542 -2920
rect 10302 -3860 10322 -2940
rect 10522 -3860 10542 -2940
rect 10702 -3152 11602 -3052
rect 10702 -3552 10802 -3152
rect 11502 -3552 11602 -3152
rect 10702 -3652 11602 -3552
rect 12002 -3340 14802 -3200
rect 10302 -4052 10542 -3860
rect 2600 -4120 7000 -4100
rect 2600 -4280 2620 -4120
rect 2700 -4280 7000 -4120
rect 2600 -4300 7000 -4280
rect 6800 -5400 7000 -4300
rect 10302 -4192 11602 -4052
rect 6800 -5420 8300 -5400
rect 6800 -5580 8120 -5420
rect 8280 -5580 8300 -5420
rect 6800 -5600 8300 -5580
rect 5000 -6340 5600 -6310
rect 0 -6600 100 -6400
rect 200 -6600 300 -6400
rect 0 -6700 300 -6600
rect 400 -6700 500 -6400
rect 600 -6700 700 -6400
rect 800 -6600 1100 -6400
rect 5000 -6420 5030 -6340
rect 5000 -6580 5020 -6420
rect 5570 -6420 5600 -6340
rect 5580 -6580 5600 -6420
rect 5000 -6600 5600 -6580
rect 800 -6700 900 -6600
rect 1000 -6700 1100 -6600
rect 6000 -6650 6130 -6640
rect 6000 -6700 6010 -6650
rect 5000 -6740 6010 -6700
rect 6120 -6740 6130 -6650
rect 5000 -6750 6130 -6740
rect 5000 -6920 5050 -6750
rect -360 -7080 5050 -6920
rect 5000 -9350 5050 -7080
rect 5750 -6760 6130 -6750
rect 5750 -9350 5800 -6760
rect 5000 -9400 5800 -9350
rect 6402 -9300 9802 -9200
rect 3400 -9800 4600 -9600
rect 6402 -9800 6502 -9300
rect 9702 -9800 9802 -9300
rect 10302 -9512 10442 -4192
rect 11462 -9512 11602 -4192
rect 10302 -9652 11602 -9512
rect 12002 -9460 12142 -3340
rect 14662 -9100 14802 -3340
rect 15537 -6680 15597 -1371
rect 15877 -771 15931 -440
rect 16251 -440 16645 -380
rect 16251 -771 16311 -440
rect 15877 -1371 16311 -771
rect 15877 -6680 15931 -1371
rect 15537 -6740 15931 -6680
rect 16251 -6680 16311 -1371
rect 16591 -771 16645 -440
rect 16965 -440 17359 -380
rect 16965 -771 17025 -440
rect 16591 -1371 17025 -771
rect 16591 -6680 16645 -1371
rect 16251 -6740 16645 -6680
rect 16965 -6680 17025 -1371
rect 17305 -771 17359 -440
rect 17679 -440 18073 -380
rect 17679 -771 17739 -440
rect 17305 -1371 17739 -771
rect 17305 -6680 17359 -1371
rect 16965 -6740 17359 -6680
rect 17679 -6680 17739 -1371
rect 18019 -771 18073 -440
rect 18393 -440 18787 -380
rect 18393 -771 18453 -440
rect 18019 -1371 18453 -771
rect 18019 -6680 18073 -1371
rect 17679 -6740 18073 -6680
rect 18393 -6680 18453 -1371
rect 18733 -771 18787 -440
rect 19107 -440 19501 -380
rect 19107 -771 19167 -440
rect 18733 -1371 19167 -771
rect 18733 -6680 18787 -1371
rect 18393 -6740 18787 -6680
rect 19107 -6680 19167 -1371
rect 19447 -771 19501 -440
rect 19821 -440 20215 -380
rect 19821 -771 19881 -440
rect 19447 -1371 19881 -771
rect 19447 -6680 19501 -1371
rect 19107 -6740 19501 -6680
rect 19821 -6680 19881 -1371
rect 20161 -771 20215 -440
rect 20535 -440 20929 -380
rect 20535 -771 20595 -440
rect 20161 -1371 20595 -771
rect 20161 -6680 20215 -1371
rect 19821 -6740 20215 -6680
rect 20535 -6680 20595 -1371
rect 20875 -771 20929 -440
rect 21249 -440 21643 -380
rect 21249 -771 21309 -440
rect 20875 -1371 21309 -771
rect 20875 -6680 20929 -1371
rect 20535 -6740 20929 -6680
rect 21249 -6680 21309 -1371
rect 21589 -771 21643 -440
rect 21963 -440 22357 -380
rect 21963 -771 22023 -440
rect 21589 -1371 22023 -771
rect 21589 -6680 21643 -1371
rect 21249 -6740 21643 -6680
rect 21963 -6680 22023 -1371
rect 22303 -771 22357 -440
rect 22677 -440 23071 -380
rect 22677 -771 22737 -440
rect 22303 -1371 22737 -771
rect 22303 -6680 22357 -1371
rect 21963 -6740 22357 -6680
rect 22677 -6680 22737 -1371
rect 23017 -771 23071 -440
rect 23391 -440 23785 -380
rect 23391 -771 23451 -440
rect 23017 -1371 23451 -771
rect 23017 -6680 23071 -1371
rect 22677 -6740 23071 -6680
rect 23391 -6680 23451 -1371
rect 23731 -771 23785 -440
rect 24105 -440 24499 -380
rect 24105 -771 24165 -440
rect 23731 -1371 24165 -771
rect 23731 -6680 23785 -1371
rect 23391 -6740 23785 -6680
rect 24105 -6680 24165 -1371
rect 24445 -771 24499 -440
rect 24819 -440 25213 -380
rect 24819 -771 24879 -440
rect 24445 -1371 24879 -771
rect 24445 -6680 24499 -1371
rect 24105 -6740 24499 -6680
rect 24819 -6680 24879 -1371
rect 25159 -771 25213 -440
rect 25533 -440 25927 -380
rect 25533 -771 25593 -440
rect 25159 -1371 25593 -771
rect 25159 -6680 25213 -1371
rect 24819 -6740 25213 -6680
rect 25533 -6680 25593 -1371
rect 25873 -771 25927 -440
rect 26247 -440 26641 -380
rect 26247 -771 26307 -440
rect 25873 -1371 26307 -771
rect 25873 -6680 25927 -1371
rect 25533 -6740 25927 -6680
rect 26247 -6680 26307 -1371
rect 26587 -771 26641 -440
rect 26961 -440 27355 -380
rect 26961 -771 27021 -440
rect 26587 -1371 27021 -771
rect 26587 -6680 26641 -1371
rect 26247 -6740 26641 -6680
rect 26961 -6680 27021 -1371
rect 27301 -771 27355 -440
rect 27675 -440 28069 -380
rect 27675 -771 27735 -440
rect 27301 -1371 27735 -771
rect 27301 -6680 27355 -1371
rect 26961 -6740 27355 -6680
rect 27675 -6680 27735 -1371
rect 28015 -771 28069 -440
rect 28389 -440 28783 -380
rect 28389 -771 28449 -440
rect 28015 -1371 28449 -771
rect 28015 -6680 28069 -1371
rect 27675 -6740 28069 -6680
rect 28389 -6680 28449 -1371
rect 28729 -771 28783 -440
rect 29103 -440 29497 -380
rect 29103 -771 29163 -440
rect 28729 -1371 29163 -771
rect 28729 -6680 28783 -1371
rect 28389 -6740 28783 -6680
rect 29103 -6680 29163 -1371
rect 29443 -771 29497 -440
rect 29817 -440 30211 -380
rect 29817 -771 29877 -440
rect 29443 -1371 29877 -771
rect 29443 -6680 29497 -1371
rect 29103 -6740 29497 -6680
rect 29817 -6680 29877 -1371
rect 30157 -771 30211 -440
rect 30531 -440 30925 -380
rect 30531 -771 30591 -440
rect 30157 -1371 30591 -771
rect 30157 -6680 30211 -1371
rect 29817 -6740 30211 -6680
rect 30531 -6680 30591 -1371
rect 30871 -771 30925 -440
rect 31245 -440 31639 -380
rect 31245 -771 31305 -440
rect 30871 -1371 31305 -771
rect 30871 -6680 30925 -1371
rect 30531 -6740 30925 -6680
rect 31245 -6680 31305 -1371
rect 31585 -771 31639 -440
rect 31959 -440 32353 -380
rect 31959 -771 32019 -440
rect 31585 -1371 32019 -771
rect 31585 -6680 31639 -1371
rect 31245 -6740 31639 -6680
rect 31959 -6680 32019 -1371
rect 32299 -771 32353 -440
rect 32673 -440 33067 -380
rect 32673 -771 32733 -440
rect 32299 -1371 32733 -771
rect 32299 -6680 32353 -1371
rect 31959 -6740 32353 -6680
rect 32673 -6680 32733 -1371
rect 33013 -771 33067 -440
rect 33387 -440 33781 -380
rect 33387 -771 33447 -440
rect 33013 -1371 33447 -771
rect 33013 -6680 33067 -1371
rect 32673 -6740 33067 -6680
rect 33387 -6680 33447 -1371
rect 33727 -771 33781 -440
rect 34101 -440 34495 -380
rect 34101 -771 34161 -440
rect 33727 -1371 34161 -771
rect 33727 -6680 33781 -1371
rect 33387 -6740 33781 -6680
rect 34101 -6680 34161 -1371
rect 34441 -771 34495 -440
rect 34815 -440 35209 -380
rect 34815 -771 34875 -440
rect 34441 -1371 34875 -771
rect 34441 -6680 34495 -1371
rect 34101 -6740 34495 -6680
rect 34815 -6680 34875 -1371
rect 35155 -771 35209 -440
rect 35529 -440 35923 -380
rect 35529 -771 35589 -440
rect 35155 -1371 35589 -771
rect 35155 -6680 35209 -1371
rect 34815 -6740 35209 -6680
rect 35529 -6680 35589 -1371
rect 35869 -771 35923 -440
rect 36243 -440 36637 -380
rect 36243 -771 36303 -440
rect 35869 -1371 36303 -771
rect 35869 -6680 35923 -1371
rect 35529 -6740 35923 -6680
rect 36243 -6680 36303 -1371
rect 36583 -771 36637 -440
rect 36957 -440 37351 -380
rect 36957 -771 37017 -440
rect 36583 -1371 37017 -771
rect 36583 -6680 36637 -1371
rect 36243 -6740 36637 -6680
rect 36957 -6680 37017 -1371
rect 37297 -771 37351 -440
rect 37671 -440 38065 -380
rect 37671 -771 37731 -440
rect 37297 -1371 37731 -771
rect 37297 -6680 37351 -1371
rect 36957 -6740 37351 -6680
rect 37671 -6680 37731 -1371
rect 38011 -771 38065 -440
rect 38385 -440 38779 -380
rect 38385 -771 38445 -440
rect 38011 -1371 38445 -771
rect 38011 -6680 38065 -1371
rect 37671 -6740 38065 -6680
rect 38385 -6680 38445 -1371
rect 38725 -6680 38779 -440
rect 40000 -900 40600 -800
rect 40000 -1300 40100 -900
rect 40500 -1300 40600 -900
rect 40000 -1400 40600 -1300
rect 38385 -6740 38779 -6680
rect 14662 -9200 44200 -9100
rect 14662 -9460 43100 -9200
rect 12002 -9600 43100 -9460
rect 3400 -10400 3600 -9800
rect 4400 -9900 9802 -9800
rect 12202 -9900 43100 -9600
rect 4400 -10300 43100 -9900
rect 44100 -10300 44200 -9200
rect 4400 -10400 44200 -10300
rect 3400 -10600 4600 -10400
<< via4 >>
rect 3600 13200 4400 13800
rect 5030 9740 5570 9980
rect 10802 6552 11502 6952
rect 43100 12600 44100 13700
rect 12102 5500 14702 6100
rect 3228 3995 3468 4315
rect 4374 3995 4614 4315
rect 8640 3960 9560 4260
rect 3228 3281 3468 3601
rect 4374 3281 4614 3601
rect 3941 225 4181 545
rect 3941 -489 4181 -169
rect 9920 -740 10040 -420
rect 10040 -740 10160 -420
rect 40100 1900 40500 2100
rect 40100 1700 40500 1900
rect 15577 902 15897 1142
rect 16291 902 16611 1142
rect 17005 902 17325 1142
rect 17719 902 18039 1142
rect 18433 902 18753 1142
rect 19147 902 19467 1142
rect 19861 902 20181 1142
rect 20575 902 20895 1142
rect 21289 902 21609 1142
rect 22003 902 22323 1142
rect 22717 902 23037 1142
rect 23431 902 23751 1142
rect 24145 902 24465 1142
rect 24859 902 25179 1142
rect 25573 902 25893 1142
rect 26287 902 26607 1142
rect 27001 902 27321 1142
rect 27715 902 28035 1142
rect 28429 902 28749 1142
rect 29143 902 29463 1142
rect 29857 902 30177 1142
rect 30571 902 30891 1142
rect 31285 902 31605 1142
rect 31999 902 32319 1142
rect 32713 902 33033 1142
rect 33427 902 33747 1142
rect 34141 902 34461 1142
rect 34855 902 35175 1142
rect 35569 902 35889 1142
rect 36283 902 36603 1142
rect 36997 902 37317 1142
rect 37711 902 38031 1142
rect 38425 902 38745 1142
rect 12020 -180 12780 100
rect 15577 -280 15897 -40
rect 16291 -280 16611 -40
rect 17005 -280 17325 -40
rect 17719 -280 18039 -40
rect 18433 -280 18753 -40
rect 19147 -280 19467 -40
rect 19861 -280 20181 -40
rect 20575 -280 20895 -40
rect 21289 -280 21609 -40
rect 22003 -280 22323 -40
rect 22717 -280 23037 -40
rect 23431 -280 23751 -40
rect 24145 -280 24465 -40
rect 24859 -280 25179 -40
rect 25573 -280 25893 -40
rect 26287 -280 26607 -40
rect 27001 -280 27321 -40
rect 27715 -280 28035 -40
rect 28429 -280 28749 -40
rect 29143 -280 29463 -40
rect 29857 -280 30177 -40
rect 30571 -280 30891 -40
rect 31285 -280 31605 -40
rect 31999 -280 32319 -40
rect 32713 -280 33033 -40
rect 33427 -280 33747 -40
rect 34141 -280 34461 -40
rect 34855 -280 35175 -40
rect 35569 -280 35889 -40
rect 36283 -280 36603 -40
rect 36997 -280 37317 -40
rect 37711 -280 38031 -40
rect 38425 -280 38745 -40
rect 12102 -2700 14702 -2100
rect 10802 -3552 11502 -3152
rect 5030 -6580 5570 -6340
rect 40100 -1100 40500 -900
rect 40100 -1300 40500 -1100
rect 3600 -10400 4400 -9800
rect 43100 -10300 44100 -9200
<< mimcap2 >>
rect 10402 12912 11502 12952
rect 5030 12750 5770 12770
rect 5030 10150 5050 12750
rect 5750 10150 5770 12750
rect 5030 10130 5770 10150
rect 10402 7592 10442 12912
rect 11462 7592 11502 12912
rect 10402 7552 11502 7592
rect 12102 12860 14702 12900
rect 12102 6740 12142 12860
rect 14662 6740 14702 12860
rect 12102 6700 14702 6740
rect 15577 7542 15897 7562
rect 1518 4295 3088 4315
rect 1518 4015 1538 4295
rect 3068 4015 3088 4295
rect 1518 3995 3088 4015
rect 4754 4295 6324 4315
rect 4754 4015 4774 4295
rect 6304 4015 6324 4295
rect 4754 3995 6324 4015
rect -52 3581 3088 3601
rect -52 3301 -32 3581
rect 3068 3301 3088 3581
rect -52 3281 3088 3301
rect 4754 3581 7894 3601
rect 4754 3301 4774 3581
rect 7874 3301 7894 3581
rect 4754 3281 7894 3301
rect 15577 1302 15597 7542
rect 15877 1302 15897 7542
rect 15577 1282 15897 1302
rect 16291 7542 16611 7562
rect 16291 1302 16311 7542
rect 16591 1302 16611 7542
rect 16291 1282 16611 1302
rect 17005 7542 17325 7562
rect 17005 1302 17025 7542
rect 17305 1302 17325 7542
rect 17005 1282 17325 1302
rect 17719 7542 18039 7562
rect 17719 1302 17739 7542
rect 18019 1302 18039 7542
rect 17719 1282 18039 1302
rect 18433 7542 18753 7562
rect 18433 1302 18453 7542
rect 18733 1302 18753 7542
rect 18433 1282 18753 1302
rect 19147 7542 19467 7562
rect 19147 1302 19167 7542
rect 19447 1302 19467 7542
rect 19147 1282 19467 1302
rect 19861 7542 20181 7562
rect 19861 1302 19881 7542
rect 20161 1302 20181 7542
rect 19861 1282 20181 1302
rect 20575 7542 20895 7562
rect 20575 1302 20595 7542
rect 20875 1302 20895 7542
rect 20575 1282 20895 1302
rect 21289 7542 21609 7562
rect 21289 1302 21309 7542
rect 21589 1302 21609 7542
rect 21289 1282 21609 1302
rect 22003 7542 22323 7562
rect 22003 1302 22023 7542
rect 22303 1302 22323 7542
rect 22003 1282 22323 1302
rect 22717 7542 23037 7562
rect 22717 1302 22737 7542
rect 23017 1302 23037 7542
rect 22717 1282 23037 1302
rect 23431 7542 23751 7562
rect 23431 1302 23451 7542
rect 23731 1302 23751 7542
rect 23431 1282 23751 1302
rect 24145 7542 24465 7562
rect 24145 1302 24165 7542
rect 24445 1302 24465 7542
rect 24145 1282 24465 1302
rect 24859 7542 25179 7562
rect 24859 1302 24879 7542
rect 25159 1302 25179 7542
rect 24859 1282 25179 1302
rect 25573 7542 25893 7562
rect 25573 1302 25593 7542
rect 25873 1302 25893 7542
rect 25573 1282 25893 1302
rect 26287 7542 26607 7562
rect 26287 1302 26307 7542
rect 26587 1302 26607 7542
rect 26287 1282 26607 1302
rect 27001 7542 27321 7562
rect 27001 1302 27021 7542
rect 27301 1302 27321 7542
rect 27001 1282 27321 1302
rect 27715 7542 28035 7562
rect 27715 1302 27735 7542
rect 28015 1302 28035 7542
rect 27715 1282 28035 1302
rect 28429 7542 28749 7562
rect 28429 1302 28449 7542
rect 28729 1302 28749 7542
rect 28429 1282 28749 1302
rect 29143 7542 29463 7562
rect 29143 1302 29163 7542
rect 29443 1302 29463 7542
rect 29143 1282 29463 1302
rect 29857 7542 30177 7562
rect 29857 1302 29877 7542
rect 30157 1302 30177 7542
rect 29857 1282 30177 1302
rect 30571 7542 30891 7562
rect 30571 1302 30591 7542
rect 30871 1302 30891 7542
rect 30571 1282 30891 1302
rect 31285 7542 31605 7562
rect 31285 1302 31305 7542
rect 31585 1302 31605 7542
rect 31285 1282 31605 1302
rect 31999 7542 32319 7562
rect 31999 1302 32019 7542
rect 32299 1302 32319 7542
rect 31999 1282 32319 1302
rect 32713 7542 33033 7562
rect 32713 1302 32733 7542
rect 33013 1302 33033 7542
rect 32713 1282 33033 1302
rect 33427 7542 33747 7562
rect 33427 1302 33447 7542
rect 33727 1302 33747 7542
rect 33427 1282 33747 1302
rect 34141 7542 34461 7562
rect 34141 1302 34161 7542
rect 34441 1302 34461 7542
rect 34141 1282 34461 1302
rect 34855 7542 35175 7562
rect 34855 1302 34875 7542
rect 35155 1302 35175 7542
rect 34855 1282 35175 1302
rect 35569 7542 35889 7562
rect 35569 1302 35589 7542
rect 35869 1302 35889 7542
rect 35569 1282 35889 1302
rect 36283 7542 36603 7562
rect 36283 1302 36303 7542
rect 36583 1302 36603 7542
rect 36283 1282 36603 1302
rect 36997 7542 37317 7562
rect 36997 1302 37017 7542
rect 37297 1302 37317 7542
rect 36997 1282 37317 1302
rect 37711 4402 38031 4422
rect 37711 1302 37731 4402
rect 38011 1302 38031 4402
rect 37711 1282 38031 1302
rect 38425 2832 38745 2852
rect 38425 1302 38445 2832
rect 38725 1302 38745 2832
rect 38425 1282 38745 1302
rect 4321 525 5891 545
rect 4321 245 4341 525
rect 5871 245 5891 525
rect 4321 225 5891 245
rect 4321 -189 7461 -169
rect 4321 -469 4341 -189
rect 7441 -469 7461 -189
rect 4321 -489 7461 -469
rect 15577 -440 15897 -420
rect 12102 -3340 14702 -3300
rect 10402 -4192 11502 -4152
rect 5030 -6750 5770 -6730
rect 5030 -9350 5050 -6750
rect 5750 -9350 5770 -6750
rect 5030 -9370 5770 -9350
rect 10402 -9512 10442 -4192
rect 11462 -9512 11502 -4192
rect 12102 -9460 12142 -3340
rect 14662 -9460 14702 -3340
rect 15577 -6680 15597 -440
rect 15877 -6680 15897 -440
rect 15577 -6700 15897 -6680
rect 16291 -440 16611 -420
rect 16291 -6680 16311 -440
rect 16591 -6680 16611 -440
rect 16291 -6700 16611 -6680
rect 17005 -440 17325 -420
rect 17005 -6680 17025 -440
rect 17305 -6680 17325 -440
rect 17005 -6700 17325 -6680
rect 17719 -440 18039 -420
rect 17719 -6680 17739 -440
rect 18019 -6680 18039 -440
rect 17719 -6700 18039 -6680
rect 18433 -440 18753 -420
rect 18433 -6680 18453 -440
rect 18733 -6680 18753 -440
rect 18433 -6700 18753 -6680
rect 19147 -440 19467 -420
rect 19147 -6680 19167 -440
rect 19447 -6680 19467 -440
rect 19147 -6700 19467 -6680
rect 19861 -440 20181 -420
rect 19861 -6680 19881 -440
rect 20161 -6680 20181 -440
rect 19861 -6700 20181 -6680
rect 20575 -440 20895 -420
rect 20575 -6680 20595 -440
rect 20875 -6680 20895 -440
rect 20575 -6700 20895 -6680
rect 21289 -440 21609 -420
rect 21289 -6680 21309 -440
rect 21589 -6680 21609 -440
rect 21289 -6700 21609 -6680
rect 22003 -440 22323 -420
rect 22003 -6680 22023 -440
rect 22303 -6680 22323 -440
rect 22003 -6700 22323 -6680
rect 22717 -440 23037 -420
rect 22717 -6680 22737 -440
rect 23017 -6680 23037 -440
rect 22717 -6700 23037 -6680
rect 23431 -440 23751 -420
rect 23431 -6680 23451 -440
rect 23731 -6680 23751 -440
rect 23431 -6700 23751 -6680
rect 24145 -440 24465 -420
rect 24145 -6680 24165 -440
rect 24445 -6680 24465 -440
rect 24145 -6700 24465 -6680
rect 24859 -440 25179 -420
rect 24859 -6680 24879 -440
rect 25159 -6680 25179 -440
rect 24859 -6700 25179 -6680
rect 25573 -440 25893 -420
rect 25573 -6680 25593 -440
rect 25873 -6680 25893 -440
rect 25573 -6700 25893 -6680
rect 26287 -440 26607 -420
rect 26287 -6680 26307 -440
rect 26587 -6680 26607 -440
rect 26287 -6700 26607 -6680
rect 27001 -440 27321 -420
rect 27001 -6680 27021 -440
rect 27301 -6680 27321 -440
rect 27001 -6700 27321 -6680
rect 27715 -440 28035 -420
rect 27715 -6680 27735 -440
rect 28015 -6680 28035 -440
rect 27715 -6700 28035 -6680
rect 28429 -440 28749 -420
rect 28429 -6680 28449 -440
rect 28729 -6680 28749 -440
rect 28429 -6700 28749 -6680
rect 29143 -440 29463 -420
rect 29143 -6680 29163 -440
rect 29443 -6680 29463 -440
rect 29143 -6700 29463 -6680
rect 29857 -440 30177 -420
rect 29857 -6680 29877 -440
rect 30157 -6680 30177 -440
rect 29857 -6700 30177 -6680
rect 30571 -440 30891 -420
rect 30571 -6680 30591 -440
rect 30871 -6680 30891 -440
rect 30571 -6700 30891 -6680
rect 31285 -440 31605 -420
rect 31285 -6680 31305 -440
rect 31585 -6680 31605 -440
rect 31285 -6700 31605 -6680
rect 31999 -440 32319 -420
rect 31999 -6680 32019 -440
rect 32299 -6680 32319 -440
rect 31999 -6700 32319 -6680
rect 32713 -440 33033 -420
rect 32713 -6680 32733 -440
rect 33013 -6680 33033 -440
rect 32713 -6700 33033 -6680
rect 33427 -440 33747 -420
rect 33427 -6680 33447 -440
rect 33727 -6680 33747 -440
rect 33427 -6700 33747 -6680
rect 34141 -440 34461 -420
rect 34141 -6680 34161 -440
rect 34441 -6680 34461 -440
rect 34141 -6700 34461 -6680
rect 34855 -440 35175 -420
rect 34855 -6680 34875 -440
rect 35155 -6680 35175 -440
rect 34855 -6700 35175 -6680
rect 35569 -440 35889 -420
rect 35569 -6680 35589 -440
rect 35869 -6680 35889 -440
rect 35569 -6700 35889 -6680
rect 36283 -440 36603 -420
rect 36283 -6680 36303 -440
rect 36583 -6680 36603 -440
rect 36283 -6700 36603 -6680
rect 36997 -440 37317 -420
rect 36997 -6680 37017 -440
rect 37297 -6680 37317 -440
rect 36997 -6700 37317 -6680
rect 37711 -440 38031 -420
rect 37711 -6680 37731 -440
rect 38011 -6680 38031 -440
rect 37711 -6700 38031 -6680
rect 38425 -440 38745 -420
rect 38425 -6680 38445 -440
rect 38725 -6680 38745 -440
rect 38425 -6700 38745 -6680
rect 12102 -9500 14702 -9460
rect 10402 -9552 11502 -9512
<< mimcap2contact >>
rect 5050 10150 5750 12750
rect 10442 7592 11462 12912
rect 12142 6740 14662 12860
rect 1538 4015 3068 4295
rect 4774 4015 6304 4295
rect -32 3301 3068 3581
rect 4774 3301 7874 3581
rect 15597 1302 15877 7542
rect 16311 1302 16591 7542
rect 17025 1302 17305 7542
rect 17739 1302 18019 7542
rect 18453 1302 18733 7542
rect 19167 1302 19447 7542
rect 19881 1302 20161 7542
rect 20595 1302 20875 7542
rect 21309 1302 21589 7542
rect 22023 1302 22303 7542
rect 22737 1302 23017 7542
rect 23451 1302 23731 7542
rect 24165 1302 24445 7542
rect 24879 1302 25159 7542
rect 25593 1302 25873 7542
rect 26307 1302 26587 7542
rect 27021 1302 27301 7542
rect 27735 1302 28015 7542
rect 28449 1302 28729 7542
rect 29163 1302 29443 7542
rect 29877 1302 30157 7542
rect 30591 1302 30871 7542
rect 31305 1302 31585 7542
rect 32019 1302 32299 7542
rect 32733 1302 33013 7542
rect 33447 1302 33727 7542
rect 34161 1302 34441 7542
rect 34875 1302 35155 7542
rect 35589 1302 35869 7542
rect 36303 1302 36583 7542
rect 37017 1302 37297 7542
rect 37731 1302 38011 4402
rect 38445 1302 38725 2832
rect 4341 245 5871 525
rect 4341 -469 7441 -189
rect 5050 -9350 5750 -6750
rect 10442 -9512 11462 -4192
rect 12142 -9460 14662 -3340
rect 15597 -6680 15877 -440
rect 16311 -6680 16591 -440
rect 17025 -6680 17305 -440
rect 17739 -6680 18019 -440
rect 18453 -6680 18733 -440
rect 19167 -6680 19447 -440
rect 19881 -6680 20161 -440
rect 20595 -6680 20875 -440
rect 21309 -6680 21589 -440
rect 22023 -6680 22303 -440
rect 22737 -6680 23017 -440
rect 23451 -6680 23731 -440
rect 24165 -6680 24445 -440
rect 24879 -6680 25159 -440
rect 25593 -6680 25873 -440
rect 26307 -6680 26587 -440
rect 27021 -6680 27301 -440
rect 27735 -6680 28015 -440
rect 28449 -6680 28729 -440
rect 29163 -6680 29443 -440
rect 29877 -6680 30157 -440
rect 30591 -6680 30871 -440
rect 31305 -6680 31585 -440
rect 32019 -6680 32299 -440
rect 32733 -6680 33013 -440
rect 33447 -6680 33727 -440
rect 34161 -6680 34441 -440
rect 34875 -6680 35155 -440
rect 35589 -6680 35869 -440
rect 36303 -6680 36583 -440
rect 37017 -6680 37297 -440
rect 37731 -6680 38011 -440
rect 38445 -6680 38725 -440
<< metal5 >>
rect 3400 13800 4600 15000
rect 3400 13200 3600 13800
rect 4400 13200 4600 13800
rect 3400 5400 4600 13200
rect 10302 12912 11602 13052
rect 5000 12750 5800 12800
rect 5000 10150 5050 12750
rect 5750 10150 5800 12750
rect 5000 10100 5800 10150
rect 5000 9980 5600 10100
rect 5000 9740 5030 9980
rect 5570 9740 5600 9980
rect 5000 9710 5600 9740
rect 10302 7592 10442 12912
rect 11462 7592 11602 12912
rect 10302 7452 11602 7592
rect 10702 6952 11602 7452
rect 10702 6552 10802 6952
rect 11502 6552 11602 6952
rect 10702 6452 11602 6552
rect 12000 13000 13200 15000
rect 12000 12860 14802 13000
rect 12000 6740 12142 12860
rect 14662 6740 14802 12860
rect 12000 6100 14802 6740
rect 12000 5500 12102 6100
rect 14702 5500 14802 6100
rect 12000 5400 14802 5500
rect 15537 7542 15931 7602
rect 3400 4800 9600 5400
rect 1478 4315 3508 4355
rect 1478 4295 3228 4315
rect 1478 4015 1538 4295
rect 3068 4015 3228 4295
rect 1478 3995 3228 4015
rect 3468 3995 3508 4315
rect 1478 3961 3508 3995
rect 4334 4315 6364 4355
rect 4334 3995 4374 4315
rect 4614 4295 6364 4315
rect 4614 4015 4774 4295
rect 6304 4015 6364 4295
rect 4614 3995 6364 4015
rect 4334 3961 6364 3995
rect 8600 4260 9600 4800
rect 8600 3960 8640 4260
rect 9560 3960 9600 4260
rect -92 3601 3508 3641
rect -92 3581 3228 3601
rect -92 3301 -32 3581
rect 3068 3301 3228 3581
rect -92 3281 3228 3301
rect 3468 3281 3508 3601
rect -92 3247 3508 3281
rect 4334 3601 7934 3641
rect 4334 3281 4374 3601
rect 4614 3581 7934 3601
rect 4614 3301 4774 3581
rect 7874 3301 7934 3581
rect 4614 3281 7934 3301
rect 4334 3247 7934 3281
rect 3901 545 5931 585
rect 3901 225 3941 545
rect 4181 525 5931 545
rect 4181 245 4341 525
rect 5871 245 5931 525
rect 4181 225 5931 245
rect 3901 191 5931 225
rect 3901 -169 7501 -129
rect 3901 -489 3941 -169
rect 4181 -189 7501 -169
rect 4181 -469 4341 -189
rect 7441 -469 7501 -189
rect 4181 -489 7501 -469
rect 3901 -523 7501 -489
rect 8600 -380 9600 3960
rect 11600 5000 13200 5400
rect 11600 120 12800 5000
rect 15537 1302 15597 7542
rect 15877 1302 15931 7542
rect 15537 1142 15931 1302
rect 15537 902 15577 1142
rect 15897 902 15931 1142
rect 15537 863 15931 902
rect 16251 7542 16645 7602
rect 16251 1302 16311 7542
rect 16591 1302 16645 7542
rect 16251 1142 16645 1302
rect 16251 902 16291 1142
rect 16611 902 16645 1142
rect 16251 863 16645 902
rect 16965 7542 17359 7602
rect 16965 1302 17025 7542
rect 17305 1302 17359 7542
rect 16965 1142 17359 1302
rect 16965 902 17005 1142
rect 17325 902 17359 1142
rect 16965 863 17359 902
rect 17679 7542 18073 7602
rect 17679 1302 17739 7542
rect 18019 1302 18073 7542
rect 17679 1142 18073 1302
rect 17679 902 17719 1142
rect 18039 902 18073 1142
rect 17679 863 18073 902
rect 18393 7542 18787 7602
rect 18393 1302 18453 7542
rect 18733 1302 18787 7542
rect 18393 1142 18787 1302
rect 18393 902 18433 1142
rect 18753 902 18787 1142
rect 18393 863 18787 902
rect 19107 7542 19501 7602
rect 19107 1302 19167 7542
rect 19447 1302 19501 7542
rect 19107 1142 19501 1302
rect 19107 902 19147 1142
rect 19467 902 19501 1142
rect 19107 863 19501 902
rect 19821 7542 20215 7602
rect 19821 1302 19881 7542
rect 20161 1302 20215 7542
rect 19821 1142 20215 1302
rect 19821 902 19861 1142
rect 20181 902 20215 1142
rect 19821 863 20215 902
rect 20535 7542 20929 7602
rect 20535 1302 20595 7542
rect 20875 1302 20929 7542
rect 20535 1142 20929 1302
rect 20535 902 20575 1142
rect 20895 902 20929 1142
rect 20535 863 20929 902
rect 21249 7542 21643 7602
rect 21249 1302 21309 7542
rect 21589 1302 21643 7542
rect 21249 1142 21643 1302
rect 21249 902 21289 1142
rect 21609 902 21643 1142
rect 21249 863 21643 902
rect 21963 7542 22357 7602
rect 21963 1302 22023 7542
rect 22303 1302 22357 7542
rect 21963 1142 22357 1302
rect 21963 902 22003 1142
rect 22323 902 22357 1142
rect 21963 863 22357 902
rect 22677 7542 23071 7602
rect 22677 1302 22737 7542
rect 23017 1302 23071 7542
rect 22677 1142 23071 1302
rect 22677 902 22717 1142
rect 23037 902 23071 1142
rect 22677 863 23071 902
rect 23391 7542 23785 7602
rect 23391 1302 23451 7542
rect 23731 1302 23785 7542
rect 23391 1142 23785 1302
rect 23391 902 23431 1142
rect 23751 902 23785 1142
rect 23391 863 23785 902
rect 24105 7542 24499 7602
rect 24105 1302 24165 7542
rect 24445 1302 24499 7542
rect 24105 1142 24499 1302
rect 24105 902 24145 1142
rect 24465 902 24499 1142
rect 24105 863 24499 902
rect 24819 7542 25213 7602
rect 24819 1302 24879 7542
rect 25159 1302 25213 7542
rect 24819 1142 25213 1302
rect 24819 902 24859 1142
rect 25179 902 25213 1142
rect 24819 863 25213 902
rect 25533 7542 25927 7602
rect 25533 1302 25593 7542
rect 25873 1302 25927 7542
rect 25533 1142 25927 1302
rect 25533 902 25573 1142
rect 25893 902 25927 1142
rect 25533 863 25927 902
rect 26247 7542 26641 7602
rect 26247 1302 26307 7542
rect 26587 1302 26641 7542
rect 26247 1142 26641 1302
rect 26247 902 26287 1142
rect 26607 902 26641 1142
rect 26247 863 26641 902
rect 26961 7542 27355 7602
rect 26961 1302 27021 7542
rect 27301 1302 27355 7542
rect 26961 1142 27355 1302
rect 26961 902 27001 1142
rect 27321 902 27355 1142
rect 26961 863 27355 902
rect 27675 7542 28069 7602
rect 27675 1302 27735 7542
rect 28015 1302 28069 7542
rect 27675 1142 28069 1302
rect 27675 902 27715 1142
rect 28035 902 28069 1142
rect 27675 863 28069 902
rect 28389 7542 28783 7602
rect 28389 1302 28449 7542
rect 28729 1302 28783 7542
rect 28389 1142 28783 1302
rect 28389 902 28429 1142
rect 28749 902 28783 1142
rect 28389 863 28783 902
rect 29103 7542 29497 7602
rect 29103 1302 29163 7542
rect 29443 1302 29497 7542
rect 29103 1142 29497 1302
rect 29103 902 29143 1142
rect 29463 902 29497 1142
rect 29103 863 29497 902
rect 29817 7542 30211 7602
rect 29817 1302 29877 7542
rect 30157 1302 30211 7542
rect 29817 1142 30211 1302
rect 29817 902 29857 1142
rect 30177 902 30211 1142
rect 29817 863 30211 902
rect 30531 7542 30925 7602
rect 30531 1302 30591 7542
rect 30871 1302 30925 7542
rect 30531 1142 30925 1302
rect 30531 902 30571 1142
rect 30891 902 30925 1142
rect 30531 863 30925 902
rect 31245 7542 31639 7602
rect 31245 1302 31305 7542
rect 31585 1302 31639 7542
rect 31245 1142 31639 1302
rect 31245 902 31285 1142
rect 31605 902 31639 1142
rect 31245 863 31639 902
rect 31959 7542 32353 7602
rect 31959 1302 32019 7542
rect 32299 1302 32353 7542
rect 31959 1142 32353 1302
rect 31959 902 31999 1142
rect 32319 902 32353 1142
rect 31959 863 32353 902
rect 32673 7542 33067 7602
rect 32673 1302 32733 7542
rect 33013 1302 33067 7542
rect 32673 1142 33067 1302
rect 32673 902 32713 1142
rect 33033 902 33067 1142
rect 32673 863 33067 902
rect 33387 7542 33781 7602
rect 33387 1302 33447 7542
rect 33727 1302 33781 7542
rect 33387 1142 33781 1302
rect 33387 902 33427 1142
rect 33747 902 33781 1142
rect 33387 863 33781 902
rect 34101 7542 34495 7602
rect 34101 1302 34161 7542
rect 34441 1302 34495 7542
rect 34101 1142 34495 1302
rect 34101 902 34141 1142
rect 34461 902 34495 1142
rect 34101 863 34495 902
rect 34815 7542 35209 7602
rect 34815 1302 34875 7542
rect 35155 1302 35209 7542
rect 34815 1142 35209 1302
rect 34815 902 34855 1142
rect 35175 902 35209 1142
rect 34815 863 35209 902
rect 35529 7542 35923 7602
rect 35529 1302 35589 7542
rect 35869 1302 35923 7542
rect 35529 1142 35923 1302
rect 35529 902 35569 1142
rect 35889 902 35923 1142
rect 35529 863 35923 902
rect 36243 7542 36637 7602
rect 36243 1302 36303 7542
rect 36583 1302 36637 7542
rect 36243 1142 36637 1302
rect 36243 902 36283 1142
rect 36603 902 36637 1142
rect 36243 863 36637 902
rect 36957 7542 37351 7602
rect 36957 1302 37017 7542
rect 37297 1302 37351 7542
rect 36957 1142 37351 1302
rect 36957 902 36997 1142
rect 37317 902 37351 1142
rect 36957 863 37351 902
rect 37671 4402 38065 4462
rect 37671 1302 37731 4402
rect 38011 1302 38065 4402
rect 37671 1142 38065 1302
rect 37671 902 37711 1142
rect 38031 902 38065 1142
rect 37671 862 38065 902
rect 38385 2832 38779 2892
rect 38385 1302 38445 2832
rect 38725 1302 38779 2832
rect 38385 1142 38779 1302
rect 38385 902 38425 1142
rect 38745 902 38779 1142
rect 38385 862 38779 902
rect 40000 2100 41200 15000
rect 40000 1700 40100 2100
rect 40500 1700 41200 2100
rect 11600 100 12820 120
rect 11600 -180 12020 100
rect 12780 -180 12820 100
rect 11600 -200 12820 -180
rect 15537 -40 15931 -1
rect 8600 -420 10200 -380
rect 8600 -740 9920 -420
rect 10160 -740 10200 -420
rect 8600 -780 10200 -740
rect 8600 -1000 9600 -780
rect 3400 -1600 9600 -1000
rect 11600 -1600 12800 -200
rect 15537 -280 15577 -40
rect 15897 -280 15931 -40
rect 15537 -440 15931 -280
rect 3400 -9800 4600 -1600
rect 11600 -2000 13200 -1600
rect 12000 -2100 14802 -2000
rect 12000 -2700 12102 -2100
rect 14702 -2700 14802 -2100
rect 10702 -3152 11602 -3052
rect 10702 -3552 10802 -3152
rect 11502 -3552 11602 -3152
rect 10702 -4052 11602 -3552
rect 10302 -4192 11602 -4052
rect 5000 -6340 5600 -6310
rect 5000 -6580 5030 -6340
rect 5570 -6580 5600 -6340
rect 5000 -6700 5600 -6580
rect 5000 -6750 5800 -6700
rect 5000 -9350 5050 -6750
rect 5750 -9350 5800 -6750
rect 5000 -9400 5800 -9350
rect 10302 -9512 10442 -4192
rect 11462 -9512 11602 -4192
rect 10302 -9652 11602 -9512
rect 12000 -3340 14802 -2700
rect 12000 -9460 12142 -3340
rect 14662 -9460 14802 -3340
rect 15537 -6680 15597 -440
rect 15877 -6680 15931 -440
rect 15537 -6740 15931 -6680
rect 16251 -40 16645 -1
rect 16251 -280 16291 -40
rect 16611 -280 16645 -40
rect 16251 -440 16645 -280
rect 16251 -6680 16311 -440
rect 16591 -6680 16645 -440
rect 16251 -6740 16645 -6680
rect 16965 -40 17359 -1
rect 16965 -280 17005 -40
rect 17325 -280 17359 -40
rect 16965 -440 17359 -280
rect 16965 -6680 17025 -440
rect 17305 -6680 17359 -440
rect 16965 -6740 17359 -6680
rect 17679 -40 18073 -1
rect 17679 -280 17719 -40
rect 18039 -280 18073 -40
rect 17679 -440 18073 -280
rect 17679 -6680 17739 -440
rect 18019 -6680 18073 -440
rect 17679 -6740 18073 -6680
rect 18393 -40 18787 -1
rect 18393 -280 18433 -40
rect 18753 -280 18787 -40
rect 18393 -440 18787 -280
rect 18393 -6680 18453 -440
rect 18733 -6680 18787 -440
rect 18393 -6740 18787 -6680
rect 19107 -40 19501 -1
rect 19107 -280 19147 -40
rect 19467 -280 19501 -40
rect 19107 -440 19501 -280
rect 19107 -6680 19167 -440
rect 19447 -6680 19501 -440
rect 19107 -6740 19501 -6680
rect 19821 -40 20215 -1
rect 19821 -280 19861 -40
rect 20181 -280 20215 -40
rect 19821 -440 20215 -280
rect 19821 -6680 19881 -440
rect 20161 -6680 20215 -440
rect 19821 -6740 20215 -6680
rect 20535 -40 20929 -1
rect 20535 -280 20575 -40
rect 20895 -280 20929 -40
rect 20535 -440 20929 -280
rect 20535 -6680 20595 -440
rect 20875 -6680 20929 -440
rect 20535 -6740 20929 -6680
rect 21249 -40 21643 -1
rect 21249 -280 21289 -40
rect 21609 -280 21643 -40
rect 21249 -440 21643 -280
rect 21249 -6680 21309 -440
rect 21589 -6680 21643 -440
rect 21249 -6740 21643 -6680
rect 21963 -40 22357 -1
rect 21963 -280 22003 -40
rect 22323 -280 22357 -40
rect 21963 -440 22357 -280
rect 21963 -6680 22023 -440
rect 22303 -6680 22357 -440
rect 21963 -6740 22357 -6680
rect 22677 -40 23071 -1
rect 22677 -280 22717 -40
rect 23037 -280 23071 -40
rect 22677 -440 23071 -280
rect 22677 -6680 22737 -440
rect 23017 -6680 23071 -440
rect 22677 -6740 23071 -6680
rect 23391 -40 23785 -1
rect 23391 -280 23431 -40
rect 23751 -280 23785 -40
rect 23391 -440 23785 -280
rect 23391 -6680 23451 -440
rect 23731 -6680 23785 -440
rect 23391 -6740 23785 -6680
rect 24105 -40 24499 -1
rect 24105 -280 24145 -40
rect 24465 -280 24499 -40
rect 24105 -440 24499 -280
rect 24105 -6680 24165 -440
rect 24445 -6680 24499 -440
rect 24105 -6740 24499 -6680
rect 24819 -40 25213 -1
rect 24819 -280 24859 -40
rect 25179 -280 25213 -40
rect 24819 -440 25213 -280
rect 24819 -6680 24879 -440
rect 25159 -6680 25213 -440
rect 24819 -6740 25213 -6680
rect 25533 -40 25927 -1
rect 25533 -280 25573 -40
rect 25893 -280 25927 -40
rect 25533 -440 25927 -280
rect 25533 -6680 25593 -440
rect 25873 -6680 25927 -440
rect 25533 -6740 25927 -6680
rect 26247 -40 26641 -1
rect 26247 -280 26287 -40
rect 26607 -280 26641 -40
rect 26247 -440 26641 -280
rect 26247 -6680 26307 -440
rect 26587 -6680 26641 -440
rect 26247 -6740 26641 -6680
rect 26961 -40 27355 -1
rect 26961 -280 27001 -40
rect 27321 -280 27355 -40
rect 26961 -440 27355 -280
rect 26961 -6680 27021 -440
rect 27301 -6680 27355 -440
rect 26961 -6740 27355 -6680
rect 27675 -40 28069 -1
rect 27675 -280 27715 -40
rect 28035 -280 28069 -40
rect 27675 -440 28069 -280
rect 27675 -6680 27735 -440
rect 28015 -6680 28069 -440
rect 27675 -6740 28069 -6680
rect 28389 -40 28783 -1
rect 28389 -280 28429 -40
rect 28749 -280 28783 -40
rect 28389 -440 28783 -280
rect 28389 -6680 28449 -440
rect 28729 -6680 28783 -440
rect 28389 -6740 28783 -6680
rect 29103 -40 29497 -1
rect 29103 -280 29143 -40
rect 29463 -280 29497 -40
rect 29103 -440 29497 -280
rect 29103 -6680 29163 -440
rect 29443 -6680 29497 -440
rect 29103 -6740 29497 -6680
rect 29817 -40 30211 -1
rect 29817 -280 29857 -40
rect 30177 -280 30211 -40
rect 29817 -440 30211 -280
rect 29817 -6680 29877 -440
rect 30157 -6680 30211 -440
rect 29817 -6740 30211 -6680
rect 30531 -40 30925 -1
rect 30531 -280 30571 -40
rect 30891 -280 30925 -40
rect 30531 -440 30925 -280
rect 30531 -6680 30591 -440
rect 30871 -6680 30925 -440
rect 30531 -6740 30925 -6680
rect 31245 -40 31639 -1
rect 31245 -280 31285 -40
rect 31605 -280 31639 -40
rect 31245 -440 31639 -280
rect 31245 -6680 31305 -440
rect 31585 -6680 31639 -440
rect 31245 -6740 31639 -6680
rect 31959 -40 32353 -1
rect 31959 -280 31999 -40
rect 32319 -280 32353 -40
rect 31959 -440 32353 -280
rect 31959 -6680 32019 -440
rect 32299 -6680 32353 -440
rect 31959 -6740 32353 -6680
rect 32673 -40 33067 -1
rect 32673 -280 32713 -40
rect 33033 -280 33067 -40
rect 32673 -440 33067 -280
rect 32673 -6680 32733 -440
rect 33013 -6680 33067 -440
rect 32673 -6740 33067 -6680
rect 33387 -40 33781 -1
rect 33387 -280 33427 -40
rect 33747 -280 33781 -40
rect 33387 -440 33781 -280
rect 33387 -6680 33447 -440
rect 33727 -6680 33781 -440
rect 33387 -6740 33781 -6680
rect 34101 -40 34495 -1
rect 34101 -280 34141 -40
rect 34461 -280 34495 -40
rect 34101 -440 34495 -280
rect 34101 -6680 34161 -440
rect 34441 -6680 34495 -440
rect 34101 -6740 34495 -6680
rect 34815 -40 35209 -1
rect 34815 -280 34855 -40
rect 35175 -280 35209 -40
rect 34815 -440 35209 -280
rect 34815 -6680 34875 -440
rect 35155 -6680 35209 -440
rect 34815 -6740 35209 -6680
rect 35529 -40 35923 -1
rect 35529 -280 35569 -40
rect 35889 -280 35923 -40
rect 35529 -440 35923 -280
rect 35529 -6680 35589 -440
rect 35869 -6680 35923 -440
rect 35529 -6740 35923 -6680
rect 36243 -40 36637 -1
rect 36243 -280 36283 -40
rect 36603 -280 36637 -40
rect 36243 -440 36637 -280
rect 36243 -6680 36303 -440
rect 36583 -6680 36637 -440
rect 36243 -6740 36637 -6680
rect 36957 -40 37351 -1
rect 36957 -280 36997 -40
rect 37317 -280 37351 -40
rect 36957 -440 37351 -280
rect 36957 -6680 37017 -440
rect 37297 -6680 37351 -440
rect 36957 -6740 37351 -6680
rect 37671 -40 38065 -1
rect 37671 -280 37711 -40
rect 38031 -280 38065 -40
rect 37671 -440 38065 -280
rect 37671 -6680 37731 -440
rect 38011 -6680 38065 -440
rect 37671 -6740 38065 -6680
rect 38385 -40 38779 -1
rect 38385 -280 38425 -40
rect 38745 -280 38779 -40
rect 38385 -440 38779 -280
rect 38385 -6680 38445 -440
rect 38725 -6680 38779 -440
rect 38385 -6740 38779 -6680
rect 40000 -900 41200 1700
rect 40000 -1300 40100 -900
rect 40500 -1300 41200 -900
rect 12000 -9600 14802 -9460
rect 3400 -10400 3600 -9800
rect 4400 -10400 4600 -9800
rect 3400 -13000 4600 -10400
rect 12000 -13000 13200 -9600
rect 40000 -13000 41200 -1300
rect 43000 13700 44200 15000
rect 43000 12600 43100 13700
rect 44100 12600 44200 13700
rect 43000 -9200 44200 12600
rect 43000 -10300 43100 -9200
rect 44100 -10300 44200 -9200
rect 43000 -13000 44200 -10300
<< comment >>
rect 7997 8100 8000 12640
rect 7997 -9240 8000 -4700
<< res0p35 >>
rect 39793 973 39897 1047
rect 39793 807 39897 881
rect 39793 641 39897 715
rect 39793 475 39897 549
rect 39793 309 39897 383
rect 39793 143 39897 217
rect 39793 -23 39897 51
rect 39793 -189 39897 -115
<< res1p41 >>
rect 3121 2345 3225 2631
rect 3121 1793 3225 2079
rect 4273 1013 4377 1299
<< labels >>
rlabel metal3 1900 -9060 2000 -8860 1 CLKIN
port 6 n
rlabel metal3 1400 -9060 1520 -8860 1 LLIM
port 7 n
rlabel metal3 40500 980 40530 1040 1 B0
port 8 n
rlabel metal3 40500 820 40530 880 1 B1
port 9 n
rlabel metal3 40500 650 40530 710 1 B2
port 10 n
rlabel metal3 40500 480 40530 540 1 B3
port 11 n
rlabel metal3 40500 310 40530 370 1 B4
port 12 n
rlabel metal3 40500 150 40530 210 1 B5
port 13 n
rlabel metal3 40500 -10 40530 50 1 B6
port 14 n
rlabel metal3 40500 -180 40530 -120 1 B7
port 15 n
rlabel metal5 3400 -13000 4600 -12400 1 VHI
port 16 n
rlabel metal5 12000 -13000 13200 -12400 1 VLO
port 17 n
rlabel metal4 14800 1700 15100 2200 1 VOUT
port 18 n
rlabel metal3 12810 1600 13180 1700 1 VREFP
port 19 n
rlabel metal4 12810 1350 13180 1450 1 VREFN
port 20 n
rlabel metal3 2420 -9060 2540 -8860 1 C50
port 4 n
rlabel metal3 2240 -9060 2360 -8860 1 C100
port 5 n
rlabel metal3 2780 -9060 2900 -8860 1 IREF
port 2 n
rlabel metal3 2600 -9060 2720 -8860 1 ULIM
port 3 n
rlabel metal3 2960 -9060 3080 -8860 1 OPAEN
port 21 n
rlabel metal3 10360 1890 10450 1960 1 GP
port 22 n
rlabel metal3 10390 1150 10440 1200 1 GN
port 23 n
<< end >>
