* NGSPICE file created from sarcon_sync_flat_1.ext - technology: sky130A

.subckt sarcon_sync_flat_1 clk comp dq[0] dq[1] dq[2] dq[3] dq[4] dq[5] dq[6] dq[7]
+ last_cycle rst_n valid vccd1 vssd1
X0 a_12283_4726# _31_.A0 a_12283_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 _54_.CLK a_9494_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.1892e+14p ps=1.17526e+09u w=1e+06u l=150000u
X2 a_5322_2741# a_5172_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X3 vccd1 a_6700_5175# _43_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 vssd1 a_4043_4373# _52_.RESET_B vssd1 sky130_fd_pr__nfet_01v8 ad=8.07775e+13p pd=8.5953e+08u as=0p ps=0u w=420000u l=150000u
X5 a_4680_2223# _45_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 vssd1 a_9494_2767# _54_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 vssd1 a_9034_3855# clkbuf_0_clk.X vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 output6.A a_15175_4159# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_7458_2899# a_7775_3009# a_7733_3133# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X10 _29_.A a_5742_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_5436_3133# a_5322_2741# a_5364_3133# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 _32_.X a_12856_5737# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 vssd1 a_16727_4564# _30_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X14 vssd1 hold1.X a_2235_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X15 vccd1 a_2764_2223# a_2939_2197# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 a_2997_3133# a_2618_2767# a_2925_3133# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X18 a_14085_3861# a_13919_3861# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 a_5280_2767# a_4333_2773# a_5172_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X21 a_2489_3133# a_2011_2741# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X23 a_11650_5737# _35_.B a_11568_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 _41_.B a_7867_5814# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_11760_5175# _40_.A1 a_11902_5309# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 vssd1 a_12189_5241# a_12123_5309# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X28 vccd1 clkbuf_0_clk.X a_4605_3285# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 vssd1 a_4605_3285# _63_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 a_12715_2460# a_12559_2365# a_12860_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X31 vccd1 _63_.CLK a_4259_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X32 a_5340_2223# a_4259_2223# a_4993_2465# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X33 vccd1 a_9494_2767# _54_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 vccd1 a_9034_3855# clkbuf_0_clk.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 a_12242_3563# a_12520_3579# a_12476_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X36 a_2104_2223# _26_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X37 a_4702_2767# a_4167_2773# a_4616_3145# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X38 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X39 vccd1 fanout13.A a_9135_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X40 clkbuf_0_clk.X a_9034_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X41 a_9258_4649# _47_.B a_9176_4649# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X42 vccd1 _26_.A a_10638_4649# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X43 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X44 a_15248_4649# _28_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X45 a_13278_2589# a_12520_2491# a_12715_2460# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X46 a_1849_2223# a_1683_2223# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X47 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X48 vssd1 _63_.CLK a_1683_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X49 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X50 vccd1 a_8928_5321# a_9103_5247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X51 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X52 _63_.CLK a_4605_3285# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X53 vssd1 fanout13.A a_9135_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X54 a_7355_3311# a_6909_3311# a_7259_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X55 a_9794_2589# a_9668_2491# a_9390_2475# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X56 a_9034_3855# clk vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X57 a_13231_4564# _35_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X58 _63_.CLK a_4605_3285# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X59 a_12283_3009# _54_.CLK vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X60 a_5172_2767# a_4167_2773# a_5096_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X61 vssd1 _63_.RESET_B a_12277_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X62 vccd1 a_12559_2365# a_12520_2491# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X63 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X64 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X65 a_7692_2767# a_7255_2741# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X66 _54_.CLK a_9494_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X67 vssd1 a_9034_3855# clkbuf_0_clk.X vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X68 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X69 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X70 a_4069_4233# a_2879_3861# a_3960_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X71 a_12646_2589# a_12520_2491# a_12242_2475# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X72 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X73 vssd1 _25_.S a_13919_2775# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X74 vccd1 _40_.S a_8081_5814# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X75 a_2926_3677# a_1849_3311# a_2764_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X76 a_6791_5652# _45_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X77 a_6909_3311# a_6743_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X78 a_9863_2460# a_9707_2365# a_10008_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X79 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X80 vssd1 _63_.CLK a_6743_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X81 a_7477_3553# a_7259_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X82 dq[5] a_14471_7127# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X83 a_8013_4949# a_7847_4949# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X84 a_3300_4221# _39_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X85 a_8178_3311# _52_.RESET_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X86 vssd1 a_12715_2460# a_12646_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X87 a_5515_2197# a_5340_2223# a_5694_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X88 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X89 a_8081_5814# output6.A a_7867_5814# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X90 vccd1 a_7129_5241# a_7159_4982# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X91 vccd1 a_9034_3855# clkbuf_0_clk.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X92 a_14543_3855# _52_.RESET_B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X93 vccd1 a_10103_3476# _48_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X94 _63_.RESET_B a_9135_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X95 a_10351_4982# output3.A a_10351_5309# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X96 a_8268_5309# _40_.S vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X97 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X98 a_10426_2589# a_9668_2491# a_9863_2460# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X99 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X100 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X101 vssd1 a_15175_4159# a_15109_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X102 vccd1 a_9494_2767# _54_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X103 a_7775_3009# _54_.CLK vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X104 vccd1 _63_.RESET_B a_7255_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X105 a_2687_2741# a_2531_3009# a_2832_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X106 _52_.RESET_B a_4043_4373# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X107 a_5172_2767# a_4333_2773# a_5196_3133# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X108 vssd1 a_2531_3009# a_2492_2883# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X109 _28_.X a_13203_4982# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X110 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X111 a_12584_3855# a_12370_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X112 a_2939_2197# a_2764_2223# a_3118_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X113 dq[7] a_18059_7127# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X114 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X115 vccd1 _29_.A a_15330_4649# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X116 vccd1 a_9707_2365# a_9668_2491# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X117 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X118 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X119 a_12211_4726# a_12029_4726# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X120 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X121 a_3250_2767# a_2492_2883# a_2687_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X122 vssd1 a_5172_2767# a_5742_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X123 vccd1 a_7900_7093# dq[3] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X124 a_14653_3829# a_14435_4233# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X125 _31_.A0 a_2939_3285# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X126 vccd1 a_15015_2460# a_14946_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X127 a_11568_5737# _35_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X128 a_5502_2589# a_4425_2223# a_5340_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
R0 vccd1 _60__15.HI sky130_fd_pr__res_generic_po w=480000u l=45000u
X129 clkbuf_0_clk.X a_9034_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X130 _54_.CLK a_9494_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X131 vssd1 a_9034_3855# clkbuf_0_clk.X vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X132 a_4993_2465# a_4775_2223# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X133 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X134 a_8325_4373# _41_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X135 a_4333_2773# a_4167_2773# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X136 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X137 a_15015_2460# a_14859_2365# a_15160_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X138 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X139 dq[3] a_7900_7093# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X140 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X141 a_12200_3855# a_11763_3829# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X142 vccd1 a_9135_3311# _63_.RESET_B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X143 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X144 vccd1 clkbuf_0_clk.X a_4605_3285# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X145 vssd1 a_4605_3285# _63_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X146 vccd1 _35_.A a_13278_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X147 vssd1 _52_.RESET_B a_2461_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X148 a_15578_2589# a_14820_2491# a_15015_2460# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X149 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X150 vccd1 clk a_9034_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X151 vccd1 a_4993_2465# a_4883_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X152 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X153 vccd1 a_4605_3285# _63_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X154 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X155 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X156 a_3657_4221# a_3613_3829# a_3491_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X157 a_12039_3285# a_12242_3563# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X158 vccd1 a_4036_7093# dq[1] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X159 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X160 a_6085_4551# _34_.S vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X161 vccd1 a_2489_4551# hold1.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X162 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X163 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X164 vssd1 _63_.RESET_B a_14577_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X165 vccd1 a_14859_2365# a_14820_2491# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X166 a_7795_5814# a_7613_5814# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X167 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X168 _63_.CLK a_4605_3285# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X169 vccd1 _63_.RESET_B a_12860_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X170 dq[1] a_4036_7093# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X171 a_6700_5175# output5.A a_6842_4982# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X172 a_12504_4399# _40_.A1 a_12283_4726# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X173 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X174 a_13278_3677# a_12559_3453# a_12715_3548# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X175 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X176 a_6791_5652# _45_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X177 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X178 vccd1 _52_.RESET_B a_11763_3829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X179 a_12283_4097# _54_.CLK vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X180 a_15175_4159# a_15000_4233# a_15354_4221# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X181 a_14946_2589# a_14820_2491# a_14542_2475# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X182 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X183 a_4043_4373# fanout13.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X184 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X185 a_12476_2589# a_12039_2197# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X186 a_6842_4982# _63_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X187 vssd1 _52_.RESET_B a_5037_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X188 vssd1 a_5692_7093# dq[2] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X189 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X190 _47_.B a_7959_3894# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X191 clkbuf_0_clk.X a_9034_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X192 vssd1 a_10103_3476# _48_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X193 a_12189_5241# _34_.S vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X194 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X195 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X196 vccd1 a_5322_2741# a_5280_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X197 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X198 _54_.CLK a_9494_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X199 a_2687_2741# a_2492_2883# a_2997_3133# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X200 vccd1 _54_.CLK a_13919_3861# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X201 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X202 vssd1 a_4043_4373# _52_.RESET_B vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X203 vccd1 a_15000_4233# a_15175_4159# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X204 a_11966_2899# a_12244_2883# a_12200_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X205 a_13417_4982# _28_.A0 a_13203_4982# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X206 a_4122_3855# a_3045_3861# a_3960_4233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X207 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X208 a_4521_2767# _60__15.LO vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X209 dq[0] a_1644_7093# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X210 a_12953_2223# _63_.RESET_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X211 a_2214_2899# a_2531_3009# a_2489_3133# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X212 vssd1 a_4605_3285# _63_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X213 a_3521_4917# a_3303_5321# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X214 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X215 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X216 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X217 vccd1 a_2417_3553# a_2307_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X218 a_12559_3453# _54_.CLK vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X219 vssd1 a_8325_4373# a_8259_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X220 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X221 vssd1 _35_.A a_13278_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X222 vccd1 _63_.RESET_B a_12039_2197# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X223 a_8154_6147# _41_.B a_8072_6147# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X224 vccd1 a_4792_2741# a_4702_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X225 _52_.RESET_B a_4043_4373# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X226 _63_.CLK a_4605_3285# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X227 vssd1 _48_.X a_8494_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X228 clkbuf_0_clk.X a_9034_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X229 a_2417_2465# a_2199_2223# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X230 _42_.X a_11343_4399# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X231 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X232 vccd1 a_12715_3548# a_12646_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X233 a_2873_3311# a_1683_3311# a_2764_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X234 _49_.D a_10975_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X235 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X236 a_2764_2223# a_1849_2223# a_2417_2465# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
D0 vssd1 rst_n sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
X237 a_4605_3285# clkbuf_0_clk.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X238 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X239 a_8241_3133# a_7862_2767# a_8169_3133# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X240 vssd1 _32_.A a_13424_5309# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X241 vssd1 a_7255_2741# output4.A vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X242 a_7999_3285# _52_.RESET_B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X243 _35_.X a_11568_5737# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X244 a_4043_5247# _52_.RESET_B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X245 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X246 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X247 vssd1 a_9034_3855# clkbuf_0_clk.X vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X248 _54_.CLK a_9494_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X249 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X250 a_10572_5309# _40_.A1 a_10351_4982# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X251 vssd1 a_11760_5175# _35_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X252 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X253 a_11763_3829# a_11966_3987# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X254 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X255 a_3045_3861# a_2879_3861# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X256 a_7477_3553# a_7259_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X257 dq[2] a_5692_7093# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X258 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X259 a_3521_4917# a_3303_5321# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X260 vccd1 _26_.A a_8173_3894# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X261 vccd1 clk a_9034_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X262 a_12559_2365# _54_.CLK vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X263 a_13002_2767# a_12283_3009# a_12439_2741# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X264 _54_.CLK a_9494_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X265 vccd1 a_4605_3285# _63_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X266 a_7900_7093# output6.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X267 a_4043_5247# a_3868_5321# a_4222_5309# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X268 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X269 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X270 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X271 _25_.X a_10351_4982# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X272 a_12219_4982# _40_.A1 a_11760_5175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X273 a_7824_3311# a_6909_3311# a_7477_3553# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X274 vccd1 a_12039_2197# _41_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X275 _63_.Q a_9103_5247# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X276 vccd1 a_16727_4564# _30_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X277 a_8173_3894# output4.A a_7959_3894# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X278 vccd1 a_9034_3855# clkbuf_0_clk.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X279 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X280 _63_.CLK a_4605_3285# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X281 a_3868_5321# a_2787_4949# a_3521_4917# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X282 vccd1 a_4043_5247# a_4030_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X283 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X284 a_12283_4726# _40_.A1 a_12211_4726# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X285 a_14776_2589# a_14339_2197# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X286 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X287 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X288 vccd1 _63_.RESET_B a_10008_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X289 vccd1 _26_.A a_17507_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X290 a_4871_2223# a_4425_2223# a_4775_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X291 a_12001_3133# a_11966_2899# a_11763_2741# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X292 vccd1 _52_.RESET_B a_2011_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X293 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X294 a_12677_3133# _63_.RESET_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X295 a_12370_2767# a_12283_3009# a_11966_2899# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X296 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X297 a_12277_2223# a_12242_2475# a_12039_2197# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X298 a_16083_4564# _32_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X299 vssd1 _49_.D a_13002_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X300 a_4605_3285# clkbuf_0_clk.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X301 vccd1 a_13919_2775# valid vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X302 a_8013_4949# a_7847_4949# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X303 vssd1 _26_.A a_17507_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X304 a_12370_2767# a_12244_2883# a_11966_2899# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X305 clkbuf_0_clk.X a_9034_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X306 a_6085_4551# _37_.X a_6248_4649# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X307 a_9494_2767# clkbuf_0_clk.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X308 a_2295_2223# a_1849_2223# a_2199_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X309 vccd1 _32_.A a_13002_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X310 vssd1 a_7931_2741# a_7862_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X311 vssd1 a_14471_7127# dq[5] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X312 a_7259_3311# a_6743_3311# a_7164_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X313 a_7775_3009# _54_.CLK vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X314 a_13231_4564# _35_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X315 vccd1 a_4605_3285# _63_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X316 a_3960_4233# a_3045_3861# a_3613_3829# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X317 vccd1 _63_.RESET_B a_14339_2197# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X318 a_5694_2223# _52_.RESET_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X319 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X320 _49_.D a_10975_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X321 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X322 vssd1 a_10055_7119# _40_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X323 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X324 a_4792_2741# a_4616_3145# a_4936_3133# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X325 _41_.X a_8072_6147# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X326 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X327 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X328 vccd1 _63_.RESET_B a_12584_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X329 a_7867_5814# _40_.A1 a_7795_5814# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X330 a_13203_4982# _28_.A0 a_13203_5309# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X331 vccd1 a_11763_3829# output3.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X332 vccd1 a_12439_3829# a_12370_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X333 vssd1 _63_.RESET_B a_9425_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X334 vccd1 _63_.RESET_B a_15160_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X335 a_3303_5321# a_2787_4949# a_3208_5309# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X336 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X337 a_3118_2223# _52_.RESET_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X338 vccd1 a_9494_2767# _54_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X339 last_cycle a_17507_2223# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X340 a_4726_3145# a_4333_2773# a_4616_3145# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X341 a_5692_7093# output5.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X342 vccd1 a_2764_3311# a_2939_3285# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X343 vssd1 a_9494_2767# _54_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X344 a_9037_5321# a_7847_4949# a_8928_5321# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X345 _52_.RESET_B a_4043_4373# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X346 _26_.X a_10556_4649# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X347 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X348 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X349 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X350 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X351 a_7887_3894# a_7705_3894# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X352 dq[6] a_16863_7127# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X353 a_12715_3548# a_12559_3453# a_12860_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X354 vssd1 _40_.S a_8088_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X355 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X356 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X357 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X358 vssd1 _26_.A a_8180_4221# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X359 a_7867_5814# output6.A a_7867_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X360 a_8459_5321# a_8013_4949# a_8363_5321# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X361 a_14653_3829# a_14435_4233# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X362 a_2104_3311# _33_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X363 valid a_13919_2775# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X364 vccd1 _34_.A0 a_14471_7127# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X365 a_8268_5309# _40_.S vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X366 vssd1 clkbuf_0_clk.X a_4605_3285# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X367 _28_.A0 a_7999_3285# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X368 _54_.CLK a_9494_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X369 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X370 a_14859_2365# _54_.CLK vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X371 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X372 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X373 vccd1 _35_.A a_12029_4726# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X374 a_1849_3311# a_1683_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X375 vssd1 _63_.CLK a_1683_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X376 a_2417_3553# a_2199_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X377 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X378 a_13278_3677# a_12520_3579# a_12715_3548# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X379 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X380 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X381 a_2953_4949# a_2787_4949# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X382 a_16727_4564# _30_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X383 vccd1 a_14339_2197# _32_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X384 a_8625_5309# a_8581_4917# a_8459_5321# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X385 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X386 vccd1 a_8325_4373# a_8355_4726# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X387 a_3491_4233# a_3045_3861# a_3395_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X388 a_9390_2475# a_9707_2365# a_9665_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X389 a_12283_4097# _54_.CLK vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X390 vccd1 a_17507_2223# last_cycle vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X391 vccd1 a_12559_3453# a_12520_3579# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X392 vssd1 _63_.RESET_B a_12277_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X393 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X394 vccd1 a_18059_7127# dq[7] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X395 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X396 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X397 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X398 _63_.CLK a_4605_3285# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X399 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X400 vccd1 _63_.CLK a_4167_2773# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X401 vssd1 a_2687_2741# a_2618_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X402 a_12715_2460# a_12520_2491# a_13025_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X403 a_14577_2223# a_14542_2475# a_14339_2197# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X404 vccd1 a_6085_4551# _38_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X405 vssd1 clkbuf_0_clk.X a_9494_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X406 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X407 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X408 a_12856_5737# _32_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X409 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X410 vssd1 _54_.CLK a_13919_3861# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X411 a_12646_3677# a_12520_3579# a_12242_3563# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X412 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X413 vccd1 _40_.S a_6958_4649# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X414 a_12242_2475# a_12559_2365# a_12517_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X415 vssd1 _63_.Q a_3250_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X416 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X417 a_15354_4221# _52_.RESET_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X418 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X419 a_7259_3311# a_6909_3311# a_7164_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X420 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X421 a_8325_4373# _41_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X422 a_3303_5321# a_2953_4949# a_3208_5309# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X423 vssd1 _63_.CLK a_4259_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X424 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X425 _29_.A a_5742_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X426 vssd1 a_12715_3548# a_12646_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X427 _30_.A a_15248_4649# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X428 output6.A a_15175_4159# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X429 a_9494_2767# clkbuf_0_clk.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X430 vccd1 _40_.S a_7613_5814# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X431 clkbuf_0_clk.X a_9034_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X432 a_8076_2767# a_7862_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X433 vccd1 a_4605_3285# _63_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X434 a_7367_3677# a_6743_3311# a_7259_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X435 vssd1 a_2011_2741# _26_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X436 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X437 a_1849_2223# a_1683_2223# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X438 a_12439_2741# a_12283_3009# a_12584_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X439 a_3411_4943# a_2787_4949# a_3303_5321# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X440 a_10279_4982# a_10097_4982# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X441 vccd1 a_12263_7127# dq[4] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X442 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X443 a_9176_4649# _47_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X444 a_2939_3285# a_2764_3311# a_3118_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X445 vccd1 a_2939_2197# a_2926_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X446 _32_.B a_12283_4726# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X447 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X448 vccd1 a_4043_4373# _52_.RESET_B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X449 a_10638_4649# _25_.X a_10556_4649# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X450 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X451 a_13002_2767# a_12244_2883# a_12439_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X452 vssd1 a_12559_2365# a_12520_2491# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X453 vssd1 _63_.RESET_B a_12001_3133# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X454 a_7458_2899# a_7736_2883# a_7692_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X455 _34_.A0 a_4043_5247# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X456 a_9624_2589# a_9187_2197# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X457 dq[4] a_12263_7127# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X458 a_12749_3133# a_12370_2767# a_12677_3133# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X459 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X460 vccd1 a_9494_2767# _54_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X461 _45_.A a_6876_4649# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X462 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X463 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X464 _52_.RESET_B a_4043_4373# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X465 a_8259_4399# _37_.A0 a_7896_4551# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X466 a_3300_4221# _39_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X467 a_6909_3311# a_6743_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X468 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X469 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X470 a_3045_3861# a_2879_3861# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X471 a_5515_2197# _52_.RESET_B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X472 vccd1 _32_.A a_12938_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X473 a_9090_4943# a_8013_4949# a_8928_5321# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X474 vccd1 a_7896_4551# _37_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X475 a_4792_2741# _52_.RESET_B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X476 vssd1 a_9135_3311# _63_.RESET_B vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X477 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X478 vssd1 a_9103_5247# a_9037_5321# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X479 _42_.X a_11343_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X480 a_9034_3855# clk vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X481 vssd1 clkbuf_0_clk.X a_4605_3285# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X482 _54_.CLK a_9494_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X483 vccd1 _35_.A a_11650_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X484 vccd1 _32_.A a_13417_4982# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X485 vssd1 a_4605_3285# _63_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X486 vccd1 _63_.RESET_B a_9187_2197# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X487 a_2307_2589# _52_.RESET_B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X488 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X489 vssd1 _28_.A0 a_18059_7127# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X490 a_13424_5309# _40_.A1 a_13203_4982# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X491 vssd1 a_2843_4373# a_2585_4373# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X492 a_2939_2197# _52_.RESET_B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X493 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X494 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X495 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X496 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X497 a_9707_2365# _54_.CLK vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X498 a_4222_5309# _52_.RESET_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X499 vccd1 a_8581_4917# a_8471_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X500 vssd1 a_9707_2365# a_9668_2491# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X501 a_15015_2460# a_14820_2491# a_15325_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X502 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X503 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X504 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X505 a_12497_4726# _31_.A0 a_12283_4726# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X506 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X507 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X508 a_12476_3677# a_12039_3285# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X509 vccd1 a_5515_2197# a_5502_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X510 vssd1 a_2939_2197# a_2873_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X511 a_4616_3145# a_4333_2773# a_4521_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X512 a_2832_2767# a_2618_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X513 vccd1 _63_.Q a_9258_4649# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X514 a_14340_4221# _42_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X515 a_14542_2475# a_14859_2365# a_14817_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X516 _28_.X a_13203_4982# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X517 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X518 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X519 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X520 vssd1 a_9494_2767# _54_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X521 vssd1 clkbuf_0_clk.X a_9494_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X522 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X523 vssd1 a_9034_3855# clkbuf_0_clk.X vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X524 a_2489_4551# a_2585_4373# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X525 a_12439_2741# a_12244_2883# a_12749_3133# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X526 a_7959_3894# _40_.A1 a_7887_3894# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X527 _63_.CLK a_4605_3285# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X528 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X529 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X530 a_7367_3677# _52_.RESET_B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X531 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X532 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X533 fanout13.A a_2235_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X534 a_11966_3987# a_12244_3971# a_12200_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X535 a_15000_4233# a_13919_3861# a_14653_3829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X536 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X537 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X538 a_12953_3311# _63_.RESET_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X539 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X540 vssd1 _37_.A0 a_12263_7127# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X541 a_6700_5175# _40_.A1 a_6842_5309# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X542 vssd1 a_7129_5241# a_7063_5309# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X543 a_3977_5321# a_2787_4949# a_3868_5321# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X544 clkbuf_0_clk.X a_9034_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X545 clkbuf_0_clk.X a_9034_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X546 a_12860_2589# a_12646_2589# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X547 a_3503_3855# _52_.RESET_B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X548 a_4775_2223# a_4259_2223# a_4680_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X549 a_7862_2767# a_7775_3009# a_7458_2899# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X550 vccd1 _63_.RESET_B a_12039_3285# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X551 vssd1 _63_.RESET_B a_8625_5309# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X552 vccd1 a_9187_2197# _40_.S vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X553 vssd1 a_4135_4159# a_4069_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X554 a_4135_4159# _52_.RESET_B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X555 vssd1 a_7999_3285# a_7933_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X556 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X557 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X558 a_16083_4564# _32_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X559 a_2417_3553# a_2199_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X560 a_7862_2767# a_7736_2883# a_7458_2899# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X561 vssd1 a_14859_2365# a_14820_2491# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X562 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X563 vccd1 a_7931_2741# a_7862_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X564 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X565 vccd1 a_4043_4373# _52_.RESET_B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X566 vssd1 a_13231_4564# _52_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X567 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X568 vccd1 _48_.X a_8494_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X569 a_5322_2741# a_5172_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=540000u l=150000u
X570 vccd1 _63_.CLK a_7847_4949# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X571 a_2199_2223# a_1683_2223# a_2104_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X572 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X573 _47_.X a_9176_4649# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X574 a_12283_4399# a_12029_4726# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X575 a_2764_3311# a_1849_3311# a_2417_3553# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X576 a_9425_2223# a_9390_2475# a_9187_2197# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X577 vccd1 _52_.RESET_B a_5172_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X578 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X579 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X580 vssd1 a_16863_7127# dq[6] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X581 a_3613_3829# a_3395_4233# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X582 a_7164_3311# _30_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X583 _41_.B a_7867_5814# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X584 vccd1 a_9034_3855# clkbuf_0_clk.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X585 a_4605_3285# clkbuf_0_clk.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X586 vccd1 a_9494_2767# _54_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X587 vssd1 a_9494_2767# _54_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X588 dq[7] a_18059_7127# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X589 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X590 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X591 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X592 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X593 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X594 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X595 a_8038_4726# _41_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X596 vccd1 a_7999_3285# a_7986_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X597 a_2531_3009# _63_.CLK vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X598 a_4521_2767# _60__15.LO vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X599 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X600 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X601 a_8928_5321# a_8013_4949# a_8581_4917# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X602 a_12123_5309# _34_.A0 a_11760_5175# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X603 vccd1 a_6791_5652# _45_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X604 a_11902_5309# _34_.S vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X605 vccd1 a_4135_4159# a_4122_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X606 vssd1 a_1644_7093# dq[0] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X607 vssd1 a_15015_2460# a_14946_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X608 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X609 a_2953_4949# a_2787_4949# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X610 _47_.B a_7959_3894# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X611 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X612 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X613 a_10008_2589# a_9794_2589# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X614 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X615 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X616 a_13002_3855# a_12283_4097# a_12439_3829# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X617 a_4993_2465# a_4775_2223# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X618 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X619 a_12559_3453# _54_.CLK vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X620 output5.A a_5515_2197# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X621 clkbuf_0_clk.X a_9034_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X622 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X623 dq[3] a_7900_7093# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X624 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X625 vssd1 a_4605_3285# _63_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X626 vccd1 a_12039_3285# _34_.S vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X627 vssd1 _63_.CLK a_4167_2773# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X628 a_7896_4551# _40_.A1 a_8038_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X629 a_5340_2223# a_4425_2223# a_4993_2465# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X630 _54_.CLK a_9494_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X631 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X632 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X633 vssd1 a_12039_2197# _41_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X634 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X635 a_8088_5487# _40_.A1 a_7867_5814# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X636 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X637 a_12001_4221# a_11966_3987# a_11763_3829# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X638 a_7867_5487# a_7613_5814# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X639 vssd1 _52_.RESET_B a_3657_4221# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X640 a_12677_4221# _52_.RESET_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X641 _25_.S a_2939_2197# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X642 a_7959_4221# a_7705_3894# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X643 a_12370_3855# a_12283_4097# a_11966_3987# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X644 a_15162_3855# a_14085_3861# a_15000_4233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X645 vccd1 a_12283_3009# a_12244_2883# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X646 a_12277_3311# a_12242_3563# a_12039_3285# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X647 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X648 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X649 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X650 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X651 _32_.X a_12856_5737# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X652 a_12370_3855# a_12244_3971# a_11966_3987# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X653 vccd1 a_3868_5321# a_4043_5247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X654 a_6699_4074# _38_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X655 vssd1 a_9034_3855# clkbuf_0_clk.X vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X656 vccd1 a_9034_3855# clkbuf_0_clk.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X657 a_11966_2899# a_12283_3009# a_12241_3133# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X658 vssd1 a_9494_2767# _54_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X659 dq[1] a_4036_7093# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X660 a_16727_4564# _30_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
R1 _60__15.LO vssd1 sky130_fd_pr__res_generic_po w=480000u l=45000u
X661 a_2295_3311# a_1849_3311# a_2199_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X662 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X663 a_2214_2899# a_2492_2883# a_2448_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X664 vccd1 _49_.D a_13002_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X665 a_3395_4233# a_2879_3861# a_3300_4221# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X666 vccd1 _63_.CLK a_2879_3861# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X667 _63_.CLK a_4605_3285# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X668 a_9665_2223# a_9187_2197# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X669 a_15160_2589# a_14946_2589# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X670 a_4775_2223# a_4425_2223# a_4680_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X671 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X672 vccd1 a_14653_3829# a_14543_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X673 vccd1 a_5692_7093# dq[2] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X674 vssd1 a_4605_3285# _63_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X675 a_10101_2223# _63_.RESET_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X676 vccd1 a_7255_2741# output4.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X677 a_10351_5309# a_10097_4982# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X678 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X679 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X680 vssd1 _35_.A a_12029_4726# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X681 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X682 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X683 vccd1 _25_.S a_13919_2775# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X684 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X685 vssd1 _26_.A a_10556_4649# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X686 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X687 a_9034_3855# clk vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X688 a_12646_2589# a_12559_2365# a_12242_2475# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X689 vssd1 _41_.A a_8072_6147# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X690 vccd1 _52_.RESET_B a_12584_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X691 a_7986_3677# a_6909_3311# a_7824_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X692 a_13025_2223# a_12646_2589# a_12953_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X693 a_4883_2589# a_4259_2223# a_4775_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X694 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X695 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X696 vccd1 a_11760_5175# _35_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X697 a_12517_2223# a_12039_2197# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X698 a_2199_2223# a_1849_2223# a_2104_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X699 dq[0] a_1644_7093# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X700 vccd1 a_10055_7119# _40_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X701 _54_.CLK a_9494_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X702 a_3565_5309# a_3521_4917# a_3399_5321# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X703 a_3118_3311# _52_.RESET_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X704 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X705 vccd1 _41_.A a_8154_6147# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X706 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X707 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X708 vssd1 a_6791_5652# _45_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X709 vccd1 a_5172_2767# a_5742_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X710 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X711 a_3208_5309# _52_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X712 a_13131_4982# a_12949_4982# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X713 fanout13.A a_2235_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X714 a_2307_2589# a_1683_2223# a_2199_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X715 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X716 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X717 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X718 vssd1 _32_.A a_12949_4982# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X719 vssd1 a_9034_3855# clkbuf_0_clk.X vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X720 vccd1 a_9034_3855# clkbuf_0_clk.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X721 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X722 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X723 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X724 a_15253_2223# _63_.RESET_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X725 vssd1 _63_.RESET_B a_7493_3133# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X726 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X727 _28_.A0 a_7999_3285# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X728 vssd1 a_9494_2767# _54_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X729 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X730 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X731 a_5692_7093# output5.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X732 vssd1 _40_.S a_7613_5814# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X733 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X734 a_6248_4649# _34_.S vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X735 a_6958_4649# _43_.X a_6876_4649# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X736 a_4425_2223# a_4259_2223# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X737 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X738 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X739 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X740 vccd1 a_2843_4373# a_2585_4373# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X741 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X742 vssd1 a_14339_2197# _32_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X743 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X744 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X745 a_2618_2767# a_2531_3009# a_2214_2899# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X746 a_4036_7093# output4.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X747 a_3395_4233# a_3045_3861# a_3300_4221# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X748 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X749 _54_.CLK a_9494_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X750 clkbuf_0_clk.X a_9034_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X751 a_12715_3548# a_12520_3579# a_13025_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X752 vssd1 _41_.X a_11343_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X753 vssd1 a_17507_2223# last_cycle vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X754 vssd1 _29_.A a_15248_4649# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X755 vccd1 _41_.A a_10426_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X756 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X757 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X758 a_3503_3855# a_2879_3861# a_3395_4233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X759 vccd1 _26_.X a_10975_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X760 vccd1 a_2687_2741# a_2618_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X761 a_12242_3563# a_12559_3453# a_12517_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X762 a_7129_5241# _63_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X763 vssd1 _25_.S a_10097_4982# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X764 a_2489_4551# a_2585_4373# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X765 vccd1 a_12189_5241# a_12219_4982# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X766 vssd1 _31_.A0 a_16863_7127# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X767 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X768 vssd1 _52_.RESET_B a_5436_3133# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X769 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X770 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X771 vssd1 clk a_9034_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X772 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X773 vccd1 _63_.Q a_3250_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X774 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X775 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X776 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X777 _54_.CLK a_9494_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X778 a_1644_7093# output3.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X779 _37_.A0 a_4135_4159# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X780 a_7959_3894# output4.A a_7959_4221# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X781 a_12241_3133# a_11763_2741# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X782 vssd1 a_11763_2741# _35_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X783 a_12439_3829# a_12283_4097# a_12584_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X784 a_1849_3311# a_1683_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X785 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X786 a_2011_2741# a_2214_2899# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X787 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X788 _63_.CLK a_4605_3285# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X789 a_14946_2589# a_14859_2365# a_14542_2475# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X790 vssd1 a_6700_5175# _43_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X791 vssd1 a_4605_3285# _63_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X792 a_10426_2589# a_9707_2365# a_9863_2460# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X793 a_4030_4943# a_2953_4949# a_3868_5321# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X794 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X795 vccd1 a_2939_3285# a_2926_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X796 a_14817_2223# a_14339_2197# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X797 vssd1 comp a_10055_7119# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X798 a_2843_4373# rst_n vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X799 valid a_13919_2775# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X800 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X801 vssd1 _63_.CLK a_7847_4949# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X802 a_13002_3855# a_12244_3971# a_12439_3829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X803 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X804 vccd1 a_14471_7127# dq[5] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X805 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X806 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X807 vssd1 a_2489_4551# hold1.X vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X808 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X809 vssd1 _52_.RESET_B a_12001_4221# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X810 vssd1 a_12559_3453# a_12520_3579# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X811 a_5096_2767# a_4616_3145# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X812 clkbuf_0_clk.X a_9034_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X813 a_12749_4221# a_12370_3855# a_12677_4221# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X814 dq[5] a_14471_7127# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X815 a_7159_4982# _40_.A1 a_6700_5175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X816 a_6699_4074# _38_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X817 clkbuf_0_clk.X a_9034_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X818 vccd1 a_4605_3285# _63_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X819 vccd1 a_12715_2460# a_12646_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X820 a_15109_4233# a_13919_3861# a_15000_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X821 a_2531_3009# _63_.CLK vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X822 vccd1 a_3521_4917# a_3411_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X823 _41_.X a_8072_6147# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X824 _35_.X a_11568_5737# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X825 a_4043_4373# fanout13.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X826 vccd1 _35_.A a_12497_4726# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X827 a_3250_2767# a_2531_3009# a_2687_2741# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X828 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X829 vssd1 a_16083_4564# _33_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X830 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X831 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X832 a_4680_2223# _45_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X833 vssd1 _41_.A a_10426_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X834 vccd1 a_9034_3855# clkbuf_0_clk.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X835 a_14531_4233# a_14085_3861# a_14435_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X836 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X837 _40_.A1 a_10055_7119# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X838 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X839 a_8471_4943# _63_.RESET_B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X840 a_3613_3829# a_3395_4233# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X841 a_7933_3311# a_6743_3311# a_7824_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X842 a_2461_2223# a_2417_2465# a_2295_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X843 vssd1 a_7900_7093# dq[3] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X844 vccd1 a_13231_4564# _52_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X845 a_10173_2223# a_9794_2589# a_10101_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X846 a_2307_3677# _52_.RESET_B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X847 vssd1 a_4792_2741# a_4726_3145# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X848 a_2249_3133# a_2214_2899# a_2011_2741# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X849 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X850 a_15330_4649# _28_.X a_15248_4649# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X851 vccd1 _63_.CLK a_1683_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X852 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X853 a_11760_5175# _34_.A0 a_11902_4982# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X854 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X855 a_2104_2223# _26_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X856 a_2939_3285# _52_.RESET_B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X857 a_9103_5247# _63_.RESET_B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X858 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X859 vssd1 _26_.X a_10975_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X860 vssd1 a_12439_2741# a_12370_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X861 _54_.CLK a_9494_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X862 a_2764_2223# a_1683_2223# a_2417_2465# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X863 a_11902_4982# _34_.S vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X864 vssd1 a_12283_3009# a_12244_2883# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X865 vccd1 a_2011_2741# _26_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X866 vssd1 _52_.RESET_B a_3565_5309# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X867 a_9390_2475# a_9668_2491# a_9624_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X868 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X869 vssd1 a_2939_3285# a_2873_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X870 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X871 vccd1 a_6699_4074# _39_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X872 a_9103_5247# a_8928_5321# a_9282_5309# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X873 vssd1 _37_.X a_6085_4551# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X874 _54_.CLK a_9494_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X875 vccd1 _28_.A0 a_18059_7127# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X876 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X877 a_12439_3829# a_12244_3971# a_12749_4221# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X878 vccd1 _63_.CLK a_2787_4949# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X879 vssd1 _63_.CLK a_2879_3861# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X880 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X881 vccd1 a_4605_3285# _63_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X882 a_7521_3311# a_7477_3553# a_7355_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X883 vssd1 a_4036_7093# dq[1] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X884 vccd1 _63_.CLK a_6743_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X885 _63_.CLK a_4605_3285# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X886 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X887 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X888 _34_.A0 a_4043_5247# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X889 vccd1 a_5340_2223# a_5515_2197# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X890 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X891 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X892 vssd1 _25_.S a_10572_5309# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X893 vccd1 a_9103_5247# a_9090_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X894 a_8038_4399# _41_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X895 vssd1 clk a_9034_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X896 a_12242_2475# a_12520_2491# a_12476_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X897 a_7896_4551# _37_.A0 a_8038_4726# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X898 a_7824_3311# a_6743_3311# a_7477_3553# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X899 a_9494_2767# clkbuf_0_clk.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X900 a_12860_3677# a_12646_3677# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X901 a_14697_4221# a_14653_3829# a_14531_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X902 a_3868_5321# a_2953_4949# a_3521_4917# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X903 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X904 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X905 vccd1 a_7775_3009# a_7736_2883# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X906 a_7255_2741# a_7458_2899# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X907 a_12938_5737# _32_.B a_12856_5737# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X908 vssd1 a_9034_3855# clkbuf_0_clk.X vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X909 _63_.CLK a_4605_3285# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X910 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X911 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X912 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X913 vssd1 a_5515_2197# a_5449_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X914 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X915 vssd1 a_9187_2197# _40_.S vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X916 a_5037_2223# a_4993_2465# a_4871_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X917 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X918 a_9707_2365# _54_.CLK vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X919 vssd1 _52_.RESET_B a_2249_3133# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X920 a_13203_5309# a_12949_4982# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X921 a_14340_4221# _42_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X922 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X923 a_2199_3311# a_1683_3311# a_2104_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X924 vccd1 _37_.A0 a_12263_7127# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X925 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X926 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X927 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X928 a_10351_4982# _40_.A1 a_10279_4982# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X929 clkbuf_0_clk.X a_9034_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X930 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X931 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X932 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X933 vccd1 a_9494_2767# _54_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X934 a_8494_2767# a_7775_3009# a_7931_2741# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X935 vccd1 _26_.A a_7705_3894# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X936 a_2926_2589# a_1849_2223# a_2764_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X937 dq[4] a_12263_7127# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X938 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X939 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X940 a_8363_5321# a_7847_4949# a_8268_5309# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X941 a_4135_4159# a_3960_4233# a_4314_4221# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X942 a_8180_4221# _40_.A1 a_7959_3894# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X943 _63_.RESET_B a_9135_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X944 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X945 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X946 a_2417_2465# a_2199_2223# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X947 vccd1 a_7824_3311# a_7999_3285# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X948 vssd1 a_9863_2460# a_9794_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X949 a_9794_2589# a_9707_2365# a_9390_2475# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X950 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X951 output5.A a_5515_2197# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X952 a_8169_3133# _63_.RESET_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X953 a_7493_3133# a_7458_2899# a_7255_2741# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X954 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X955 vccd1 a_3960_4233# a_4135_4159# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X956 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X957 vccd1 _32_.A a_12949_4982# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X958 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X959 a_7164_3311# _30_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X960 vssd1 a_12039_3285# _34_.S vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X961 a_12584_2767# a_12370_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X962 vssd1 a_9494_2767# _54_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X963 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X964 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X965 a_3399_5321# a_2953_4949# a_3303_5321# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X966 a_3208_5309# _52_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X967 _31_.A0 a_2939_3285# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X968 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X969 vccd1 a_12283_4097# a_12244_3971# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X970 _25_.S a_2939_2197# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X971 dq[2] a_5692_7093# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X972 vccd1 clkbuf_0_clk.X a_9494_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X973 a_11966_3987# a_12283_4097# a_12241_4221# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X974 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X975 _54_.CLK a_9494_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X976 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X977 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X978 _26_.X a_10556_4649# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X979 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X980 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X981 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X982 a_15175_4159# _52_.RESET_B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X983 vccd1 a_4605_3285# _63_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X984 a_14542_2475# a_14820_2491# a_14776_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X985 a_9187_2197# a_9390_2475# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X986 a_14085_3861# a_13919_3861# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X987 a_12200_2767# a_11763_2741# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X988 a_4616_3145# a_4167_2773# a_4521_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X989 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X990 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X991 vccd1 _63_.RESET_B a_8076_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X992 a_3960_4233# a_2879_3861# a_3613_3829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X993 vccd1 _34_.S a_13278_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X994 vssd1 _52_.RESET_B a_2461_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X995 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X996 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X997 vccd1 _41_.X a_11343_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X998 _63_.CLK a_4605_3285# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X999 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1000 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1001 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X1002 a_9494_2767# clkbuf_0_clk.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1003 a_7129_5241# _63_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1004 a_12646_3677# a_12559_3453# a_12242_3563# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1005 vccd1 _25_.S a_10097_4982# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1006 _32_.B a_12283_4726# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1007 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1008 a_13025_3311# a_12646_3677# a_12953_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1009 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1010 a_2843_4373# rst_n vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1011 a_12039_2197# a_12242_2475# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1012 a_12517_3311# a_12039_3285# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1013 vssd1 a_6699_4074# _39_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1014 _63_.CLK a_4605_3285# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1015 a_2199_3311# a_1849_3311# a_2104_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1016 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1017 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1018 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1019 a_8363_5321# a_8013_4949# a_8268_5309# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1020 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1021 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1022 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1023 vccd1 _63_.RESET_B a_12860_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1024 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1025 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1026 a_13278_2589# a_12559_2365# a_12715_2460# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
D1 vssd1 comp sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
X1027 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1028 _45_.A a_6876_4649# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1029 vccd1 a_15175_4159# a_15162_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1030 a_7733_3133# a_7255_2741# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1031 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X1032 vssd1 _26_.A a_7705_3894# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1033 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1034 a_2307_3677# a_1683_3311# a_2199_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1035 a_12283_3009# _54_.CLK vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1036 vccd1 _63_.RESET_B a_11763_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1037 a_5364_3133# a_4167_2773# a_5172_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1038 a_8471_4943# a_7847_4949# a_8363_5321# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1039 vssd1 a_6085_4551# _38_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1040 a_2925_3133# _52_.RESET_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1041 vssd1 _52_.RESET_B a_7521_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1042 a_7999_3285# a_7824_3311# a_8178_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1043 a_9863_2460# a_9668_2491# a_10173_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1044 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1045 vssd1 _40_.S a_6876_4649# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1046 clkbuf_0_clk.X a_9034_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1047 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1048 a_15000_4233# a_14085_3861# a_14653_3829# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1049 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1050 _63_.Q a_9103_5247# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1051 _25_.X a_10351_4982# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1052 vccd1 a_4605_3285# _63_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1053 a_4936_3133# _52_.RESET_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1054 a_2618_2767# a_2492_2883# a_2214_2899# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1055 vccd1 hold1.X a_2235_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1056 vccd1 a_16863_7127# dq[6] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1057 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X1058 vssd1 _52_.RESET_B a_14697_4221# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1059 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1060 _30_.A a_15248_4649# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1061 a_12559_2365# _54_.CLK vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1062 vccd1 a_2417_2465# a_2307_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1063 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1064 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1065 a_9034_3855# clk vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1066 a_10103_3476# _47_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1067 vssd1 _34_.S a_13278_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1068 _63_.CLK a_4605_3285# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1069 vssd1 a_13919_2775# valid vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1070 vccd1 a_1644_7093# dq[0] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1071 vccd1 a_2531_3009# a_2492_2883# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1072 dq[6] a_16863_7127# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1073 vccd1 a_16083_4564# _33_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1074 vccd1 a_9863_2460# a_9794_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1075 vssd1 a_9494_2767# _54_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1076 vssd1 a_4043_5247# a_3977_5321# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1077 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1078 vccd1 _52_.RESET_B a_2832_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1079 vssd1 _63_.CLK a_2787_4949# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1080 a_14435_4233# a_13919_3861# a_14340_4221# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1081 a_2873_2223# a_1683_2223# a_2764_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1082 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1083 a_7900_7093# output6.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1084 a_7931_2741# a_7775_3009# a_8076_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1085 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1086 a_8581_4917# a_8363_5321# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1087 vssd1 _35_.A a_12504_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1088 vccd1 a_9034_3855# clkbuf_0_clk.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1089 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X1090 vccd1 a_9494_2767# _54_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1091 vccd1 clkbuf_0_clk.X a_9494_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1092 a_4036_7093# output4.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1093 a_9282_5309# _63_.RESET_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1094 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X1095 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1096 vccd1 a_7477_3553# a_7367_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1097 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1098 vccd1 _29_.A a_15578_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1099 _54_.CLK a_9494_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1100 a_4333_2773# a_4167_2773# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1101 vssd1 a_11763_3829# output3.A vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1102 a_12241_4221# a_11763_3829# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1103 vssd1 a_7775_3009# a_7736_2883# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1104 vssd1 a_18059_7127# dq[7] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1105 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1106 a_8494_2767# a_7736_2883# a_7931_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1107 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1108 vssd1 _32_.A a_12856_5737# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1109 a_8355_4726# _40_.A1 a_7896_4551# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1110 a_11763_2741# a_11966_2899# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1111 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1112 a_6842_5309# _63_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1113 a_7063_5309# output5.A a_6700_5175# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1114 vssd1 a_7896_4551# _37_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1115 a_14339_2197# a_14542_2475# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1116 a_4425_2223# a_4259_2223# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1117 vccd1 a_3613_3829# a_3503_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1118 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1119 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1120 _63_.CLK a_4605_3285# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1121 a_5196_3133# a_4616_3145# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1122 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1123 vccd1 _31_.A0 a_16863_7127# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1124 a_3411_4943# _52_.RESET_B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1125 a_12189_5241# _34_.S vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1126 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1127 vssd1 _35_.A a_11568_5737# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1128 a_6876_4649# _43_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1129 clkbuf_0_clk.X a_9034_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1130 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1131 _63_.CLK a_4605_3285# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1132 a_15578_2589# a_14859_2365# a_15015_2460# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1133 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X1134 vccd1 comp a_10055_7119# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1135 vccd1 _25_.S a_10565_4982# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1136 _47_.X a_9176_4649# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
D2 vssd1 clk sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
X1137 a_1644_7093# output3.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1138 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1139 a_2448_2767# a_2011_2741# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1140 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1141 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1142 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1143 a_4605_3285# clkbuf_0_clk.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1144 a_10565_4982# output3.A a_10351_4982# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1145 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X1146 vssd1 a_4605_3285# _63_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1147 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1148 vssd1 _63_.Q a_9176_4649# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1149 vssd1 _32_.A a_13002_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1150 vssd1 a_12263_7127# dq[4] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1151 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1152 a_10556_4649# _25_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1153 a_10103_3476# _47_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1154 a_8581_4917# a_8363_5321# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1155 a_5449_2223# a_4259_2223# a_5340_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1156 vccd1 a_9494_2767# _54_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1157 a_13203_4982# _40_.A1 a_13131_4982# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1158 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1159 clkbuf_0_clk.X a_9034_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1160 a_14435_4233# a_14085_3861# a_14340_4221# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1161 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X1162 a_8072_6147# _41_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1163 a_2461_3311# a_2417_3553# a_2295_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1164 a_14859_2365# _54_.CLK vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1165 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1166 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1167 vccd1 _63_.CLK a_1683_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1168 vssd1 _29_.A a_15578_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1169 _40_.A1 a_10055_7119# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1170 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1171 a_4314_4221# _52_.RESET_B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1172 a_2104_3311# _33_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1173 a_8928_5321# a_7847_4949# a_8581_4917# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1174 a_4883_2589# _52_.RESET_B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1175 vssd1 a_12439_3829# a_12370_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1176 a_14543_3855# a_13919_3861# a_14435_4233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1177 a_15325_2223# a_14946_2589# a_15253_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1178 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1179 a_2764_3311# a_1683_3311# a_2417_3553# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1180 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1181 _37_.A0 a_4135_4159# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1182 vccd1 a_4616_3145# a_4792_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1183 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1184 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1185 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X1186 vssd1 a_12283_4097# a_12244_3971# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1187 last_cycle a_17507_2223# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1188 vccd1 a_12439_2741# a_12370_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1189 vccd1 a_11763_2741# _35_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1190 a_7931_2741# a_7736_2883# a_8241_3133# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1191 vssd1 _34_.A0 a_14471_7127# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
C0 clkbuf_0_clk.X vccd1 2.86fF
C1 _26_.A vccd1 2.64fF
C2 _29_.A vccd1 3.13fF
C3 _52_.RESET_B vccd1 4.20fF
C4 vccd1 output3.A 6.20fF
C5 _54_.CLK vccd1 3.22fF
C6 vccd1 _25_.S 5.14fF
C7 vccd1 fanout13.A 3.09fF
C8 _63_.CLK vccd1 7.82fF
C9 vccd1 _40_.A1 2.44fF
C10 _41_.X vccd1 2.33fF
C11 vccd1 _28_.A0 3.94fF
C12 vccd1 _33_.X 7.83fF
C13 vccd1 _63_.Q 3.73fF
C14 output6.A vccd1 3.43fF
C15 vccd1 _31_.A0 3.40fF
C16 clk vccd1 2.17fF
C17 _52_.D vccd1 6.36fF
C18 vccd1 _32_.A 2.06fF
C19 _52_.RESET_B _26_.A 2.05fF
C20 _40_.S vccd1 2.01fF
C21 clkbuf_0_clk.X vssd1 2.22fF $ **FLOATING
C22 _54_.CLK vssd1 4.22fF $ **FLOATING
C23 _30_.X vssd1 3.46fF $ **FLOATING
C24 _26_.A vssd1 9.30fF $ **FLOATING
C25 fanout13.A vssd1 2.14fF $ **FLOATING
C26 _34_.S vssd1 2.89fF $ **FLOATING
C27 _63_.RESET_B vssd1 4.91fF $ **FLOATING
C28 _52_.RESET_B vssd1 6.77fF $ **FLOATING
C29 _63_.CLK vssd1 2.50fF $ **FLOATING
C30 _40_.A1 vssd1 3.49fF $ **FLOATING
C31 _31_.A0 vssd1 4.04fF $ **FLOATING
C32 _34_.A0 vssd1 3.65fF $ **FLOATING
C33 _37_.A0 vssd1 2.77fF $ **FLOATING
C34 output3.A vssd1 2.16fF $ **FLOATING
C35 vccd1 vssd1 443.17fF
.ends
