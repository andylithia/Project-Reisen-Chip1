** sch_path: /home/andylithia/openmpw/Project-Reisen-Chip1/xschem/shn_test.sch
**.subckt shn_test
C1 vout GND 1p m=1
V1 vin GND 0.9 AC 1
.save i(v1)
XM1 vin net1 vout GND sky130_fd_pr__nfet_01v8 L=0.15 W=40 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
V2 net1 GND 1.8
.save i(v2)
**** begin user architecture code
.lib /home/andylithia/openmpw/pdk_1/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.include /home/andylithia/openmpw/pdk_1/sky130A/libs.ref/sky130_fd_sc_hs/spice/sky130_fd_sc_hs.spice



.noise v(vout) V1 dec 100 1 1e9
* .tran 0.1ns 100ns
.save onoise_spectrum inoise_spectrum
.control
run
setplot noise1
plot inoise_spectrum
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
