magic
tech sky130A
timestamp 1671334348
<< pwell >>
rect -142 -283 142 283
<< psubdiff >>
rect -124 248 -76 265
rect 76 248 124 265
rect -124 217 -107 248
rect 107 217 124 248
rect -124 -248 -107 -217
rect 107 -248 124 -217
rect -124 -265 -76 -248
rect 76 -265 124 -248
<< psubdiffcont >>
rect -76 248 76 265
rect -124 -217 -107 217
rect 107 -217 124 217
rect -76 -265 76 -248
<< xpolycontact >>
rect -59 -200 -24 16
rect 24 -200 59 16
<< ppolyres >>
rect -59 165 59 200
rect -59 16 -24 165
rect 24 16 59 165
<< locali >>
rect -124 248 -76 265
rect 76 248 124 265
rect -124 217 -107 248
rect 107 217 124 248
rect -124 -248 -107 -217
rect 107 -248 124 -217
rect -124 -265 -76 -248
rect 76 -265 124 -248
<< properties >>
string FIXED_BBOX -115 -256 115 256
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.35 l 4 m 1 nx 2 wmin 0.350 lmin 0.50 rho 319.8 val 8.742k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 1 full_metal 1 wmax 0.350 vias 1 n_guard 0 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
