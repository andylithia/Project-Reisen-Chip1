magic
tech sky130A
magscale 1 2
timestamp 1671210538
<< pwell >>
rect -201 -104954 201 104954
<< psubdiff >>
rect -165 104884 -69 104918
rect 69 104884 165 104918
rect -165 104822 -131 104884
rect 131 104822 165 104884
rect -165 -104884 -131 -104822
rect 131 -104884 165 -104822
rect -165 -104918 -69 -104884
rect 69 -104918 165 -104884
<< psubdiffcont >>
rect -69 104884 69 104918
rect -165 -104822 -131 104822
rect 131 -104822 165 104822
rect -69 -104918 69 -104884
<< xpolycontact >>
rect -35 104356 35 104788
rect -35 83924 35 84356
rect -35 83388 35 83820
rect -35 62956 35 63388
rect -35 62420 35 62852
rect -35 41988 35 42420
rect -35 41452 35 41884
rect -35 21020 35 21452
rect -35 20484 35 20916
rect -35 52 35 484
rect -35 -484 35 -52
rect -35 -20916 35 -20484
rect -35 -21452 35 -21020
rect -35 -41884 35 -41452
rect -35 -42420 35 -41988
rect -35 -62852 35 -62420
rect -35 -63388 35 -62956
rect -35 -83820 35 -83388
rect -35 -84356 35 -83924
rect -35 -104788 35 -104356
<< xpolyres >>
rect -35 84356 35 104356
rect -35 63388 35 83388
rect -35 42420 35 62420
rect -35 21452 35 41452
rect -35 484 35 20484
rect -35 -20484 35 -484
rect -35 -41452 35 -21452
rect -35 -62420 35 -42420
rect -35 -83388 35 -63388
rect -35 -104356 35 -84356
<< locali >>
rect -165 104884 -69 104918
rect 69 104884 165 104918
rect -165 104822 -131 104884
rect 131 104822 165 104884
rect -165 -104884 -131 -104822
rect 131 -104884 165 -104822
rect -165 -104918 -69 -104884
rect 69 -104918 165 -104884
<< viali >>
rect -19 104373 19 104770
rect -19 83942 19 84339
rect -19 83405 19 83802
rect -19 62974 19 63371
rect -19 62437 19 62834
rect -19 42006 19 42403
rect -19 41469 19 41866
rect -19 21038 19 21435
rect -19 20501 19 20898
rect -19 70 19 467
rect -19 -467 19 -70
rect -19 -20898 19 -20501
rect -19 -21435 19 -21038
rect -19 -41866 19 -41469
rect -19 -42403 19 -42006
rect -19 -62834 19 -62437
rect -19 -63371 19 -62974
rect -19 -83802 19 -83405
rect -19 -84339 19 -83942
rect -19 -104770 19 -104373
<< metal1 >>
rect -25 104770 25 104782
rect -25 104373 -19 104770
rect 19 104373 25 104770
rect -25 104361 25 104373
rect -25 84339 25 84351
rect -25 83942 -19 84339
rect 19 83942 25 84339
rect -25 83930 25 83942
rect -25 83802 25 83814
rect -25 83405 -19 83802
rect 19 83405 25 83802
rect -25 83393 25 83405
rect -25 63371 25 63383
rect -25 62974 -19 63371
rect 19 62974 25 63371
rect -25 62962 25 62974
rect -25 62834 25 62846
rect -25 62437 -19 62834
rect 19 62437 25 62834
rect -25 62425 25 62437
rect -25 42403 25 42415
rect -25 42006 -19 42403
rect 19 42006 25 42403
rect -25 41994 25 42006
rect -25 41866 25 41878
rect -25 41469 -19 41866
rect 19 41469 25 41866
rect -25 41457 25 41469
rect -25 21435 25 21447
rect -25 21038 -19 21435
rect 19 21038 25 21435
rect -25 21026 25 21038
rect -25 20898 25 20910
rect -25 20501 -19 20898
rect 19 20501 25 20898
rect -25 20489 25 20501
rect -25 467 25 479
rect -25 70 -19 467
rect 19 70 25 467
rect -25 58 25 70
rect -25 -70 25 -58
rect -25 -467 -19 -70
rect 19 -467 25 -70
rect -25 -479 25 -467
rect -25 -20501 25 -20489
rect -25 -20898 -19 -20501
rect 19 -20898 25 -20501
rect -25 -20910 25 -20898
rect -25 -21038 25 -21026
rect -25 -21435 -19 -21038
rect 19 -21435 25 -21038
rect -25 -21447 25 -21435
rect -25 -41469 25 -41457
rect -25 -41866 -19 -41469
rect 19 -41866 25 -41469
rect -25 -41878 25 -41866
rect -25 -42006 25 -41994
rect -25 -42403 -19 -42006
rect 19 -42403 25 -42006
rect -25 -42415 25 -42403
rect -25 -62437 25 -62425
rect -25 -62834 -19 -62437
rect 19 -62834 25 -62437
rect -25 -62846 25 -62834
rect -25 -62974 25 -62962
rect -25 -63371 -19 -62974
rect 19 -63371 25 -62974
rect -25 -63383 25 -63371
rect -25 -83405 25 -83393
rect -25 -83802 -19 -83405
rect 19 -83802 25 -83405
rect -25 -83814 25 -83802
rect -25 -83942 25 -83930
rect -25 -84339 -19 -83942
rect 19 -84339 25 -83942
rect -25 -84351 25 -84339
rect -25 -104373 25 -104361
rect -25 -104770 -19 -104373
rect 19 -104770 25 -104373
rect -25 -104782 25 -104770
<< res0p35 >>
rect -37 84354 37 104358
rect -37 63386 37 83390
rect -37 42418 37 62422
rect -37 21450 37 41454
rect -37 482 37 20486
rect -37 -20486 37 -482
rect -37 -41454 37 -21450
rect -37 -62422 37 -42418
rect -37 -83390 37 -63386
rect -37 -104358 37 -84354
<< properties >>
string FIXED_BBOX -148 -104901 148 104901
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.35 l 100 m 10 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 572.504k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 1 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
