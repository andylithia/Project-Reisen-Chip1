magic
tech sky130A
magscale 1 2
timestamp 1672341375
<< pwell >>
rect -191 10502 191 10588
rect -191 -10502 -105 10502
rect 105 -10502 191 10502
rect -191 -10588 191 -10502
<< psubdiff >>
rect -165 10528 -51 10562
rect -17 10528 17 10562
rect 51 10528 165 10562
rect -165 10455 -131 10528
rect 131 10455 165 10528
rect -165 10387 -131 10421
rect -165 10319 -131 10353
rect -165 10251 -131 10285
rect -165 10183 -131 10217
rect -165 10115 -131 10149
rect -165 10047 -131 10081
rect -165 9979 -131 10013
rect -165 9911 -131 9945
rect -165 9843 -131 9877
rect -165 9775 -131 9809
rect -165 9707 -131 9741
rect -165 9639 -131 9673
rect -165 9571 -131 9605
rect -165 9503 -131 9537
rect -165 9435 -131 9469
rect -165 9367 -131 9401
rect -165 9299 -131 9333
rect -165 9231 -131 9265
rect -165 9163 -131 9197
rect -165 9095 -131 9129
rect -165 9027 -131 9061
rect -165 8959 -131 8993
rect -165 8891 -131 8925
rect -165 8823 -131 8857
rect -165 8755 -131 8789
rect -165 8687 -131 8721
rect -165 8619 -131 8653
rect -165 8551 -131 8585
rect -165 8483 -131 8517
rect -165 8415 -131 8449
rect -165 8347 -131 8381
rect -165 8279 -131 8313
rect -165 8211 -131 8245
rect -165 8143 -131 8177
rect -165 8075 -131 8109
rect -165 8007 -131 8041
rect -165 7939 -131 7973
rect -165 7871 -131 7905
rect -165 7803 -131 7837
rect -165 7735 -131 7769
rect -165 7667 -131 7701
rect -165 7599 -131 7633
rect -165 7531 -131 7565
rect -165 7463 -131 7497
rect -165 7395 -131 7429
rect -165 7327 -131 7361
rect -165 7259 -131 7293
rect -165 7191 -131 7225
rect -165 7123 -131 7157
rect -165 7055 -131 7089
rect -165 6987 -131 7021
rect -165 6919 -131 6953
rect -165 6851 -131 6885
rect -165 6783 -131 6817
rect -165 6715 -131 6749
rect -165 6647 -131 6681
rect -165 6579 -131 6613
rect -165 6511 -131 6545
rect -165 6443 -131 6477
rect -165 6375 -131 6409
rect -165 6307 -131 6341
rect -165 6239 -131 6273
rect -165 6171 -131 6205
rect -165 6103 -131 6137
rect -165 6035 -131 6069
rect -165 5967 -131 6001
rect -165 5899 -131 5933
rect -165 5831 -131 5865
rect -165 5763 -131 5797
rect -165 5695 -131 5729
rect -165 5627 -131 5661
rect -165 5559 -131 5593
rect -165 5491 -131 5525
rect -165 5423 -131 5457
rect -165 5355 -131 5389
rect -165 5287 -131 5321
rect -165 5219 -131 5253
rect -165 5151 -131 5185
rect -165 5083 -131 5117
rect -165 5015 -131 5049
rect -165 4947 -131 4981
rect -165 4879 -131 4913
rect -165 4811 -131 4845
rect -165 4743 -131 4777
rect -165 4675 -131 4709
rect -165 4607 -131 4641
rect -165 4539 -131 4573
rect -165 4471 -131 4505
rect -165 4403 -131 4437
rect -165 4335 -131 4369
rect -165 4267 -131 4301
rect -165 4199 -131 4233
rect -165 4131 -131 4165
rect -165 4063 -131 4097
rect -165 3995 -131 4029
rect -165 3927 -131 3961
rect -165 3859 -131 3893
rect -165 3791 -131 3825
rect -165 3723 -131 3757
rect -165 3655 -131 3689
rect -165 3587 -131 3621
rect -165 3519 -131 3553
rect -165 3451 -131 3485
rect -165 3383 -131 3417
rect -165 3315 -131 3349
rect -165 3247 -131 3281
rect -165 3179 -131 3213
rect -165 3111 -131 3145
rect -165 3043 -131 3077
rect -165 2975 -131 3009
rect -165 2907 -131 2941
rect -165 2839 -131 2873
rect -165 2771 -131 2805
rect -165 2703 -131 2737
rect -165 2635 -131 2669
rect -165 2567 -131 2601
rect -165 2499 -131 2533
rect -165 2431 -131 2465
rect -165 2363 -131 2397
rect -165 2295 -131 2329
rect -165 2227 -131 2261
rect -165 2159 -131 2193
rect -165 2091 -131 2125
rect -165 2023 -131 2057
rect -165 1955 -131 1989
rect -165 1887 -131 1921
rect -165 1819 -131 1853
rect -165 1751 -131 1785
rect -165 1683 -131 1717
rect -165 1615 -131 1649
rect -165 1547 -131 1581
rect -165 1479 -131 1513
rect -165 1411 -131 1445
rect -165 1343 -131 1377
rect -165 1275 -131 1309
rect -165 1207 -131 1241
rect -165 1139 -131 1173
rect -165 1071 -131 1105
rect -165 1003 -131 1037
rect -165 935 -131 969
rect -165 867 -131 901
rect -165 799 -131 833
rect -165 731 -131 765
rect -165 663 -131 697
rect -165 595 -131 629
rect -165 527 -131 561
rect -165 459 -131 493
rect -165 391 -131 425
rect -165 323 -131 357
rect -165 255 -131 289
rect -165 187 -131 221
rect -165 119 -131 153
rect -165 51 -131 85
rect -165 -17 -131 17
rect -165 -85 -131 -51
rect -165 -153 -131 -119
rect -165 -221 -131 -187
rect -165 -289 -131 -255
rect -165 -357 -131 -323
rect -165 -425 -131 -391
rect -165 -493 -131 -459
rect -165 -561 -131 -527
rect -165 -629 -131 -595
rect -165 -697 -131 -663
rect -165 -765 -131 -731
rect -165 -833 -131 -799
rect -165 -901 -131 -867
rect -165 -969 -131 -935
rect -165 -1037 -131 -1003
rect -165 -1105 -131 -1071
rect -165 -1173 -131 -1139
rect -165 -1241 -131 -1207
rect -165 -1309 -131 -1275
rect -165 -1377 -131 -1343
rect -165 -1445 -131 -1411
rect -165 -1513 -131 -1479
rect -165 -1581 -131 -1547
rect -165 -1649 -131 -1615
rect -165 -1717 -131 -1683
rect -165 -1785 -131 -1751
rect -165 -1853 -131 -1819
rect -165 -1921 -131 -1887
rect -165 -1989 -131 -1955
rect -165 -2057 -131 -2023
rect -165 -2125 -131 -2091
rect -165 -2193 -131 -2159
rect -165 -2261 -131 -2227
rect -165 -2329 -131 -2295
rect -165 -2397 -131 -2363
rect -165 -2465 -131 -2431
rect -165 -2533 -131 -2499
rect -165 -2601 -131 -2567
rect -165 -2669 -131 -2635
rect -165 -2737 -131 -2703
rect -165 -2805 -131 -2771
rect -165 -2873 -131 -2839
rect -165 -2941 -131 -2907
rect -165 -3009 -131 -2975
rect -165 -3077 -131 -3043
rect -165 -3145 -131 -3111
rect -165 -3213 -131 -3179
rect -165 -3281 -131 -3247
rect -165 -3349 -131 -3315
rect -165 -3417 -131 -3383
rect -165 -3485 -131 -3451
rect -165 -3553 -131 -3519
rect -165 -3621 -131 -3587
rect -165 -3689 -131 -3655
rect -165 -3757 -131 -3723
rect -165 -3825 -131 -3791
rect -165 -3893 -131 -3859
rect -165 -3961 -131 -3927
rect -165 -4029 -131 -3995
rect -165 -4097 -131 -4063
rect -165 -4165 -131 -4131
rect -165 -4233 -131 -4199
rect -165 -4301 -131 -4267
rect -165 -4369 -131 -4335
rect -165 -4437 -131 -4403
rect -165 -4505 -131 -4471
rect -165 -4573 -131 -4539
rect -165 -4641 -131 -4607
rect -165 -4709 -131 -4675
rect -165 -4777 -131 -4743
rect -165 -4845 -131 -4811
rect -165 -4913 -131 -4879
rect -165 -4981 -131 -4947
rect -165 -5049 -131 -5015
rect -165 -5117 -131 -5083
rect -165 -5185 -131 -5151
rect -165 -5253 -131 -5219
rect -165 -5321 -131 -5287
rect -165 -5389 -131 -5355
rect -165 -5457 -131 -5423
rect -165 -5525 -131 -5491
rect -165 -5593 -131 -5559
rect -165 -5661 -131 -5627
rect -165 -5729 -131 -5695
rect -165 -5797 -131 -5763
rect -165 -5865 -131 -5831
rect -165 -5933 -131 -5899
rect -165 -6001 -131 -5967
rect -165 -6069 -131 -6035
rect -165 -6137 -131 -6103
rect -165 -6205 -131 -6171
rect -165 -6273 -131 -6239
rect -165 -6341 -131 -6307
rect -165 -6409 -131 -6375
rect -165 -6477 -131 -6443
rect -165 -6545 -131 -6511
rect -165 -6613 -131 -6579
rect -165 -6681 -131 -6647
rect -165 -6749 -131 -6715
rect -165 -6817 -131 -6783
rect -165 -6885 -131 -6851
rect -165 -6953 -131 -6919
rect -165 -7021 -131 -6987
rect -165 -7089 -131 -7055
rect -165 -7157 -131 -7123
rect -165 -7225 -131 -7191
rect -165 -7293 -131 -7259
rect -165 -7361 -131 -7327
rect -165 -7429 -131 -7395
rect -165 -7497 -131 -7463
rect -165 -7565 -131 -7531
rect -165 -7633 -131 -7599
rect -165 -7701 -131 -7667
rect -165 -7769 -131 -7735
rect -165 -7837 -131 -7803
rect -165 -7905 -131 -7871
rect -165 -7973 -131 -7939
rect -165 -8041 -131 -8007
rect -165 -8109 -131 -8075
rect -165 -8177 -131 -8143
rect -165 -8245 -131 -8211
rect -165 -8313 -131 -8279
rect -165 -8381 -131 -8347
rect -165 -8449 -131 -8415
rect -165 -8517 -131 -8483
rect -165 -8585 -131 -8551
rect -165 -8653 -131 -8619
rect -165 -8721 -131 -8687
rect -165 -8789 -131 -8755
rect -165 -8857 -131 -8823
rect -165 -8925 -131 -8891
rect -165 -8993 -131 -8959
rect -165 -9061 -131 -9027
rect -165 -9129 -131 -9095
rect -165 -9197 -131 -9163
rect -165 -9265 -131 -9231
rect -165 -9333 -131 -9299
rect -165 -9401 -131 -9367
rect -165 -9469 -131 -9435
rect -165 -9537 -131 -9503
rect -165 -9605 -131 -9571
rect -165 -9673 -131 -9639
rect -165 -9741 -131 -9707
rect -165 -9809 -131 -9775
rect -165 -9877 -131 -9843
rect -165 -9945 -131 -9911
rect -165 -10013 -131 -9979
rect -165 -10081 -131 -10047
rect -165 -10149 -131 -10115
rect -165 -10217 -131 -10183
rect -165 -10285 -131 -10251
rect -165 -10353 -131 -10319
rect -165 -10421 -131 -10387
rect 131 10387 165 10421
rect 131 10319 165 10353
rect 131 10251 165 10285
rect 131 10183 165 10217
rect 131 10115 165 10149
rect 131 10047 165 10081
rect 131 9979 165 10013
rect 131 9911 165 9945
rect 131 9843 165 9877
rect 131 9775 165 9809
rect 131 9707 165 9741
rect 131 9639 165 9673
rect 131 9571 165 9605
rect 131 9503 165 9537
rect 131 9435 165 9469
rect 131 9367 165 9401
rect 131 9299 165 9333
rect 131 9231 165 9265
rect 131 9163 165 9197
rect 131 9095 165 9129
rect 131 9027 165 9061
rect 131 8959 165 8993
rect 131 8891 165 8925
rect 131 8823 165 8857
rect 131 8755 165 8789
rect 131 8687 165 8721
rect 131 8619 165 8653
rect 131 8551 165 8585
rect 131 8483 165 8517
rect 131 8415 165 8449
rect 131 8347 165 8381
rect 131 8279 165 8313
rect 131 8211 165 8245
rect 131 8143 165 8177
rect 131 8075 165 8109
rect 131 8007 165 8041
rect 131 7939 165 7973
rect 131 7871 165 7905
rect 131 7803 165 7837
rect 131 7735 165 7769
rect 131 7667 165 7701
rect 131 7599 165 7633
rect 131 7531 165 7565
rect 131 7463 165 7497
rect 131 7395 165 7429
rect 131 7327 165 7361
rect 131 7259 165 7293
rect 131 7191 165 7225
rect 131 7123 165 7157
rect 131 7055 165 7089
rect 131 6987 165 7021
rect 131 6919 165 6953
rect 131 6851 165 6885
rect 131 6783 165 6817
rect 131 6715 165 6749
rect 131 6647 165 6681
rect 131 6579 165 6613
rect 131 6511 165 6545
rect 131 6443 165 6477
rect 131 6375 165 6409
rect 131 6307 165 6341
rect 131 6239 165 6273
rect 131 6171 165 6205
rect 131 6103 165 6137
rect 131 6035 165 6069
rect 131 5967 165 6001
rect 131 5899 165 5933
rect 131 5831 165 5865
rect 131 5763 165 5797
rect 131 5695 165 5729
rect 131 5627 165 5661
rect 131 5559 165 5593
rect 131 5491 165 5525
rect 131 5423 165 5457
rect 131 5355 165 5389
rect 131 5287 165 5321
rect 131 5219 165 5253
rect 131 5151 165 5185
rect 131 5083 165 5117
rect 131 5015 165 5049
rect 131 4947 165 4981
rect 131 4879 165 4913
rect 131 4811 165 4845
rect 131 4743 165 4777
rect 131 4675 165 4709
rect 131 4607 165 4641
rect 131 4539 165 4573
rect 131 4471 165 4505
rect 131 4403 165 4437
rect 131 4335 165 4369
rect 131 4267 165 4301
rect 131 4199 165 4233
rect 131 4131 165 4165
rect 131 4063 165 4097
rect 131 3995 165 4029
rect 131 3927 165 3961
rect 131 3859 165 3893
rect 131 3791 165 3825
rect 131 3723 165 3757
rect 131 3655 165 3689
rect 131 3587 165 3621
rect 131 3519 165 3553
rect 131 3451 165 3485
rect 131 3383 165 3417
rect 131 3315 165 3349
rect 131 3247 165 3281
rect 131 3179 165 3213
rect 131 3111 165 3145
rect 131 3043 165 3077
rect 131 2975 165 3009
rect 131 2907 165 2941
rect 131 2839 165 2873
rect 131 2771 165 2805
rect 131 2703 165 2737
rect 131 2635 165 2669
rect 131 2567 165 2601
rect 131 2499 165 2533
rect 131 2431 165 2465
rect 131 2363 165 2397
rect 131 2295 165 2329
rect 131 2227 165 2261
rect 131 2159 165 2193
rect 131 2091 165 2125
rect 131 2023 165 2057
rect 131 1955 165 1989
rect 131 1887 165 1921
rect 131 1819 165 1853
rect 131 1751 165 1785
rect 131 1683 165 1717
rect 131 1615 165 1649
rect 131 1547 165 1581
rect 131 1479 165 1513
rect 131 1411 165 1445
rect 131 1343 165 1377
rect 131 1275 165 1309
rect 131 1207 165 1241
rect 131 1139 165 1173
rect 131 1071 165 1105
rect 131 1003 165 1037
rect 131 935 165 969
rect 131 867 165 901
rect 131 799 165 833
rect 131 731 165 765
rect 131 663 165 697
rect 131 595 165 629
rect 131 527 165 561
rect 131 459 165 493
rect 131 391 165 425
rect 131 323 165 357
rect 131 255 165 289
rect 131 187 165 221
rect 131 119 165 153
rect 131 51 165 85
rect 131 -17 165 17
rect 131 -85 165 -51
rect 131 -153 165 -119
rect 131 -221 165 -187
rect 131 -289 165 -255
rect 131 -357 165 -323
rect 131 -425 165 -391
rect 131 -493 165 -459
rect 131 -561 165 -527
rect 131 -629 165 -595
rect 131 -697 165 -663
rect 131 -765 165 -731
rect 131 -833 165 -799
rect 131 -901 165 -867
rect 131 -969 165 -935
rect 131 -1037 165 -1003
rect 131 -1105 165 -1071
rect 131 -1173 165 -1139
rect 131 -1241 165 -1207
rect 131 -1309 165 -1275
rect 131 -1377 165 -1343
rect 131 -1445 165 -1411
rect 131 -1513 165 -1479
rect 131 -1581 165 -1547
rect 131 -1649 165 -1615
rect 131 -1717 165 -1683
rect 131 -1785 165 -1751
rect 131 -1853 165 -1819
rect 131 -1921 165 -1887
rect 131 -1989 165 -1955
rect 131 -2057 165 -2023
rect 131 -2125 165 -2091
rect 131 -2193 165 -2159
rect 131 -2261 165 -2227
rect 131 -2329 165 -2295
rect 131 -2397 165 -2363
rect 131 -2465 165 -2431
rect 131 -2533 165 -2499
rect 131 -2601 165 -2567
rect 131 -2669 165 -2635
rect 131 -2737 165 -2703
rect 131 -2805 165 -2771
rect 131 -2873 165 -2839
rect 131 -2941 165 -2907
rect 131 -3009 165 -2975
rect 131 -3077 165 -3043
rect 131 -3145 165 -3111
rect 131 -3213 165 -3179
rect 131 -3281 165 -3247
rect 131 -3349 165 -3315
rect 131 -3417 165 -3383
rect 131 -3485 165 -3451
rect 131 -3553 165 -3519
rect 131 -3621 165 -3587
rect 131 -3689 165 -3655
rect 131 -3757 165 -3723
rect 131 -3825 165 -3791
rect 131 -3893 165 -3859
rect 131 -3961 165 -3927
rect 131 -4029 165 -3995
rect 131 -4097 165 -4063
rect 131 -4165 165 -4131
rect 131 -4233 165 -4199
rect 131 -4301 165 -4267
rect 131 -4369 165 -4335
rect 131 -4437 165 -4403
rect 131 -4505 165 -4471
rect 131 -4573 165 -4539
rect 131 -4641 165 -4607
rect 131 -4709 165 -4675
rect 131 -4777 165 -4743
rect 131 -4845 165 -4811
rect 131 -4913 165 -4879
rect 131 -4981 165 -4947
rect 131 -5049 165 -5015
rect 131 -5117 165 -5083
rect 131 -5185 165 -5151
rect 131 -5253 165 -5219
rect 131 -5321 165 -5287
rect 131 -5389 165 -5355
rect 131 -5457 165 -5423
rect 131 -5525 165 -5491
rect 131 -5593 165 -5559
rect 131 -5661 165 -5627
rect 131 -5729 165 -5695
rect 131 -5797 165 -5763
rect 131 -5865 165 -5831
rect 131 -5933 165 -5899
rect 131 -6001 165 -5967
rect 131 -6069 165 -6035
rect 131 -6137 165 -6103
rect 131 -6205 165 -6171
rect 131 -6273 165 -6239
rect 131 -6341 165 -6307
rect 131 -6409 165 -6375
rect 131 -6477 165 -6443
rect 131 -6545 165 -6511
rect 131 -6613 165 -6579
rect 131 -6681 165 -6647
rect 131 -6749 165 -6715
rect 131 -6817 165 -6783
rect 131 -6885 165 -6851
rect 131 -6953 165 -6919
rect 131 -7021 165 -6987
rect 131 -7089 165 -7055
rect 131 -7157 165 -7123
rect 131 -7225 165 -7191
rect 131 -7293 165 -7259
rect 131 -7361 165 -7327
rect 131 -7429 165 -7395
rect 131 -7497 165 -7463
rect 131 -7565 165 -7531
rect 131 -7633 165 -7599
rect 131 -7701 165 -7667
rect 131 -7769 165 -7735
rect 131 -7837 165 -7803
rect 131 -7905 165 -7871
rect 131 -7973 165 -7939
rect 131 -8041 165 -8007
rect 131 -8109 165 -8075
rect 131 -8177 165 -8143
rect 131 -8245 165 -8211
rect 131 -8313 165 -8279
rect 131 -8381 165 -8347
rect 131 -8449 165 -8415
rect 131 -8517 165 -8483
rect 131 -8585 165 -8551
rect 131 -8653 165 -8619
rect 131 -8721 165 -8687
rect 131 -8789 165 -8755
rect 131 -8857 165 -8823
rect 131 -8925 165 -8891
rect 131 -8993 165 -8959
rect 131 -9061 165 -9027
rect 131 -9129 165 -9095
rect 131 -9197 165 -9163
rect 131 -9265 165 -9231
rect 131 -9333 165 -9299
rect 131 -9401 165 -9367
rect 131 -9469 165 -9435
rect 131 -9537 165 -9503
rect 131 -9605 165 -9571
rect 131 -9673 165 -9639
rect 131 -9741 165 -9707
rect 131 -9809 165 -9775
rect 131 -9877 165 -9843
rect 131 -9945 165 -9911
rect 131 -10013 165 -9979
rect 131 -10081 165 -10047
rect 131 -10149 165 -10115
rect 131 -10217 165 -10183
rect 131 -10285 165 -10251
rect 131 -10353 165 -10319
rect 131 -10421 165 -10387
rect -165 -10528 -131 -10455
rect 131 -10528 165 -10455
rect -165 -10562 -51 -10528
rect -17 -10562 17 -10528
rect 51 -10562 165 -10528
<< psubdiffcont >>
rect -51 10528 -17 10562
rect 17 10528 51 10562
rect -165 10421 -131 10455
rect -165 10353 -131 10387
rect -165 10285 -131 10319
rect -165 10217 -131 10251
rect -165 10149 -131 10183
rect -165 10081 -131 10115
rect -165 10013 -131 10047
rect -165 9945 -131 9979
rect -165 9877 -131 9911
rect -165 9809 -131 9843
rect -165 9741 -131 9775
rect -165 9673 -131 9707
rect -165 9605 -131 9639
rect -165 9537 -131 9571
rect -165 9469 -131 9503
rect -165 9401 -131 9435
rect -165 9333 -131 9367
rect -165 9265 -131 9299
rect -165 9197 -131 9231
rect -165 9129 -131 9163
rect -165 9061 -131 9095
rect -165 8993 -131 9027
rect -165 8925 -131 8959
rect -165 8857 -131 8891
rect -165 8789 -131 8823
rect -165 8721 -131 8755
rect -165 8653 -131 8687
rect -165 8585 -131 8619
rect -165 8517 -131 8551
rect -165 8449 -131 8483
rect -165 8381 -131 8415
rect -165 8313 -131 8347
rect -165 8245 -131 8279
rect -165 8177 -131 8211
rect -165 8109 -131 8143
rect -165 8041 -131 8075
rect -165 7973 -131 8007
rect -165 7905 -131 7939
rect -165 7837 -131 7871
rect -165 7769 -131 7803
rect -165 7701 -131 7735
rect -165 7633 -131 7667
rect -165 7565 -131 7599
rect -165 7497 -131 7531
rect -165 7429 -131 7463
rect -165 7361 -131 7395
rect -165 7293 -131 7327
rect -165 7225 -131 7259
rect -165 7157 -131 7191
rect -165 7089 -131 7123
rect -165 7021 -131 7055
rect -165 6953 -131 6987
rect -165 6885 -131 6919
rect -165 6817 -131 6851
rect -165 6749 -131 6783
rect -165 6681 -131 6715
rect -165 6613 -131 6647
rect -165 6545 -131 6579
rect -165 6477 -131 6511
rect -165 6409 -131 6443
rect -165 6341 -131 6375
rect -165 6273 -131 6307
rect -165 6205 -131 6239
rect -165 6137 -131 6171
rect -165 6069 -131 6103
rect -165 6001 -131 6035
rect -165 5933 -131 5967
rect -165 5865 -131 5899
rect -165 5797 -131 5831
rect -165 5729 -131 5763
rect -165 5661 -131 5695
rect -165 5593 -131 5627
rect -165 5525 -131 5559
rect -165 5457 -131 5491
rect -165 5389 -131 5423
rect -165 5321 -131 5355
rect -165 5253 -131 5287
rect -165 5185 -131 5219
rect -165 5117 -131 5151
rect -165 5049 -131 5083
rect -165 4981 -131 5015
rect -165 4913 -131 4947
rect -165 4845 -131 4879
rect -165 4777 -131 4811
rect -165 4709 -131 4743
rect -165 4641 -131 4675
rect -165 4573 -131 4607
rect -165 4505 -131 4539
rect -165 4437 -131 4471
rect -165 4369 -131 4403
rect -165 4301 -131 4335
rect -165 4233 -131 4267
rect -165 4165 -131 4199
rect -165 4097 -131 4131
rect -165 4029 -131 4063
rect -165 3961 -131 3995
rect -165 3893 -131 3927
rect -165 3825 -131 3859
rect -165 3757 -131 3791
rect -165 3689 -131 3723
rect -165 3621 -131 3655
rect -165 3553 -131 3587
rect -165 3485 -131 3519
rect -165 3417 -131 3451
rect -165 3349 -131 3383
rect -165 3281 -131 3315
rect -165 3213 -131 3247
rect -165 3145 -131 3179
rect -165 3077 -131 3111
rect -165 3009 -131 3043
rect -165 2941 -131 2975
rect -165 2873 -131 2907
rect -165 2805 -131 2839
rect -165 2737 -131 2771
rect -165 2669 -131 2703
rect -165 2601 -131 2635
rect -165 2533 -131 2567
rect -165 2465 -131 2499
rect -165 2397 -131 2431
rect -165 2329 -131 2363
rect -165 2261 -131 2295
rect -165 2193 -131 2227
rect -165 2125 -131 2159
rect -165 2057 -131 2091
rect -165 1989 -131 2023
rect -165 1921 -131 1955
rect -165 1853 -131 1887
rect -165 1785 -131 1819
rect -165 1717 -131 1751
rect -165 1649 -131 1683
rect -165 1581 -131 1615
rect -165 1513 -131 1547
rect -165 1445 -131 1479
rect -165 1377 -131 1411
rect -165 1309 -131 1343
rect -165 1241 -131 1275
rect -165 1173 -131 1207
rect -165 1105 -131 1139
rect -165 1037 -131 1071
rect -165 969 -131 1003
rect -165 901 -131 935
rect -165 833 -131 867
rect -165 765 -131 799
rect -165 697 -131 731
rect -165 629 -131 663
rect -165 561 -131 595
rect -165 493 -131 527
rect -165 425 -131 459
rect -165 357 -131 391
rect -165 289 -131 323
rect -165 221 -131 255
rect -165 153 -131 187
rect -165 85 -131 119
rect -165 17 -131 51
rect -165 -51 -131 -17
rect -165 -119 -131 -85
rect -165 -187 -131 -153
rect -165 -255 -131 -221
rect -165 -323 -131 -289
rect -165 -391 -131 -357
rect -165 -459 -131 -425
rect -165 -527 -131 -493
rect -165 -595 -131 -561
rect -165 -663 -131 -629
rect -165 -731 -131 -697
rect -165 -799 -131 -765
rect -165 -867 -131 -833
rect -165 -935 -131 -901
rect -165 -1003 -131 -969
rect -165 -1071 -131 -1037
rect -165 -1139 -131 -1105
rect -165 -1207 -131 -1173
rect -165 -1275 -131 -1241
rect -165 -1343 -131 -1309
rect -165 -1411 -131 -1377
rect -165 -1479 -131 -1445
rect -165 -1547 -131 -1513
rect -165 -1615 -131 -1581
rect -165 -1683 -131 -1649
rect -165 -1751 -131 -1717
rect -165 -1819 -131 -1785
rect -165 -1887 -131 -1853
rect -165 -1955 -131 -1921
rect -165 -2023 -131 -1989
rect -165 -2091 -131 -2057
rect -165 -2159 -131 -2125
rect -165 -2227 -131 -2193
rect -165 -2295 -131 -2261
rect -165 -2363 -131 -2329
rect -165 -2431 -131 -2397
rect -165 -2499 -131 -2465
rect -165 -2567 -131 -2533
rect -165 -2635 -131 -2601
rect -165 -2703 -131 -2669
rect -165 -2771 -131 -2737
rect -165 -2839 -131 -2805
rect -165 -2907 -131 -2873
rect -165 -2975 -131 -2941
rect -165 -3043 -131 -3009
rect -165 -3111 -131 -3077
rect -165 -3179 -131 -3145
rect -165 -3247 -131 -3213
rect -165 -3315 -131 -3281
rect -165 -3383 -131 -3349
rect -165 -3451 -131 -3417
rect -165 -3519 -131 -3485
rect -165 -3587 -131 -3553
rect -165 -3655 -131 -3621
rect -165 -3723 -131 -3689
rect -165 -3791 -131 -3757
rect -165 -3859 -131 -3825
rect -165 -3927 -131 -3893
rect -165 -3995 -131 -3961
rect -165 -4063 -131 -4029
rect -165 -4131 -131 -4097
rect -165 -4199 -131 -4165
rect -165 -4267 -131 -4233
rect -165 -4335 -131 -4301
rect -165 -4403 -131 -4369
rect -165 -4471 -131 -4437
rect -165 -4539 -131 -4505
rect -165 -4607 -131 -4573
rect -165 -4675 -131 -4641
rect -165 -4743 -131 -4709
rect -165 -4811 -131 -4777
rect -165 -4879 -131 -4845
rect -165 -4947 -131 -4913
rect -165 -5015 -131 -4981
rect -165 -5083 -131 -5049
rect -165 -5151 -131 -5117
rect -165 -5219 -131 -5185
rect -165 -5287 -131 -5253
rect -165 -5355 -131 -5321
rect -165 -5423 -131 -5389
rect -165 -5491 -131 -5457
rect -165 -5559 -131 -5525
rect -165 -5627 -131 -5593
rect -165 -5695 -131 -5661
rect -165 -5763 -131 -5729
rect -165 -5831 -131 -5797
rect -165 -5899 -131 -5865
rect -165 -5967 -131 -5933
rect -165 -6035 -131 -6001
rect -165 -6103 -131 -6069
rect -165 -6171 -131 -6137
rect -165 -6239 -131 -6205
rect -165 -6307 -131 -6273
rect -165 -6375 -131 -6341
rect -165 -6443 -131 -6409
rect -165 -6511 -131 -6477
rect -165 -6579 -131 -6545
rect -165 -6647 -131 -6613
rect -165 -6715 -131 -6681
rect -165 -6783 -131 -6749
rect -165 -6851 -131 -6817
rect -165 -6919 -131 -6885
rect -165 -6987 -131 -6953
rect -165 -7055 -131 -7021
rect -165 -7123 -131 -7089
rect -165 -7191 -131 -7157
rect -165 -7259 -131 -7225
rect -165 -7327 -131 -7293
rect -165 -7395 -131 -7361
rect -165 -7463 -131 -7429
rect -165 -7531 -131 -7497
rect -165 -7599 -131 -7565
rect -165 -7667 -131 -7633
rect -165 -7735 -131 -7701
rect -165 -7803 -131 -7769
rect -165 -7871 -131 -7837
rect -165 -7939 -131 -7905
rect -165 -8007 -131 -7973
rect -165 -8075 -131 -8041
rect -165 -8143 -131 -8109
rect -165 -8211 -131 -8177
rect -165 -8279 -131 -8245
rect -165 -8347 -131 -8313
rect -165 -8415 -131 -8381
rect -165 -8483 -131 -8449
rect -165 -8551 -131 -8517
rect -165 -8619 -131 -8585
rect -165 -8687 -131 -8653
rect -165 -8755 -131 -8721
rect -165 -8823 -131 -8789
rect -165 -8891 -131 -8857
rect -165 -8959 -131 -8925
rect -165 -9027 -131 -8993
rect -165 -9095 -131 -9061
rect -165 -9163 -131 -9129
rect -165 -9231 -131 -9197
rect -165 -9299 -131 -9265
rect -165 -9367 -131 -9333
rect -165 -9435 -131 -9401
rect -165 -9503 -131 -9469
rect -165 -9571 -131 -9537
rect -165 -9639 -131 -9605
rect -165 -9707 -131 -9673
rect -165 -9775 -131 -9741
rect -165 -9843 -131 -9809
rect -165 -9911 -131 -9877
rect -165 -9979 -131 -9945
rect -165 -10047 -131 -10013
rect -165 -10115 -131 -10081
rect -165 -10183 -131 -10149
rect -165 -10251 -131 -10217
rect -165 -10319 -131 -10285
rect -165 -10387 -131 -10353
rect -165 -10455 -131 -10421
rect 131 10421 165 10455
rect 131 10353 165 10387
rect 131 10285 165 10319
rect 131 10217 165 10251
rect 131 10149 165 10183
rect 131 10081 165 10115
rect 131 10013 165 10047
rect 131 9945 165 9979
rect 131 9877 165 9911
rect 131 9809 165 9843
rect 131 9741 165 9775
rect 131 9673 165 9707
rect 131 9605 165 9639
rect 131 9537 165 9571
rect 131 9469 165 9503
rect 131 9401 165 9435
rect 131 9333 165 9367
rect 131 9265 165 9299
rect 131 9197 165 9231
rect 131 9129 165 9163
rect 131 9061 165 9095
rect 131 8993 165 9027
rect 131 8925 165 8959
rect 131 8857 165 8891
rect 131 8789 165 8823
rect 131 8721 165 8755
rect 131 8653 165 8687
rect 131 8585 165 8619
rect 131 8517 165 8551
rect 131 8449 165 8483
rect 131 8381 165 8415
rect 131 8313 165 8347
rect 131 8245 165 8279
rect 131 8177 165 8211
rect 131 8109 165 8143
rect 131 8041 165 8075
rect 131 7973 165 8007
rect 131 7905 165 7939
rect 131 7837 165 7871
rect 131 7769 165 7803
rect 131 7701 165 7735
rect 131 7633 165 7667
rect 131 7565 165 7599
rect 131 7497 165 7531
rect 131 7429 165 7463
rect 131 7361 165 7395
rect 131 7293 165 7327
rect 131 7225 165 7259
rect 131 7157 165 7191
rect 131 7089 165 7123
rect 131 7021 165 7055
rect 131 6953 165 6987
rect 131 6885 165 6919
rect 131 6817 165 6851
rect 131 6749 165 6783
rect 131 6681 165 6715
rect 131 6613 165 6647
rect 131 6545 165 6579
rect 131 6477 165 6511
rect 131 6409 165 6443
rect 131 6341 165 6375
rect 131 6273 165 6307
rect 131 6205 165 6239
rect 131 6137 165 6171
rect 131 6069 165 6103
rect 131 6001 165 6035
rect 131 5933 165 5967
rect 131 5865 165 5899
rect 131 5797 165 5831
rect 131 5729 165 5763
rect 131 5661 165 5695
rect 131 5593 165 5627
rect 131 5525 165 5559
rect 131 5457 165 5491
rect 131 5389 165 5423
rect 131 5321 165 5355
rect 131 5253 165 5287
rect 131 5185 165 5219
rect 131 5117 165 5151
rect 131 5049 165 5083
rect 131 4981 165 5015
rect 131 4913 165 4947
rect 131 4845 165 4879
rect 131 4777 165 4811
rect 131 4709 165 4743
rect 131 4641 165 4675
rect 131 4573 165 4607
rect 131 4505 165 4539
rect 131 4437 165 4471
rect 131 4369 165 4403
rect 131 4301 165 4335
rect 131 4233 165 4267
rect 131 4165 165 4199
rect 131 4097 165 4131
rect 131 4029 165 4063
rect 131 3961 165 3995
rect 131 3893 165 3927
rect 131 3825 165 3859
rect 131 3757 165 3791
rect 131 3689 165 3723
rect 131 3621 165 3655
rect 131 3553 165 3587
rect 131 3485 165 3519
rect 131 3417 165 3451
rect 131 3349 165 3383
rect 131 3281 165 3315
rect 131 3213 165 3247
rect 131 3145 165 3179
rect 131 3077 165 3111
rect 131 3009 165 3043
rect 131 2941 165 2975
rect 131 2873 165 2907
rect 131 2805 165 2839
rect 131 2737 165 2771
rect 131 2669 165 2703
rect 131 2601 165 2635
rect 131 2533 165 2567
rect 131 2465 165 2499
rect 131 2397 165 2431
rect 131 2329 165 2363
rect 131 2261 165 2295
rect 131 2193 165 2227
rect 131 2125 165 2159
rect 131 2057 165 2091
rect 131 1989 165 2023
rect 131 1921 165 1955
rect 131 1853 165 1887
rect 131 1785 165 1819
rect 131 1717 165 1751
rect 131 1649 165 1683
rect 131 1581 165 1615
rect 131 1513 165 1547
rect 131 1445 165 1479
rect 131 1377 165 1411
rect 131 1309 165 1343
rect 131 1241 165 1275
rect 131 1173 165 1207
rect 131 1105 165 1139
rect 131 1037 165 1071
rect 131 969 165 1003
rect 131 901 165 935
rect 131 833 165 867
rect 131 765 165 799
rect 131 697 165 731
rect 131 629 165 663
rect 131 561 165 595
rect 131 493 165 527
rect 131 425 165 459
rect 131 357 165 391
rect 131 289 165 323
rect 131 221 165 255
rect 131 153 165 187
rect 131 85 165 119
rect 131 17 165 51
rect 131 -51 165 -17
rect 131 -119 165 -85
rect 131 -187 165 -153
rect 131 -255 165 -221
rect 131 -323 165 -289
rect 131 -391 165 -357
rect 131 -459 165 -425
rect 131 -527 165 -493
rect 131 -595 165 -561
rect 131 -663 165 -629
rect 131 -731 165 -697
rect 131 -799 165 -765
rect 131 -867 165 -833
rect 131 -935 165 -901
rect 131 -1003 165 -969
rect 131 -1071 165 -1037
rect 131 -1139 165 -1105
rect 131 -1207 165 -1173
rect 131 -1275 165 -1241
rect 131 -1343 165 -1309
rect 131 -1411 165 -1377
rect 131 -1479 165 -1445
rect 131 -1547 165 -1513
rect 131 -1615 165 -1581
rect 131 -1683 165 -1649
rect 131 -1751 165 -1717
rect 131 -1819 165 -1785
rect 131 -1887 165 -1853
rect 131 -1955 165 -1921
rect 131 -2023 165 -1989
rect 131 -2091 165 -2057
rect 131 -2159 165 -2125
rect 131 -2227 165 -2193
rect 131 -2295 165 -2261
rect 131 -2363 165 -2329
rect 131 -2431 165 -2397
rect 131 -2499 165 -2465
rect 131 -2567 165 -2533
rect 131 -2635 165 -2601
rect 131 -2703 165 -2669
rect 131 -2771 165 -2737
rect 131 -2839 165 -2805
rect 131 -2907 165 -2873
rect 131 -2975 165 -2941
rect 131 -3043 165 -3009
rect 131 -3111 165 -3077
rect 131 -3179 165 -3145
rect 131 -3247 165 -3213
rect 131 -3315 165 -3281
rect 131 -3383 165 -3349
rect 131 -3451 165 -3417
rect 131 -3519 165 -3485
rect 131 -3587 165 -3553
rect 131 -3655 165 -3621
rect 131 -3723 165 -3689
rect 131 -3791 165 -3757
rect 131 -3859 165 -3825
rect 131 -3927 165 -3893
rect 131 -3995 165 -3961
rect 131 -4063 165 -4029
rect 131 -4131 165 -4097
rect 131 -4199 165 -4165
rect 131 -4267 165 -4233
rect 131 -4335 165 -4301
rect 131 -4403 165 -4369
rect 131 -4471 165 -4437
rect 131 -4539 165 -4505
rect 131 -4607 165 -4573
rect 131 -4675 165 -4641
rect 131 -4743 165 -4709
rect 131 -4811 165 -4777
rect 131 -4879 165 -4845
rect 131 -4947 165 -4913
rect 131 -5015 165 -4981
rect 131 -5083 165 -5049
rect 131 -5151 165 -5117
rect 131 -5219 165 -5185
rect 131 -5287 165 -5253
rect 131 -5355 165 -5321
rect 131 -5423 165 -5389
rect 131 -5491 165 -5457
rect 131 -5559 165 -5525
rect 131 -5627 165 -5593
rect 131 -5695 165 -5661
rect 131 -5763 165 -5729
rect 131 -5831 165 -5797
rect 131 -5899 165 -5865
rect 131 -5967 165 -5933
rect 131 -6035 165 -6001
rect 131 -6103 165 -6069
rect 131 -6171 165 -6137
rect 131 -6239 165 -6205
rect 131 -6307 165 -6273
rect 131 -6375 165 -6341
rect 131 -6443 165 -6409
rect 131 -6511 165 -6477
rect 131 -6579 165 -6545
rect 131 -6647 165 -6613
rect 131 -6715 165 -6681
rect 131 -6783 165 -6749
rect 131 -6851 165 -6817
rect 131 -6919 165 -6885
rect 131 -6987 165 -6953
rect 131 -7055 165 -7021
rect 131 -7123 165 -7089
rect 131 -7191 165 -7157
rect 131 -7259 165 -7225
rect 131 -7327 165 -7293
rect 131 -7395 165 -7361
rect 131 -7463 165 -7429
rect 131 -7531 165 -7497
rect 131 -7599 165 -7565
rect 131 -7667 165 -7633
rect 131 -7735 165 -7701
rect 131 -7803 165 -7769
rect 131 -7871 165 -7837
rect 131 -7939 165 -7905
rect 131 -8007 165 -7973
rect 131 -8075 165 -8041
rect 131 -8143 165 -8109
rect 131 -8211 165 -8177
rect 131 -8279 165 -8245
rect 131 -8347 165 -8313
rect 131 -8415 165 -8381
rect 131 -8483 165 -8449
rect 131 -8551 165 -8517
rect 131 -8619 165 -8585
rect 131 -8687 165 -8653
rect 131 -8755 165 -8721
rect 131 -8823 165 -8789
rect 131 -8891 165 -8857
rect 131 -8959 165 -8925
rect 131 -9027 165 -8993
rect 131 -9095 165 -9061
rect 131 -9163 165 -9129
rect 131 -9231 165 -9197
rect 131 -9299 165 -9265
rect 131 -9367 165 -9333
rect 131 -9435 165 -9401
rect 131 -9503 165 -9469
rect 131 -9571 165 -9537
rect 131 -9639 165 -9605
rect 131 -9707 165 -9673
rect 131 -9775 165 -9741
rect 131 -9843 165 -9809
rect 131 -9911 165 -9877
rect 131 -9979 165 -9945
rect 131 -10047 165 -10013
rect 131 -10115 165 -10081
rect 131 -10183 165 -10149
rect 131 -10251 165 -10217
rect 131 -10319 165 -10285
rect 131 -10387 165 -10353
rect 131 -10455 165 -10421
rect -51 -10562 -17 -10528
rect 17 -10562 51 -10528
<< xpolycontact >>
rect -35 10000 35 10432
rect -35 -10432 35 -10000
<< xpolyres >>
rect -35 -10000 35 10000
<< locali >>
rect -165 10528 -51 10562
rect -17 10528 17 10562
rect 51 10528 165 10562
rect -165 10455 -131 10528
rect 131 10455 165 10528
rect -165 10387 -131 10421
rect -165 10319 -131 10353
rect -165 10251 -131 10285
rect -165 10183 -131 10217
rect -165 10115 -131 10149
rect -165 10047 -131 10081
rect -165 9979 -131 10013
rect 131 10387 165 10421
rect 131 10319 165 10353
rect 131 10251 165 10285
rect 131 10183 165 10217
rect 131 10115 165 10149
rect 131 10047 165 10081
rect -165 9911 -131 9945
rect -165 9843 -131 9877
rect -165 9775 -131 9809
rect -165 9707 -131 9741
rect -165 9639 -131 9673
rect -165 9571 -131 9605
rect -165 9503 -131 9537
rect -165 9435 -131 9469
rect -165 9367 -131 9401
rect -165 9299 -131 9333
rect -165 9231 -131 9265
rect -165 9163 -131 9197
rect -165 9095 -131 9129
rect -165 9027 -131 9061
rect -165 8959 -131 8993
rect -165 8891 -131 8925
rect -165 8823 -131 8857
rect -165 8755 -131 8789
rect -165 8687 -131 8721
rect -165 8619 -131 8653
rect -165 8551 -131 8585
rect -165 8483 -131 8517
rect -165 8415 -131 8449
rect -165 8347 -131 8381
rect -165 8279 -131 8313
rect -165 8211 -131 8245
rect -165 8143 -131 8177
rect -165 8075 -131 8109
rect -165 8007 -131 8041
rect -165 7939 -131 7973
rect -165 7871 -131 7905
rect -165 7803 -131 7837
rect -165 7735 -131 7769
rect -165 7667 -131 7701
rect -165 7599 -131 7633
rect -165 7531 -131 7565
rect -165 7463 -131 7497
rect -165 7395 -131 7429
rect -165 7327 -131 7361
rect -165 7259 -131 7293
rect -165 7191 -131 7225
rect -165 7123 -131 7157
rect -165 7055 -131 7089
rect -165 6987 -131 7021
rect -165 6919 -131 6953
rect -165 6851 -131 6885
rect -165 6783 -131 6817
rect -165 6715 -131 6749
rect -165 6647 -131 6681
rect -165 6579 -131 6613
rect -165 6511 -131 6545
rect -165 6443 -131 6477
rect -165 6375 -131 6409
rect -165 6307 -131 6341
rect -165 6239 -131 6273
rect -165 6171 -131 6205
rect -165 6103 -131 6137
rect -165 6035 -131 6069
rect -165 5967 -131 6001
rect -165 5899 -131 5933
rect -165 5831 -131 5865
rect -165 5763 -131 5797
rect -165 5695 -131 5729
rect -165 5627 -131 5661
rect -165 5559 -131 5593
rect -165 5491 -131 5525
rect -165 5423 -131 5457
rect -165 5355 -131 5389
rect -165 5287 -131 5321
rect -165 5219 -131 5253
rect -165 5151 -131 5185
rect -165 5083 -131 5117
rect -165 5015 -131 5049
rect -165 4947 -131 4981
rect -165 4879 -131 4913
rect -165 4811 -131 4845
rect -165 4743 -131 4777
rect -165 4675 -131 4709
rect -165 4607 -131 4641
rect -165 4539 -131 4573
rect -165 4471 -131 4505
rect -165 4403 -131 4437
rect -165 4335 -131 4369
rect -165 4267 -131 4301
rect -165 4199 -131 4233
rect -165 4131 -131 4165
rect -165 4063 -131 4097
rect -165 3995 -131 4029
rect -165 3927 -131 3961
rect -165 3859 -131 3893
rect -165 3791 -131 3825
rect -165 3723 -131 3757
rect -165 3655 -131 3689
rect -165 3587 -131 3621
rect -165 3519 -131 3553
rect -165 3451 -131 3485
rect -165 3383 -131 3417
rect -165 3315 -131 3349
rect -165 3247 -131 3281
rect -165 3179 -131 3213
rect -165 3111 -131 3145
rect -165 3043 -131 3077
rect -165 2975 -131 3009
rect -165 2907 -131 2941
rect -165 2839 -131 2873
rect -165 2771 -131 2805
rect -165 2703 -131 2737
rect -165 2635 -131 2669
rect -165 2567 -131 2601
rect -165 2499 -131 2533
rect -165 2431 -131 2465
rect -165 2363 -131 2397
rect -165 2295 -131 2329
rect -165 2227 -131 2261
rect -165 2159 -131 2193
rect -165 2091 -131 2125
rect -165 2023 -131 2057
rect -165 1955 -131 1989
rect -165 1887 -131 1921
rect -165 1819 -131 1853
rect -165 1751 -131 1785
rect -165 1683 -131 1717
rect -165 1615 -131 1649
rect -165 1547 -131 1581
rect -165 1479 -131 1513
rect -165 1411 -131 1445
rect -165 1343 -131 1377
rect -165 1275 -131 1309
rect -165 1207 -131 1241
rect -165 1139 -131 1173
rect -165 1071 -131 1105
rect -165 1003 -131 1037
rect -165 935 -131 969
rect -165 867 -131 901
rect -165 799 -131 833
rect -165 731 -131 765
rect -165 663 -131 697
rect -165 595 -131 629
rect -165 527 -131 561
rect -165 459 -131 493
rect -165 391 -131 425
rect -165 323 -131 357
rect -165 255 -131 289
rect -165 187 -131 221
rect -165 119 -131 153
rect -165 51 -131 85
rect -165 -17 -131 17
rect -165 -85 -131 -51
rect -165 -153 -131 -119
rect -165 -221 -131 -187
rect -165 -289 -131 -255
rect -165 -357 -131 -323
rect -165 -425 -131 -391
rect -165 -493 -131 -459
rect -165 -561 -131 -527
rect -165 -629 -131 -595
rect -165 -697 -131 -663
rect -165 -765 -131 -731
rect -165 -833 -131 -799
rect -165 -901 -131 -867
rect -165 -969 -131 -935
rect -165 -1037 -131 -1003
rect -165 -1105 -131 -1071
rect -165 -1173 -131 -1139
rect -165 -1241 -131 -1207
rect -165 -1309 -131 -1275
rect -165 -1377 -131 -1343
rect -165 -1445 -131 -1411
rect -165 -1513 -131 -1479
rect -165 -1581 -131 -1547
rect -165 -1649 -131 -1615
rect -165 -1717 -131 -1683
rect -165 -1785 -131 -1751
rect -165 -1853 -131 -1819
rect -165 -1921 -131 -1887
rect -165 -1989 -131 -1955
rect -165 -2057 -131 -2023
rect -165 -2125 -131 -2091
rect -165 -2193 -131 -2159
rect -165 -2261 -131 -2227
rect -165 -2329 -131 -2295
rect -165 -2397 -131 -2363
rect -165 -2465 -131 -2431
rect -165 -2533 -131 -2499
rect -165 -2601 -131 -2567
rect -165 -2669 -131 -2635
rect -165 -2737 -131 -2703
rect -165 -2805 -131 -2771
rect -165 -2873 -131 -2839
rect -165 -2941 -131 -2907
rect -165 -3009 -131 -2975
rect -165 -3077 -131 -3043
rect -165 -3145 -131 -3111
rect -165 -3213 -131 -3179
rect -165 -3281 -131 -3247
rect -165 -3349 -131 -3315
rect -165 -3417 -131 -3383
rect -165 -3485 -131 -3451
rect -165 -3553 -131 -3519
rect -165 -3621 -131 -3587
rect -165 -3689 -131 -3655
rect -165 -3757 -131 -3723
rect -165 -3825 -131 -3791
rect -165 -3893 -131 -3859
rect -165 -3961 -131 -3927
rect -165 -4029 -131 -3995
rect -165 -4097 -131 -4063
rect -165 -4165 -131 -4131
rect -165 -4233 -131 -4199
rect -165 -4301 -131 -4267
rect -165 -4369 -131 -4335
rect -165 -4437 -131 -4403
rect -165 -4505 -131 -4471
rect -165 -4573 -131 -4539
rect -165 -4641 -131 -4607
rect -165 -4709 -131 -4675
rect -165 -4777 -131 -4743
rect -165 -4845 -131 -4811
rect -165 -4913 -131 -4879
rect -165 -4981 -131 -4947
rect -165 -5049 -131 -5015
rect -165 -5117 -131 -5083
rect -165 -5185 -131 -5151
rect -165 -5253 -131 -5219
rect -165 -5321 -131 -5287
rect -165 -5389 -131 -5355
rect -165 -5457 -131 -5423
rect -165 -5525 -131 -5491
rect -165 -5593 -131 -5559
rect -165 -5661 -131 -5627
rect -165 -5729 -131 -5695
rect -165 -5797 -131 -5763
rect -165 -5865 -131 -5831
rect -165 -5933 -131 -5899
rect -165 -6001 -131 -5967
rect -165 -6069 -131 -6035
rect -165 -6137 -131 -6103
rect -165 -6205 -131 -6171
rect -165 -6273 -131 -6239
rect -165 -6341 -131 -6307
rect -165 -6409 -131 -6375
rect -165 -6477 -131 -6443
rect -165 -6545 -131 -6511
rect -165 -6613 -131 -6579
rect -165 -6681 -131 -6647
rect -165 -6749 -131 -6715
rect -165 -6817 -131 -6783
rect -165 -6885 -131 -6851
rect -165 -6953 -131 -6919
rect -165 -7021 -131 -6987
rect -165 -7089 -131 -7055
rect -165 -7157 -131 -7123
rect -165 -7225 -131 -7191
rect -165 -7293 -131 -7259
rect -165 -7361 -131 -7327
rect -165 -7429 -131 -7395
rect -165 -7497 -131 -7463
rect -165 -7565 -131 -7531
rect -165 -7633 -131 -7599
rect -165 -7701 -131 -7667
rect -165 -7769 -131 -7735
rect -165 -7837 -131 -7803
rect -165 -7905 -131 -7871
rect -165 -7973 -131 -7939
rect -165 -8041 -131 -8007
rect -165 -8109 -131 -8075
rect -165 -8177 -131 -8143
rect -165 -8245 -131 -8211
rect -165 -8313 -131 -8279
rect -165 -8381 -131 -8347
rect -165 -8449 -131 -8415
rect -165 -8517 -131 -8483
rect -165 -8585 -131 -8551
rect -165 -8653 -131 -8619
rect -165 -8721 -131 -8687
rect -165 -8789 -131 -8755
rect -165 -8857 -131 -8823
rect -165 -8925 -131 -8891
rect -165 -8993 -131 -8959
rect -165 -9061 -131 -9027
rect -165 -9129 -131 -9095
rect -165 -9197 -131 -9163
rect -165 -9265 -131 -9231
rect -165 -9333 -131 -9299
rect -165 -9401 -131 -9367
rect -165 -9469 -131 -9435
rect -165 -9537 -131 -9503
rect -165 -9605 -131 -9571
rect -165 -9673 -131 -9639
rect -165 -9741 -131 -9707
rect -165 -9809 -131 -9775
rect -165 -9877 -131 -9843
rect -165 -9945 -131 -9911
rect -165 -10013 -131 -9979
rect 131 9979 165 10013
rect 131 9911 165 9945
rect 131 9843 165 9877
rect 131 9775 165 9809
rect 131 9707 165 9741
rect 131 9639 165 9673
rect 131 9571 165 9605
rect 131 9503 165 9537
rect 131 9435 165 9469
rect 131 9367 165 9401
rect 131 9299 165 9333
rect 131 9231 165 9265
rect 131 9163 165 9197
rect 131 9095 165 9129
rect 131 9027 165 9061
rect 131 8959 165 8993
rect 131 8891 165 8925
rect 131 8823 165 8857
rect 131 8755 165 8789
rect 131 8687 165 8721
rect 131 8619 165 8653
rect 131 8551 165 8585
rect 131 8483 165 8517
rect 131 8415 165 8449
rect 131 8347 165 8381
rect 131 8279 165 8313
rect 131 8211 165 8245
rect 131 8143 165 8177
rect 131 8075 165 8109
rect 131 8007 165 8041
rect 131 7939 165 7973
rect 131 7871 165 7905
rect 131 7803 165 7837
rect 131 7735 165 7769
rect 131 7667 165 7701
rect 131 7599 165 7633
rect 131 7531 165 7565
rect 131 7463 165 7497
rect 131 7395 165 7429
rect 131 7327 165 7361
rect 131 7259 165 7293
rect 131 7191 165 7225
rect 131 7123 165 7157
rect 131 7055 165 7089
rect 131 6987 165 7021
rect 131 6919 165 6953
rect 131 6851 165 6885
rect 131 6783 165 6817
rect 131 6715 165 6749
rect 131 6647 165 6681
rect 131 6579 165 6613
rect 131 6511 165 6545
rect 131 6443 165 6477
rect 131 6375 165 6409
rect 131 6307 165 6341
rect 131 6239 165 6273
rect 131 6171 165 6205
rect 131 6103 165 6137
rect 131 6035 165 6069
rect 131 5967 165 6001
rect 131 5899 165 5933
rect 131 5831 165 5865
rect 131 5763 165 5797
rect 131 5695 165 5729
rect 131 5627 165 5661
rect 131 5559 165 5593
rect 131 5491 165 5525
rect 131 5423 165 5457
rect 131 5355 165 5389
rect 131 5287 165 5321
rect 131 5219 165 5253
rect 131 5151 165 5185
rect 131 5083 165 5117
rect 131 5015 165 5049
rect 131 4947 165 4981
rect 131 4879 165 4913
rect 131 4811 165 4845
rect 131 4743 165 4777
rect 131 4675 165 4709
rect 131 4607 165 4641
rect 131 4539 165 4573
rect 131 4471 165 4505
rect 131 4403 165 4437
rect 131 4335 165 4369
rect 131 4267 165 4301
rect 131 4199 165 4233
rect 131 4131 165 4165
rect 131 4063 165 4097
rect 131 3995 165 4029
rect 131 3927 165 3961
rect 131 3859 165 3893
rect 131 3791 165 3825
rect 131 3723 165 3757
rect 131 3655 165 3689
rect 131 3587 165 3621
rect 131 3519 165 3553
rect 131 3451 165 3485
rect 131 3383 165 3417
rect 131 3315 165 3349
rect 131 3247 165 3281
rect 131 3179 165 3213
rect 131 3111 165 3145
rect 131 3043 165 3077
rect 131 2975 165 3009
rect 131 2907 165 2941
rect 131 2839 165 2873
rect 131 2771 165 2805
rect 131 2703 165 2737
rect 131 2635 165 2669
rect 131 2567 165 2601
rect 131 2499 165 2533
rect 131 2431 165 2465
rect 131 2363 165 2397
rect 131 2295 165 2329
rect 131 2227 165 2261
rect 131 2159 165 2193
rect 131 2091 165 2125
rect 131 2023 165 2057
rect 131 1955 165 1989
rect 131 1887 165 1921
rect 131 1819 165 1853
rect 131 1751 165 1785
rect 131 1683 165 1717
rect 131 1615 165 1649
rect 131 1547 165 1581
rect 131 1479 165 1513
rect 131 1411 165 1445
rect 131 1343 165 1377
rect 131 1275 165 1309
rect 131 1207 165 1241
rect 131 1139 165 1173
rect 131 1071 165 1105
rect 131 1003 165 1037
rect 131 935 165 969
rect 131 867 165 901
rect 131 799 165 833
rect 131 731 165 765
rect 131 663 165 697
rect 131 595 165 629
rect 131 527 165 561
rect 131 459 165 493
rect 131 391 165 425
rect 131 323 165 357
rect 131 255 165 289
rect 131 187 165 221
rect 131 119 165 153
rect 131 51 165 85
rect 131 -17 165 17
rect 131 -85 165 -51
rect 131 -153 165 -119
rect 131 -221 165 -187
rect 131 -289 165 -255
rect 131 -357 165 -323
rect 131 -425 165 -391
rect 131 -493 165 -459
rect 131 -561 165 -527
rect 131 -629 165 -595
rect 131 -697 165 -663
rect 131 -765 165 -731
rect 131 -833 165 -799
rect 131 -901 165 -867
rect 131 -969 165 -935
rect 131 -1037 165 -1003
rect 131 -1105 165 -1071
rect 131 -1173 165 -1139
rect 131 -1241 165 -1207
rect 131 -1309 165 -1275
rect 131 -1377 165 -1343
rect 131 -1445 165 -1411
rect 131 -1513 165 -1479
rect 131 -1581 165 -1547
rect 131 -1649 165 -1615
rect 131 -1717 165 -1683
rect 131 -1785 165 -1751
rect 131 -1853 165 -1819
rect 131 -1921 165 -1887
rect 131 -1989 165 -1955
rect 131 -2057 165 -2023
rect 131 -2125 165 -2091
rect 131 -2193 165 -2159
rect 131 -2261 165 -2227
rect 131 -2329 165 -2295
rect 131 -2397 165 -2363
rect 131 -2465 165 -2431
rect 131 -2533 165 -2499
rect 131 -2601 165 -2567
rect 131 -2669 165 -2635
rect 131 -2737 165 -2703
rect 131 -2805 165 -2771
rect 131 -2873 165 -2839
rect 131 -2941 165 -2907
rect 131 -3009 165 -2975
rect 131 -3077 165 -3043
rect 131 -3145 165 -3111
rect 131 -3213 165 -3179
rect 131 -3281 165 -3247
rect 131 -3349 165 -3315
rect 131 -3417 165 -3383
rect 131 -3485 165 -3451
rect 131 -3553 165 -3519
rect 131 -3621 165 -3587
rect 131 -3689 165 -3655
rect 131 -3757 165 -3723
rect 131 -3825 165 -3791
rect 131 -3893 165 -3859
rect 131 -3961 165 -3927
rect 131 -4029 165 -3995
rect 131 -4097 165 -4063
rect 131 -4165 165 -4131
rect 131 -4233 165 -4199
rect 131 -4301 165 -4267
rect 131 -4369 165 -4335
rect 131 -4437 165 -4403
rect 131 -4505 165 -4471
rect 131 -4573 165 -4539
rect 131 -4641 165 -4607
rect 131 -4709 165 -4675
rect 131 -4777 165 -4743
rect 131 -4845 165 -4811
rect 131 -4913 165 -4879
rect 131 -4981 165 -4947
rect 131 -5049 165 -5015
rect 131 -5117 165 -5083
rect 131 -5185 165 -5151
rect 131 -5253 165 -5219
rect 131 -5321 165 -5287
rect 131 -5389 165 -5355
rect 131 -5457 165 -5423
rect 131 -5525 165 -5491
rect 131 -5593 165 -5559
rect 131 -5661 165 -5627
rect 131 -5729 165 -5695
rect 131 -5797 165 -5763
rect 131 -5865 165 -5831
rect 131 -5933 165 -5899
rect 131 -6001 165 -5967
rect 131 -6069 165 -6035
rect 131 -6137 165 -6103
rect 131 -6205 165 -6171
rect 131 -6273 165 -6239
rect 131 -6341 165 -6307
rect 131 -6409 165 -6375
rect 131 -6477 165 -6443
rect 131 -6545 165 -6511
rect 131 -6613 165 -6579
rect 131 -6681 165 -6647
rect 131 -6749 165 -6715
rect 131 -6817 165 -6783
rect 131 -6885 165 -6851
rect 131 -6953 165 -6919
rect 131 -7021 165 -6987
rect 131 -7089 165 -7055
rect 131 -7157 165 -7123
rect 131 -7225 165 -7191
rect 131 -7293 165 -7259
rect 131 -7361 165 -7327
rect 131 -7429 165 -7395
rect 131 -7497 165 -7463
rect 131 -7565 165 -7531
rect 131 -7633 165 -7599
rect 131 -7701 165 -7667
rect 131 -7769 165 -7735
rect 131 -7837 165 -7803
rect 131 -7905 165 -7871
rect 131 -7973 165 -7939
rect 131 -8041 165 -8007
rect 131 -8109 165 -8075
rect 131 -8177 165 -8143
rect 131 -8245 165 -8211
rect 131 -8313 165 -8279
rect 131 -8381 165 -8347
rect 131 -8449 165 -8415
rect 131 -8517 165 -8483
rect 131 -8585 165 -8551
rect 131 -8653 165 -8619
rect 131 -8721 165 -8687
rect 131 -8789 165 -8755
rect 131 -8857 165 -8823
rect 131 -8925 165 -8891
rect 131 -8993 165 -8959
rect 131 -9061 165 -9027
rect 131 -9129 165 -9095
rect 131 -9197 165 -9163
rect 131 -9265 165 -9231
rect 131 -9333 165 -9299
rect 131 -9401 165 -9367
rect 131 -9469 165 -9435
rect 131 -9537 165 -9503
rect 131 -9605 165 -9571
rect 131 -9673 165 -9639
rect 131 -9741 165 -9707
rect 131 -9809 165 -9775
rect 131 -9877 165 -9843
rect 131 -9945 165 -9911
rect -165 -10081 -131 -10047
rect -165 -10149 -131 -10115
rect -165 -10217 -131 -10183
rect -165 -10285 -131 -10251
rect -165 -10353 -131 -10319
rect -165 -10421 -131 -10387
rect 131 -10013 165 -9979
rect 131 -10081 165 -10047
rect 131 -10149 165 -10115
rect 131 -10217 165 -10183
rect 131 -10285 165 -10251
rect 131 -10353 165 -10319
rect 131 -10421 165 -10387
rect -165 -10528 -131 -10455
rect 131 -10528 165 -10455
rect -165 -10562 -51 -10528
rect -17 -10562 17 -10528
rect 51 -10562 165 -10528
<< viali >>
rect -17 10378 17 10412
rect -17 10306 17 10340
rect -17 10234 17 10268
rect -17 10162 17 10196
rect -17 10090 17 10124
rect -17 10018 17 10052
rect -17 -10053 17 -10019
rect -17 -10125 17 -10091
rect -17 -10197 17 -10163
rect -17 -10269 17 -10235
rect -17 -10341 17 -10307
rect -17 -10413 17 -10379
<< metal1 >>
rect -25 10412 25 10426
rect -25 10378 -17 10412
rect 17 10378 25 10412
rect -25 10340 25 10378
rect -25 10306 -17 10340
rect 17 10306 25 10340
rect -25 10268 25 10306
rect -25 10234 -17 10268
rect 17 10234 25 10268
rect -25 10196 25 10234
rect -25 10162 -17 10196
rect 17 10162 25 10196
rect -25 10124 25 10162
rect -25 10090 -17 10124
rect 17 10090 25 10124
rect -25 10052 25 10090
rect -25 10018 -17 10052
rect 17 10018 25 10052
rect -25 10005 25 10018
rect -25 -10019 25 -10005
rect -25 -10053 -17 -10019
rect 17 -10053 25 -10019
rect -25 -10091 25 -10053
rect -25 -10125 -17 -10091
rect 17 -10125 25 -10091
rect -25 -10163 25 -10125
rect -25 -10197 -17 -10163
rect 17 -10197 25 -10163
rect -25 -10235 25 -10197
rect -25 -10269 -17 -10235
rect 17 -10269 25 -10235
rect -25 -10307 25 -10269
rect -25 -10341 -17 -10307
rect 17 -10341 25 -10307
rect -25 -10379 25 -10341
rect -25 -10413 -17 -10379
rect 17 -10413 25 -10379
rect -25 -10426 25 -10413
<< properties >>
string FIXED_BBOX -148 -10545 148 10545
<< end >>
