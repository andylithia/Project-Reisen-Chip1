magic
tech sky130B
timestamp 1668125106
<< metal4 >>
rect 1860 4420 2140 4520
rect 1860 -160 1920 4420
rect 1950 -160 2050 4390
rect 2080 -160 2140 4420
<< fillblock >>
rect 1860 -160 2140 4520
<< labels >>
rlabel metal4 1950 -160 2050 -100 1 TOP
rlabel metal4 1920 4420 2080 4520 1 BOT
<< end >>
