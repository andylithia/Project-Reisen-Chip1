magic
tech sky130A
magscale 1 2
timestamp 1671207568
<< error_p >>
rect -383 172 -325 178
rect -265 172 -207 178
rect -147 172 -89 178
rect -29 172 29 178
rect 89 172 147 178
rect 207 172 265 178
rect 325 172 383 178
rect -383 138 -371 172
rect -265 138 -253 172
rect -147 138 -135 172
rect -29 138 -17 172
rect 89 138 101 172
rect 207 138 219 172
rect 325 138 337 172
rect -383 132 -325 138
rect -265 132 -207 138
rect -147 132 -89 138
rect -29 132 29 138
rect 89 132 147 138
rect 207 132 265 138
rect 325 132 383 138
rect -383 -138 -325 -132
rect -265 -138 -207 -132
rect -147 -138 -89 -132
rect -29 -138 29 -132
rect 89 -138 147 -132
rect 207 -138 265 -132
rect 325 -138 383 -132
rect -383 -172 -371 -138
rect -265 -172 -253 -138
rect -147 -172 -135 -138
rect -29 -172 -17 -138
rect 89 -172 101 -138
rect 207 -172 219 -138
rect 325 -172 337 -138
rect -383 -178 -325 -172
rect -265 -178 -207 -172
rect -147 -178 -89 -172
rect -29 -178 29 -172
rect 89 -178 147 -172
rect 207 -178 265 -172
rect 325 -178 383 -172
<< pwell >>
rect -580 -310 580 310
<< nmos >>
rect -384 -100 -324 100
rect -266 -100 -206 100
rect -148 -100 -88 100
rect -30 -100 30 100
rect 88 -100 148 100
rect 206 -100 266 100
rect 324 -100 384 100
<< ndiff >>
rect -442 88 -384 100
rect -442 -88 -430 88
rect -396 -88 -384 88
rect -442 -100 -384 -88
rect -324 88 -266 100
rect -324 -88 -312 88
rect -278 -88 -266 88
rect -324 -100 -266 -88
rect -206 88 -148 100
rect -206 -88 -194 88
rect -160 -88 -148 88
rect -206 -100 -148 -88
rect -88 88 -30 100
rect -88 -88 -76 88
rect -42 -88 -30 88
rect -88 -100 -30 -88
rect 30 88 88 100
rect 30 -88 42 88
rect 76 -88 88 88
rect 30 -100 88 -88
rect 148 88 206 100
rect 148 -88 160 88
rect 194 -88 206 88
rect 148 -100 206 -88
rect 266 88 324 100
rect 266 -88 278 88
rect 312 -88 324 88
rect 266 -100 324 -88
rect 384 88 442 100
rect 384 -88 396 88
rect 430 -88 442 88
rect 384 -100 442 -88
<< ndiffc >>
rect -430 -88 -396 88
rect -312 -88 -278 88
rect -194 -88 -160 88
rect -76 -88 -42 88
rect 42 -88 76 88
rect 160 -88 194 88
rect 278 -88 312 88
rect 396 -88 430 88
<< psubdiff >>
rect -544 240 -448 274
rect 448 240 544 274
rect -544 178 -510 240
rect 510 178 544 240
rect -544 -240 -510 -178
rect 510 -240 544 -178
rect -544 -274 -448 -240
rect 448 -274 544 -240
<< psubdiffcont >>
rect -448 240 448 274
rect -544 -178 -510 178
rect 510 -178 544 178
rect -448 -274 448 -240
<< poly >>
rect -387 172 -321 188
rect -387 138 -371 172
rect -337 138 -321 172
rect -387 122 -321 138
rect -269 172 -203 188
rect -269 138 -253 172
rect -219 138 -203 172
rect -269 122 -203 138
rect -151 172 -85 188
rect -151 138 -135 172
rect -101 138 -85 172
rect -151 122 -85 138
rect -33 172 33 188
rect -33 138 -17 172
rect 17 138 33 172
rect -33 122 33 138
rect 85 172 151 188
rect 85 138 101 172
rect 135 138 151 172
rect 85 122 151 138
rect 203 172 269 188
rect 203 138 219 172
rect 253 138 269 172
rect 203 122 269 138
rect 321 172 387 188
rect 321 138 337 172
rect 371 138 387 172
rect 321 122 387 138
rect -384 100 -324 122
rect -266 100 -206 122
rect -148 100 -88 122
rect -30 100 30 122
rect 88 100 148 122
rect 206 100 266 122
rect 324 100 384 122
rect -384 -122 -324 -100
rect -266 -122 -206 -100
rect -148 -122 -88 -100
rect -30 -122 30 -100
rect 88 -122 148 -100
rect 206 -122 266 -100
rect 324 -122 384 -100
rect -387 -138 -321 -122
rect -387 -172 -371 -138
rect -337 -172 -321 -138
rect -387 -188 -321 -172
rect -269 -138 -203 -122
rect -269 -172 -253 -138
rect -219 -172 -203 -138
rect -269 -188 -203 -172
rect -151 -138 -85 -122
rect -151 -172 -135 -138
rect -101 -172 -85 -138
rect -151 -188 -85 -172
rect -33 -138 33 -122
rect -33 -172 -17 -138
rect 17 -172 33 -138
rect -33 -188 33 -172
rect 85 -138 151 -122
rect 85 -172 101 -138
rect 135 -172 151 -138
rect 85 -188 151 -172
rect 203 -138 269 -122
rect 203 -172 219 -138
rect 253 -172 269 -138
rect 203 -188 269 -172
rect 321 -138 387 -122
rect 321 -172 337 -138
rect 371 -172 387 -138
rect 321 -188 387 -172
<< polycont >>
rect -371 138 -337 172
rect -253 138 -219 172
rect -135 138 -101 172
rect -17 138 17 172
rect 101 138 135 172
rect 219 138 253 172
rect 337 138 371 172
rect -371 -172 -337 -138
rect -253 -172 -219 -138
rect -135 -172 -101 -138
rect -17 -172 17 -138
rect 101 -172 135 -138
rect 219 -172 253 -138
rect 337 -172 371 -138
<< locali >>
rect -544 240 -448 274
rect 448 240 544 274
rect -544 178 -510 240
rect 510 178 544 240
rect -387 138 -371 172
rect -337 138 -321 172
rect -269 138 -253 172
rect -219 138 -203 172
rect -151 138 -135 172
rect -101 138 -85 172
rect -33 138 -17 172
rect 17 138 33 172
rect 85 138 101 172
rect 135 138 151 172
rect 203 138 219 172
rect 253 138 269 172
rect 321 138 337 172
rect 371 138 387 172
rect -430 88 -396 104
rect -430 -104 -396 -88
rect -312 88 -278 104
rect -312 -104 -278 -88
rect -194 88 -160 104
rect -194 -104 -160 -88
rect -76 88 -42 104
rect -76 -104 -42 -88
rect 42 88 76 104
rect 42 -104 76 -88
rect 160 88 194 104
rect 160 -104 194 -88
rect 278 88 312 104
rect 278 -104 312 -88
rect 396 88 430 104
rect 396 -104 430 -88
rect -387 -172 -371 -138
rect -337 -172 -321 -138
rect -269 -172 -253 -138
rect -219 -172 -203 -138
rect -151 -172 -135 -138
rect -101 -172 -85 -138
rect -33 -172 -17 -138
rect 17 -172 33 -138
rect 85 -172 101 -138
rect 135 -172 151 -138
rect 203 -172 219 -138
rect 253 -172 269 -138
rect 321 -172 337 -138
rect 371 -172 387 -138
rect -544 -240 -510 -178
rect 510 -240 544 -178
rect -544 -274 -448 -240
rect 448 -274 544 -240
<< viali >>
rect -371 138 -337 172
rect -253 138 -219 172
rect -135 138 -101 172
rect -17 138 17 172
rect 101 138 135 172
rect 219 138 253 172
rect 337 138 371 172
rect -430 -88 -396 88
rect -312 -88 -278 88
rect -194 -88 -160 88
rect -76 -88 -42 88
rect 42 -88 76 88
rect 160 -88 194 88
rect 278 -88 312 88
rect 396 -88 430 88
rect -371 -172 -337 -138
rect -253 -172 -219 -138
rect -135 -172 -101 -138
rect -17 -172 17 -138
rect 101 -172 135 -138
rect 219 -172 253 -138
rect 337 -172 371 -138
<< metal1 >>
rect -383 172 -325 178
rect -383 138 -371 172
rect -337 138 -325 172
rect -383 132 -325 138
rect -265 172 -207 178
rect -265 138 -253 172
rect -219 138 -207 172
rect -265 132 -207 138
rect -147 172 -89 178
rect -147 138 -135 172
rect -101 138 -89 172
rect -147 132 -89 138
rect -29 172 29 178
rect -29 138 -17 172
rect 17 138 29 172
rect -29 132 29 138
rect 89 172 147 178
rect 89 138 101 172
rect 135 138 147 172
rect 89 132 147 138
rect 207 172 265 178
rect 207 138 219 172
rect 253 138 265 172
rect 207 132 265 138
rect 325 172 383 178
rect 325 138 337 172
rect 371 138 383 172
rect 325 132 383 138
rect -436 88 -390 100
rect -436 -88 -430 88
rect -396 -88 -390 88
rect -436 -100 -390 -88
rect -318 88 -272 100
rect -318 -88 -312 88
rect -278 -88 -272 88
rect -318 -100 -272 -88
rect -200 88 -154 100
rect -200 -88 -194 88
rect -160 -88 -154 88
rect -200 -100 -154 -88
rect -82 88 -36 100
rect -82 -88 -76 88
rect -42 -88 -36 88
rect -82 -100 -36 -88
rect 36 88 82 100
rect 36 -88 42 88
rect 76 -88 82 88
rect 36 -100 82 -88
rect 154 88 200 100
rect 154 -88 160 88
rect 194 -88 200 88
rect 154 -100 200 -88
rect 272 88 318 100
rect 272 -88 278 88
rect 312 -88 318 88
rect 272 -100 318 -88
rect 390 88 436 100
rect 390 -88 396 88
rect 430 -88 436 88
rect 390 -100 436 -88
rect -383 -138 -325 -132
rect -383 -172 -371 -138
rect -337 -172 -325 -138
rect -383 -178 -325 -172
rect -265 -138 -207 -132
rect -265 -172 -253 -138
rect -219 -172 -207 -138
rect -265 -178 -207 -172
rect -147 -138 -89 -132
rect -147 -172 -135 -138
rect -101 -172 -89 -138
rect -147 -178 -89 -172
rect -29 -138 29 -132
rect -29 -172 -17 -138
rect 17 -172 29 -138
rect -29 -178 29 -172
rect 89 -138 147 -132
rect 89 -172 101 -138
rect 135 -172 147 -138
rect 89 -178 147 -172
rect 207 -138 265 -132
rect 207 -172 219 -138
rect 253 -172 265 -138
rect 207 -178 265 -172
rect 325 -138 383 -132
rect 325 -172 337 -138
rect 371 -172 383 -138
rect 325 -178 383 -172
<< properties >>
string FIXED_BBOX -527 -257 527 257
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 0.3 m 1 nf 7 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
