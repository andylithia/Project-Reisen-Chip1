magic
tech sky130A
timestamp 1671334348
<< pwell >>
rect -142 -242 142 242
<< psubdiff >>
rect -124 207 -76 224
rect 76 207 124 224
rect -124 176 -107 207
rect 107 176 124 207
rect -124 -207 -107 -176
rect 107 -207 124 -176
rect -124 -224 -76 -207
rect 76 -224 124 -207
<< psubdiffcont >>
rect -76 207 76 224
rect -124 -176 -107 176
rect 107 -176 124 176
rect -76 -224 76 -207
<< xpolycontact >>
rect -59 -159 -24 57
rect 24 -159 59 57
<< xpolyres >>
rect -59 124 59 159
rect -59 57 -24 124
rect 24 57 59 124
<< locali >>
rect -124 207 -76 224
rect 76 207 124 224
rect -124 176 -107 207
rect 107 176 124 207
rect -124 -207 -107 -176
rect 107 -207 124 -176
rect -124 -224 -76 -207
rect 76 -224 124 -207
<< properties >>
string FIXED_BBOX -115 -215 115 215
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.35 l 0.5 m 1 nx 2 wmin 0.350 lmin 0.50 rho 2000 val 8.789k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 1 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
