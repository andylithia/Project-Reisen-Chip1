magic
tech sky130A
magscale 1 2
timestamp 1671152619
<< error_p >>
rect -2684 1081 -2626 1087
rect -2566 1081 -2508 1087
rect -2448 1081 -2390 1087
rect -2330 1081 -2272 1087
rect -2212 1081 -2154 1087
rect -2094 1081 -2036 1087
rect -1976 1081 -1918 1087
rect -1858 1081 -1800 1087
rect -1740 1081 -1682 1087
rect -1622 1081 -1564 1087
rect -1504 1081 -1446 1087
rect -1386 1081 -1328 1087
rect -1268 1081 -1210 1087
rect -1150 1081 -1092 1087
rect -1032 1081 -974 1087
rect -914 1081 -856 1087
rect -796 1081 -738 1087
rect -678 1081 -620 1087
rect -560 1081 -502 1087
rect -442 1081 -384 1087
rect -324 1081 -266 1087
rect -206 1081 -148 1087
rect -88 1081 -30 1087
rect 30 1081 88 1087
rect 148 1081 206 1087
rect 266 1081 324 1087
rect 384 1081 442 1087
rect 502 1081 560 1087
rect 620 1081 678 1087
rect 738 1081 796 1087
rect 856 1081 914 1087
rect 974 1081 1032 1087
rect 1092 1081 1150 1087
rect 1210 1081 1268 1087
rect 1328 1081 1386 1087
rect 1446 1081 1504 1087
rect 1564 1081 1622 1087
rect 1682 1081 1740 1087
rect 1800 1081 1858 1087
rect 1918 1081 1976 1087
rect 2036 1081 2094 1087
rect 2154 1081 2212 1087
rect 2272 1081 2330 1087
rect 2390 1081 2448 1087
rect 2508 1081 2566 1087
rect 2626 1081 2684 1087
rect -2684 1047 -2672 1081
rect -2566 1047 -2554 1081
rect -2448 1047 -2436 1081
rect -2330 1047 -2318 1081
rect -2212 1047 -2200 1081
rect -2094 1047 -2082 1081
rect -1976 1047 -1964 1081
rect -1858 1047 -1846 1081
rect -1740 1047 -1728 1081
rect -1622 1047 -1610 1081
rect -1504 1047 -1492 1081
rect -1386 1047 -1374 1081
rect -1268 1047 -1256 1081
rect -1150 1047 -1138 1081
rect -1032 1047 -1020 1081
rect -914 1047 -902 1081
rect -796 1047 -784 1081
rect -678 1047 -666 1081
rect -560 1047 -548 1081
rect -442 1047 -430 1081
rect -324 1047 -312 1081
rect -206 1047 -194 1081
rect -88 1047 -76 1081
rect 30 1047 42 1081
rect 148 1047 160 1081
rect 266 1047 278 1081
rect 384 1047 396 1081
rect 502 1047 514 1081
rect 620 1047 632 1081
rect 738 1047 750 1081
rect 856 1047 868 1081
rect 974 1047 986 1081
rect 1092 1047 1104 1081
rect 1210 1047 1222 1081
rect 1328 1047 1340 1081
rect 1446 1047 1458 1081
rect 1564 1047 1576 1081
rect 1682 1047 1694 1081
rect 1800 1047 1812 1081
rect 1918 1047 1930 1081
rect 2036 1047 2048 1081
rect 2154 1047 2166 1081
rect 2272 1047 2284 1081
rect 2390 1047 2402 1081
rect 2508 1047 2520 1081
rect 2626 1047 2638 1081
rect -2684 1041 -2626 1047
rect -2566 1041 -2508 1047
rect -2448 1041 -2390 1047
rect -2330 1041 -2272 1047
rect -2212 1041 -2154 1047
rect -2094 1041 -2036 1047
rect -1976 1041 -1918 1047
rect -1858 1041 -1800 1047
rect -1740 1041 -1682 1047
rect -1622 1041 -1564 1047
rect -1504 1041 -1446 1047
rect -1386 1041 -1328 1047
rect -1268 1041 -1210 1047
rect -1150 1041 -1092 1047
rect -1032 1041 -974 1047
rect -914 1041 -856 1047
rect -796 1041 -738 1047
rect -678 1041 -620 1047
rect -560 1041 -502 1047
rect -442 1041 -384 1047
rect -324 1041 -266 1047
rect -206 1041 -148 1047
rect -88 1041 -30 1047
rect 30 1041 88 1047
rect 148 1041 206 1047
rect 266 1041 324 1047
rect 384 1041 442 1047
rect 502 1041 560 1047
rect 620 1041 678 1047
rect 738 1041 796 1047
rect 856 1041 914 1047
rect 974 1041 1032 1047
rect 1092 1041 1150 1047
rect 1210 1041 1268 1047
rect 1328 1041 1386 1047
rect 1446 1041 1504 1047
rect 1564 1041 1622 1047
rect 1682 1041 1740 1047
rect 1800 1041 1858 1047
rect 1918 1041 1976 1047
rect 2036 1041 2094 1047
rect 2154 1041 2212 1047
rect 2272 1041 2330 1047
rect 2390 1041 2448 1047
rect 2508 1041 2566 1047
rect 2626 1041 2684 1047
rect -2684 -1047 -2626 -1041
rect -2566 -1047 -2508 -1041
rect -2448 -1047 -2390 -1041
rect -2330 -1047 -2272 -1041
rect -2212 -1047 -2154 -1041
rect -2094 -1047 -2036 -1041
rect -1976 -1047 -1918 -1041
rect -1858 -1047 -1800 -1041
rect -1740 -1047 -1682 -1041
rect -1622 -1047 -1564 -1041
rect -1504 -1047 -1446 -1041
rect -1386 -1047 -1328 -1041
rect -1268 -1047 -1210 -1041
rect -1150 -1047 -1092 -1041
rect -1032 -1047 -974 -1041
rect -914 -1047 -856 -1041
rect -796 -1047 -738 -1041
rect -678 -1047 -620 -1041
rect -560 -1047 -502 -1041
rect -442 -1047 -384 -1041
rect -324 -1047 -266 -1041
rect -206 -1047 -148 -1041
rect -88 -1047 -30 -1041
rect 30 -1047 88 -1041
rect 148 -1047 206 -1041
rect 266 -1047 324 -1041
rect 384 -1047 442 -1041
rect 502 -1047 560 -1041
rect 620 -1047 678 -1041
rect 738 -1047 796 -1041
rect 856 -1047 914 -1041
rect 974 -1047 1032 -1041
rect 1092 -1047 1150 -1041
rect 1210 -1047 1268 -1041
rect 1328 -1047 1386 -1041
rect 1446 -1047 1504 -1041
rect 1564 -1047 1622 -1041
rect 1682 -1047 1740 -1041
rect 1800 -1047 1858 -1041
rect 1918 -1047 1976 -1041
rect 2036 -1047 2094 -1041
rect 2154 -1047 2212 -1041
rect 2272 -1047 2330 -1041
rect 2390 -1047 2448 -1041
rect 2508 -1047 2566 -1041
rect 2626 -1047 2684 -1041
rect -2684 -1081 -2672 -1047
rect -2566 -1081 -2554 -1047
rect -2448 -1081 -2436 -1047
rect -2330 -1081 -2318 -1047
rect -2212 -1081 -2200 -1047
rect -2094 -1081 -2082 -1047
rect -1976 -1081 -1964 -1047
rect -1858 -1081 -1846 -1047
rect -1740 -1081 -1728 -1047
rect -1622 -1081 -1610 -1047
rect -1504 -1081 -1492 -1047
rect -1386 -1081 -1374 -1047
rect -1268 -1081 -1256 -1047
rect -1150 -1081 -1138 -1047
rect -1032 -1081 -1020 -1047
rect -914 -1081 -902 -1047
rect -796 -1081 -784 -1047
rect -678 -1081 -666 -1047
rect -560 -1081 -548 -1047
rect -442 -1081 -430 -1047
rect -324 -1081 -312 -1047
rect -206 -1081 -194 -1047
rect -88 -1081 -76 -1047
rect 30 -1081 42 -1047
rect 148 -1081 160 -1047
rect 266 -1081 278 -1047
rect 384 -1081 396 -1047
rect 502 -1081 514 -1047
rect 620 -1081 632 -1047
rect 738 -1081 750 -1047
rect 856 -1081 868 -1047
rect 974 -1081 986 -1047
rect 1092 -1081 1104 -1047
rect 1210 -1081 1222 -1047
rect 1328 -1081 1340 -1047
rect 1446 -1081 1458 -1047
rect 1564 -1081 1576 -1047
rect 1682 -1081 1694 -1047
rect 1800 -1081 1812 -1047
rect 1918 -1081 1930 -1047
rect 2036 -1081 2048 -1047
rect 2154 -1081 2166 -1047
rect 2272 -1081 2284 -1047
rect 2390 -1081 2402 -1047
rect 2508 -1081 2520 -1047
rect 2626 -1081 2638 -1047
rect -2684 -1087 -2626 -1081
rect -2566 -1087 -2508 -1081
rect -2448 -1087 -2390 -1081
rect -2330 -1087 -2272 -1081
rect -2212 -1087 -2154 -1081
rect -2094 -1087 -2036 -1081
rect -1976 -1087 -1918 -1081
rect -1858 -1087 -1800 -1081
rect -1740 -1087 -1682 -1081
rect -1622 -1087 -1564 -1081
rect -1504 -1087 -1446 -1081
rect -1386 -1087 -1328 -1081
rect -1268 -1087 -1210 -1081
rect -1150 -1087 -1092 -1081
rect -1032 -1087 -974 -1081
rect -914 -1087 -856 -1081
rect -796 -1087 -738 -1081
rect -678 -1087 -620 -1081
rect -560 -1087 -502 -1081
rect -442 -1087 -384 -1081
rect -324 -1087 -266 -1081
rect -206 -1087 -148 -1081
rect -88 -1087 -30 -1081
rect 30 -1087 88 -1081
rect 148 -1087 206 -1081
rect 266 -1087 324 -1081
rect 384 -1087 442 -1081
rect 502 -1087 560 -1081
rect 620 -1087 678 -1081
rect 738 -1087 796 -1081
rect 856 -1087 914 -1081
rect 974 -1087 1032 -1081
rect 1092 -1087 1150 -1081
rect 1210 -1087 1268 -1081
rect 1328 -1087 1386 -1081
rect 1446 -1087 1504 -1081
rect 1564 -1087 1622 -1081
rect 1682 -1087 1740 -1081
rect 1800 -1087 1858 -1081
rect 1918 -1087 1976 -1081
rect 2036 -1087 2094 -1081
rect 2154 -1087 2212 -1081
rect 2272 -1087 2330 -1081
rect 2390 -1087 2448 -1081
rect 2508 -1087 2566 -1081
rect 2626 -1087 2684 -1081
<< nwell >>
rect -2881 -1219 2881 1219
<< pmos >>
rect -2685 -1000 -2625 1000
rect -2567 -1000 -2507 1000
rect -2449 -1000 -2389 1000
rect -2331 -1000 -2271 1000
rect -2213 -1000 -2153 1000
rect -2095 -1000 -2035 1000
rect -1977 -1000 -1917 1000
rect -1859 -1000 -1799 1000
rect -1741 -1000 -1681 1000
rect -1623 -1000 -1563 1000
rect -1505 -1000 -1445 1000
rect -1387 -1000 -1327 1000
rect -1269 -1000 -1209 1000
rect -1151 -1000 -1091 1000
rect -1033 -1000 -973 1000
rect -915 -1000 -855 1000
rect -797 -1000 -737 1000
rect -679 -1000 -619 1000
rect -561 -1000 -501 1000
rect -443 -1000 -383 1000
rect -325 -1000 -265 1000
rect -207 -1000 -147 1000
rect -89 -1000 -29 1000
rect 29 -1000 89 1000
rect 147 -1000 207 1000
rect 265 -1000 325 1000
rect 383 -1000 443 1000
rect 501 -1000 561 1000
rect 619 -1000 679 1000
rect 737 -1000 797 1000
rect 855 -1000 915 1000
rect 973 -1000 1033 1000
rect 1091 -1000 1151 1000
rect 1209 -1000 1269 1000
rect 1327 -1000 1387 1000
rect 1445 -1000 1505 1000
rect 1563 -1000 1623 1000
rect 1681 -1000 1741 1000
rect 1799 -1000 1859 1000
rect 1917 -1000 1977 1000
rect 2035 -1000 2095 1000
rect 2153 -1000 2213 1000
rect 2271 -1000 2331 1000
rect 2389 -1000 2449 1000
rect 2507 -1000 2567 1000
rect 2625 -1000 2685 1000
<< pdiff >>
rect -2743 988 -2685 1000
rect -2743 -988 -2731 988
rect -2697 -988 -2685 988
rect -2743 -1000 -2685 -988
rect -2625 988 -2567 1000
rect -2625 -988 -2613 988
rect -2579 -988 -2567 988
rect -2625 -1000 -2567 -988
rect -2507 988 -2449 1000
rect -2507 -988 -2495 988
rect -2461 -988 -2449 988
rect -2507 -1000 -2449 -988
rect -2389 988 -2331 1000
rect -2389 -988 -2377 988
rect -2343 -988 -2331 988
rect -2389 -1000 -2331 -988
rect -2271 988 -2213 1000
rect -2271 -988 -2259 988
rect -2225 -988 -2213 988
rect -2271 -1000 -2213 -988
rect -2153 988 -2095 1000
rect -2153 -988 -2141 988
rect -2107 -988 -2095 988
rect -2153 -1000 -2095 -988
rect -2035 988 -1977 1000
rect -2035 -988 -2023 988
rect -1989 -988 -1977 988
rect -2035 -1000 -1977 -988
rect -1917 988 -1859 1000
rect -1917 -988 -1905 988
rect -1871 -988 -1859 988
rect -1917 -1000 -1859 -988
rect -1799 988 -1741 1000
rect -1799 -988 -1787 988
rect -1753 -988 -1741 988
rect -1799 -1000 -1741 -988
rect -1681 988 -1623 1000
rect -1681 -988 -1669 988
rect -1635 -988 -1623 988
rect -1681 -1000 -1623 -988
rect -1563 988 -1505 1000
rect -1563 -988 -1551 988
rect -1517 -988 -1505 988
rect -1563 -1000 -1505 -988
rect -1445 988 -1387 1000
rect -1445 -988 -1433 988
rect -1399 -988 -1387 988
rect -1445 -1000 -1387 -988
rect -1327 988 -1269 1000
rect -1327 -988 -1315 988
rect -1281 -988 -1269 988
rect -1327 -1000 -1269 -988
rect -1209 988 -1151 1000
rect -1209 -988 -1197 988
rect -1163 -988 -1151 988
rect -1209 -1000 -1151 -988
rect -1091 988 -1033 1000
rect -1091 -988 -1079 988
rect -1045 -988 -1033 988
rect -1091 -1000 -1033 -988
rect -973 988 -915 1000
rect -973 -988 -961 988
rect -927 -988 -915 988
rect -973 -1000 -915 -988
rect -855 988 -797 1000
rect -855 -988 -843 988
rect -809 -988 -797 988
rect -855 -1000 -797 -988
rect -737 988 -679 1000
rect -737 -988 -725 988
rect -691 -988 -679 988
rect -737 -1000 -679 -988
rect -619 988 -561 1000
rect -619 -988 -607 988
rect -573 -988 -561 988
rect -619 -1000 -561 -988
rect -501 988 -443 1000
rect -501 -988 -489 988
rect -455 -988 -443 988
rect -501 -1000 -443 -988
rect -383 988 -325 1000
rect -383 -988 -371 988
rect -337 -988 -325 988
rect -383 -1000 -325 -988
rect -265 988 -207 1000
rect -265 -988 -253 988
rect -219 -988 -207 988
rect -265 -1000 -207 -988
rect -147 988 -89 1000
rect -147 -988 -135 988
rect -101 -988 -89 988
rect -147 -1000 -89 -988
rect -29 988 29 1000
rect -29 -988 -17 988
rect 17 -988 29 988
rect -29 -1000 29 -988
rect 89 988 147 1000
rect 89 -988 101 988
rect 135 -988 147 988
rect 89 -1000 147 -988
rect 207 988 265 1000
rect 207 -988 219 988
rect 253 -988 265 988
rect 207 -1000 265 -988
rect 325 988 383 1000
rect 325 -988 337 988
rect 371 -988 383 988
rect 325 -1000 383 -988
rect 443 988 501 1000
rect 443 -988 455 988
rect 489 -988 501 988
rect 443 -1000 501 -988
rect 561 988 619 1000
rect 561 -988 573 988
rect 607 -988 619 988
rect 561 -1000 619 -988
rect 679 988 737 1000
rect 679 -988 691 988
rect 725 -988 737 988
rect 679 -1000 737 -988
rect 797 988 855 1000
rect 797 -988 809 988
rect 843 -988 855 988
rect 797 -1000 855 -988
rect 915 988 973 1000
rect 915 -988 927 988
rect 961 -988 973 988
rect 915 -1000 973 -988
rect 1033 988 1091 1000
rect 1033 -988 1045 988
rect 1079 -988 1091 988
rect 1033 -1000 1091 -988
rect 1151 988 1209 1000
rect 1151 -988 1163 988
rect 1197 -988 1209 988
rect 1151 -1000 1209 -988
rect 1269 988 1327 1000
rect 1269 -988 1281 988
rect 1315 -988 1327 988
rect 1269 -1000 1327 -988
rect 1387 988 1445 1000
rect 1387 -988 1399 988
rect 1433 -988 1445 988
rect 1387 -1000 1445 -988
rect 1505 988 1563 1000
rect 1505 -988 1517 988
rect 1551 -988 1563 988
rect 1505 -1000 1563 -988
rect 1623 988 1681 1000
rect 1623 -988 1635 988
rect 1669 -988 1681 988
rect 1623 -1000 1681 -988
rect 1741 988 1799 1000
rect 1741 -988 1753 988
rect 1787 -988 1799 988
rect 1741 -1000 1799 -988
rect 1859 988 1917 1000
rect 1859 -988 1871 988
rect 1905 -988 1917 988
rect 1859 -1000 1917 -988
rect 1977 988 2035 1000
rect 1977 -988 1989 988
rect 2023 -988 2035 988
rect 1977 -1000 2035 -988
rect 2095 988 2153 1000
rect 2095 -988 2107 988
rect 2141 -988 2153 988
rect 2095 -1000 2153 -988
rect 2213 988 2271 1000
rect 2213 -988 2225 988
rect 2259 -988 2271 988
rect 2213 -1000 2271 -988
rect 2331 988 2389 1000
rect 2331 -988 2343 988
rect 2377 -988 2389 988
rect 2331 -1000 2389 -988
rect 2449 988 2507 1000
rect 2449 -988 2461 988
rect 2495 -988 2507 988
rect 2449 -1000 2507 -988
rect 2567 988 2625 1000
rect 2567 -988 2579 988
rect 2613 -988 2625 988
rect 2567 -1000 2625 -988
rect 2685 988 2743 1000
rect 2685 -988 2697 988
rect 2731 -988 2743 988
rect 2685 -1000 2743 -988
<< pdiffc >>
rect -2731 -988 -2697 988
rect -2613 -988 -2579 988
rect -2495 -988 -2461 988
rect -2377 -988 -2343 988
rect -2259 -988 -2225 988
rect -2141 -988 -2107 988
rect -2023 -988 -1989 988
rect -1905 -988 -1871 988
rect -1787 -988 -1753 988
rect -1669 -988 -1635 988
rect -1551 -988 -1517 988
rect -1433 -988 -1399 988
rect -1315 -988 -1281 988
rect -1197 -988 -1163 988
rect -1079 -988 -1045 988
rect -961 -988 -927 988
rect -843 -988 -809 988
rect -725 -988 -691 988
rect -607 -988 -573 988
rect -489 -988 -455 988
rect -371 -988 -337 988
rect -253 -988 -219 988
rect -135 -988 -101 988
rect -17 -988 17 988
rect 101 -988 135 988
rect 219 -988 253 988
rect 337 -988 371 988
rect 455 -988 489 988
rect 573 -988 607 988
rect 691 -988 725 988
rect 809 -988 843 988
rect 927 -988 961 988
rect 1045 -988 1079 988
rect 1163 -988 1197 988
rect 1281 -988 1315 988
rect 1399 -988 1433 988
rect 1517 -988 1551 988
rect 1635 -988 1669 988
rect 1753 -988 1787 988
rect 1871 -988 1905 988
rect 1989 -988 2023 988
rect 2107 -988 2141 988
rect 2225 -988 2259 988
rect 2343 -988 2377 988
rect 2461 -988 2495 988
rect 2579 -988 2613 988
rect 2697 -988 2731 988
<< nsubdiff >>
rect -2845 1149 -2749 1183
rect 2749 1149 2845 1183
rect -2845 1087 -2811 1149
rect 2811 1087 2845 1149
rect -2845 -1149 -2811 -1087
rect 2811 -1149 2845 -1087
rect -2845 -1183 -2749 -1149
rect 2749 -1183 2845 -1149
<< nsubdiffcont >>
rect -2749 1149 2749 1183
rect -2845 -1087 -2811 1087
rect 2811 -1087 2845 1087
rect -2749 -1183 2749 -1149
<< poly >>
rect -2688 1081 -2622 1097
rect -2688 1047 -2672 1081
rect -2638 1047 -2622 1081
rect -2688 1031 -2622 1047
rect -2570 1081 -2504 1097
rect -2570 1047 -2554 1081
rect -2520 1047 -2504 1081
rect -2570 1031 -2504 1047
rect -2452 1081 -2386 1097
rect -2452 1047 -2436 1081
rect -2402 1047 -2386 1081
rect -2452 1031 -2386 1047
rect -2334 1081 -2268 1097
rect -2334 1047 -2318 1081
rect -2284 1047 -2268 1081
rect -2334 1031 -2268 1047
rect -2216 1081 -2150 1097
rect -2216 1047 -2200 1081
rect -2166 1047 -2150 1081
rect -2216 1031 -2150 1047
rect -2098 1081 -2032 1097
rect -2098 1047 -2082 1081
rect -2048 1047 -2032 1081
rect -2098 1031 -2032 1047
rect -1980 1081 -1914 1097
rect -1980 1047 -1964 1081
rect -1930 1047 -1914 1081
rect -1980 1031 -1914 1047
rect -1862 1081 -1796 1097
rect -1862 1047 -1846 1081
rect -1812 1047 -1796 1081
rect -1862 1031 -1796 1047
rect -1744 1081 -1678 1097
rect -1744 1047 -1728 1081
rect -1694 1047 -1678 1081
rect -1744 1031 -1678 1047
rect -1626 1081 -1560 1097
rect -1626 1047 -1610 1081
rect -1576 1047 -1560 1081
rect -1626 1031 -1560 1047
rect -1508 1081 -1442 1097
rect -1508 1047 -1492 1081
rect -1458 1047 -1442 1081
rect -1508 1031 -1442 1047
rect -1390 1081 -1324 1097
rect -1390 1047 -1374 1081
rect -1340 1047 -1324 1081
rect -1390 1031 -1324 1047
rect -1272 1081 -1206 1097
rect -1272 1047 -1256 1081
rect -1222 1047 -1206 1081
rect -1272 1031 -1206 1047
rect -1154 1081 -1088 1097
rect -1154 1047 -1138 1081
rect -1104 1047 -1088 1081
rect -1154 1031 -1088 1047
rect -1036 1081 -970 1097
rect -1036 1047 -1020 1081
rect -986 1047 -970 1081
rect -1036 1031 -970 1047
rect -918 1081 -852 1097
rect -918 1047 -902 1081
rect -868 1047 -852 1081
rect -918 1031 -852 1047
rect -800 1081 -734 1097
rect -800 1047 -784 1081
rect -750 1047 -734 1081
rect -800 1031 -734 1047
rect -682 1081 -616 1097
rect -682 1047 -666 1081
rect -632 1047 -616 1081
rect -682 1031 -616 1047
rect -564 1081 -498 1097
rect -564 1047 -548 1081
rect -514 1047 -498 1081
rect -564 1031 -498 1047
rect -446 1081 -380 1097
rect -446 1047 -430 1081
rect -396 1047 -380 1081
rect -446 1031 -380 1047
rect -328 1081 -262 1097
rect -328 1047 -312 1081
rect -278 1047 -262 1081
rect -328 1031 -262 1047
rect -210 1081 -144 1097
rect -210 1047 -194 1081
rect -160 1047 -144 1081
rect -210 1031 -144 1047
rect -92 1081 -26 1097
rect -92 1047 -76 1081
rect -42 1047 -26 1081
rect -92 1031 -26 1047
rect 26 1081 92 1097
rect 26 1047 42 1081
rect 76 1047 92 1081
rect 26 1031 92 1047
rect 144 1081 210 1097
rect 144 1047 160 1081
rect 194 1047 210 1081
rect 144 1031 210 1047
rect 262 1081 328 1097
rect 262 1047 278 1081
rect 312 1047 328 1081
rect 262 1031 328 1047
rect 380 1081 446 1097
rect 380 1047 396 1081
rect 430 1047 446 1081
rect 380 1031 446 1047
rect 498 1081 564 1097
rect 498 1047 514 1081
rect 548 1047 564 1081
rect 498 1031 564 1047
rect 616 1081 682 1097
rect 616 1047 632 1081
rect 666 1047 682 1081
rect 616 1031 682 1047
rect 734 1081 800 1097
rect 734 1047 750 1081
rect 784 1047 800 1081
rect 734 1031 800 1047
rect 852 1081 918 1097
rect 852 1047 868 1081
rect 902 1047 918 1081
rect 852 1031 918 1047
rect 970 1081 1036 1097
rect 970 1047 986 1081
rect 1020 1047 1036 1081
rect 970 1031 1036 1047
rect 1088 1081 1154 1097
rect 1088 1047 1104 1081
rect 1138 1047 1154 1081
rect 1088 1031 1154 1047
rect 1206 1081 1272 1097
rect 1206 1047 1222 1081
rect 1256 1047 1272 1081
rect 1206 1031 1272 1047
rect 1324 1081 1390 1097
rect 1324 1047 1340 1081
rect 1374 1047 1390 1081
rect 1324 1031 1390 1047
rect 1442 1081 1508 1097
rect 1442 1047 1458 1081
rect 1492 1047 1508 1081
rect 1442 1031 1508 1047
rect 1560 1081 1626 1097
rect 1560 1047 1576 1081
rect 1610 1047 1626 1081
rect 1560 1031 1626 1047
rect 1678 1081 1744 1097
rect 1678 1047 1694 1081
rect 1728 1047 1744 1081
rect 1678 1031 1744 1047
rect 1796 1081 1862 1097
rect 1796 1047 1812 1081
rect 1846 1047 1862 1081
rect 1796 1031 1862 1047
rect 1914 1081 1980 1097
rect 1914 1047 1930 1081
rect 1964 1047 1980 1081
rect 1914 1031 1980 1047
rect 2032 1081 2098 1097
rect 2032 1047 2048 1081
rect 2082 1047 2098 1081
rect 2032 1031 2098 1047
rect 2150 1081 2216 1097
rect 2150 1047 2166 1081
rect 2200 1047 2216 1081
rect 2150 1031 2216 1047
rect 2268 1081 2334 1097
rect 2268 1047 2284 1081
rect 2318 1047 2334 1081
rect 2268 1031 2334 1047
rect 2386 1081 2452 1097
rect 2386 1047 2402 1081
rect 2436 1047 2452 1081
rect 2386 1031 2452 1047
rect 2504 1081 2570 1097
rect 2504 1047 2520 1081
rect 2554 1047 2570 1081
rect 2504 1031 2570 1047
rect 2622 1081 2688 1097
rect 2622 1047 2638 1081
rect 2672 1047 2688 1081
rect 2622 1031 2688 1047
rect -2685 1000 -2625 1031
rect -2567 1000 -2507 1031
rect -2449 1000 -2389 1031
rect -2331 1000 -2271 1031
rect -2213 1000 -2153 1031
rect -2095 1000 -2035 1031
rect -1977 1000 -1917 1031
rect -1859 1000 -1799 1031
rect -1741 1000 -1681 1031
rect -1623 1000 -1563 1031
rect -1505 1000 -1445 1031
rect -1387 1000 -1327 1031
rect -1269 1000 -1209 1031
rect -1151 1000 -1091 1031
rect -1033 1000 -973 1031
rect -915 1000 -855 1031
rect -797 1000 -737 1031
rect -679 1000 -619 1031
rect -561 1000 -501 1031
rect -443 1000 -383 1031
rect -325 1000 -265 1031
rect -207 1000 -147 1031
rect -89 1000 -29 1031
rect 29 1000 89 1031
rect 147 1000 207 1031
rect 265 1000 325 1031
rect 383 1000 443 1031
rect 501 1000 561 1031
rect 619 1000 679 1031
rect 737 1000 797 1031
rect 855 1000 915 1031
rect 973 1000 1033 1031
rect 1091 1000 1151 1031
rect 1209 1000 1269 1031
rect 1327 1000 1387 1031
rect 1445 1000 1505 1031
rect 1563 1000 1623 1031
rect 1681 1000 1741 1031
rect 1799 1000 1859 1031
rect 1917 1000 1977 1031
rect 2035 1000 2095 1031
rect 2153 1000 2213 1031
rect 2271 1000 2331 1031
rect 2389 1000 2449 1031
rect 2507 1000 2567 1031
rect 2625 1000 2685 1031
rect -2685 -1031 -2625 -1000
rect -2567 -1031 -2507 -1000
rect -2449 -1031 -2389 -1000
rect -2331 -1031 -2271 -1000
rect -2213 -1031 -2153 -1000
rect -2095 -1031 -2035 -1000
rect -1977 -1031 -1917 -1000
rect -1859 -1031 -1799 -1000
rect -1741 -1031 -1681 -1000
rect -1623 -1031 -1563 -1000
rect -1505 -1031 -1445 -1000
rect -1387 -1031 -1327 -1000
rect -1269 -1031 -1209 -1000
rect -1151 -1031 -1091 -1000
rect -1033 -1031 -973 -1000
rect -915 -1031 -855 -1000
rect -797 -1031 -737 -1000
rect -679 -1031 -619 -1000
rect -561 -1031 -501 -1000
rect -443 -1031 -383 -1000
rect -325 -1031 -265 -1000
rect -207 -1031 -147 -1000
rect -89 -1031 -29 -1000
rect 29 -1031 89 -1000
rect 147 -1031 207 -1000
rect 265 -1031 325 -1000
rect 383 -1031 443 -1000
rect 501 -1031 561 -1000
rect 619 -1031 679 -1000
rect 737 -1031 797 -1000
rect 855 -1031 915 -1000
rect 973 -1031 1033 -1000
rect 1091 -1031 1151 -1000
rect 1209 -1031 1269 -1000
rect 1327 -1031 1387 -1000
rect 1445 -1031 1505 -1000
rect 1563 -1031 1623 -1000
rect 1681 -1031 1741 -1000
rect 1799 -1031 1859 -1000
rect 1917 -1031 1977 -1000
rect 2035 -1031 2095 -1000
rect 2153 -1031 2213 -1000
rect 2271 -1031 2331 -1000
rect 2389 -1031 2449 -1000
rect 2507 -1031 2567 -1000
rect 2625 -1031 2685 -1000
rect -2688 -1047 -2622 -1031
rect -2688 -1081 -2672 -1047
rect -2638 -1081 -2622 -1047
rect -2688 -1097 -2622 -1081
rect -2570 -1047 -2504 -1031
rect -2570 -1081 -2554 -1047
rect -2520 -1081 -2504 -1047
rect -2570 -1097 -2504 -1081
rect -2452 -1047 -2386 -1031
rect -2452 -1081 -2436 -1047
rect -2402 -1081 -2386 -1047
rect -2452 -1097 -2386 -1081
rect -2334 -1047 -2268 -1031
rect -2334 -1081 -2318 -1047
rect -2284 -1081 -2268 -1047
rect -2334 -1097 -2268 -1081
rect -2216 -1047 -2150 -1031
rect -2216 -1081 -2200 -1047
rect -2166 -1081 -2150 -1047
rect -2216 -1097 -2150 -1081
rect -2098 -1047 -2032 -1031
rect -2098 -1081 -2082 -1047
rect -2048 -1081 -2032 -1047
rect -2098 -1097 -2032 -1081
rect -1980 -1047 -1914 -1031
rect -1980 -1081 -1964 -1047
rect -1930 -1081 -1914 -1047
rect -1980 -1097 -1914 -1081
rect -1862 -1047 -1796 -1031
rect -1862 -1081 -1846 -1047
rect -1812 -1081 -1796 -1047
rect -1862 -1097 -1796 -1081
rect -1744 -1047 -1678 -1031
rect -1744 -1081 -1728 -1047
rect -1694 -1081 -1678 -1047
rect -1744 -1097 -1678 -1081
rect -1626 -1047 -1560 -1031
rect -1626 -1081 -1610 -1047
rect -1576 -1081 -1560 -1047
rect -1626 -1097 -1560 -1081
rect -1508 -1047 -1442 -1031
rect -1508 -1081 -1492 -1047
rect -1458 -1081 -1442 -1047
rect -1508 -1097 -1442 -1081
rect -1390 -1047 -1324 -1031
rect -1390 -1081 -1374 -1047
rect -1340 -1081 -1324 -1047
rect -1390 -1097 -1324 -1081
rect -1272 -1047 -1206 -1031
rect -1272 -1081 -1256 -1047
rect -1222 -1081 -1206 -1047
rect -1272 -1097 -1206 -1081
rect -1154 -1047 -1088 -1031
rect -1154 -1081 -1138 -1047
rect -1104 -1081 -1088 -1047
rect -1154 -1097 -1088 -1081
rect -1036 -1047 -970 -1031
rect -1036 -1081 -1020 -1047
rect -986 -1081 -970 -1047
rect -1036 -1097 -970 -1081
rect -918 -1047 -852 -1031
rect -918 -1081 -902 -1047
rect -868 -1081 -852 -1047
rect -918 -1097 -852 -1081
rect -800 -1047 -734 -1031
rect -800 -1081 -784 -1047
rect -750 -1081 -734 -1047
rect -800 -1097 -734 -1081
rect -682 -1047 -616 -1031
rect -682 -1081 -666 -1047
rect -632 -1081 -616 -1047
rect -682 -1097 -616 -1081
rect -564 -1047 -498 -1031
rect -564 -1081 -548 -1047
rect -514 -1081 -498 -1047
rect -564 -1097 -498 -1081
rect -446 -1047 -380 -1031
rect -446 -1081 -430 -1047
rect -396 -1081 -380 -1047
rect -446 -1097 -380 -1081
rect -328 -1047 -262 -1031
rect -328 -1081 -312 -1047
rect -278 -1081 -262 -1047
rect -328 -1097 -262 -1081
rect -210 -1047 -144 -1031
rect -210 -1081 -194 -1047
rect -160 -1081 -144 -1047
rect -210 -1097 -144 -1081
rect -92 -1047 -26 -1031
rect -92 -1081 -76 -1047
rect -42 -1081 -26 -1047
rect -92 -1097 -26 -1081
rect 26 -1047 92 -1031
rect 26 -1081 42 -1047
rect 76 -1081 92 -1047
rect 26 -1097 92 -1081
rect 144 -1047 210 -1031
rect 144 -1081 160 -1047
rect 194 -1081 210 -1047
rect 144 -1097 210 -1081
rect 262 -1047 328 -1031
rect 262 -1081 278 -1047
rect 312 -1081 328 -1047
rect 262 -1097 328 -1081
rect 380 -1047 446 -1031
rect 380 -1081 396 -1047
rect 430 -1081 446 -1047
rect 380 -1097 446 -1081
rect 498 -1047 564 -1031
rect 498 -1081 514 -1047
rect 548 -1081 564 -1047
rect 498 -1097 564 -1081
rect 616 -1047 682 -1031
rect 616 -1081 632 -1047
rect 666 -1081 682 -1047
rect 616 -1097 682 -1081
rect 734 -1047 800 -1031
rect 734 -1081 750 -1047
rect 784 -1081 800 -1047
rect 734 -1097 800 -1081
rect 852 -1047 918 -1031
rect 852 -1081 868 -1047
rect 902 -1081 918 -1047
rect 852 -1097 918 -1081
rect 970 -1047 1036 -1031
rect 970 -1081 986 -1047
rect 1020 -1081 1036 -1047
rect 970 -1097 1036 -1081
rect 1088 -1047 1154 -1031
rect 1088 -1081 1104 -1047
rect 1138 -1081 1154 -1047
rect 1088 -1097 1154 -1081
rect 1206 -1047 1272 -1031
rect 1206 -1081 1222 -1047
rect 1256 -1081 1272 -1047
rect 1206 -1097 1272 -1081
rect 1324 -1047 1390 -1031
rect 1324 -1081 1340 -1047
rect 1374 -1081 1390 -1047
rect 1324 -1097 1390 -1081
rect 1442 -1047 1508 -1031
rect 1442 -1081 1458 -1047
rect 1492 -1081 1508 -1047
rect 1442 -1097 1508 -1081
rect 1560 -1047 1626 -1031
rect 1560 -1081 1576 -1047
rect 1610 -1081 1626 -1047
rect 1560 -1097 1626 -1081
rect 1678 -1047 1744 -1031
rect 1678 -1081 1694 -1047
rect 1728 -1081 1744 -1047
rect 1678 -1097 1744 -1081
rect 1796 -1047 1862 -1031
rect 1796 -1081 1812 -1047
rect 1846 -1081 1862 -1047
rect 1796 -1097 1862 -1081
rect 1914 -1047 1980 -1031
rect 1914 -1081 1930 -1047
rect 1964 -1081 1980 -1047
rect 1914 -1097 1980 -1081
rect 2032 -1047 2098 -1031
rect 2032 -1081 2048 -1047
rect 2082 -1081 2098 -1047
rect 2032 -1097 2098 -1081
rect 2150 -1047 2216 -1031
rect 2150 -1081 2166 -1047
rect 2200 -1081 2216 -1047
rect 2150 -1097 2216 -1081
rect 2268 -1047 2334 -1031
rect 2268 -1081 2284 -1047
rect 2318 -1081 2334 -1047
rect 2268 -1097 2334 -1081
rect 2386 -1047 2452 -1031
rect 2386 -1081 2402 -1047
rect 2436 -1081 2452 -1047
rect 2386 -1097 2452 -1081
rect 2504 -1047 2570 -1031
rect 2504 -1081 2520 -1047
rect 2554 -1081 2570 -1047
rect 2504 -1097 2570 -1081
rect 2622 -1047 2688 -1031
rect 2622 -1081 2638 -1047
rect 2672 -1081 2688 -1047
rect 2622 -1097 2688 -1081
<< polycont >>
rect -2672 1047 -2638 1081
rect -2554 1047 -2520 1081
rect -2436 1047 -2402 1081
rect -2318 1047 -2284 1081
rect -2200 1047 -2166 1081
rect -2082 1047 -2048 1081
rect -1964 1047 -1930 1081
rect -1846 1047 -1812 1081
rect -1728 1047 -1694 1081
rect -1610 1047 -1576 1081
rect -1492 1047 -1458 1081
rect -1374 1047 -1340 1081
rect -1256 1047 -1222 1081
rect -1138 1047 -1104 1081
rect -1020 1047 -986 1081
rect -902 1047 -868 1081
rect -784 1047 -750 1081
rect -666 1047 -632 1081
rect -548 1047 -514 1081
rect -430 1047 -396 1081
rect -312 1047 -278 1081
rect -194 1047 -160 1081
rect -76 1047 -42 1081
rect 42 1047 76 1081
rect 160 1047 194 1081
rect 278 1047 312 1081
rect 396 1047 430 1081
rect 514 1047 548 1081
rect 632 1047 666 1081
rect 750 1047 784 1081
rect 868 1047 902 1081
rect 986 1047 1020 1081
rect 1104 1047 1138 1081
rect 1222 1047 1256 1081
rect 1340 1047 1374 1081
rect 1458 1047 1492 1081
rect 1576 1047 1610 1081
rect 1694 1047 1728 1081
rect 1812 1047 1846 1081
rect 1930 1047 1964 1081
rect 2048 1047 2082 1081
rect 2166 1047 2200 1081
rect 2284 1047 2318 1081
rect 2402 1047 2436 1081
rect 2520 1047 2554 1081
rect 2638 1047 2672 1081
rect -2672 -1081 -2638 -1047
rect -2554 -1081 -2520 -1047
rect -2436 -1081 -2402 -1047
rect -2318 -1081 -2284 -1047
rect -2200 -1081 -2166 -1047
rect -2082 -1081 -2048 -1047
rect -1964 -1081 -1930 -1047
rect -1846 -1081 -1812 -1047
rect -1728 -1081 -1694 -1047
rect -1610 -1081 -1576 -1047
rect -1492 -1081 -1458 -1047
rect -1374 -1081 -1340 -1047
rect -1256 -1081 -1222 -1047
rect -1138 -1081 -1104 -1047
rect -1020 -1081 -986 -1047
rect -902 -1081 -868 -1047
rect -784 -1081 -750 -1047
rect -666 -1081 -632 -1047
rect -548 -1081 -514 -1047
rect -430 -1081 -396 -1047
rect -312 -1081 -278 -1047
rect -194 -1081 -160 -1047
rect -76 -1081 -42 -1047
rect 42 -1081 76 -1047
rect 160 -1081 194 -1047
rect 278 -1081 312 -1047
rect 396 -1081 430 -1047
rect 514 -1081 548 -1047
rect 632 -1081 666 -1047
rect 750 -1081 784 -1047
rect 868 -1081 902 -1047
rect 986 -1081 1020 -1047
rect 1104 -1081 1138 -1047
rect 1222 -1081 1256 -1047
rect 1340 -1081 1374 -1047
rect 1458 -1081 1492 -1047
rect 1576 -1081 1610 -1047
rect 1694 -1081 1728 -1047
rect 1812 -1081 1846 -1047
rect 1930 -1081 1964 -1047
rect 2048 -1081 2082 -1047
rect 2166 -1081 2200 -1047
rect 2284 -1081 2318 -1047
rect 2402 -1081 2436 -1047
rect 2520 -1081 2554 -1047
rect 2638 -1081 2672 -1047
<< locali >>
rect -2845 1149 -2749 1183
rect 2749 1149 2845 1183
rect -2845 1087 -2811 1149
rect 2811 1087 2845 1149
rect -2688 1047 -2672 1081
rect -2638 1047 -2622 1081
rect -2570 1047 -2554 1081
rect -2520 1047 -2504 1081
rect -2452 1047 -2436 1081
rect -2402 1047 -2386 1081
rect -2334 1047 -2318 1081
rect -2284 1047 -2268 1081
rect -2216 1047 -2200 1081
rect -2166 1047 -2150 1081
rect -2098 1047 -2082 1081
rect -2048 1047 -2032 1081
rect -1980 1047 -1964 1081
rect -1930 1047 -1914 1081
rect -1862 1047 -1846 1081
rect -1812 1047 -1796 1081
rect -1744 1047 -1728 1081
rect -1694 1047 -1678 1081
rect -1626 1047 -1610 1081
rect -1576 1047 -1560 1081
rect -1508 1047 -1492 1081
rect -1458 1047 -1442 1081
rect -1390 1047 -1374 1081
rect -1340 1047 -1324 1081
rect -1272 1047 -1256 1081
rect -1222 1047 -1206 1081
rect -1154 1047 -1138 1081
rect -1104 1047 -1088 1081
rect -1036 1047 -1020 1081
rect -986 1047 -970 1081
rect -918 1047 -902 1081
rect -868 1047 -852 1081
rect -800 1047 -784 1081
rect -750 1047 -734 1081
rect -682 1047 -666 1081
rect -632 1047 -616 1081
rect -564 1047 -548 1081
rect -514 1047 -498 1081
rect -446 1047 -430 1081
rect -396 1047 -380 1081
rect -328 1047 -312 1081
rect -278 1047 -262 1081
rect -210 1047 -194 1081
rect -160 1047 -144 1081
rect -92 1047 -76 1081
rect -42 1047 -26 1081
rect 26 1047 42 1081
rect 76 1047 92 1081
rect 144 1047 160 1081
rect 194 1047 210 1081
rect 262 1047 278 1081
rect 312 1047 328 1081
rect 380 1047 396 1081
rect 430 1047 446 1081
rect 498 1047 514 1081
rect 548 1047 564 1081
rect 616 1047 632 1081
rect 666 1047 682 1081
rect 734 1047 750 1081
rect 784 1047 800 1081
rect 852 1047 868 1081
rect 902 1047 918 1081
rect 970 1047 986 1081
rect 1020 1047 1036 1081
rect 1088 1047 1104 1081
rect 1138 1047 1154 1081
rect 1206 1047 1222 1081
rect 1256 1047 1272 1081
rect 1324 1047 1340 1081
rect 1374 1047 1390 1081
rect 1442 1047 1458 1081
rect 1492 1047 1508 1081
rect 1560 1047 1576 1081
rect 1610 1047 1626 1081
rect 1678 1047 1694 1081
rect 1728 1047 1744 1081
rect 1796 1047 1812 1081
rect 1846 1047 1862 1081
rect 1914 1047 1930 1081
rect 1964 1047 1980 1081
rect 2032 1047 2048 1081
rect 2082 1047 2098 1081
rect 2150 1047 2166 1081
rect 2200 1047 2216 1081
rect 2268 1047 2284 1081
rect 2318 1047 2334 1081
rect 2386 1047 2402 1081
rect 2436 1047 2452 1081
rect 2504 1047 2520 1081
rect 2554 1047 2570 1081
rect 2622 1047 2638 1081
rect 2672 1047 2688 1081
rect -2731 988 -2697 1004
rect -2731 -1004 -2697 -988
rect -2613 988 -2579 1004
rect -2613 -1004 -2579 -988
rect -2495 988 -2461 1004
rect -2495 -1004 -2461 -988
rect -2377 988 -2343 1004
rect -2377 -1004 -2343 -988
rect -2259 988 -2225 1004
rect -2259 -1004 -2225 -988
rect -2141 988 -2107 1004
rect -2141 -1004 -2107 -988
rect -2023 988 -1989 1004
rect -2023 -1004 -1989 -988
rect -1905 988 -1871 1004
rect -1905 -1004 -1871 -988
rect -1787 988 -1753 1004
rect -1787 -1004 -1753 -988
rect -1669 988 -1635 1004
rect -1669 -1004 -1635 -988
rect -1551 988 -1517 1004
rect -1551 -1004 -1517 -988
rect -1433 988 -1399 1004
rect -1433 -1004 -1399 -988
rect -1315 988 -1281 1004
rect -1315 -1004 -1281 -988
rect -1197 988 -1163 1004
rect -1197 -1004 -1163 -988
rect -1079 988 -1045 1004
rect -1079 -1004 -1045 -988
rect -961 988 -927 1004
rect -961 -1004 -927 -988
rect -843 988 -809 1004
rect -843 -1004 -809 -988
rect -725 988 -691 1004
rect -725 -1004 -691 -988
rect -607 988 -573 1004
rect -607 -1004 -573 -988
rect -489 988 -455 1004
rect -489 -1004 -455 -988
rect -371 988 -337 1004
rect -371 -1004 -337 -988
rect -253 988 -219 1004
rect -253 -1004 -219 -988
rect -135 988 -101 1004
rect -135 -1004 -101 -988
rect -17 988 17 1004
rect -17 -1004 17 -988
rect 101 988 135 1004
rect 101 -1004 135 -988
rect 219 988 253 1004
rect 219 -1004 253 -988
rect 337 988 371 1004
rect 337 -1004 371 -988
rect 455 988 489 1004
rect 455 -1004 489 -988
rect 573 988 607 1004
rect 573 -1004 607 -988
rect 691 988 725 1004
rect 691 -1004 725 -988
rect 809 988 843 1004
rect 809 -1004 843 -988
rect 927 988 961 1004
rect 927 -1004 961 -988
rect 1045 988 1079 1004
rect 1045 -1004 1079 -988
rect 1163 988 1197 1004
rect 1163 -1004 1197 -988
rect 1281 988 1315 1004
rect 1281 -1004 1315 -988
rect 1399 988 1433 1004
rect 1399 -1004 1433 -988
rect 1517 988 1551 1004
rect 1517 -1004 1551 -988
rect 1635 988 1669 1004
rect 1635 -1004 1669 -988
rect 1753 988 1787 1004
rect 1753 -1004 1787 -988
rect 1871 988 1905 1004
rect 1871 -1004 1905 -988
rect 1989 988 2023 1004
rect 1989 -1004 2023 -988
rect 2107 988 2141 1004
rect 2107 -1004 2141 -988
rect 2225 988 2259 1004
rect 2225 -1004 2259 -988
rect 2343 988 2377 1004
rect 2343 -1004 2377 -988
rect 2461 988 2495 1004
rect 2461 -1004 2495 -988
rect 2579 988 2613 1004
rect 2579 -1004 2613 -988
rect 2697 988 2731 1004
rect 2697 -1004 2731 -988
rect -2688 -1081 -2672 -1047
rect -2638 -1081 -2622 -1047
rect -2570 -1081 -2554 -1047
rect -2520 -1081 -2504 -1047
rect -2452 -1081 -2436 -1047
rect -2402 -1081 -2386 -1047
rect -2334 -1081 -2318 -1047
rect -2284 -1081 -2268 -1047
rect -2216 -1081 -2200 -1047
rect -2166 -1081 -2150 -1047
rect -2098 -1081 -2082 -1047
rect -2048 -1081 -2032 -1047
rect -1980 -1081 -1964 -1047
rect -1930 -1081 -1914 -1047
rect -1862 -1081 -1846 -1047
rect -1812 -1081 -1796 -1047
rect -1744 -1081 -1728 -1047
rect -1694 -1081 -1678 -1047
rect -1626 -1081 -1610 -1047
rect -1576 -1081 -1560 -1047
rect -1508 -1081 -1492 -1047
rect -1458 -1081 -1442 -1047
rect -1390 -1081 -1374 -1047
rect -1340 -1081 -1324 -1047
rect -1272 -1081 -1256 -1047
rect -1222 -1081 -1206 -1047
rect -1154 -1081 -1138 -1047
rect -1104 -1081 -1088 -1047
rect -1036 -1081 -1020 -1047
rect -986 -1081 -970 -1047
rect -918 -1081 -902 -1047
rect -868 -1081 -852 -1047
rect -800 -1081 -784 -1047
rect -750 -1081 -734 -1047
rect -682 -1081 -666 -1047
rect -632 -1081 -616 -1047
rect -564 -1081 -548 -1047
rect -514 -1081 -498 -1047
rect -446 -1081 -430 -1047
rect -396 -1081 -380 -1047
rect -328 -1081 -312 -1047
rect -278 -1081 -262 -1047
rect -210 -1081 -194 -1047
rect -160 -1081 -144 -1047
rect -92 -1081 -76 -1047
rect -42 -1081 -26 -1047
rect 26 -1081 42 -1047
rect 76 -1081 92 -1047
rect 144 -1081 160 -1047
rect 194 -1081 210 -1047
rect 262 -1081 278 -1047
rect 312 -1081 328 -1047
rect 380 -1081 396 -1047
rect 430 -1081 446 -1047
rect 498 -1081 514 -1047
rect 548 -1081 564 -1047
rect 616 -1081 632 -1047
rect 666 -1081 682 -1047
rect 734 -1081 750 -1047
rect 784 -1081 800 -1047
rect 852 -1081 868 -1047
rect 902 -1081 918 -1047
rect 970 -1081 986 -1047
rect 1020 -1081 1036 -1047
rect 1088 -1081 1104 -1047
rect 1138 -1081 1154 -1047
rect 1206 -1081 1222 -1047
rect 1256 -1081 1272 -1047
rect 1324 -1081 1340 -1047
rect 1374 -1081 1390 -1047
rect 1442 -1081 1458 -1047
rect 1492 -1081 1508 -1047
rect 1560 -1081 1576 -1047
rect 1610 -1081 1626 -1047
rect 1678 -1081 1694 -1047
rect 1728 -1081 1744 -1047
rect 1796 -1081 1812 -1047
rect 1846 -1081 1862 -1047
rect 1914 -1081 1930 -1047
rect 1964 -1081 1980 -1047
rect 2032 -1081 2048 -1047
rect 2082 -1081 2098 -1047
rect 2150 -1081 2166 -1047
rect 2200 -1081 2216 -1047
rect 2268 -1081 2284 -1047
rect 2318 -1081 2334 -1047
rect 2386 -1081 2402 -1047
rect 2436 -1081 2452 -1047
rect 2504 -1081 2520 -1047
rect 2554 -1081 2570 -1047
rect 2622 -1081 2638 -1047
rect 2672 -1081 2688 -1047
rect -2845 -1149 -2811 -1087
rect 2811 -1149 2845 -1087
rect -2845 -1183 -2749 -1149
rect 2749 -1183 2845 -1149
<< viali >>
rect -2672 1047 -2638 1081
rect -2554 1047 -2520 1081
rect -2436 1047 -2402 1081
rect -2318 1047 -2284 1081
rect -2200 1047 -2166 1081
rect -2082 1047 -2048 1081
rect -1964 1047 -1930 1081
rect -1846 1047 -1812 1081
rect -1728 1047 -1694 1081
rect -1610 1047 -1576 1081
rect -1492 1047 -1458 1081
rect -1374 1047 -1340 1081
rect -1256 1047 -1222 1081
rect -1138 1047 -1104 1081
rect -1020 1047 -986 1081
rect -902 1047 -868 1081
rect -784 1047 -750 1081
rect -666 1047 -632 1081
rect -548 1047 -514 1081
rect -430 1047 -396 1081
rect -312 1047 -278 1081
rect -194 1047 -160 1081
rect -76 1047 -42 1081
rect 42 1047 76 1081
rect 160 1047 194 1081
rect 278 1047 312 1081
rect 396 1047 430 1081
rect 514 1047 548 1081
rect 632 1047 666 1081
rect 750 1047 784 1081
rect 868 1047 902 1081
rect 986 1047 1020 1081
rect 1104 1047 1138 1081
rect 1222 1047 1256 1081
rect 1340 1047 1374 1081
rect 1458 1047 1492 1081
rect 1576 1047 1610 1081
rect 1694 1047 1728 1081
rect 1812 1047 1846 1081
rect 1930 1047 1964 1081
rect 2048 1047 2082 1081
rect 2166 1047 2200 1081
rect 2284 1047 2318 1081
rect 2402 1047 2436 1081
rect 2520 1047 2554 1081
rect 2638 1047 2672 1081
rect -2731 -988 -2697 988
rect -2613 -988 -2579 988
rect -2495 -988 -2461 988
rect -2377 -988 -2343 988
rect -2259 -988 -2225 988
rect -2141 -988 -2107 988
rect -2023 -988 -1989 988
rect -1905 -988 -1871 988
rect -1787 -988 -1753 988
rect -1669 -988 -1635 988
rect -1551 -988 -1517 988
rect -1433 -988 -1399 988
rect -1315 -988 -1281 988
rect -1197 -988 -1163 988
rect -1079 -988 -1045 988
rect -961 -988 -927 988
rect -843 -988 -809 988
rect -725 -988 -691 988
rect -607 -988 -573 988
rect -489 -988 -455 988
rect -371 -988 -337 988
rect -253 -988 -219 988
rect -135 -988 -101 988
rect -17 -988 17 988
rect 101 -988 135 988
rect 219 -988 253 988
rect 337 -988 371 988
rect 455 -988 489 988
rect 573 -988 607 988
rect 691 -988 725 988
rect 809 -988 843 988
rect 927 -988 961 988
rect 1045 -988 1079 988
rect 1163 -988 1197 988
rect 1281 -988 1315 988
rect 1399 -988 1433 988
rect 1517 -988 1551 988
rect 1635 -988 1669 988
rect 1753 -988 1787 988
rect 1871 -988 1905 988
rect 1989 -988 2023 988
rect 2107 -988 2141 988
rect 2225 -988 2259 988
rect 2343 -988 2377 988
rect 2461 -988 2495 988
rect 2579 -988 2613 988
rect 2697 -988 2731 988
rect -2672 -1081 -2638 -1047
rect -2554 -1081 -2520 -1047
rect -2436 -1081 -2402 -1047
rect -2318 -1081 -2284 -1047
rect -2200 -1081 -2166 -1047
rect -2082 -1081 -2048 -1047
rect -1964 -1081 -1930 -1047
rect -1846 -1081 -1812 -1047
rect -1728 -1081 -1694 -1047
rect -1610 -1081 -1576 -1047
rect -1492 -1081 -1458 -1047
rect -1374 -1081 -1340 -1047
rect -1256 -1081 -1222 -1047
rect -1138 -1081 -1104 -1047
rect -1020 -1081 -986 -1047
rect -902 -1081 -868 -1047
rect -784 -1081 -750 -1047
rect -666 -1081 -632 -1047
rect -548 -1081 -514 -1047
rect -430 -1081 -396 -1047
rect -312 -1081 -278 -1047
rect -194 -1081 -160 -1047
rect -76 -1081 -42 -1047
rect 42 -1081 76 -1047
rect 160 -1081 194 -1047
rect 278 -1081 312 -1047
rect 396 -1081 430 -1047
rect 514 -1081 548 -1047
rect 632 -1081 666 -1047
rect 750 -1081 784 -1047
rect 868 -1081 902 -1047
rect 986 -1081 1020 -1047
rect 1104 -1081 1138 -1047
rect 1222 -1081 1256 -1047
rect 1340 -1081 1374 -1047
rect 1458 -1081 1492 -1047
rect 1576 -1081 1610 -1047
rect 1694 -1081 1728 -1047
rect 1812 -1081 1846 -1047
rect 1930 -1081 1964 -1047
rect 2048 -1081 2082 -1047
rect 2166 -1081 2200 -1047
rect 2284 -1081 2318 -1047
rect 2402 -1081 2436 -1047
rect 2520 -1081 2554 -1047
rect 2638 -1081 2672 -1047
<< metal1 >>
rect -2684 1081 -2626 1087
rect -2684 1047 -2672 1081
rect -2638 1047 -2626 1081
rect -2684 1041 -2626 1047
rect -2566 1081 -2508 1087
rect -2566 1047 -2554 1081
rect -2520 1047 -2508 1081
rect -2566 1041 -2508 1047
rect -2448 1081 -2390 1087
rect -2448 1047 -2436 1081
rect -2402 1047 -2390 1081
rect -2448 1041 -2390 1047
rect -2330 1081 -2272 1087
rect -2330 1047 -2318 1081
rect -2284 1047 -2272 1081
rect -2330 1041 -2272 1047
rect -2212 1081 -2154 1087
rect -2212 1047 -2200 1081
rect -2166 1047 -2154 1081
rect -2212 1041 -2154 1047
rect -2094 1081 -2036 1087
rect -2094 1047 -2082 1081
rect -2048 1047 -2036 1081
rect -2094 1041 -2036 1047
rect -1976 1081 -1918 1087
rect -1976 1047 -1964 1081
rect -1930 1047 -1918 1081
rect -1976 1041 -1918 1047
rect -1858 1081 -1800 1087
rect -1858 1047 -1846 1081
rect -1812 1047 -1800 1081
rect -1858 1041 -1800 1047
rect -1740 1081 -1682 1087
rect -1740 1047 -1728 1081
rect -1694 1047 -1682 1081
rect -1740 1041 -1682 1047
rect -1622 1081 -1564 1087
rect -1622 1047 -1610 1081
rect -1576 1047 -1564 1081
rect -1622 1041 -1564 1047
rect -1504 1081 -1446 1087
rect -1504 1047 -1492 1081
rect -1458 1047 -1446 1081
rect -1504 1041 -1446 1047
rect -1386 1081 -1328 1087
rect -1386 1047 -1374 1081
rect -1340 1047 -1328 1081
rect -1386 1041 -1328 1047
rect -1268 1081 -1210 1087
rect -1268 1047 -1256 1081
rect -1222 1047 -1210 1081
rect -1268 1041 -1210 1047
rect -1150 1081 -1092 1087
rect -1150 1047 -1138 1081
rect -1104 1047 -1092 1081
rect -1150 1041 -1092 1047
rect -1032 1081 -974 1087
rect -1032 1047 -1020 1081
rect -986 1047 -974 1081
rect -1032 1041 -974 1047
rect -914 1081 -856 1087
rect -914 1047 -902 1081
rect -868 1047 -856 1081
rect -914 1041 -856 1047
rect -796 1081 -738 1087
rect -796 1047 -784 1081
rect -750 1047 -738 1081
rect -796 1041 -738 1047
rect -678 1081 -620 1087
rect -678 1047 -666 1081
rect -632 1047 -620 1081
rect -678 1041 -620 1047
rect -560 1081 -502 1087
rect -560 1047 -548 1081
rect -514 1047 -502 1081
rect -560 1041 -502 1047
rect -442 1081 -384 1087
rect -442 1047 -430 1081
rect -396 1047 -384 1081
rect -442 1041 -384 1047
rect -324 1081 -266 1087
rect -324 1047 -312 1081
rect -278 1047 -266 1081
rect -324 1041 -266 1047
rect -206 1081 -148 1087
rect -206 1047 -194 1081
rect -160 1047 -148 1081
rect -206 1041 -148 1047
rect -88 1081 -30 1087
rect -88 1047 -76 1081
rect -42 1047 -30 1081
rect -88 1041 -30 1047
rect 30 1081 88 1087
rect 30 1047 42 1081
rect 76 1047 88 1081
rect 30 1041 88 1047
rect 148 1081 206 1087
rect 148 1047 160 1081
rect 194 1047 206 1081
rect 148 1041 206 1047
rect 266 1081 324 1087
rect 266 1047 278 1081
rect 312 1047 324 1081
rect 266 1041 324 1047
rect 384 1081 442 1087
rect 384 1047 396 1081
rect 430 1047 442 1081
rect 384 1041 442 1047
rect 502 1081 560 1087
rect 502 1047 514 1081
rect 548 1047 560 1081
rect 502 1041 560 1047
rect 620 1081 678 1087
rect 620 1047 632 1081
rect 666 1047 678 1081
rect 620 1041 678 1047
rect 738 1081 796 1087
rect 738 1047 750 1081
rect 784 1047 796 1081
rect 738 1041 796 1047
rect 856 1081 914 1087
rect 856 1047 868 1081
rect 902 1047 914 1081
rect 856 1041 914 1047
rect 974 1081 1032 1087
rect 974 1047 986 1081
rect 1020 1047 1032 1081
rect 974 1041 1032 1047
rect 1092 1081 1150 1087
rect 1092 1047 1104 1081
rect 1138 1047 1150 1081
rect 1092 1041 1150 1047
rect 1210 1081 1268 1087
rect 1210 1047 1222 1081
rect 1256 1047 1268 1081
rect 1210 1041 1268 1047
rect 1328 1081 1386 1087
rect 1328 1047 1340 1081
rect 1374 1047 1386 1081
rect 1328 1041 1386 1047
rect 1446 1081 1504 1087
rect 1446 1047 1458 1081
rect 1492 1047 1504 1081
rect 1446 1041 1504 1047
rect 1564 1081 1622 1087
rect 1564 1047 1576 1081
rect 1610 1047 1622 1081
rect 1564 1041 1622 1047
rect 1682 1081 1740 1087
rect 1682 1047 1694 1081
rect 1728 1047 1740 1081
rect 1682 1041 1740 1047
rect 1800 1081 1858 1087
rect 1800 1047 1812 1081
rect 1846 1047 1858 1081
rect 1800 1041 1858 1047
rect 1918 1081 1976 1087
rect 1918 1047 1930 1081
rect 1964 1047 1976 1081
rect 1918 1041 1976 1047
rect 2036 1081 2094 1087
rect 2036 1047 2048 1081
rect 2082 1047 2094 1081
rect 2036 1041 2094 1047
rect 2154 1081 2212 1087
rect 2154 1047 2166 1081
rect 2200 1047 2212 1081
rect 2154 1041 2212 1047
rect 2272 1081 2330 1087
rect 2272 1047 2284 1081
rect 2318 1047 2330 1081
rect 2272 1041 2330 1047
rect 2390 1081 2448 1087
rect 2390 1047 2402 1081
rect 2436 1047 2448 1081
rect 2390 1041 2448 1047
rect 2508 1081 2566 1087
rect 2508 1047 2520 1081
rect 2554 1047 2566 1081
rect 2508 1041 2566 1047
rect 2626 1081 2684 1087
rect 2626 1047 2638 1081
rect 2672 1047 2684 1081
rect 2626 1041 2684 1047
rect -2737 988 -2691 1000
rect -2737 -988 -2731 988
rect -2697 -988 -2691 988
rect -2737 -1000 -2691 -988
rect -2619 988 -2573 1000
rect -2619 -988 -2613 988
rect -2579 -988 -2573 988
rect -2619 -1000 -2573 -988
rect -2501 988 -2455 1000
rect -2501 -988 -2495 988
rect -2461 -988 -2455 988
rect -2501 -1000 -2455 -988
rect -2383 988 -2337 1000
rect -2383 -988 -2377 988
rect -2343 -988 -2337 988
rect -2383 -1000 -2337 -988
rect -2265 988 -2219 1000
rect -2265 -988 -2259 988
rect -2225 -988 -2219 988
rect -2265 -1000 -2219 -988
rect -2147 988 -2101 1000
rect -2147 -988 -2141 988
rect -2107 -988 -2101 988
rect -2147 -1000 -2101 -988
rect -2029 988 -1983 1000
rect -2029 -988 -2023 988
rect -1989 -988 -1983 988
rect -2029 -1000 -1983 -988
rect -1911 988 -1865 1000
rect -1911 -988 -1905 988
rect -1871 -988 -1865 988
rect -1911 -1000 -1865 -988
rect -1793 988 -1747 1000
rect -1793 -988 -1787 988
rect -1753 -988 -1747 988
rect -1793 -1000 -1747 -988
rect -1675 988 -1629 1000
rect -1675 -988 -1669 988
rect -1635 -988 -1629 988
rect -1675 -1000 -1629 -988
rect -1557 988 -1511 1000
rect -1557 -988 -1551 988
rect -1517 -988 -1511 988
rect -1557 -1000 -1511 -988
rect -1439 988 -1393 1000
rect -1439 -988 -1433 988
rect -1399 -988 -1393 988
rect -1439 -1000 -1393 -988
rect -1321 988 -1275 1000
rect -1321 -988 -1315 988
rect -1281 -988 -1275 988
rect -1321 -1000 -1275 -988
rect -1203 988 -1157 1000
rect -1203 -988 -1197 988
rect -1163 -988 -1157 988
rect -1203 -1000 -1157 -988
rect -1085 988 -1039 1000
rect -1085 -988 -1079 988
rect -1045 -988 -1039 988
rect -1085 -1000 -1039 -988
rect -967 988 -921 1000
rect -967 -988 -961 988
rect -927 -988 -921 988
rect -967 -1000 -921 -988
rect -849 988 -803 1000
rect -849 -988 -843 988
rect -809 -988 -803 988
rect -849 -1000 -803 -988
rect -731 988 -685 1000
rect -731 -988 -725 988
rect -691 -988 -685 988
rect -731 -1000 -685 -988
rect -613 988 -567 1000
rect -613 -988 -607 988
rect -573 -988 -567 988
rect -613 -1000 -567 -988
rect -495 988 -449 1000
rect -495 -988 -489 988
rect -455 -988 -449 988
rect -495 -1000 -449 -988
rect -377 988 -331 1000
rect -377 -988 -371 988
rect -337 -988 -331 988
rect -377 -1000 -331 -988
rect -259 988 -213 1000
rect -259 -988 -253 988
rect -219 -988 -213 988
rect -259 -1000 -213 -988
rect -141 988 -95 1000
rect -141 -988 -135 988
rect -101 -988 -95 988
rect -141 -1000 -95 -988
rect -23 988 23 1000
rect -23 -988 -17 988
rect 17 -988 23 988
rect -23 -1000 23 -988
rect 95 988 141 1000
rect 95 -988 101 988
rect 135 -988 141 988
rect 95 -1000 141 -988
rect 213 988 259 1000
rect 213 -988 219 988
rect 253 -988 259 988
rect 213 -1000 259 -988
rect 331 988 377 1000
rect 331 -988 337 988
rect 371 -988 377 988
rect 331 -1000 377 -988
rect 449 988 495 1000
rect 449 -988 455 988
rect 489 -988 495 988
rect 449 -1000 495 -988
rect 567 988 613 1000
rect 567 -988 573 988
rect 607 -988 613 988
rect 567 -1000 613 -988
rect 685 988 731 1000
rect 685 -988 691 988
rect 725 -988 731 988
rect 685 -1000 731 -988
rect 803 988 849 1000
rect 803 -988 809 988
rect 843 -988 849 988
rect 803 -1000 849 -988
rect 921 988 967 1000
rect 921 -988 927 988
rect 961 -988 967 988
rect 921 -1000 967 -988
rect 1039 988 1085 1000
rect 1039 -988 1045 988
rect 1079 -988 1085 988
rect 1039 -1000 1085 -988
rect 1157 988 1203 1000
rect 1157 -988 1163 988
rect 1197 -988 1203 988
rect 1157 -1000 1203 -988
rect 1275 988 1321 1000
rect 1275 -988 1281 988
rect 1315 -988 1321 988
rect 1275 -1000 1321 -988
rect 1393 988 1439 1000
rect 1393 -988 1399 988
rect 1433 -988 1439 988
rect 1393 -1000 1439 -988
rect 1511 988 1557 1000
rect 1511 -988 1517 988
rect 1551 -988 1557 988
rect 1511 -1000 1557 -988
rect 1629 988 1675 1000
rect 1629 -988 1635 988
rect 1669 -988 1675 988
rect 1629 -1000 1675 -988
rect 1747 988 1793 1000
rect 1747 -988 1753 988
rect 1787 -988 1793 988
rect 1747 -1000 1793 -988
rect 1865 988 1911 1000
rect 1865 -988 1871 988
rect 1905 -988 1911 988
rect 1865 -1000 1911 -988
rect 1983 988 2029 1000
rect 1983 -988 1989 988
rect 2023 -988 2029 988
rect 1983 -1000 2029 -988
rect 2101 988 2147 1000
rect 2101 -988 2107 988
rect 2141 -988 2147 988
rect 2101 -1000 2147 -988
rect 2219 988 2265 1000
rect 2219 -988 2225 988
rect 2259 -988 2265 988
rect 2219 -1000 2265 -988
rect 2337 988 2383 1000
rect 2337 -988 2343 988
rect 2377 -988 2383 988
rect 2337 -1000 2383 -988
rect 2455 988 2501 1000
rect 2455 -988 2461 988
rect 2495 -988 2501 988
rect 2455 -1000 2501 -988
rect 2573 988 2619 1000
rect 2573 -988 2579 988
rect 2613 -988 2619 988
rect 2573 -1000 2619 -988
rect 2691 988 2737 1000
rect 2691 -988 2697 988
rect 2731 -988 2737 988
rect 2691 -1000 2737 -988
rect -2684 -1047 -2626 -1041
rect -2684 -1081 -2672 -1047
rect -2638 -1081 -2626 -1047
rect -2684 -1087 -2626 -1081
rect -2566 -1047 -2508 -1041
rect -2566 -1081 -2554 -1047
rect -2520 -1081 -2508 -1047
rect -2566 -1087 -2508 -1081
rect -2448 -1047 -2390 -1041
rect -2448 -1081 -2436 -1047
rect -2402 -1081 -2390 -1047
rect -2448 -1087 -2390 -1081
rect -2330 -1047 -2272 -1041
rect -2330 -1081 -2318 -1047
rect -2284 -1081 -2272 -1047
rect -2330 -1087 -2272 -1081
rect -2212 -1047 -2154 -1041
rect -2212 -1081 -2200 -1047
rect -2166 -1081 -2154 -1047
rect -2212 -1087 -2154 -1081
rect -2094 -1047 -2036 -1041
rect -2094 -1081 -2082 -1047
rect -2048 -1081 -2036 -1047
rect -2094 -1087 -2036 -1081
rect -1976 -1047 -1918 -1041
rect -1976 -1081 -1964 -1047
rect -1930 -1081 -1918 -1047
rect -1976 -1087 -1918 -1081
rect -1858 -1047 -1800 -1041
rect -1858 -1081 -1846 -1047
rect -1812 -1081 -1800 -1047
rect -1858 -1087 -1800 -1081
rect -1740 -1047 -1682 -1041
rect -1740 -1081 -1728 -1047
rect -1694 -1081 -1682 -1047
rect -1740 -1087 -1682 -1081
rect -1622 -1047 -1564 -1041
rect -1622 -1081 -1610 -1047
rect -1576 -1081 -1564 -1047
rect -1622 -1087 -1564 -1081
rect -1504 -1047 -1446 -1041
rect -1504 -1081 -1492 -1047
rect -1458 -1081 -1446 -1047
rect -1504 -1087 -1446 -1081
rect -1386 -1047 -1328 -1041
rect -1386 -1081 -1374 -1047
rect -1340 -1081 -1328 -1047
rect -1386 -1087 -1328 -1081
rect -1268 -1047 -1210 -1041
rect -1268 -1081 -1256 -1047
rect -1222 -1081 -1210 -1047
rect -1268 -1087 -1210 -1081
rect -1150 -1047 -1092 -1041
rect -1150 -1081 -1138 -1047
rect -1104 -1081 -1092 -1047
rect -1150 -1087 -1092 -1081
rect -1032 -1047 -974 -1041
rect -1032 -1081 -1020 -1047
rect -986 -1081 -974 -1047
rect -1032 -1087 -974 -1081
rect -914 -1047 -856 -1041
rect -914 -1081 -902 -1047
rect -868 -1081 -856 -1047
rect -914 -1087 -856 -1081
rect -796 -1047 -738 -1041
rect -796 -1081 -784 -1047
rect -750 -1081 -738 -1047
rect -796 -1087 -738 -1081
rect -678 -1047 -620 -1041
rect -678 -1081 -666 -1047
rect -632 -1081 -620 -1047
rect -678 -1087 -620 -1081
rect -560 -1047 -502 -1041
rect -560 -1081 -548 -1047
rect -514 -1081 -502 -1047
rect -560 -1087 -502 -1081
rect -442 -1047 -384 -1041
rect -442 -1081 -430 -1047
rect -396 -1081 -384 -1047
rect -442 -1087 -384 -1081
rect -324 -1047 -266 -1041
rect -324 -1081 -312 -1047
rect -278 -1081 -266 -1047
rect -324 -1087 -266 -1081
rect -206 -1047 -148 -1041
rect -206 -1081 -194 -1047
rect -160 -1081 -148 -1047
rect -206 -1087 -148 -1081
rect -88 -1047 -30 -1041
rect -88 -1081 -76 -1047
rect -42 -1081 -30 -1047
rect -88 -1087 -30 -1081
rect 30 -1047 88 -1041
rect 30 -1081 42 -1047
rect 76 -1081 88 -1047
rect 30 -1087 88 -1081
rect 148 -1047 206 -1041
rect 148 -1081 160 -1047
rect 194 -1081 206 -1047
rect 148 -1087 206 -1081
rect 266 -1047 324 -1041
rect 266 -1081 278 -1047
rect 312 -1081 324 -1047
rect 266 -1087 324 -1081
rect 384 -1047 442 -1041
rect 384 -1081 396 -1047
rect 430 -1081 442 -1047
rect 384 -1087 442 -1081
rect 502 -1047 560 -1041
rect 502 -1081 514 -1047
rect 548 -1081 560 -1047
rect 502 -1087 560 -1081
rect 620 -1047 678 -1041
rect 620 -1081 632 -1047
rect 666 -1081 678 -1047
rect 620 -1087 678 -1081
rect 738 -1047 796 -1041
rect 738 -1081 750 -1047
rect 784 -1081 796 -1047
rect 738 -1087 796 -1081
rect 856 -1047 914 -1041
rect 856 -1081 868 -1047
rect 902 -1081 914 -1047
rect 856 -1087 914 -1081
rect 974 -1047 1032 -1041
rect 974 -1081 986 -1047
rect 1020 -1081 1032 -1047
rect 974 -1087 1032 -1081
rect 1092 -1047 1150 -1041
rect 1092 -1081 1104 -1047
rect 1138 -1081 1150 -1047
rect 1092 -1087 1150 -1081
rect 1210 -1047 1268 -1041
rect 1210 -1081 1222 -1047
rect 1256 -1081 1268 -1047
rect 1210 -1087 1268 -1081
rect 1328 -1047 1386 -1041
rect 1328 -1081 1340 -1047
rect 1374 -1081 1386 -1047
rect 1328 -1087 1386 -1081
rect 1446 -1047 1504 -1041
rect 1446 -1081 1458 -1047
rect 1492 -1081 1504 -1047
rect 1446 -1087 1504 -1081
rect 1564 -1047 1622 -1041
rect 1564 -1081 1576 -1047
rect 1610 -1081 1622 -1047
rect 1564 -1087 1622 -1081
rect 1682 -1047 1740 -1041
rect 1682 -1081 1694 -1047
rect 1728 -1081 1740 -1047
rect 1682 -1087 1740 -1081
rect 1800 -1047 1858 -1041
rect 1800 -1081 1812 -1047
rect 1846 -1081 1858 -1047
rect 1800 -1087 1858 -1081
rect 1918 -1047 1976 -1041
rect 1918 -1081 1930 -1047
rect 1964 -1081 1976 -1047
rect 1918 -1087 1976 -1081
rect 2036 -1047 2094 -1041
rect 2036 -1081 2048 -1047
rect 2082 -1081 2094 -1047
rect 2036 -1087 2094 -1081
rect 2154 -1047 2212 -1041
rect 2154 -1081 2166 -1047
rect 2200 -1081 2212 -1047
rect 2154 -1087 2212 -1081
rect 2272 -1047 2330 -1041
rect 2272 -1081 2284 -1047
rect 2318 -1081 2330 -1047
rect 2272 -1087 2330 -1081
rect 2390 -1047 2448 -1041
rect 2390 -1081 2402 -1047
rect 2436 -1081 2448 -1047
rect 2390 -1087 2448 -1081
rect 2508 -1047 2566 -1041
rect 2508 -1081 2520 -1047
rect 2554 -1081 2566 -1047
rect 2508 -1087 2566 -1081
rect 2626 -1047 2684 -1041
rect 2626 -1081 2638 -1047
rect 2672 -1081 2684 -1047
rect 2626 -1087 2684 -1081
<< properties >>
string FIXED_BBOX -2828 -1166 2828 1166
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 10 l 0.3 m 1 nf 46 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
