magic
tech sky130A
magscale 1 2
timestamp 1671678338
<< pwell >>
rect -284 -748 284 748
<< psubdiff >>
rect -248 678 -152 712
rect 152 678 248 712
rect -248 616 -214 678
rect 214 616 248 678
rect -248 -678 -214 -616
rect 214 -678 248 -616
rect -248 -712 -152 -678
rect 152 -712 248 -678
<< psubdiffcont >>
rect -152 678 152 712
rect -248 -616 -214 616
rect 214 -616 248 616
rect -152 -712 152 -678
<< xpolycontact >>
rect -118 150 -48 582
rect -118 -582 -48 -150
rect 48 150 118 582
rect 48 -582 118 -150
<< xpolyres >>
rect -118 -150 -48 150
rect 48 -150 118 150
<< locali >>
rect -248 678 -152 712
rect 152 678 248 712
rect -248 616 -214 678
rect 214 616 248 678
rect -248 -678 -214 -616
rect 214 -678 248 -616
rect -248 -712 -152 -678
rect 152 -712 248 -678
<< viali >>
rect -102 167 -64 564
rect 64 167 102 564
rect -102 -564 -64 -167
rect 64 -564 102 -167
<< metal1 >>
rect -108 564 -58 576
rect -108 167 -102 564
rect -64 167 -58 564
rect -108 155 -58 167
rect 58 564 108 576
rect 58 167 64 564
rect 102 167 108 564
rect 58 155 108 167
rect -108 -167 -58 -155
rect -108 -564 -102 -167
rect -64 -564 -58 -167
rect -108 -576 -58 -564
rect 58 -167 108 -155
rect 58 -564 64 -167
rect 102 -564 108 -167
rect 58 -576 108 -564
<< res0p35 >>
rect -120 -152 -46 152
rect 46 -152 120 152
<< properties >>
string FIXED_BBOX -231 -695 231 695
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 1.5 m 1 nx 2 wmin 0.350 lmin 0.50 rho 2000 val 9.646k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
