magic
tech sky130A
magscale 1 2
timestamp 1671152619
<< error_p >>
rect -269 572 -211 578
rect -77 572 -19 578
rect 115 572 173 578
rect 307 572 365 578
rect -269 538 -257 572
rect -77 538 -65 572
rect 115 538 127 572
rect 307 538 319 572
rect -269 532 -211 538
rect -77 532 -19 538
rect 115 532 173 538
rect 307 532 365 538
rect -365 -538 -307 -532
rect -173 -538 -115 -532
rect 19 -538 77 -532
rect 211 -538 269 -532
rect -365 -572 -353 -538
rect -173 -572 -161 -538
rect 19 -572 31 -538
rect 211 -572 223 -538
rect -365 -578 -307 -572
rect -173 -578 -115 -572
rect 19 -578 77 -572
rect 211 -578 269 -572
<< pwell >>
rect -551 -710 551 710
<< nmos >>
rect -351 -500 -321 500
rect -255 -500 -225 500
rect -159 -500 -129 500
rect -63 -500 -33 500
rect 33 -500 63 500
rect 129 -500 159 500
rect 225 -500 255 500
rect 321 -500 351 500
<< ndiff >>
rect -413 488 -351 500
rect -413 -488 -401 488
rect -367 -488 -351 488
rect -413 -500 -351 -488
rect -321 488 -255 500
rect -321 -488 -305 488
rect -271 -488 -255 488
rect -321 -500 -255 -488
rect -225 488 -159 500
rect -225 -488 -209 488
rect -175 -488 -159 488
rect -225 -500 -159 -488
rect -129 488 -63 500
rect -129 -488 -113 488
rect -79 -488 -63 488
rect -129 -500 -63 -488
rect -33 488 33 500
rect -33 -488 -17 488
rect 17 -488 33 488
rect -33 -500 33 -488
rect 63 488 129 500
rect 63 -488 79 488
rect 113 -488 129 488
rect 63 -500 129 -488
rect 159 488 225 500
rect 159 -488 175 488
rect 209 -488 225 488
rect 159 -500 225 -488
rect 255 488 321 500
rect 255 -488 271 488
rect 305 -488 321 488
rect 255 -500 321 -488
rect 351 488 413 500
rect 351 -488 367 488
rect 401 -488 413 488
rect 351 -500 413 -488
<< ndiffc >>
rect -401 -488 -367 488
rect -305 -488 -271 488
rect -209 -488 -175 488
rect -113 -488 -79 488
rect -17 -488 17 488
rect 79 -488 113 488
rect 175 -488 209 488
rect 271 -488 305 488
rect 367 -488 401 488
<< psubdiff >>
rect -515 640 -419 674
rect 419 640 515 674
rect -515 578 -481 640
rect 481 578 515 640
rect -515 -640 -481 -578
rect 481 -640 515 -578
rect -515 -674 -419 -640
rect 419 -674 515 -640
<< psubdiffcont >>
rect -419 640 419 674
rect -515 -578 -481 578
rect 481 -578 515 578
rect -419 -674 419 -640
<< poly >>
rect -273 572 -207 588
rect -273 538 -257 572
rect -223 538 -207 572
rect -351 500 -321 526
rect -273 522 -207 538
rect -81 572 -15 588
rect -81 538 -65 572
rect -31 538 -15 572
rect -255 500 -225 522
rect -159 500 -129 526
rect -81 522 -15 538
rect 111 572 177 588
rect 111 538 127 572
rect 161 538 177 572
rect -63 500 -33 522
rect 33 500 63 526
rect 111 522 177 538
rect 303 572 369 588
rect 303 538 319 572
rect 353 538 369 572
rect 129 500 159 522
rect 225 500 255 526
rect 303 522 369 538
rect 321 500 351 522
rect -351 -522 -321 -500
rect -369 -538 -303 -522
rect -255 -526 -225 -500
rect -159 -522 -129 -500
rect -369 -572 -353 -538
rect -319 -572 -303 -538
rect -369 -588 -303 -572
rect -177 -538 -111 -522
rect -63 -526 -33 -500
rect 33 -522 63 -500
rect -177 -572 -161 -538
rect -127 -572 -111 -538
rect -177 -588 -111 -572
rect 15 -538 81 -522
rect 129 -526 159 -500
rect 225 -522 255 -500
rect 15 -572 31 -538
rect 65 -572 81 -538
rect 15 -588 81 -572
rect 207 -538 273 -522
rect 321 -526 351 -500
rect 207 -572 223 -538
rect 257 -572 273 -538
rect 207 -588 273 -572
<< polycont >>
rect -257 538 -223 572
rect -65 538 -31 572
rect 127 538 161 572
rect 319 538 353 572
rect -353 -572 -319 -538
rect -161 -572 -127 -538
rect 31 -572 65 -538
rect 223 -572 257 -538
<< locali >>
rect -515 640 -419 674
rect 419 640 515 674
rect -515 578 -481 640
rect 481 578 515 640
rect -273 538 -257 572
rect -223 538 -207 572
rect -81 538 -65 572
rect -31 538 -15 572
rect 111 538 127 572
rect 161 538 177 572
rect 303 538 319 572
rect 353 538 369 572
rect -401 488 -367 504
rect -401 -504 -367 -488
rect -305 488 -271 504
rect -305 -504 -271 -488
rect -209 488 -175 504
rect -209 -504 -175 -488
rect -113 488 -79 504
rect -113 -504 -79 -488
rect -17 488 17 504
rect -17 -504 17 -488
rect 79 488 113 504
rect 79 -504 113 -488
rect 175 488 209 504
rect 175 -504 209 -488
rect 271 488 305 504
rect 271 -504 305 -488
rect 367 488 401 504
rect 367 -504 401 -488
rect -369 -572 -353 -538
rect -319 -572 -303 -538
rect -177 -572 -161 -538
rect -127 -572 -111 -538
rect 15 -572 31 -538
rect 65 -572 81 -538
rect 207 -572 223 -538
rect 257 -572 273 -538
rect -515 -640 -481 -578
rect 481 -640 515 -578
rect -515 -674 -419 -640
rect 419 -674 515 -640
<< viali >>
rect -257 538 -223 572
rect -65 538 -31 572
rect 127 538 161 572
rect 319 538 353 572
rect -401 -488 -367 488
rect -305 -488 -271 488
rect -209 -488 -175 488
rect -113 -488 -79 488
rect -17 -488 17 488
rect 79 -488 113 488
rect 175 -488 209 488
rect 271 -488 305 488
rect 367 -488 401 488
rect -353 -572 -319 -538
rect -161 -572 -127 -538
rect 31 -572 65 -538
rect 223 -572 257 -538
<< metal1 >>
rect -269 572 -211 578
rect -269 538 -257 572
rect -223 538 -211 572
rect -269 532 -211 538
rect -77 572 -19 578
rect -77 538 -65 572
rect -31 538 -19 572
rect -77 532 -19 538
rect 115 572 173 578
rect 115 538 127 572
rect 161 538 173 572
rect 115 532 173 538
rect 307 572 365 578
rect 307 538 319 572
rect 353 538 365 572
rect 307 532 365 538
rect -407 488 -361 500
rect -407 -488 -401 488
rect -367 -488 -361 488
rect -407 -500 -361 -488
rect -311 488 -265 500
rect -311 -488 -305 488
rect -271 -488 -265 488
rect -311 -500 -265 -488
rect -215 488 -169 500
rect -215 -488 -209 488
rect -175 -488 -169 488
rect -215 -500 -169 -488
rect -119 488 -73 500
rect -119 -488 -113 488
rect -79 -488 -73 488
rect -119 -500 -73 -488
rect -23 488 23 500
rect -23 -488 -17 488
rect 17 -488 23 488
rect -23 -500 23 -488
rect 73 488 119 500
rect 73 -488 79 488
rect 113 -488 119 488
rect 73 -500 119 -488
rect 169 488 215 500
rect 169 -488 175 488
rect 209 -488 215 488
rect 169 -500 215 -488
rect 265 488 311 500
rect 265 -488 271 488
rect 305 -488 311 488
rect 265 -500 311 -488
rect 361 488 407 500
rect 361 -488 367 488
rect 401 -488 407 488
rect 361 -500 407 -488
rect -365 -538 -307 -532
rect -365 -572 -353 -538
rect -319 -572 -307 -538
rect -365 -578 -307 -572
rect -173 -538 -115 -532
rect -173 -572 -161 -538
rect -127 -572 -115 -538
rect -173 -578 -115 -572
rect 19 -538 77 -532
rect 19 -572 31 -538
rect 65 -572 77 -538
rect 19 -578 77 -572
rect 211 -538 269 -532
rect 211 -572 223 -538
rect 257 -572 269 -538
rect 211 -578 269 -572
<< properties >>
string FIXED_BBOX -498 -657 498 657
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 5 l 0.15 m 1 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
