magic
tech sky130A
magscale 1 2
timestamp 1671856655
<< nwell >>
rect 17947 -5634 22057 -3196
rect 23118 -7653 23838 -7332
rect 16790 -10900 17111 -10456
<< pwell >>
rect 17710 -8134 18752 -5714
rect 18875 -6810 21129 -5890
rect 21251 -6082 22293 -5714
rect 16440 -8714 17360 -8248
rect 16440 -8718 17198 -8714
rect 17244 -8718 17360 -8714
rect 16440 -9034 17360 -8718
rect 16440 -9140 17272 -9034
rect 17281 -9140 17360 -9034
rect 16440 -9382 17360 -9140
rect 18919 -9250 21085 -6830
rect 21251 -7450 22996 -6082
rect 21251 -8134 22293 -7450
rect 23159 -7876 23245 -7719
rect 23253 -7901 23431 -7711
rect 23435 -7876 23521 -7719
rect 23529 -7901 23707 -7711
rect 23711 -7876 23797 -7719
rect 23277 -7931 23311 -7901
rect 23553 -7931 23587 -7901
rect 17177 -10583 17334 -10497
rect 17169 -10615 17359 -10591
rect 17169 -10649 17389 -10615
rect 17169 -10769 17359 -10649
rect 17177 -10859 17334 -10773
<< nmos >>
rect 17906 -7924 17966 -5924
rect 18024 -7924 18084 -5924
rect 18142 -7924 18202 -5924
rect 18260 -7924 18320 -5924
rect 18378 -7924 18438 -5924
rect 18496 -7924 18556 -5924
rect 16650 -8478 17150 -8448
rect 16650 -8574 17150 -8544
rect 16650 -8670 17150 -8640
rect 16650 -8766 17150 -8736
rect 19115 -9040 19515 -7040
rect 19573 -9040 19973 -7040
rect 20031 -9040 20431 -7040
rect 20489 -9040 20889 -7040
rect 21447 -7924 21507 -5924
rect 21565 -7924 21625 -5924
rect 21683 -7924 21743 -5924
rect 21801 -7924 21861 -5924
rect 21919 -7924 21979 -5924
rect 22037 -7924 22097 -5924
<< pmos >>
rect 18143 -5415 18203 -3415
rect 18261 -5415 18321 -3415
rect 18379 -5415 18439 -3415
rect 18497 -5415 18557 -3415
rect 18615 -5415 18675 -3415
rect 18733 -5415 18793 -3415
rect 18851 -5415 18911 -3415
rect 18969 -5415 19029 -3415
rect 19087 -5415 19147 -3415
rect 19205 -5415 19265 -3415
rect 19323 -5415 19383 -3415
rect 19441 -5415 19501 -3415
rect 19559 -5415 19619 -3415
rect 19677 -5415 19737 -3415
rect 19795 -5415 19855 -3415
rect 19913 -5415 19973 -3415
rect 20031 -5415 20091 -3415
rect 20149 -5415 20209 -3415
rect 20267 -5415 20327 -3415
rect 20385 -5415 20445 -3415
rect 20503 -5415 20563 -3415
rect 20621 -5415 20681 -3415
rect 20739 -5415 20799 -3415
rect 20857 -5415 20917 -3415
rect 20975 -5415 21035 -3415
rect 21093 -5415 21153 -3415
rect 21211 -5415 21271 -3415
rect 21329 -5415 21389 -3415
rect 21447 -5415 21507 -3415
rect 21565 -5415 21625 -3415
rect 21683 -5415 21743 -3415
rect 21801 -5415 21861 -3415
<< nmoslvt >>
rect 19075 -6600 19105 -6100
rect 19171 -6600 19201 -6100
rect 19267 -6600 19297 -6100
rect 19363 -6600 19393 -6100
rect 19459 -6600 19489 -6100
rect 19555 -6600 19585 -6100
rect 19651 -6600 19681 -6100
rect 19747 -6600 19777 -6100
rect 19843 -6600 19873 -6100
rect 19939 -6600 19969 -6100
rect 20035 -6600 20065 -6100
rect 20131 -6600 20161 -6100
rect 20227 -6600 20257 -6100
rect 20323 -6600 20353 -6100
rect 20419 -6600 20449 -6100
rect 20515 -6600 20545 -6100
rect 20611 -6600 20641 -6100
rect 20707 -6600 20737 -6100
rect 20803 -6600 20833 -6100
rect 20899 -6600 20929 -6100
<< ndiff >>
rect 17848 -5936 17906 -5924
rect 17848 -7912 17860 -5936
rect 17894 -7912 17906 -5936
rect 17848 -7924 17906 -7912
rect 17966 -5936 18024 -5924
rect 17966 -7912 17978 -5936
rect 18012 -7912 18024 -5936
rect 17966 -7924 18024 -7912
rect 18084 -5936 18142 -5924
rect 18084 -7912 18096 -5936
rect 18130 -7912 18142 -5936
rect 18084 -7924 18142 -7912
rect 18202 -5936 18260 -5924
rect 18202 -7912 18214 -5936
rect 18248 -7912 18260 -5936
rect 18202 -7924 18260 -7912
rect 18320 -5936 18378 -5924
rect 18320 -7912 18332 -5936
rect 18366 -7912 18378 -5936
rect 18320 -7924 18378 -7912
rect 18438 -5936 18496 -5924
rect 18438 -7912 18450 -5936
rect 18484 -7912 18496 -5936
rect 18438 -7924 18496 -7912
rect 18556 -5936 18614 -5924
rect 18556 -7912 18568 -5936
rect 18602 -7912 18614 -5936
rect 18556 -7924 18614 -7912
rect 19013 -6112 19075 -6100
rect 19013 -6588 19025 -6112
rect 19059 -6588 19075 -6112
rect 19013 -6600 19075 -6588
rect 19105 -6112 19171 -6100
rect 19105 -6588 19121 -6112
rect 19155 -6588 19171 -6112
rect 19105 -6600 19171 -6588
rect 19201 -6112 19267 -6100
rect 19201 -6588 19217 -6112
rect 19251 -6588 19267 -6112
rect 19201 -6600 19267 -6588
rect 19297 -6112 19363 -6100
rect 19297 -6588 19313 -6112
rect 19347 -6588 19363 -6112
rect 19297 -6600 19363 -6588
rect 19393 -6112 19459 -6100
rect 19393 -6588 19409 -6112
rect 19443 -6588 19459 -6112
rect 19393 -6600 19459 -6588
rect 19489 -6112 19555 -6100
rect 19489 -6588 19505 -6112
rect 19539 -6588 19555 -6112
rect 19489 -6600 19555 -6588
rect 19585 -6112 19651 -6100
rect 19585 -6588 19601 -6112
rect 19635 -6588 19651 -6112
rect 19585 -6600 19651 -6588
rect 19681 -6112 19747 -6100
rect 19681 -6588 19697 -6112
rect 19731 -6588 19747 -6112
rect 19681 -6600 19747 -6588
rect 19777 -6112 19843 -6100
rect 19777 -6588 19793 -6112
rect 19827 -6588 19843 -6112
rect 19777 -6600 19843 -6588
rect 19873 -6112 19939 -6100
rect 19873 -6588 19889 -6112
rect 19923 -6588 19939 -6112
rect 19873 -6600 19939 -6588
rect 19969 -6112 20035 -6100
rect 19969 -6588 19985 -6112
rect 20019 -6588 20035 -6112
rect 19969 -6600 20035 -6588
rect 20065 -6112 20131 -6100
rect 20065 -6588 20081 -6112
rect 20115 -6588 20131 -6112
rect 20065 -6600 20131 -6588
rect 20161 -6112 20227 -6100
rect 20161 -6588 20177 -6112
rect 20211 -6588 20227 -6112
rect 20161 -6600 20227 -6588
rect 20257 -6112 20323 -6100
rect 20257 -6588 20273 -6112
rect 20307 -6588 20323 -6112
rect 20257 -6600 20323 -6588
rect 20353 -6112 20419 -6100
rect 20353 -6588 20369 -6112
rect 20403 -6588 20419 -6112
rect 20353 -6600 20419 -6588
rect 20449 -6112 20515 -6100
rect 20449 -6588 20465 -6112
rect 20499 -6588 20515 -6112
rect 20449 -6600 20515 -6588
rect 20545 -6112 20611 -6100
rect 20545 -6588 20561 -6112
rect 20595 -6588 20611 -6112
rect 20545 -6600 20611 -6588
rect 20641 -6112 20707 -6100
rect 20641 -6588 20657 -6112
rect 20691 -6588 20707 -6112
rect 20641 -6600 20707 -6588
rect 20737 -6112 20803 -6100
rect 20737 -6588 20753 -6112
rect 20787 -6588 20803 -6112
rect 20737 -6600 20803 -6588
rect 20833 -6112 20899 -6100
rect 20833 -6588 20849 -6112
rect 20883 -6588 20899 -6112
rect 20833 -6600 20899 -6588
rect 20929 -6112 20991 -6100
rect 20929 -6588 20945 -6112
rect 20979 -6588 20991 -6112
rect 20929 -6600 20991 -6588
rect 16650 -8398 17150 -8386
rect 16650 -8432 16662 -8398
rect 17138 -8432 17150 -8398
rect 16650 -8448 17150 -8432
rect 16650 -8494 17150 -8478
rect 16650 -8528 16662 -8494
rect 17138 -8528 17150 -8494
rect 16650 -8544 17150 -8528
rect 16650 -8590 17150 -8574
rect 16650 -8624 16662 -8590
rect 17138 -8624 17150 -8590
rect 16650 -8640 17150 -8624
rect 16650 -8686 17150 -8670
rect 16650 -8720 16662 -8686
rect 17138 -8720 17150 -8686
rect 16650 -8736 17150 -8720
rect 16650 -8782 17150 -8766
rect 16650 -8816 16662 -8782
rect 17138 -8816 17150 -8782
rect 16650 -8828 17150 -8816
rect 19057 -7052 19115 -7040
rect 19057 -9028 19069 -7052
rect 19103 -9028 19115 -7052
rect 19057 -9040 19115 -9028
rect 19515 -7052 19573 -7040
rect 19515 -9028 19527 -7052
rect 19561 -9028 19573 -7052
rect 19515 -9040 19573 -9028
rect 19973 -7052 20031 -7040
rect 19973 -9028 19985 -7052
rect 20019 -9028 20031 -7052
rect 19973 -9040 20031 -9028
rect 20431 -7052 20489 -7040
rect 20431 -9028 20443 -7052
rect 20477 -9028 20489 -7052
rect 20431 -9040 20489 -9028
rect 20889 -7052 20947 -7040
rect 20889 -9028 20901 -7052
rect 20935 -9028 20947 -7052
rect 20889 -9040 20947 -9028
rect 21389 -5936 21447 -5924
rect 21389 -7912 21401 -5936
rect 21435 -7912 21447 -5936
rect 21389 -7924 21447 -7912
rect 21507 -5936 21565 -5924
rect 21507 -7912 21519 -5936
rect 21553 -7912 21565 -5936
rect 21507 -7924 21565 -7912
rect 21625 -5936 21683 -5924
rect 21625 -7912 21637 -5936
rect 21671 -7912 21683 -5936
rect 21625 -7924 21683 -7912
rect 21743 -5936 21801 -5924
rect 21743 -7912 21755 -5936
rect 21789 -7912 21801 -5936
rect 21743 -7924 21801 -7912
rect 21861 -5936 21919 -5924
rect 21861 -7912 21873 -5936
rect 21907 -7912 21919 -5936
rect 21861 -7924 21919 -7912
rect 21979 -5936 22037 -5924
rect 21979 -7912 21991 -5936
rect 22025 -7912 22037 -5936
rect 21979 -7924 22037 -7912
rect 22097 -5936 22155 -5924
rect 22097 -7912 22109 -5936
rect 22143 -7912 22155 -5936
rect 22097 -7924 22155 -7912
<< pdiff >>
rect 18085 -3427 18143 -3415
rect 18085 -5403 18097 -3427
rect 18131 -5403 18143 -3427
rect 18085 -5415 18143 -5403
rect 18203 -3427 18261 -3415
rect 18203 -5403 18215 -3427
rect 18249 -5403 18261 -3427
rect 18203 -5415 18261 -5403
rect 18321 -3427 18379 -3415
rect 18321 -5403 18333 -3427
rect 18367 -5403 18379 -3427
rect 18321 -5415 18379 -5403
rect 18439 -3427 18497 -3415
rect 18439 -5403 18451 -3427
rect 18485 -5403 18497 -3427
rect 18439 -5415 18497 -5403
rect 18557 -3427 18615 -3415
rect 18557 -5403 18569 -3427
rect 18603 -5403 18615 -3427
rect 18557 -5415 18615 -5403
rect 18675 -3427 18733 -3415
rect 18675 -5403 18687 -3427
rect 18721 -5403 18733 -3427
rect 18675 -5415 18733 -5403
rect 18793 -3427 18851 -3415
rect 18793 -5403 18805 -3427
rect 18839 -5403 18851 -3427
rect 18793 -5415 18851 -5403
rect 18911 -3427 18969 -3415
rect 18911 -5403 18923 -3427
rect 18957 -5403 18969 -3427
rect 18911 -5415 18969 -5403
rect 19029 -3427 19087 -3415
rect 19029 -5403 19041 -3427
rect 19075 -5403 19087 -3427
rect 19029 -5415 19087 -5403
rect 19147 -3427 19205 -3415
rect 19147 -5403 19159 -3427
rect 19193 -5403 19205 -3427
rect 19147 -5415 19205 -5403
rect 19265 -3427 19323 -3415
rect 19265 -5403 19277 -3427
rect 19311 -5403 19323 -3427
rect 19265 -5415 19323 -5403
rect 19383 -3427 19441 -3415
rect 19383 -5403 19395 -3427
rect 19429 -5403 19441 -3427
rect 19383 -5415 19441 -5403
rect 19501 -3427 19559 -3415
rect 19501 -5403 19513 -3427
rect 19547 -5403 19559 -3427
rect 19501 -5415 19559 -5403
rect 19619 -3427 19677 -3415
rect 19619 -5403 19631 -3427
rect 19665 -5403 19677 -3427
rect 19619 -5415 19677 -5403
rect 19737 -3427 19795 -3415
rect 19737 -5403 19749 -3427
rect 19783 -5403 19795 -3427
rect 19737 -5415 19795 -5403
rect 19855 -3427 19913 -3415
rect 19855 -5403 19867 -3427
rect 19901 -5403 19913 -3427
rect 19855 -5415 19913 -5403
rect 19973 -3427 20031 -3415
rect 19973 -5403 19985 -3427
rect 20019 -5403 20031 -3427
rect 19973 -5415 20031 -5403
rect 20091 -3427 20149 -3415
rect 20091 -5403 20103 -3427
rect 20137 -5403 20149 -3427
rect 20091 -5415 20149 -5403
rect 20209 -3427 20267 -3415
rect 20209 -5403 20221 -3427
rect 20255 -5403 20267 -3427
rect 20209 -5415 20267 -5403
rect 20327 -3427 20385 -3415
rect 20327 -5403 20339 -3427
rect 20373 -5403 20385 -3427
rect 20327 -5415 20385 -5403
rect 20445 -3427 20503 -3415
rect 20445 -5403 20457 -3427
rect 20491 -5403 20503 -3427
rect 20445 -5415 20503 -5403
rect 20563 -3427 20621 -3415
rect 20563 -5403 20575 -3427
rect 20609 -5403 20621 -3427
rect 20563 -5415 20621 -5403
rect 20681 -3427 20739 -3415
rect 20681 -5403 20693 -3427
rect 20727 -5403 20739 -3427
rect 20681 -5415 20739 -5403
rect 20799 -3427 20857 -3415
rect 20799 -5403 20811 -3427
rect 20845 -5403 20857 -3427
rect 20799 -5415 20857 -5403
rect 20917 -3427 20975 -3415
rect 20917 -5403 20929 -3427
rect 20963 -5403 20975 -3427
rect 20917 -5415 20975 -5403
rect 21035 -3427 21093 -3415
rect 21035 -5403 21047 -3427
rect 21081 -5403 21093 -3427
rect 21035 -5415 21093 -5403
rect 21153 -3427 21211 -3415
rect 21153 -5403 21165 -3427
rect 21199 -5403 21211 -3427
rect 21153 -5415 21211 -5403
rect 21271 -3427 21329 -3415
rect 21271 -5403 21283 -3427
rect 21317 -5403 21329 -3427
rect 21271 -5415 21329 -5403
rect 21389 -3427 21447 -3415
rect 21389 -5403 21401 -3427
rect 21435 -5403 21447 -3427
rect 21389 -5415 21447 -5403
rect 21507 -3427 21565 -3415
rect 21507 -5403 21519 -3427
rect 21553 -5403 21565 -3427
rect 21507 -5415 21565 -5403
rect 21625 -3427 21683 -3415
rect 21625 -5403 21637 -3427
rect 21671 -5403 21683 -3427
rect 21625 -5415 21683 -5403
rect 21743 -3427 21801 -3415
rect 21743 -5403 21755 -3427
rect 21789 -5403 21801 -3427
rect 21743 -5415 21801 -5403
rect 21861 -3427 21919 -3415
rect 21861 -5403 21873 -3427
rect 21907 -5403 21919 -3427
rect 21861 -5415 21919 -5403
<< ndiffc >>
rect 17860 -7912 17894 -5936
rect 17978 -7912 18012 -5936
rect 18096 -7912 18130 -5936
rect 18214 -7912 18248 -5936
rect 18332 -7912 18366 -5936
rect 18450 -7912 18484 -5936
rect 18568 -7912 18602 -5936
rect 19025 -6588 19059 -6112
rect 19121 -6588 19155 -6112
rect 19217 -6588 19251 -6112
rect 19313 -6588 19347 -6112
rect 19409 -6588 19443 -6112
rect 19505 -6588 19539 -6112
rect 19601 -6588 19635 -6112
rect 19697 -6588 19731 -6112
rect 19793 -6588 19827 -6112
rect 19889 -6588 19923 -6112
rect 19985 -6588 20019 -6112
rect 20081 -6588 20115 -6112
rect 20177 -6588 20211 -6112
rect 20273 -6588 20307 -6112
rect 20369 -6588 20403 -6112
rect 20465 -6588 20499 -6112
rect 20561 -6588 20595 -6112
rect 20657 -6588 20691 -6112
rect 20753 -6588 20787 -6112
rect 20849 -6588 20883 -6112
rect 20945 -6588 20979 -6112
rect 16662 -8432 17138 -8398
rect 16662 -8528 17138 -8494
rect 16662 -8624 17138 -8590
rect 16662 -8720 17138 -8686
rect 16662 -8816 17138 -8782
rect 19069 -9028 19103 -7052
rect 19527 -9028 19561 -7052
rect 19985 -9028 20019 -7052
rect 20443 -9028 20477 -7052
rect 20901 -9028 20935 -7052
rect 21401 -7912 21435 -5936
rect 21519 -7912 21553 -5936
rect 21637 -7912 21671 -5936
rect 21755 -7912 21789 -5936
rect 21873 -7912 21907 -5936
rect 21991 -7912 22025 -5936
rect 22109 -7912 22143 -5936
<< pdiffc >>
rect 18097 -5403 18131 -3427
rect 18215 -5403 18249 -3427
rect 18333 -5403 18367 -3427
rect 18451 -5403 18485 -3427
rect 18569 -5403 18603 -3427
rect 18687 -5403 18721 -3427
rect 18805 -5403 18839 -3427
rect 18923 -5403 18957 -3427
rect 19041 -5403 19075 -3427
rect 19159 -5403 19193 -3427
rect 19277 -5403 19311 -3427
rect 19395 -5403 19429 -3427
rect 19513 -5403 19547 -3427
rect 19631 -5403 19665 -3427
rect 19749 -5403 19783 -3427
rect 19867 -5403 19901 -3427
rect 19985 -5403 20019 -3427
rect 20103 -5403 20137 -3427
rect 20221 -5403 20255 -3427
rect 20339 -5403 20373 -3427
rect 20457 -5403 20491 -3427
rect 20575 -5403 20609 -3427
rect 20693 -5403 20727 -3427
rect 20811 -5403 20845 -3427
rect 20929 -5403 20963 -3427
rect 21047 -5403 21081 -3427
rect 21165 -5403 21199 -3427
rect 21283 -5403 21317 -3427
rect 21401 -5403 21435 -3427
rect 21519 -5403 21553 -3427
rect 21637 -5403 21671 -3427
rect 21755 -5403 21789 -3427
rect 21873 -5403 21907 -3427
<< psubdiff >>
rect 17746 -5784 17842 -5750
rect 18620 -5784 18716 -5750
rect 17746 -5846 17780 -5784
rect 18682 -5846 18716 -5784
rect 17746 -8064 17780 -8002
rect 21287 -5784 21383 -5750
rect 22161 -5784 22257 -5750
rect 21287 -5846 21321 -5784
rect 18911 -5960 19007 -5926
rect 20997 -5960 21093 -5926
rect 18911 -6022 18945 -5960
rect 21059 -6022 21093 -5960
rect 18911 -6740 18945 -6678
rect 21059 -6740 21093 -6678
rect 18911 -6774 19007 -6740
rect 20997 -6774 21093 -6740
rect 18682 -8064 18716 -8002
rect 17746 -8098 17842 -8064
rect 18620 -8098 18716 -8064
rect 18955 -6900 19051 -6866
rect 20953 -6900 21049 -6866
rect 18955 -6962 18989 -6900
rect 16476 -8318 16572 -8284
rect 17228 -8318 17324 -8284
rect 16476 -8380 16510 -8318
rect 17290 -8380 17324 -8318
rect 16476 -9312 16510 -9230
rect 21015 -6962 21049 -6900
rect 18955 -9180 18989 -9118
rect 22223 -5846 22257 -5784
rect 21287 -8064 21321 -8002
rect 22328 -6152 22424 -6118
rect 22864 -6152 22960 -6118
rect 22328 -6214 22362 -6152
rect 22926 -6214 22960 -6152
rect 22328 -7380 22362 -7318
rect 22926 -7380 22960 -7318
rect 22328 -7414 22424 -7380
rect 22864 -7414 22960 -7380
rect 23185 -7769 23219 -7745
rect 23185 -7850 23219 -7803
rect 23461 -7769 23495 -7745
rect 23461 -7850 23495 -7803
rect 23737 -7769 23771 -7745
rect 23737 -7850 23771 -7803
rect 22223 -8064 22257 -8002
rect 21287 -8098 21383 -8064
rect 22161 -8098 22257 -8064
rect 21015 -9180 21049 -9118
rect 18955 -9214 19051 -9180
rect 20953 -9214 21049 -9180
rect 17290 -9312 17324 -9230
rect 16476 -9346 16572 -9312
rect 17228 -9346 17324 -9312
rect 17203 -10557 17227 -10523
rect 17261 -10557 17308 -10523
rect 17203 -10833 17227 -10799
rect 17261 -10833 17308 -10799
<< nsubdiff >>
rect 17983 -3266 18079 -3232
rect 21925 -3266 22021 -3232
rect 17983 -3328 18017 -3266
rect 21987 -3328 22021 -3266
rect 17983 -5564 18017 -5502
rect 21987 -5564 22021 -5502
rect 17983 -5598 18079 -5564
rect 21925 -5598 22021 -5564
rect 23185 -7458 23219 -7434
rect 23185 -7551 23219 -7492
rect 23185 -7609 23219 -7585
rect 23461 -7458 23495 -7434
rect 23461 -7551 23495 -7492
rect 23461 -7609 23495 -7585
rect 23737 -7458 23771 -7434
rect 23737 -7551 23771 -7492
rect 23737 -7609 23771 -7585
rect 16892 -10557 16916 -10523
rect 16950 -10557 17009 -10523
rect 17043 -10557 17067 -10523
rect 16892 -10833 16916 -10799
rect 16950 -10833 17009 -10799
rect 17043 -10833 17067 -10799
<< psubdiffcont >>
rect 17842 -5784 18620 -5750
rect 17746 -8002 17780 -5846
rect 18682 -8002 18716 -5846
rect 21383 -5784 22161 -5750
rect 19007 -5960 20997 -5926
rect 18911 -6678 18945 -6022
rect 21059 -6678 21093 -6022
rect 19007 -6774 20997 -6740
rect 17842 -8098 18620 -8064
rect 19051 -6900 20953 -6866
rect 16572 -8318 17228 -8284
rect 16476 -9230 16510 -8380
rect 17290 -9230 17324 -8380
rect 18955 -9118 18989 -6962
rect 21015 -9118 21049 -6962
rect 21287 -8002 21321 -5846
rect 22223 -8002 22257 -5846
rect 22424 -6152 22864 -6118
rect 22328 -7318 22362 -6214
rect 22926 -7318 22960 -6214
rect 22424 -7414 22864 -7380
rect 23185 -7803 23219 -7769
rect 23461 -7803 23495 -7769
rect 23737 -7803 23771 -7769
rect 21383 -8098 22161 -8064
rect 19051 -9214 20953 -9180
rect 16572 -9346 17228 -9312
rect 17227 -10557 17261 -10523
rect 17227 -10833 17261 -10799
<< nsubdiffcont >>
rect 18079 -3266 21925 -3232
rect 17983 -5502 18017 -3328
rect 21987 -5502 22021 -3328
rect 18079 -5598 21925 -5564
rect 23185 -7492 23219 -7458
rect 23185 -7585 23219 -7551
rect 23461 -7492 23495 -7458
rect 23461 -7585 23495 -7551
rect 23737 -7492 23771 -7458
rect 23737 -7585 23771 -7551
rect 16916 -10557 16950 -10523
rect 17009 -10557 17043 -10523
rect 16916 -10833 16950 -10799
rect 17009 -10833 17043 -10799
<< poly >>
rect 18140 -3334 18206 -3318
rect 18140 -3368 18156 -3334
rect 18190 -3368 18206 -3334
rect 18140 -3384 18206 -3368
rect 18258 -3334 18324 -3318
rect 18258 -3368 18274 -3334
rect 18308 -3368 18324 -3334
rect 18258 -3384 18324 -3368
rect 18376 -3334 18442 -3318
rect 18376 -3368 18392 -3334
rect 18426 -3368 18442 -3334
rect 18376 -3384 18442 -3368
rect 18494 -3334 18560 -3318
rect 18494 -3368 18510 -3334
rect 18544 -3368 18560 -3334
rect 18494 -3384 18560 -3368
rect 18612 -3334 18678 -3318
rect 18612 -3368 18628 -3334
rect 18662 -3368 18678 -3334
rect 18612 -3384 18678 -3368
rect 18730 -3334 18796 -3318
rect 18730 -3368 18746 -3334
rect 18780 -3368 18796 -3334
rect 18730 -3384 18796 -3368
rect 18848 -3334 18914 -3318
rect 18848 -3368 18864 -3334
rect 18898 -3368 18914 -3334
rect 18848 -3384 18914 -3368
rect 18966 -3334 19032 -3318
rect 18966 -3368 18982 -3334
rect 19016 -3368 19032 -3334
rect 18966 -3384 19032 -3368
rect 19084 -3334 19150 -3318
rect 19084 -3368 19100 -3334
rect 19134 -3368 19150 -3334
rect 19084 -3384 19150 -3368
rect 19202 -3334 19268 -3318
rect 19202 -3368 19218 -3334
rect 19252 -3368 19268 -3334
rect 19202 -3384 19268 -3368
rect 19320 -3334 19386 -3318
rect 19320 -3368 19336 -3334
rect 19370 -3368 19386 -3334
rect 19320 -3384 19386 -3368
rect 19438 -3334 19504 -3318
rect 19438 -3368 19454 -3334
rect 19488 -3368 19504 -3334
rect 19438 -3384 19504 -3368
rect 19556 -3384 19622 -3318
rect 19674 -3384 19740 -3318
rect 19792 -3384 19858 -3318
rect 19910 -3384 19976 -3318
rect 20028 -3384 20094 -3318
rect 20146 -3384 20212 -3318
rect 20264 -3384 20330 -3318
rect 20382 -3384 20448 -3318
rect 20500 -3334 20566 -3318
rect 20500 -3368 20516 -3334
rect 20550 -3368 20566 -3334
rect 20500 -3384 20566 -3368
rect 20618 -3334 20684 -3318
rect 20618 -3368 20634 -3334
rect 20668 -3368 20684 -3334
rect 20618 -3384 20684 -3368
rect 20736 -3334 20802 -3318
rect 20736 -3368 20752 -3334
rect 20786 -3368 20802 -3334
rect 20736 -3384 20802 -3368
rect 20854 -3334 20920 -3318
rect 20854 -3368 20870 -3334
rect 20904 -3368 20920 -3334
rect 20854 -3384 20920 -3368
rect 20972 -3334 21038 -3318
rect 20972 -3368 20988 -3334
rect 21022 -3368 21038 -3334
rect 20972 -3384 21038 -3368
rect 21090 -3334 21156 -3318
rect 21090 -3368 21106 -3334
rect 21140 -3368 21156 -3334
rect 21090 -3384 21156 -3368
rect 21208 -3334 21274 -3318
rect 21208 -3368 21224 -3334
rect 21258 -3368 21274 -3334
rect 21208 -3384 21274 -3368
rect 21326 -3334 21392 -3318
rect 21326 -3368 21342 -3334
rect 21376 -3368 21392 -3334
rect 21326 -3384 21392 -3368
rect 21444 -3334 21510 -3318
rect 21444 -3368 21460 -3334
rect 21494 -3368 21510 -3334
rect 21444 -3384 21510 -3368
rect 21562 -3334 21628 -3318
rect 21562 -3368 21578 -3334
rect 21612 -3368 21628 -3334
rect 21562 -3384 21628 -3368
rect 21680 -3334 21746 -3318
rect 21680 -3368 21696 -3334
rect 21730 -3368 21746 -3334
rect 21680 -3384 21746 -3368
rect 21798 -3334 21864 -3318
rect 21798 -3368 21814 -3334
rect 21848 -3368 21864 -3334
rect 21798 -3384 21864 -3368
rect 18143 -3415 18203 -3384
rect 18261 -3415 18321 -3384
rect 18379 -3415 18439 -3384
rect 18497 -3415 18557 -3384
rect 18615 -3415 18675 -3384
rect 18733 -3415 18793 -3384
rect 18851 -3415 18911 -3384
rect 18969 -3415 19029 -3384
rect 19087 -3415 19147 -3384
rect 19205 -3415 19265 -3384
rect 19323 -3415 19383 -3384
rect 19441 -3415 19501 -3384
rect 19559 -3415 19619 -3384
rect 19677 -3415 19737 -3384
rect 19795 -3415 19855 -3384
rect 19913 -3415 19973 -3384
rect 20031 -3415 20091 -3384
rect 20149 -3415 20209 -3384
rect 20267 -3415 20327 -3384
rect 20385 -3415 20445 -3384
rect 20503 -3415 20563 -3384
rect 20621 -3415 20681 -3384
rect 20739 -3415 20799 -3384
rect 20857 -3415 20917 -3384
rect 20975 -3415 21035 -3384
rect 21093 -3415 21153 -3384
rect 21211 -3415 21271 -3384
rect 21329 -3415 21389 -3384
rect 21447 -3415 21507 -3384
rect 21565 -3415 21625 -3384
rect 21683 -3415 21743 -3384
rect 21801 -3415 21861 -3384
rect 18143 -5446 18203 -5415
rect 18261 -5446 18321 -5415
rect 18379 -5446 18439 -5415
rect 18497 -5446 18557 -5415
rect 18615 -5446 18675 -5415
rect 18733 -5446 18793 -5415
rect 18851 -5446 18911 -5415
rect 18969 -5446 19029 -5415
rect 19087 -5446 19147 -5415
rect 19205 -5446 19265 -5415
rect 19323 -5446 19383 -5415
rect 19441 -5446 19501 -5415
rect 19559 -5446 19619 -5415
rect 19677 -5446 19737 -5415
rect 19795 -5446 19855 -5415
rect 19913 -5446 19973 -5415
rect 20031 -5446 20091 -5415
rect 20149 -5446 20209 -5415
rect 20267 -5446 20327 -5415
rect 20385 -5446 20445 -5415
rect 20503 -5446 20563 -5415
rect 20621 -5446 20681 -5415
rect 20739 -5446 20799 -5415
rect 20857 -5446 20917 -5415
rect 20975 -5446 21035 -5415
rect 21093 -5446 21153 -5415
rect 21211 -5446 21271 -5415
rect 21329 -5446 21389 -5415
rect 21447 -5446 21507 -5415
rect 21565 -5446 21625 -5415
rect 21683 -5446 21743 -5415
rect 21801 -5446 21861 -5415
rect 18140 -5462 18206 -5446
rect 18140 -5496 18156 -5462
rect 18190 -5496 18206 -5462
rect 18140 -5512 18206 -5496
rect 18258 -5462 18324 -5446
rect 18258 -5496 18274 -5462
rect 18308 -5496 18324 -5462
rect 18258 -5512 18324 -5496
rect 18376 -5462 18442 -5446
rect 18376 -5496 18392 -5462
rect 18426 -5496 18442 -5462
rect 18376 -5512 18442 -5496
rect 18494 -5462 18560 -5446
rect 18494 -5496 18510 -5462
rect 18544 -5496 18560 -5462
rect 18494 -5512 18560 -5496
rect 18612 -5462 18678 -5446
rect 18612 -5496 18628 -5462
rect 18662 -5496 18678 -5462
rect 18612 -5512 18678 -5496
rect 18730 -5462 18796 -5446
rect 18730 -5496 18746 -5462
rect 18780 -5496 18796 -5462
rect 18730 -5512 18796 -5496
rect 18848 -5462 18914 -5446
rect 18848 -5496 18864 -5462
rect 18898 -5496 18914 -5462
rect 18848 -5512 18914 -5496
rect 18966 -5462 19032 -5446
rect 18966 -5496 18982 -5462
rect 19016 -5496 19032 -5462
rect 18966 -5512 19032 -5496
rect 19084 -5462 19150 -5446
rect 19084 -5496 19100 -5462
rect 19134 -5496 19150 -5462
rect 19084 -5512 19150 -5496
rect 19202 -5462 19268 -5446
rect 19202 -5496 19218 -5462
rect 19252 -5496 19268 -5462
rect 19202 -5512 19268 -5496
rect 19320 -5462 19386 -5446
rect 19320 -5496 19336 -5462
rect 19370 -5496 19386 -5462
rect 19320 -5512 19386 -5496
rect 19438 -5462 19504 -5446
rect 19438 -5496 19454 -5462
rect 19488 -5496 19504 -5462
rect 19438 -5512 19504 -5496
rect 19556 -5462 19622 -5446
rect 19556 -5496 19572 -5462
rect 19606 -5496 19622 -5462
rect 19556 -5512 19622 -5496
rect 19674 -5462 19740 -5446
rect 19674 -5496 19690 -5462
rect 19724 -5496 19740 -5462
rect 19674 -5512 19740 -5496
rect 19792 -5462 19858 -5446
rect 19792 -5496 19808 -5462
rect 19842 -5496 19858 -5462
rect 19792 -5512 19858 -5496
rect 19910 -5462 19976 -5446
rect 19910 -5496 19926 -5462
rect 19960 -5496 19976 -5462
rect 19910 -5512 19976 -5496
rect 20028 -5462 20094 -5446
rect 20028 -5496 20044 -5462
rect 20078 -5496 20094 -5462
rect 20028 -5512 20094 -5496
rect 20146 -5462 20212 -5446
rect 20146 -5496 20162 -5462
rect 20196 -5496 20212 -5462
rect 20146 -5512 20212 -5496
rect 20264 -5462 20330 -5446
rect 20264 -5496 20280 -5462
rect 20314 -5496 20330 -5462
rect 20264 -5512 20330 -5496
rect 20382 -5462 20448 -5446
rect 20382 -5496 20398 -5462
rect 20432 -5496 20448 -5462
rect 20382 -5512 20448 -5496
rect 20500 -5462 20566 -5446
rect 20500 -5496 20516 -5462
rect 20550 -5496 20566 -5462
rect 20500 -5512 20566 -5496
rect 20618 -5462 20684 -5446
rect 20618 -5496 20634 -5462
rect 20668 -5496 20684 -5462
rect 20618 -5512 20684 -5496
rect 20736 -5462 20802 -5446
rect 20736 -5496 20752 -5462
rect 20786 -5496 20802 -5462
rect 20736 -5512 20802 -5496
rect 20854 -5462 20920 -5446
rect 20854 -5496 20870 -5462
rect 20904 -5496 20920 -5462
rect 20854 -5512 20920 -5496
rect 20972 -5462 21038 -5446
rect 20972 -5496 20988 -5462
rect 21022 -5496 21038 -5462
rect 20972 -5512 21038 -5496
rect 21090 -5462 21156 -5446
rect 21090 -5496 21106 -5462
rect 21140 -5496 21156 -5462
rect 21090 -5512 21156 -5496
rect 21208 -5462 21274 -5446
rect 21208 -5496 21224 -5462
rect 21258 -5496 21274 -5462
rect 21208 -5512 21274 -5496
rect 21326 -5462 21392 -5446
rect 21326 -5496 21342 -5462
rect 21376 -5496 21392 -5462
rect 21326 -5512 21392 -5496
rect 21444 -5462 21510 -5446
rect 21444 -5496 21460 -5462
rect 21494 -5496 21510 -5462
rect 21444 -5512 21510 -5496
rect 21562 -5462 21628 -5446
rect 21562 -5496 21578 -5462
rect 21612 -5496 21628 -5462
rect 21562 -5512 21628 -5496
rect 21680 -5462 21746 -5446
rect 21680 -5496 21696 -5462
rect 21730 -5496 21746 -5462
rect 21680 -5512 21746 -5496
rect 21798 -5462 21864 -5446
rect 21798 -5496 21814 -5462
rect 21848 -5496 21864 -5462
rect 21798 -5512 21864 -5496
rect 17903 -5852 17969 -5836
rect 17903 -5886 17919 -5852
rect 17953 -5886 17969 -5852
rect 17903 -5902 17969 -5886
rect 18021 -5852 18087 -5836
rect 18021 -5886 18037 -5852
rect 18071 -5886 18087 -5852
rect 18021 -5902 18087 -5886
rect 18139 -5852 18205 -5836
rect 18139 -5886 18155 -5852
rect 18189 -5886 18205 -5852
rect 18139 -5902 18205 -5886
rect 18257 -5852 18323 -5836
rect 18257 -5886 18273 -5852
rect 18307 -5886 18323 -5852
rect 18257 -5902 18323 -5886
rect 18375 -5852 18441 -5836
rect 18375 -5886 18391 -5852
rect 18425 -5886 18441 -5852
rect 18375 -5902 18441 -5886
rect 18493 -5852 18559 -5836
rect 18493 -5886 18509 -5852
rect 18543 -5886 18559 -5852
rect 18493 -5902 18559 -5886
rect 17906 -5924 17966 -5902
rect 18024 -5924 18084 -5902
rect 18142 -5924 18202 -5902
rect 18260 -5924 18320 -5902
rect 18378 -5924 18438 -5902
rect 18496 -5924 18556 -5902
rect 17906 -7946 17966 -7924
rect 18024 -7946 18084 -7924
rect 18142 -7946 18202 -7924
rect 18260 -7946 18320 -7924
rect 18378 -7946 18438 -7924
rect 18496 -7946 18556 -7924
rect 17903 -7962 17969 -7946
rect 17903 -7996 17919 -7962
rect 17953 -7996 17969 -7962
rect 17903 -8012 17969 -7996
rect 18021 -7962 18087 -7946
rect 18021 -7996 18037 -7962
rect 18071 -7996 18087 -7962
rect 18021 -8012 18087 -7996
rect 18139 -7962 18205 -7946
rect 18139 -7996 18155 -7962
rect 18189 -7996 18205 -7962
rect 18139 -8012 18205 -7996
rect 18257 -7962 18323 -7946
rect 18257 -7996 18273 -7962
rect 18307 -7996 18323 -7962
rect 18257 -8012 18323 -7996
rect 18375 -7962 18441 -7946
rect 18375 -7996 18391 -7962
rect 18425 -7996 18441 -7962
rect 18375 -8012 18441 -7996
rect 18493 -7962 18559 -7946
rect 18493 -7996 18509 -7962
rect 18543 -7996 18559 -7962
rect 18493 -8012 18559 -7996
rect 19075 -6024 19201 -5996
rect 19075 -6058 19121 -6024
rect 19155 -6058 19201 -6024
rect 19075 -6074 19201 -6058
rect 20803 -6024 20929 -5996
rect 20803 -6058 20849 -6024
rect 20883 -6058 20929 -6024
rect 20803 -6074 20929 -6058
rect 19075 -6100 19105 -6074
rect 19171 -6100 19201 -6074
rect 19267 -6100 19297 -6074
rect 19363 -6100 19393 -6074
rect 19459 -6100 19489 -6074
rect 19555 -6100 19585 -6074
rect 19651 -6100 19681 -6074
rect 19747 -6100 19777 -6074
rect 19843 -6100 19873 -6074
rect 19939 -6100 19969 -6074
rect 20035 -6100 20065 -6074
rect 20131 -6100 20161 -6074
rect 20227 -6100 20257 -6074
rect 20323 -6100 20353 -6074
rect 20419 -6100 20449 -6074
rect 20515 -6100 20545 -6074
rect 20611 -6100 20641 -6074
rect 20707 -6100 20737 -6074
rect 20803 -6100 20833 -6074
rect 20899 -6100 20929 -6074
rect 19075 -6626 19105 -6600
rect 19171 -6626 19201 -6600
rect 19267 -6622 19297 -6600
rect 19363 -6622 19393 -6600
rect 19267 -6650 19393 -6622
rect 19267 -6684 19313 -6650
rect 19347 -6684 19393 -6650
rect 19267 -6700 19393 -6684
rect 19459 -6622 19489 -6600
rect 19555 -6622 19585 -6600
rect 19459 -6650 19585 -6622
rect 19459 -6684 19505 -6650
rect 19539 -6684 19585 -6650
rect 19459 -6700 19585 -6684
rect 19651 -6622 19681 -6600
rect 19747 -6622 19777 -6600
rect 19651 -6650 19777 -6622
rect 19651 -6684 19697 -6650
rect 19731 -6684 19777 -6650
rect 19651 -6700 19777 -6684
rect 19843 -6622 19873 -6600
rect 19939 -6622 19969 -6600
rect 19843 -6650 19969 -6622
rect 19843 -6684 19889 -6650
rect 19923 -6684 19969 -6650
rect 19843 -6700 19969 -6684
rect 20035 -6622 20065 -6600
rect 20131 -6622 20161 -6600
rect 20035 -6650 20161 -6622
rect 20035 -6684 20081 -6650
rect 20115 -6684 20161 -6650
rect 20035 -6700 20161 -6684
rect 20227 -6622 20257 -6600
rect 20323 -6622 20353 -6600
rect 20227 -6650 20353 -6622
rect 20227 -6684 20273 -6650
rect 20307 -6684 20353 -6650
rect 20227 -6700 20353 -6684
rect 20419 -6622 20449 -6600
rect 20515 -6622 20545 -6600
rect 20419 -6650 20545 -6622
rect 20419 -6684 20465 -6650
rect 20499 -6684 20545 -6650
rect 20419 -6700 20545 -6684
rect 20611 -6622 20641 -6600
rect 20707 -6622 20737 -6600
rect 20611 -6650 20737 -6622
rect 20803 -6626 20833 -6600
rect 20899 -6626 20929 -6600
rect 20611 -6684 20657 -6650
rect 20691 -6684 20737 -6650
rect 20611 -6700 20737 -6684
rect 16562 -8464 16650 -8448
rect 16562 -8498 16578 -8464
rect 16612 -8478 16650 -8464
rect 17150 -8478 17176 -8448
rect 16612 -8498 16628 -8478
rect 16562 -8544 16628 -8498
rect 16562 -8574 16650 -8544
rect 17150 -8574 17176 -8544
rect 16562 -8656 16650 -8640
rect 16562 -8690 16578 -8656
rect 16612 -8670 16650 -8656
rect 17150 -8670 17176 -8640
rect 16612 -8690 16628 -8670
rect 16562 -8736 16628 -8690
rect 16562 -8766 16650 -8736
rect 17150 -8766 17176 -8736
rect 19115 -6968 19515 -6952
rect 19115 -7002 19131 -6968
rect 19499 -7002 19515 -6968
rect 19115 -7040 19515 -7002
rect 19573 -6968 19973 -6952
rect 19573 -7002 19589 -6968
rect 19957 -7002 19973 -6968
rect 19573 -7040 19973 -7002
rect 20031 -6968 20431 -6952
rect 20031 -7002 20047 -6968
rect 20415 -7002 20431 -6968
rect 20031 -7040 20431 -7002
rect 20489 -6968 20889 -6952
rect 20489 -7002 20505 -6968
rect 20873 -7002 20889 -6968
rect 20489 -7040 20889 -7002
rect 19115 -9078 19515 -9040
rect 19115 -9112 19131 -9078
rect 19499 -9112 19515 -9078
rect 19115 -9128 19515 -9112
rect 19573 -9078 19973 -9040
rect 19573 -9112 19589 -9078
rect 19957 -9112 19973 -9078
rect 19573 -9128 19973 -9112
rect 20031 -9078 20431 -9040
rect 20031 -9112 20047 -9078
rect 20415 -9112 20431 -9078
rect 20031 -9128 20431 -9112
rect 20489 -9078 20889 -9040
rect 20489 -9112 20505 -9078
rect 20873 -9112 20889 -9078
rect 20489 -9128 20889 -9112
rect 21444 -5852 21510 -5836
rect 21444 -5886 21460 -5852
rect 21494 -5886 21510 -5852
rect 21444 -5902 21510 -5886
rect 21562 -5852 21628 -5836
rect 21562 -5886 21578 -5852
rect 21612 -5886 21628 -5852
rect 21562 -5902 21628 -5886
rect 21680 -5852 21746 -5836
rect 21680 -5886 21696 -5852
rect 21730 -5886 21746 -5852
rect 21680 -5902 21746 -5886
rect 21798 -5852 21864 -5836
rect 21798 -5886 21814 -5852
rect 21848 -5886 21864 -5852
rect 21798 -5902 21864 -5886
rect 21916 -5852 21982 -5836
rect 21916 -5886 21932 -5852
rect 21966 -5886 21982 -5852
rect 21916 -5902 21982 -5886
rect 22034 -5852 22100 -5836
rect 22034 -5886 22050 -5852
rect 22084 -5886 22100 -5852
rect 22034 -5902 22100 -5886
rect 21447 -5924 21507 -5902
rect 21565 -5924 21625 -5902
rect 21683 -5924 21743 -5902
rect 21801 -5924 21861 -5902
rect 21919 -5924 21979 -5902
rect 22037 -5924 22097 -5902
rect 21447 -7946 21507 -7924
rect 21565 -7946 21625 -7924
rect 21683 -7946 21743 -7924
rect 21801 -7946 21861 -7924
rect 21919 -7946 21979 -7924
rect 22037 -7946 22097 -7924
rect 21444 -7962 21510 -7946
rect 21444 -7996 21460 -7962
rect 21494 -7996 21510 -7962
rect 21444 -8012 21510 -7996
rect 21562 -7962 21628 -7946
rect 21562 -7996 21578 -7962
rect 21612 -7996 21628 -7962
rect 21562 -8012 21628 -7996
rect 21680 -7962 21746 -7946
rect 21680 -7996 21696 -7962
rect 21730 -7996 21746 -7962
rect 21680 -8012 21746 -7996
rect 21798 -7962 21864 -7946
rect 21798 -7996 21814 -7962
rect 21848 -7996 21864 -7962
rect 21798 -8012 21864 -7996
rect 21916 -7962 21982 -7946
rect 21916 -7996 21932 -7962
rect 21966 -7996 21982 -7962
rect 21916 -8012 21982 -7996
rect 22034 -7962 22100 -7946
rect 22034 -7996 22050 -7962
rect 22084 -7996 22100 -7962
rect 22034 -8012 22100 -7996
<< polycont >>
rect 18156 -3368 18190 -3334
rect 18274 -3368 18308 -3334
rect 18392 -3368 18426 -3334
rect 18510 -3368 18544 -3334
rect 18628 -3368 18662 -3334
rect 18746 -3368 18780 -3334
rect 18864 -3368 18898 -3334
rect 18982 -3368 19016 -3334
rect 19100 -3368 19134 -3334
rect 19218 -3368 19252 -3334
rect 19336 -3368 19370 -3334
rect 19454 -3368 19488 -3334
rect 20516 -3368 20550 -3334
rect 20634 -3368 20668 -3334
rect 20752 -3368 20786 -3334
rect 20870 -3368 20904 -3334
rect 20988 -3368 21022 -3334
rect 21106 -3368 21140 -3334
rect 21224 -3368 21258 -3334
rect 21342 -3368 21376 -3334
rect 21460 -3368 21494 -3334
rect 21578 -3368 21612 -3334
rect 21696 -3368 21730 -3334
rect 21814 -3368 21848 -3334
rect 18156 -5496 18190 -5462
rect 18274 -5496 18308 -5462
rect 18392 -5496 18426 -5462
rect 18510 -5496 18544 -5462
rect 18628 -5496 18662 -5462
rect 18746 -5496 18780 -5462
rect 18864 -5496 18898 -5462
rect 18982 -5496 19016 -5462
rect 19100 -5496 19134 -5462
rect 19218 -5496 19252 -5462
rect 19336 -5496 19370 -5462
rect 19454 -5496 19488 -5462
rect 19572 -5496 19606 -5462
rect 19690 -5496 19724 -5462
rect 19808 -5496 19842 -5462
rect 19926 -5496 19960 -5462
rect 20044 -5496 20078 -5462
rect 20162 -5496 20196 -5462
rect 20280 -5496 20314 -5462
rect 20398 -5496 20432 -5462
rect 20516 -5496 20550 -5462
rect 20634 -5496 20668 -5462
rect 20752 -5496 20786 -5462
rect 20870 -5496 20904 -5462
rect 20988 -5496 21022 -5462
rect 21106 -5496 21140 -5462
rect 21224 -5496 21258 -5462
rect 21342 -5496 21376 -5462
rect 21460 -5496 21494 -5462
rect 21578 -5496 21612 -5462
rect 21696 -5496 21730 -5462
rect 21814 -5496 21848 -5462
rect 17919 -5886 17953 -5852
rect 18037 -5886 18071 -5852
rect 18155 -5886 18189 -5852
rect 18273 -5886 18307 -5852
rect 18391 -5886 18425 -5852
rect 18509 -5886 18543 -5852
rect 17919 -7996 17953 -7962
rect 18037 -7996 18071 -7962
rect 18155 -7996 18189 -7962
rect 18273 -7996 18307 -7962
rect 18391 -7996 18425 -7962
rect 18509 -7996 18543 -7962
rect 19121 -6058 19155 -6024
rect 20849 -6058 20883 -6024
rect 19313 -6684 19347 -6650
rect 19505 -6684 19539 -6650
rect 19697 -6684 19731 -6650
rect 19889 -6684 19923 -6650
rect 20081 -6684 20115 -6650
rect 20273 -6684 20307 -6650
rect 20465 -6684 20499 -6650
rect 20657 -6684 20691 -6650
rect 16578 -8498 16612 -8464
rect 16578 -8690 16612 -8656
rect 19131 -7002 19499 -6968
rect 19589 -7002 19957 -6968
rect 20047 -7002 20415 -6968
rect 20505 -7002 20873 -6968
rect 19131 -9112 19499 -9078
rect 19589 -9112 19957 -9078
rect 20047 -9112 20415 -9078
rect 20505 -9112 20873 -9078
rect 21460 -5886 21494 -5852
rect 21578 -5886 21612 -5852
rect 21696 -5886 21730 -5852
rect 21814 -5886 21848 -5852
rect 21932 -5886 21966 -5852
rect 22050 -5886 22084 -5852
rect 21460 -7996 21494 -7962
rect 21578 -7996 21612 -7962
rect 21696 -7996 21730 -7962
rect 21814 -7996 21848 -7962
rect 21932 -7996 21966 -7962
rect 22050 -7996 22084 -7962
<< xpolycontact >>
rect 16606 -9004 17038 -8934
rect 16606 -9170 17038 -9100
rect 22458 -6680 22596 -6248
rect 22692 -6680 22830 -6248
<< ppolyres >>
rect 22458 -7146 22596 -6680
rect 22692 -7146 22830 -6680
rect 22458 -7284 22830 -7146
<< xpolyres >>
rect 17038 -9004 17174 -8934
rect 17104 -9100 17174 -9004
rect 17038 -9170 17174 -9100
<< pdiode >>
rect 23279 -7427 23405 -7409
rect 23279 -7597 23288 -7427
rect 23396 -7597 23405 -7427
rect 23555 -7427 23681 -7409
rect 23279 -7617 23405 -7597
rect 23555 -7597 23564 -7427
rect 23672 -7597 23681 -7427
rect 23555 -7617 23681 -7597
rect 16867 -10626 17075 -10617
rect 16867 -10734 16885 -10626
rect 17055 -10734 17075 -10626
rect 16867 -10743 17075 -10734
<< ndiode >>
rect 23279 -7755 23405 -7737
rect 23279 -7857 23288 -7755
rect 23397 -7857 23405 -7755
rect 23555 -7755 23681 -7737
rect 23279 -7875 23405 -7857
rect 23555 -7857 23564 -7755
rect 23673 -7857 23681 -7755
rect 23555 -7875 23681 -7857
rect 17195 -10626 17333 -10617
rect 17195 -10735 17213 -10626
rect 17315 -10735 17333 -10626
rect 17195 -10743 17333 -10735
<< pdiodec >>
rect 23288 -7597 23396 -7427
rect 23564 -7597 23672 -7427
rect 16885 -10734 17055 -10626
<< ndiodec >>
rect 23288 -7857 23397 -7755
rect 23564 -7857 23673 -7755
rect 17213 -10735 17315 -10626
<< locali >>
rect 17983 -3266 18079 -3232
rect 21925 -3266 22021 -3232
rect 17983 -3328 18017 -3266
rect 21987 -3328 22021 -3266
rect 18140 -3368 18156 -3334
rect 18190 -3368 18206 -3334
rect 18258 -3368 18274 -3334
rect 18308 -3368 18324 -3334
rect 18376 -3368 18392 -3334
rect 18426 -3368 18442 -3334
rect 18494 -3368 18510 -3334
rect 18544 -3368 18560 -3334
rect 18612 -3368 18628 -3334
rect 18662 -3368 18678 -3334
rect 18730 -3368 18746 -3334
rect 18780 -3368 18796 -3334
rect 18848 -3368 18864 -3334
rect 18898 -3368 18914 -3334
rect 18966 -3368 18982 -3334
rect 19016 -3368 19032 -3334
rect 19084 -3368 19100 -3334
rect 19134 -3368 19150 -3334
rect 19202 -3368 19218 -3334
rect 19252 -3368 19268 -3334
rect 19320 -3368 19336 -3334
rect 19370 -3368 19386 -3334
rect 19438 -3368 19454 -3334
rect 19488 -3368 19504 -3334
rect 20500 -3368 20516 -3334
rect 20550 -3368 20566 -3334
rect 20618 -3368 20634 -3334
rect 20668 -3368 20684 -3334
rect 20736 -3368 20752 -3334
rect 20786 -3368 20802 -3334
rect 20854 -3368 20870 -3334
rect 20904 -3368 20920 -3334
rect 20972 -3368 20988 -3334
rect 21022 -3368 21038 -3334
rect 21090 -3368 21106 -3334
rect 21140 -3368 21156 -3334
rect 21208 -3368 21224 -3334
rect 21258 -3368 21274 -3334
rect 21326 -3368 21342 -3334
rect 21376 -3368 21392 -3334
rect 21444 -3368 21460 -3334
rect 21494 -3368 21510 -3334
rect 21562 -3368 21578 -3334
rect 21612 -3368 21628 -3334
rect 21680 -3368 21696 -3334
rect 21730 -3368 21746 -3334
rect 21798 -3368 21814 -3334
rect 21848 -3368 21864 -3334
rect 18097 -3427 18131 -3411
rect 18097 -5419 18131 -5403
rect 18215 -3427 18249 -3411
rect 18215 -5419 18249 -5403
rect 18333 -3427 18367 -3411
rect 18333 -5419 18367 -5403
rect 18451 -3427 18485 -3411
rect 18451 -5419 18485 -5403
rect 18569 -3427 18603 -3411
rect 18569 -5419 18603 -5403
rect 18687 -3427 18721 -3411
rect 18687 -5419 18721 -5403
rect 18805 -3427 18839 -3411
rect 18805 -5419 18839 -5403
rect 18923 -3427 18957 -3411
rect 18923 -5419 18957 -5403
rect 19041 -3427 19075 -3411
rect 19041 -5419 19075 -5403
rect 19159 -3427 19193 -3411
rect 19159 -5419 19193 -5403
rect 19277 -3427 19311 -3411
rect 19277 -5419 19311 -5403
rect 19395 -3427 19429 -3411
rect 19395 -5419 19429 -5403
rect 19513 -3427 19547 -3411
rect 19513 -5419 19547 -5403
rect 19631 -3427 19665 -3411
rect 19631 -5419 19665 -5403
rect 19749 -3427 19783 -3411
rect 19749 -5419 19783 -5403
rect 19867 -3427 19901 -3411
rect 19867 -5419 19901 -5403
rect 19985 -3427 20019 -3411
rect 19985 -5419 20019 -5403
rect 20103 -3427 20137 -3411
rect 20103 -5419 20137 -5403
rect 20221 -3427 20255 -3411
rect 20221 -5419 20255 -5403
rect 20339 -3427 20373 -3411
rect 20339 -5419 20373 -5403
rect 20457 -3427 20491 -3411
rect 20457 -5419 20491 -5403
rect 20575 -3427 20609 -3411
rect 20575 -5419 20609 -5403
rect 20693 -3427 20727 -3411
rect 20693 -5419 20727 -5403
rect 20811 -3427 20845 -3411
rect 20811 -5419 20845 -5403
rect 20929 -3427 20963 -3411
rect 20929 -5419 20963 -5403
rect 21047 -3427 21081 -3411
rect 21047 -5419 21081 -5403
rect 21165 -3427 21199 -3411
rect 21165 -5419 21199 -5403
rect 21283 -3427 21317 -3411
rect 21283 -5419 21317 -5403
rect 21401 -3427 21435 -3411
rect 21401 -5419 21435 -5403
rect 21519 -3427 21553 -3411
rect 21519 -5419 21553 -5403
rect 21637 -3427 21671 -3411
rect 21637 -5419 21671 -5403
rect 21755 -3427 21789 -3411
rect 21755 -5419 21789 -5403
rect 21873 -3427 21907 -3411
rect 21873 -5419 21907 -5403
rect 18140 -5496 18156 -5462
rect 18190 -5496 18206 -5462
rect 18258 -5496 18274 -5462
rect 18308 -5496 18324 -5462
rect 18376 -5496 18392 -5462
rect 18426 -5496 18442 -5462
rect 18494 -5496 18510 -5462
rect 18544 -5496 18560 -5462
rect 18612 -5496 18628 -5462
rect 18662 -5496 18678 -5462
rect 18730 -5496 18746 -5462
rect 18780 -5496 18796 -5462
rect 18848 -5496 18864 -5462
rect 18898 -5496 18914 -5462
rect 18966 -5496 18982 -5462
rect 19016 -5496 19032 -5462
rect 19084 -5496 19100 -5462
rect 19134 -5496 19150 -5462
rect 19202 -5496 19218 -5462
rect 19252 -5496 19268 -5462
rect 19320 -5496 19336 -5462
rect 19370 -5496 19386 -5462
rect 19438 -5496 19454 -5462
rect 19488 -5496 19504 -5462
rect 19556 -5496 19572 -5462
rect 19606 -5496 19622 -5462
rect 19674 -5496 19690 -5462
rect 19724 -5496 19740 -5462
rect 19792 -5496 19808 -5462
rect 19842 -5496 19858 -5462
rect 19910 -5496 19926 -5462
rect 19960 -5496 19976 -5462
rect 20028 -5496 20044 -5462
rect 20078 -5496 20094 -5462
rect 20146 -5496 20162 -5462
rect 20196 -5496 20212 -5462
rect 20264 -5496 20280 -5462
rect 20314 -5496 20330 -5462
rect 20382 -5496 20398 -5462
rect 20432 -5496 20448 -5462
rect 20500 -5496 20516 -5462
rect 20550 -5496 20566 -5462
rect 20618 -5496 20634 -5462
rect 20668 -5496 20684 -5462
rect 20736 -5496 20752 -5462
rect 20786 -5496 20802 -5462
rect 20854 -5496 20870 -5462
rect 20904 -5496 20920 -5462
rect 20972 -5496 20988 -5462
rect 21022 -5496 21038 -5462
rect 21090 -5496 21106 -5462
rect 21140 -5496 21156 -5462
rect 21208 -5496 21224 -5462
rect 21258 -5496 21274 -5462
rect 21326 -5496 21342 -5462
rect 21376 -5496 21392 -5462
rect 21444 -5496 21460 -5462
rect 21494 -5496 21510 -5462
rect 21562 -5496 21578 -5462
rect 21612 -5496 21628 -5462
rect 21680 -5496 21696 -5462
rect 21730 -5496 21746 -5462
rect 21798 -5496 21814 -5462
rect 21848 -5496 21864 -5462
rect 17983 -5564 18017 -5502
rect 21987 -5564 22021 -5502
rect 17983 -5598 18079 -5564
rect 21925 -5598 22021 -5564
rect 17746 -5784 17842 -5750
rect 18620 -5784 18716 -5750
rect 17746 -5846 17780 -5784
rect 18682 -5846 18716 -5784
rect 17903 -5886 17919 -5852
rect 17953 -5886 17969 -5852
rect 18021 -5886 18037 -5852
rect 18071 -5886 18087 -5852
rect 18139 -5886 18155 -5852
rect 18189 -5886 18205 -5852
rect 18257 -5886 18273 -5852
rect 18307 -5886 18323 -5852
rect 18375 -5886 18391 -5852
rect 18425 -5886 18441 -5852
rect 18493 -5886 18509 -5852
rect 18543 -5886 18559 -5852
rect 17860 -5936 17894 -5920
rect 17860 -7928 17894 -7912
rect 17978 -5936 18012 -5920
rect 17978 -7928 18012 -7912
rect 18096 -5936 18130 -5920
rect 18096 -7928 18130 -7912
rect 18214 -5936 18248 -5920
rect 18214 -7928 18248 -7912
rect 18332 -5936 18366 -5920
rect 18332 -7928 18366 -7912
rect 18450 -5936 18484 -5920
rect 18450 -7928 18484 -7912
rect 18568 -5936 18602 -5920
rect 18568 -7928 18602 -7912
rect 21287 -5784 21383 -5750
rect 22161 -5784 22257 -5750
rect 21287 -5846 21321 -5784
rect 22223 -5846 22257 -5784
rect 21444 -5886 21460 -5852
rect 21494 -5886 21510 -5852
rect 21562 -5886 21578 -5852
rect 21612 -5886 21628 -5852
rect 21680 -5886 21696 -5852
rect 21730 -5886 21746 -5852
rect 21798 -5886 21814 -5852
rect 21848 -5886 21864 -5852
rect 21916 -5886 21932 -5852
rect 21966 -5886 21982 -5852
rect 22034 -5886 22050 -5852
rect 22084 -5886 22100 -5852
rect 18911 -5960 19007 -5926
rect 20997 -5960 21093 -5926
rect 18911 -6022 18945 -5960
rect 21059 -6022 21093 -5960
rect 19105 -6058 19121 -6024
rect 19155 -6058 19171 -6024
rect 20833 -6058 20849 -6024
rect 20883 -6058 20899 -6024
rect 19025 -6112 19059 -6096
rect 19025 -6604 19059 -6588
rect 19121 -6112 19155 -6096
rect 19121 -6604 19155 -6588
rect 19217 -6112 19251 -6096
rect 19217 -6604 19251 -6588
rect 19313 -6112 19347 -6096
rect 19313 -6604 19347 -6588
rect 19409 -6112 19443 -6096
rect 19409 -6604 19443 -6588
rect 19505 -6112 19539 -6096
rect 19505 -6604 19539 -6588
rect 19601 -6112 19635 -6096
rect 19601 -6604 19635 -6588
rect 19697 -6112 19731 -6096
rect 19697 -6604 19731 -6588
rect 19793 -6112 19827 -6096
rect 19793 -6604 19827 -6588
rect 19889 -6112 19923 -6096
rect 19889 -6604 19923 -6588
rect 19985 -6112 20019 -6096
rect 19985 -6604 20019 -6588
rect 20081 -6112 20115 -6096
rect 20081 -6604 20115 -6588
rect 20177 -6112 20211 -6096
rect 20177 -6604 20211 -6588
rect 20273 -6112 20307 -6096
rect 20273 -6604 20307 -6588
rect 20369 -6112 20403 -6096
rect 20369 -6604 20403 -6588
rect 20465 -6112 20499 -6096
rect 20465 -6604 20499 -6588
rect 20561 -6112 20595 -6096
rect 20561 -6604 20595 -6588
rect 20657 -6112 20691 -6096
rect 20657 -6604 20691 -6588
rect 20753 -6112 20787 -6096
rect 20753 -6604 20787 -6588
rect 20849 -6112 20883 -6096
rect 20849 -6604 20883 -6588
rect 20945 -6112 20979 -6096
rect 20945 -6604 20979 -6588
rect 18911 -6740 18945 -6678
rect 19297 -6684 19313 -6650
rect 19347 -6684 19363 -6650
rect 19489 -6684 19505 -6650
rect 19539 -6684 19555 -6650
rect 19681 -6684 19697 -6650
rect 19731 -6684 19747 -6650
rect 19873 -6684 19889 -6650
rect 19923 -6684 19939 -6650
rect 20065 -6684 20081 -6650
rect 20115 -6684 20131 -6650
rect 20257 -6684 20273 -6650
rect 20307 -6684 20323 -6650
rect 20449 -6684 20465 -6650
rect 20499 -6684 20515 -6650
rect 20641 -6684 20657 -6650
rect 20691 -6684 20707 -6650
rect 21059 -6740 21093 -6678
rect 18911 -6774 19007 -6740
rect 20997 -6774 21093 -6740
rect 17903 -7996 17919 -7962
rect 17953 -7996 17969 -7962
rect 18021 -7996 18037 -7962
rect 18071 -7996 18087 -7962
rect 18139 -7996 18155 -7962
rect 18189 -7996 18205 -7962
rect 18257 -7996 18273 -7962
rect 18307 -7996 18323 -7962
rect 18375 -7996 18391 -7962
rect 18425 -7996 18441 -7962
rect 18493 -7996 18509 -7962
rect 18543 -7996 18559 -7962
rect 17746 -8064 17780 -8002
rect 18682 -8064 18716 -8002
rect 17746 -8098 17842 -8064
rect 18620 -8098 18716 -8064
rect 18955 -6900 19051 -6866
rect 20953 -6900 21049 -6866
rect 18955 -6962 18989 -6900
rect 21015 -6962 21049 -6900
rect 19115 -7002 19131 -6968
rect 19499 -7002 19515 -6968
rect 19573 -7002 19589 -6968
rect 19957 -7002 19973 -6968
rect 20031 -7002 20047 -6968
rect 20415 -7002 20431 -6968
rect 20489 -7002 20505 -6968
rect 20873 -7002 20889 -6968
rect 16442 -8284 17358 -8250
rect 16442 -8318 16572 -8284
rect 17228 -8318 17358 -8284
rect 16442 -8380 16510 -8318
rect 16442 -9230 16476 -8380
rect 17290 -8380 17358 -8318
rect 16646 -8432 16662 -8398
rect 17138 -8432 17154 -8398
rect 16578 -8464 16612 -8448
rect 16578 -8514 16612 -8498
rect 16646 -8528 16662 -8494
rect 17138 -8528 17154 -8494
rect 16646 -8624 16662 -8590
rect 17138 -8624 17154 -8590
rect 16578 -8656 16612 -8640
rect 16578 -8706 16612 -8690
rect 16646 -8720 16662 -8686
rect 17138 -8720 17290 -8686
rect 16567 -8816 16662 -8782
rect 17138 -8816 17154 -8782
rect 16567 -8934 16618 -8816
rect 16567 -9004 16606 -8934
rect 16567 -9108 16606 -9100
rect 16567 -9161 16590 -9108
rect 16567 -9170 16606 -9161
rect 16442 -9312 16510 -9230
rect 17324 -8420 17358 -8380
rect 17324 -8440 17480 -8420
rect 17324 -9230 17400 -8440
rect 17290 -9312 17400 -9230
rect 16442 -9346 16572 -9312
rect 17228 -9346 17400 -9312
rect 16442 -9360 17400 -9346
rect 17460 -9360 17480 -8440
rect 19069 -7052 19103 -7036
rect 19069 -9044 19103 -9028
rect 19527 -7052 19561 -7036
rect 19527 -9044 19561 -9028
rect 19985 -7052 20019 -7036
rect 19985 -9044 20019 -9028
rect 20443 -7052 20477 -7036
rect 20443 -9044 20477 -9028
rect 20901 -7052 20935 -7036
rect 20901 -9044 20935 -9028
rect 21401 -5936 21435 -5920
rect 21401 -7928 21435 -7912
rect 21519 -5936 21553 -5920
rect 21519 -7928 21553 -7912
rect 21637 -5936 21671 -5920
rect 21637 -7928 21671 -7912
rect 21755 -5936 21789 -5920
rect 21755 -7928 21789 -7912
rect 21873 -5936 21907 -5920
rect 21873 -7928 21907 -7912
rect 21991 -5936 22025 -5920
rect 21991 -7928 22025 -7912
rect 22109 -5936 22143 -5920
rect 22109 -7928 22143 -7912
rect 22328 -6140 22424 -6118
rect 22257 -6152 22424 -6140
rect 22864 -6152 22960 -6118
rect 22257 -6214 22362 -6152
rect 22257 -7318 22328 -6214
rect 22926 -6214 22960 -6152
rect 22257 -7380 22362 -7318
rect 22926 -7380 22960 -7318
rect 22328 -7414 22424 -7380
rect 22864 -7414 22960 -7380
rect 23156 -7387 23185 -7353
rect 23219 -7387 23277 -7353
rect 23311 -7387 23369 -7353
rect 23403 -7387 23461 -7353
rect 23495 -7387 23553 -7353
rect 23587 -7387 23645 -7353
rect 23679 -7387 23737 -7353
rect 23771 -7387 23800 -7353
rect 23173 -7458 23231 -7387
rect 23173 -7492 23185 -7458
rect 23219 -7492 23231 -7458
rect 23173 -7551 23231 -7492
rect 23173 -7585 23185 -7551
rect 23219 -7585 23231 -7551
rect 23173 -7620 23231 -7585
rect 23265 -7427 23415 -7421
rect 23265 -7597 23288 -7427
rect 23396 -7597 23415 -7427
rect 23265 -7662 23415 -7597
rect 23449 -7458 23507 -7387
rect 23449 -7492 23461 -7458
rect 23495 -7492 23507 -7458
rect 23449 -7551 23507 -7492
rect 23449 -7585 23461 -7551
rect 23495 -7585 23507 -7551
rect 23449 -7620 23507 -7585
rect 23541 -7427 23691 -7421
rect 23541 -7597 23564 -7427
rect 23672 -7597 23691 -7427
rect 23265 -7702 23280 -7662
rect 23400 -7702 23415 -7662
rect 23173 -7769 23231 -7752
rect 23173 -7803 23185 -7769
rect 23219 -7803 23231 -7769
rect 23173 -7897 23231 -7803
rect 23265 -7755 23415 -7702
rect 23541 -7662 23691 -7597
rect 23725 -7458 23783 -7387
rect 23725 -7492 23737 -7458
rect 23771 -7492 23783 -7458
rect 23725 -7551 23783 -7492
rect 23725 -7585 23737 -7551
rect 23771 -7585 23783 -7551
rect 23725 -7620 23783 -7585
rect 23541 -7702 23556 -7662
rect 23676 -7702 23691 -7662
rect 23265 -7857 23288 -7755
rect 23397 -7857 23415 -7755
rect 23265 -7863 23415 -7857
rect 23449 -7769 23507 -7752
rect 23449 -7803 23461 -7769
rect 23495 -7803 23507 -7769
rect 23449 -7897 23507 -7803
rect 23541 -7755 23691 -7702
rect 23541 -7857 23564 -7755
rect 23673 -7857 23691 -7755
rect 23541 -7863 23691 -7857
rect 23725 -7769 23783 -7752
rect 23725 -7803 23737 -7769
rect 23771 -7803 23783 -7769
rect 23725 -7897 23783 -7803
rect 21444 -7996 21460 -7962
rect 21494 -7996 21510 -7962
rect 21562 -7996 21578 -7962
rect 21612 -7996 21628 -7962
rect 21680 -7996 21696 -7962
rect 21730 -7996 21746 -7962
rect 21798 -7996 21814 -7962
rect 21848 -7996 21864 -7962
rect 21916 -7996 21932 -7962
rect 21966 -7996 21982 -7962
rect 22034 -7996 22050 -7962
rect 22084 -7996 22100 -7962
rect 21287 -8064 21321 -8002
rect 23156 -7931 23185 -7897
rect 23219 -7931 23277 -7897
rect 23311 -7931 23369 -7897
rect 23403 -7931 23461 -7897
rect 23495 -7931 23553 -7897
rect 23587 -7931 23645 -7897
rect 23679 -7931 23737 -7897
rect 23771 -7931 23800 -7897
rect 22223 -8064 22257 -8002
rect 21287 -8098 21383 -8064
rect 22161 -8098 22257 -8064
rect 19115 -9112 19131 -9078
rect 19499 -9112 19515 -9078
rect 19573 -9112 19589 -9078
rect 19957 -9112 19973 -9078
rect 20031 -9112 20047 -9078
rect 20415 -9112 20431 -9078
rect 20489 -9112 20505 -9078
rect 20873 -9112 20889 -9078
rect 18955 -9180 18989 -9118
rect 21015 -9180 21049 -9118
rect 18955 -9214 19051 -9180
rect 20953 -9214 21049 -9180
rect 16442 -9380 17480 -9360
rect 16811 -10511 16845 -10494
rect 17355 -10511 17389 -10494
rect 16811 -10523 17078 -10511
rect 16845 -10557 16916 -10523
rect 16950 -10557 17009 -10523
rect 17043 -10557 17078 -10523
rect 16811 -10569 17078 -10557
rect 17210 -10523 17389 -10511
rect 17210 -10557 17227 -10523
rect 17261 -10557 17355 -10523
rect 17210 -10569 17389 -10557
rect 16811 -10615 16845 -10569
rect 16811 -10707 16845 -10649
rect 16811 -10787 16845 -10741
rect 16879 -10618 17321 -10603
rect 16879 -10626 17120 -10618
rect 16879 -10734 16885 -10626
rect 17055 -10734 17120 -10626
rect 16879 -10738 17120 -10734
rect 17160 -10626 17321 -10618
rect 17160 -10735 17213 -10626
rect 17315 -10735 17321 -10626
rect 17160 -10738 17321 -10735
rect 16879 -10753 17321 -10738
rect 17355 -10615 17389 -10569
rect 17355 -10707 17389 -10649
rect 17355 -10787 17389 -10741
rect 16811 -10799 17078 -10787
rect 16845 -10833 16916 -10799
rect 16950 -10833 17009 -10799
rect 17043 -10833 17078 -10799
rect 16811 -10845 17078 -10833
rect 17210 -10799 17389 -10787
rect 17210 -10833 17227 -10799
rect 17261 -10833 17355 -10799
rect 17210 -10845 17389 -10833
rect 16811 -10862 16845 -10845
rect 17355 -10862 17389 -10845
<< viali >>
rect 18156 -3368 18190 -3334
rect 18274 -3368 18308 -3334
rect 18392 -3368 18426 -3334
rect 18510 -3368 18544 -3334
rect 18628 -3368 18662 -3334
rect 18746 -3368 18780 -3334
rect 18864 -3368 18898 -3334
rect 18982 -3368 19016 -3334
rect 19100 -3368 19134 -3334
rect 19218 -3368 19252 -3334
rect 19336 -3368 19370 -3334
rect 19454 -3368 19488 -3334
rect 20516 -3368 20550 -3334
rect 20634 -3368 20668 -3334
rect 20752 -3368 20786 -3334
rect 20870 -3368 20904 -3334
rect 20988 -3368 21022 -3334
rect 21106 -3368 21140 -3334
rect 21224 -3368 21258 -3334
rect 21342 -3368 21376 -3334
rect 21460 -3368 21494 -3334
rect 21578 -3368 21612 -3334
rect 21696 -3368 21730 -3334
rect 21814 -3368 21848 -3334
rect 17983 -3815 18017 -3415
rect 17983 -5415 18017 -5015
rect 18097 -5403 18131 -3427
rect 18215 -5403 18249 -3427
rect 18333 -5403 18367 -3427
rect 18451 -5403 18485 -3427
rect 18569 -5403 18603 -3427
rect 18687 -5403 18721 -3427
rect 18805 -5403 18839 -3427
rect 18923 -5403 18957 -3427
rect 19041 -5403 19075 -3427
rect 19159 -5403 19193 -3427
rect 19277 -5403 19311 -3427
rect 19395 -5403 19429 -3427
rect 19513 -5403 19547 -3427
rect 19631 -5403 19665 -3427
rect 19749 -5403 19783 -3427
rect 19867 -5403 19901 -3427
rect 19985 -5403 20019 -3427
rect 20103 -5403 20137 -3427
rect 20221 -5403 20255 -3427
rect 20339 -5403 20373 -3427
rect 20457 -5403 20491 -3427
rect 20575 -5403 20609 -3427
rect 20693 -5403 20727 -3427
rect 20811 -5403 20845 -3427
rect 20929 -5403 20963 -3427
rect 21047 -5403 21081 -3427
rect 21165 -5403 21199 -3427
rect 21283 -5403 21317 -3427
rect 21401 -5403 21435 -3427
rect 21519 -5403 21553 -3427
rect 21637 -5403 21671 -3427
rect 21755 -5403 21789 -3427
rect 21873 -5403 21907 -3427
rect 21987 -3815 22021 -3415
rect 21987 -5415 22021 -5015
rect 18156 -5496 18190 -5462
rect 18274 -5496 18308 -5462
rect 18392 -5496 18426 -5462
rect 18510 -5496 18544 -5462
rect 18628 -5496 18662 -5462
rect 18746 -5496 18780 -5462
rect 18864 -5496 18898 -5462
rect 18982 -5496 19016 -5462
rect 19100 -5496 19134 -5462
rect 19218 -5496 19252 -5462
rect 19336 -5496 19370 -5462
rect 19454 -5496 19488 -5462
rect 19572 -5496 19606 -5462
rect 19690 -5496 19724 -5462
rect 19808 -5496 19842 -5462
rect 19926 -5496 19960 -5462
rect 20044 -5496 20078 -5462
rect 20162 -5496 20196 -5462
rect 20280 -5496 20314 -5462
rect 20398 -5496 20432 -5462
rect 20516 -5496 20550 -5462
rect 20634 -5496 20668 -5462
rect 20752 -5496 20786 -5462
rect 20870 -5496 20904 -5462
rect 20988 -5496 21022 -5462
rect 21106 -5496 21140 -5462
rect 21224 -5496 21258 -5462
rect 21342 -5496 21376 -5462
rect 21460 -5496 21494 -5462
rect 21578 -5496 21612 -5462
rect 21696 -5496 21730 -5462
rect 21814 -5496 21848 -5462
rect 17919 -5886 17953 -5852
rect 18037 -5886 18071 -5852
rect 18155 -5886 18189 -5852
rect 18273 -5886 18307 -5852
rect 18391 -5886 18425 -5852
rect 18509 -5886 18543 -5852
rect 17746 -6324 17780 -5924
rect 17746 -7924 17780 -7524
rect 17860 -7912 17894 -5936
rect 17978 -7912 18012 -5936
rect 18096 -7912 18130 -5936
rect 18214 -7912 18248 -5936
rect 18332 -7912 18366 -5936
rect 18450 -7912 18484 -5936
rect 18568 -7912 18602 -5936
rect 18682 -6324 18716 -5924
rect 21460 -5886 21494 -5852
rect 21578 -5886 21612 -5852
rect 21696 -5886 21730 -5852
rect 21814 -5886 21848 -5852
rect 21932 -5886 21966 -5852
rect 22050 -5886 22084 -5852
rect 19121 -6058 19155 -6024
rect 20849 -6058 20883 -6024
rect 18911 -6600 18945 -6100
rect 19025 -6588 19059 -6112
rect 19121 -6588 19155 -6112
rect 19217 -6588 19251 -6112
rect 19313 -6588 19347 -6112
rect 19409 -6588 19443 -6112
rect 19505 -6588 19539 -6112
rect 19601 -6588 19635 -6112
rect 19697 -6588 19731 -6112
rect 19793 -6588 19827 -6112
rect 19889 -6588 19923 -6112
rect 19985 -6588 20019 -6112
rect 20081 -6588 20115 -6112
rect 20177 -6588 20211 -6112
rect 20273 -6588 20307 -6112
rect 20369 -6588 20403 -6112
rect 20465 -6588 20499 -6112
rect 20561 -6588 20595 -6112
rect 20657 -6588 20691 -6112
rect 20753 -6588 20787 -6112
rect 20849 -6588 20883 -6112
rect 20945 -6588 20979 -6112
rect 21059 -6600 21093 -6100
rect 19313 -6684 19347 -6650
rect 19505 -6684 19539 -6650
rect 19697 -6684 19731 -6650
rect 19889 -6684 19923 -6650
rect 20081 -6684 20115 -6650
rect 20273 -6684 20307 -6650
rect 20465 -6684 20499 -6650
rect 20657 -6684 20691 -6650
rect 21287 -6324 21321 -5924
rect 18682 -7924 18716 -7524
rect 17919 -7996 17953 -7962
rect 18037 -7996 18071 -7962
rect 18155 -7996 18189 -7962
rect 18273 -7996 18307 -7962
rect 18391 -7996 18425 -7962
rect 18509 -7996 18543 -7962
rect 19131 -7002 19499 -6968
rect 19589 -7002 19957 -6968
rect 20047 -7002 20415 -6968
rect 20505 -7002 20873 -6968
rect 18955 -7440 18989 -7040
rect 16662 -8432 17138 -8398
rect 16578 -8498 16612 -8464
rect 16662 -8528 17138 -8494
rect 16662 -8624 17138 -8590
rect 16578 -8690 16612 -8656
rect 16662 -8720 17138 -8686
rect 16662 -8816 17138 -8782
rect 16590 -9161 16606 -9108
rect 16606 -9161 17022 -9108
rect 17400 -9360 17460 -8440
rect 18955 -9040 18989 -8640
rect 19069 -9028 19103 -7052
rect 19527 -9028 19561 -7052
rect 19985 -9028 20019 -7052
rect 20443 -9028 20477 -7052
rect 20901 -9028 20935 -7052
rect 21015 -7440 21049 -7040
rect 21287 -7924 21321 -7524
rect 21401 -7912 21435 -5936
rect 21519 -7912 21553 -5936
rect 21637 -7912 21671 -5936
rect 21755 -7912 21789 -5936
rect 21873 -7912 21907 -5936
rect 21991 -7912 22025 -5936
rect 22109 -7912 22143 -5936
rect 22223 -6324 22257 -5924
rect 22472 -6660 22582 -6270
rect 22702 -6660 22812 -6270
rect 23185 -7387 23219 -7353
rect 23277 -7387 23311 -7353
rect 23369 -7387 23403 -7353
rect 23461 -7387 23495 -7353
rect 23553 -7387 23587 -7353
rect 23645 -7387 23679 -7353
rect 23737 -7387 23771 -7353
rect 22223 -7924 22257 -7524
rect 23280 -7702 23400 -7662
rect 23556 -7702 23676 -7662
rect 21460 -7996 21494 -7962
rect 21578 -7996 21612 -7962
rect 21696 -7996 21730 -7962
rect 21814 -7996 21848 -7962
rect 21932 -7996 21966 -7962
rect 22050 -7996 22084 -7962
rect 23185 -7931 23219 -7897
rect 23277 -7931 23311 -7897
rect 23369 -7931 23403 -7897
rect 23461 -7931 23495 -7897
rect 23553 -7931 23587 -7897
rect 23645 -7931 23679 -7897
rect 23737 -7931 23771 -7897
rect 21015 -9040 21049 -8640
rect 19131 -9112 19499 -9078
rect 19589 -9112 19957 -9078
rect 20047 -9112 20415 -9078
rect 20505 -9112 20873 -9078
rect 16811 -10557 16845 -10523
rect 17355 -10557 17389 -10523
rect 16811 -10649 16845 -10615
rect 16811 -10741 16845 -10707
rect 17120 -10738 17160 -10618
rect 17355 -10649 17389 -10615
rect 17355 -10741 17389 -10707
rect 16811 -10833 16845 -10799
rect 17355 -10833 17389 -10799
<< metal1 >>
rect 18088 -3334 18206 -3328
rect 18088 -3368 18156 -3334
rect 18190 -3368 18206 -3334
rect 18088 -3374 18206 -3368
rect 18258 -3334 19504 -3328
rect 18258 -3368 18274 -3334
rect 18308 -3368 18392 -3334
rect 18426 -3368 18510 -3334
rect 18544 -3368 18628 -3334
rect 18662 -3368 18746 -3334
rect 18780 -3368 18864 -3334
rect 18898 -3368 18982 -3334
rect 19016 -3368 19100 -3334
rect 19134 -3368 19218 -3334
rect 19252 -3368 19336 -3334
rect 19370 -3368 19454 -3334
rect 19488 -3368 19504 -3334
rect 18258 -3374 19504 -3368
rect 20500 -3334 21746 -3328
rect 20500 -3368 20516 -3334
rect 20550 -3368 20634 -3334
rect 20668 -3368 20752 -3334
rect 20786 -3368 20870 -3334
rect 20904 -3368 20988 -3334
rect 21022 -3368 21106 -3334
rect 21140 -3368 21224 -3334
rect 21258 -3368 21342 -3334
rect 21376 -3368 21460 -3334
rect 21494 -3368 21578 -3334
rect 21612 -3368 21696 -3334
rect 21730 -3368 21746 -3334
rect 20500 -3374 21746 -3368
rect 21798 -3334 21916 -3328
rect 21798 -3368 21814 -3334
rect 21848 -3368 21916 -3334
rect 21798 -3374 21916 -3368
rect 17977 -3415 18023 -3403
rect 18088 -3415 18140 -3374
rect 17977 -3815 17983 -3415
rect 18017 -3427 18140 -3415
rect 18017 -3815 18088 -3427
rect 17977 -3827 18023 -3815
rect 17977 -5015 18023 -5003
rect 17977 -5415 17983 -5015
rect 18017 -5403 18088 -5015
rect 18017 -5415 18140 -5403
rect 17977 -5427 18023 -5415
rect 18088 -5456 18140 -5415
rect 18206 -3427 18258 -3415
rect 18206 -5416 18258 -5403
rect 18324 -3427 18376 -3415
rect 18324 -5415 18376 -5403
rect 18442 -3427 18494 -3415
rect 18442 -5415 18494 -5403
rect 18560 -3427 18612 -3415
rect 18560 -5415 18612 -5403
rect 18678 -3427 18730 -3415
rect 18678 -5415 18730 -5403
rect 18796 -3427 18848 -3415
rect 18796 -5415 18848 -5403
rect 18914 -3427 18966 -3415
rect 18914 -5415 18966 -5403
rect 19032 -3427 19084 -3415
rect 19032 -5415 19084 -5403
rect 19150 -3427 19202 -3415
rect 19150 -5415 19202 -5403
rect 19268 -3427 19320 -3415
rect 19268 -5415 19320 -5403
rect 19386 -3427 19438 -3374
rect 19386 -5456 19438 -5403
rect 19504 -3427 19556 -3415
rect 19504 -5415 19556 -5403
rect 19622 -3427 19674 -3414
rect 19622 -5415 19674 -5403
rect 19740 -3427 19792 -3415
rect 19740 -5415 19792 -5403
rect 19858 -3427 19910 -3415
rect 19858 -5415 19910 -5403
rect 19976 -3427 20028 -3415
rect 19976 -5415 20028 -5403
rect 20094 -3427 20146 -3415
rect 20094 -5415 20146 -5403
rect 20212 -3427 20264 -3415
rect 20212 -5415 20264 -5403
rect 20330 -3427 20382 -3414
rect 20330 -5415 20382 -5403
rect 20448 -3427 20500 -3415
rect 20448 -5415 20500 -5403
rect 20566 -3427 20618 -3374
rect 21864 -3415 21916 -3374
rect 21981 -3415 22027 -3403
rect 19910 -5456 19976 -5450
rect 20566 -5456 20618 -5403
rect 20684 -3427 20736 -3415
rect 20684 -5415 20736 -5403
rect 20802 -3427 20854 -3415
rect 20802 -5415 20854 -5403
rect 20920 -3427 20972 -3415
rect 20920 -5415 20972 -5403
rect 21038 -3427 21090 -3415
rect 21038 -5415 21090 -5403
rect 21156 -3427 21208 -3415
rect 21156 -5415 21208 -5403
rect 21274 -3427 21326 -3415
rect 21274 -5415 21326 -5403
rect 21392 -3427 21444 -3415
rect 21392 -5415 21444 -5403
rect 21510 -3427 21562 -3415
rect 21510 -5415 21562 -5403
rect 21628 -3427 21680 -3415
rect 21628 -5415 21680 -5403
rect 21746 -3427 21798 -3415
rect 21746 -5415 21798 -5403
rect 21864 -3427 21987 -3415
rect 21916 -3815 21987 -3427
rect 22021 -3815 22027 -3415
rect 21981 -3827 22027 -3815
rect 21981 -5015 22027 -5003
rect 21916 -5403 21987 -5015
rect 21864 -5415 21987 -5403
rect 22021 -5415 22027 -5015
rect 21864 -5456 21916 -5415
rect 21981 -5427 22027 -5415
rect 18088 -5462 18206 -5456
rect 18088 -5496 18156 -5462
rect 18190 -5496 18206 -5462
rect 18088 -5502 18206 -5496
rect 18258 -5462 19504 -5456
rect 18258 -5496 18274 -5462
rect 18308 -5496 18392 -5462
rect 18426 -5496 18510 -5462
rect 18544 -5496 18628 -5462
rect 18662 -5496 18746 -5462
rect 18780 -5496 18864 -5462
rect 18898 -5496 18982 -5462
rect 19016 -5496 19100 -5462
rect 19134 -5496 19218 -5462
rect 19252 -5496 19336 -5462
rect 19370 -5496 19454 -5462
rect 19488 -5496 19504 -5462
rect 18258 -5502 19504 -5496
rect 19556 -5462 19918 -5456
rect 19556 -5496 19572 -5462
rect 19606 -5496 19690 -5462
rect 19724 -5496 19808 -5462
rect 19842 -5496 19918 -5462
rect 19556 -5502 19918 -5496
rect 19910 -5508 19918 -5502
rect 19970 -5508 19976 -5456
rect 20032 -5462 20448 -5456
rect 20032 -5496 20044 -5462
rect 20078 -5496 20162 -5462
rect 20196 -5496 20280 -5462
rect 20314 -5496 20398 -5462
rect 20432 -5496 20448 -5462
rect 20032 -5500 20448 -5496
rect 19910 -5519 19976 -5508
rect 20027 -5552 20033 -5500
rect 20085 -5502 20448 -5500
rect 20500 -5462 21746 -5456
rect 20500 -5496 20516 -5462
rect 20550 -5496 20634 -5462
rect 20668 -5496 20752 -5462
rect 20786 -5496 20870 -5462
rect 20904 -5496 20988 -5462
rect 21022 -5496 21106 -5462
rect 21140 -5496 21224 -5462
rect 21258 -5496 21342 -5462
rect 21376 -5496 21460 -5462
rect 21494 -5496 21578 -5462
rect 21612 -5496 21696 -5462
rect 21730 -5496 21746 -5462
rect 20500 -5502 21746 -5496
rect 21798 -5462 21916 -5456
rect 21798 -5496 21814 -5462
rect 21848 -5496 21916 -5462
rect 21798 -5502 21916 -5496
rect 20085 -5552 20091 -5502
rect 18205 -5742 18257 -5736
rect 18205 -5846 18257 -5794
rect 21746 -5742 21798 -5736
rect 21746 -5846 21798 -5794
rect 17851 -5852 17969 -5846
rect 17851 -5886 17919 -5852
rect 17953 -5886 17969 -5852
rect 17851 -5892 17969 -5886
rect 18021 -5852 18437 -5846
rect 18021 -5886 18037 -5852
rect 18071 -5886 18155 -5852
rect 18189 -5886 18273 -5852
rect 18307 -5886 18391 -5852
rect 18425 -5886 18437 -5852
rect 18021 -5892 18437 -5886
rect 18497 -5852 18611 -5846
rect 18497 -5886 18509 -5852
rect 18543 -5886 18611 -5852
rect 18497 -5892 18611 -5886
rect 17740 -5924 17786 -5912
rect 17851 -5924 17903 -5892
rect 18559 -5924 18611 -5892
rect 21392 -5852 21506 -5846
rect 21392 -5886 21460 -5852
rect 21494 -5886 21506 -5852
rect 21392 -5892 21506 -5886
rect 21566 -5852 21982 -5846
rect 21566 -5886 21578 -5852
rect 21612 -5886 21696 -5852
rect 21730 -5886 21814 -5852
rect 21848 -5886 21932 -5852
rect 21966 -5886 21982 -5852
rect 21566 -5892 21982 -5886
rect 22038 -5852 22152 -5846
rect 22038 -5886 22050 -5852
rect 22084 -5886 22152 -5852
rect 22038 -5892 22152 -5886
rect 18702 -5912 18802 -5900
rect 18676 -5924 18802 -5912
rect 17740 -6324 17746 -5924
rect 17780 -5936 17903 -5924
rect 17780 -6324 17851 -5936
rect 17740 -6336 17786 -6324
rect 17740 -7524 17786 -7512
rect 17740 -7924 17746 -7524
rect 17780 -7912 17851 -7524
rect 17780 -7924 17903 -7912
rect 17969 -5936 18021 -5924
rect 17969 -7924 18021 -7912
rect 18087 -5936 18139 -5924
rect 18087 -7924 18139 -7912
rect 18205 -5936 18257 -5924
rect 18205 -7924 18257 -7912
rect 18323 -5936 18375 -5924
rect 18323 -7924 18375 -7912
rect 18441 -5936 18493 -5924
rect 18441 -7924 18493 -7912
rect 18559 -5936 18682 -5924
rect 18611 -6324 18682 -5936
rect 18716 -6000 18802 -5924
rect 21202 -5912 21302 -5900
rect 21202 -5924 21327 -5912
rect 21392 -5924 21444 -5892
rect 22100 -5924 22152 -5892
rect 22217 -5924 22263 -5912
rect 21202 -6000 21287 -5924
rect 18716 -6100 18962 -6000
rect 19019 -6024 19171 -6018
rect 19019 -6058 19121 -6024
rect 19155 -6058 19171 -6024
rect 19019 -6064 19171 -6058
rect 20833 -6024 20985 -6018
rect 20833 -6058 20849 -6024
rect 20883 -6058 20985 -6024
rect 20833 -6064 20985 -6058
rect 19019 -6100 19065 -6064
rect 19115 -6100 19161 -6064
rect 20843 -6100 20889 -6064
rect 20939 -6100 20985 -6064
rect 21042 -6100 21287 -6000
rect 18716 -6324 18911 -6100
rect 18676 -6336 18911 -6324
rect 18702 -6500 18911 -6336
rect 18802 -6600 18911 -6500
rect 18945 -6600 19015 -6100
rect 19069 -6600 19075 -6100
rect 19105 -6600 19111 -6100
rect 19165 -6600 19171 -6100
rect 19201 -6600 19207 -6100
rect 19261 -6600 19267 -6100
rect 19297 -6600 19303 -6100
rect 19357 -6600 19363 -6100
rect 19393 -6600 19399 -6100
rect 19453 -6600 19459 -6100
rect 19489 -6600 19495 -6100
rect 19549 -6600 19555 -6100
rect 19585 -6600 19591 -6100
rect 19645 -6600 19651 -6100
rect 19681 -6600 19687 -6100
rect 19741 -6600 19747 -6100
rect 19777 -6600 19783 -6100
rect 19837 -6600 19843 -6100
rect 19873 -6600 19879 -6100
rect 19933 -6600 19939 -6100
rect 19969 -6600 19975 -6100
rect 20029 -6600 20035 -6100
rect 20065 -6600 20071 -6100
rect 20125 -6600 20131 -6100
rect 20161 -6600 20167 -6100
rect 20221 -6600 20227 -6100
rect 20257 -6600 20263 -6100
rect 20317 -6600 20323 -6100
rect 20353 -6600 20359 -6100
rect 20413 -6600 20419 -6100
rect 20449 -6600 20455 -6100
rect 20509 -6600 20515 -6100
rect 20545 -6600 20551 -6100
rect 20605 -6600 20611 -6100
rect 20641 -6600 20647 -6100
rect 20701 -6600 20707 -6100
rect 20737 -6600 20743 -6100
rect 20797 -6600 20803 -6100
rect 20833 -6600 20839 -6100
rect 20893 -6600 20899 -6100
rect 20929 -6600 20935 -6100
rect 20989 -6600 21059 -6100
rect 21093 -6324 21287 -6100
rect 21321 -5936 21444 -5924
rect 21321 -6324 21392 -5936
rect 21093 -6336 21327 -6324
rect 21093 -6500 21302 -6336
rect 21093 -6600 21202 -6500
rect 18802 -6900 18962 -6600
rect 19291 -6700 19297 -6644
rect 19363 -6700 19369 -6644
rect 19483 -6700 19489 -6644
rect 19555 -6700 19561 -6644
rect 19675 -6700 19681 -6644
rect 19747 -6700 19753 -6644
rect 19867 -6700 19873 -6644
rect 19939 -6700 19945 -6644
rect 20059 -6700 20065 -6644
rect 20131 -6700 20137 -6644
rect 20251 -6700 20257 -6644
rect 20323 -6700 20329 -6644
rect 20443 -6700 20449 -6644
rect 20515 -6700 20521 -6644
rect 20635 -6700 20641 -6644
rect 20707 -6700 20713 -6644
rect 18802 -7040 19002 -6900
rect 19058 -6938 19122 -6930
rect 19122 -6968 20885 -6962
rect 19122 -7002 19131 -6968
rect 19499 -7002 19589 -6968
rect 19957 -7002 20047 -6968
rect 20415 -7002 20505 -6968
rect 20873 -7002 20885 -6968
rect 19058 -7008 20885 -7002
rect 19058 -7010 19122 -7008
rect 21042 -7028 21202 -6600
rect 21009 -7040 21202 -7028
rect 18802 -7400 18955 -7040
rect 18702 -7440 18955 -7400
rect 18989 -7052 19112 -7040
rect 18989 -7440 19060 -7052
rect 18702 -7500 19002 -7440
rect 18702 -7512 18962 -7500
rect 18676 -7524 18962 -7512
rect 18611 -7912 18682 -7524
rect 18559 -7924 18682 -7912
rect 18716 -7924 18962 -7524
rect 17740 -7936 17786 -7924
rect 17851 -7956 17903 -7924
rect 18559 -7956 18611 -7924
rect 18676 -7936 18962 -7924
rect 17851 -7962 17969 -7956
rect 17851 -7996 17919 -7962
rect 17953 -7996 17969 -7962
rect 17851 -8002 17969 -7996
rect 18021 -7962 18437 -7956
rect 18021 -7996 18037 -7962
rect 18071 -7996 18155 -7962
rect 18189 -7996 18273 -7962
rect 18307 -7996 18391 -7962
rect 18425 -7996 18437 -7962
rect 18021 -8002 18437 -7996
rect 18497 -7962 18611 -7956
rect 18497 -7996 18509 -7962
rect 18543 -7996 18611 -7962
rect 18497 -8002 18611 -7996
rect 18702 -8000 18962 -7936
rect 18802 -8060 18962 -8000
rect 16650 -8398 17258 -8392
rect 16650 -8432 16662 -8398
rect 17138 -8432 17258 -8398
rect 16650 -8438 17258 -8432
rect 16572 -8464 16618 -8448
rect 16572 -8494 16578 -8464
rect 16437 -8498 16578 -8494
rect 16612 -8498 16618 -8464
rect 16437 -8528 16618 -8498
rect 16649 -8494 16666 -8485
rect 17135 -8494 17150 -8485
rect 16649 -8528 16662 -8494
rect 17138 -8528 17150 -8494
rect 16437 -9384 16471 -8528
rect 16649 -8537 16666 -8528
rect 17135 -8537 17150 -8528
rect 17218 -8584 17258 -8438
rect 16650 -8590 17258 -8584
rect 16650 -8624 16662 -8590
rect 17138 -8624 17258 -8590
rect 16650 -8630 17258 -8624
rect 16572 -8656 16618 -8640
rect 16572 -8686 16578 -8656
rect 16431 -9510 16471 -9384
rect 16390 -9520 16471 -9510
rect 16390 -9580 16400 -9520
rect 16460 -9580 16471 -9520
rect 16390 -9584 16471 -9580
rect 16499 -8690 16578 -8686
rect 16612 -8690 16618 -8656
rect 16499 -8720 16618 -8690
rect 16650 -8686 17150 -8680
rect 16650 -8720 16662 -8686
rect 17138 -8720 17150 -8686
rect 16499 -9384 16533 -8720
rect 16650 -8726 17150 -8720
rect 17218 -8776 17258 -8630
rect 16650 -8782 17258 -8776
rect 16650 -8816 16662 -8782
rect 17138 -8816 17258 -8782
rect 16650 -8822 17258 -8816
rect 17380 -8440 17620 -8420
rect 16567 -9170 16590 -9100
rect 17019 -9108 17038 -9100
rect 17022 -9161 17038 -9108
rect 17019 -9170 17038 -9161
rect 17380 -9360 17400 -8440
rect 17600 -9360 17620 -8440
rect 18802 -9280 18822 -8060
rect 18882 -8628 18962 -8060
rect 18882 -8640 18995 -8628
rect 18882 -9040 18955 -8640
rect 18989 -9028 19060 -8640
rect 18989 -9040 19112 -9028
rect 19518 -7052 19570 -7040
rect 19518 -9040 19570 -9028
rect 19976 -7052 20028 -7040
rect 19976 -9040 20028 -9028
rect 20434 -7052 20486 -7040
rect 20434 -9040 20486 -9028
rect 20892 -7052 21015 -7040
rect 20944 -7440 21015 -7052
rect 21049 -7400 21202 -7040
rect 21049 -7440 21302 -7400
rect 21009 -7452 21302 -7440
rect 21042 -7512 21302 -7452
rect 21042 -7524 21327 -7512
rect 21042 -7924 21287 -7524
rect 21321 -7912 21392 -7524
rect 21321 -7924 21444 -7912
rect 21510 -5936 21562 -5924
rect 21510 -7924 21562 -7912
rect 21628 -5936 21680 -5924
rect 21628 -7924 21680 -7912
rect 21746 -5936 21798 -5924
rect 21746 -7924 21798 -7912
rect 21864 -5936 21916 -5924
rect 21864 -7924 21916 -7912
rect 21982 -5936 22034 -5924
rect 21982 -7924 22034 -7912
rect 22100 -5936 22223 -5924
rect 22152 -6324 22223 -5936
rect 22257 -6324 22263 -5924
rect 22217 -6336 22263 -6324
rect 22452 -6270 22602 -6250
rect 22452 -6660 22472 -6270
rect 22582 -6660 22602 -6270
rect 22452 -6680 22602 -6660
rect 22682 -6270 22832 -6250
rect 22682 -6660 22702 -6270
rect 22812 -6660 22832 -6270
rect 22682 -6680 22832 -6660
rect 23200 -7322 23300 -7200
rect 23156 -7353 23300 -7322
rect 23500 -7322 23600 -7200
rect 23500 -7353 23800 -7322
rect 23156 -7387 23185 -7353
rect 23219 -7387 23277 -7353
rect 23500 -7387 23553 -7353
rect 23587 -7387 23645 -7353
rect 23679 -7387 23737 -7353
rect 23771 -7387 23800 -7353
rect 23156 -7400 23300 -7387
rect 23500 -7400 23800 -7387
rect 23156 -7418 23800 -7400
rect 22217 -7524 22263 -7512
rect 22152 -7912 22223 -7524
rect 22100 -7924 22223 -7912
rect 22257 -7924 22263 -7524
rect 23260 -7720 23270 -7640
rect 23410 -7720 23420 -7640
rect 23540 -7720 23550 -7640
rect 23690 -7720 23700 -7640
rect 21042 -7936 21327 -7924
rect 21042 -8000 21302 -7936
rect 21392 -7956 21444 -7924
rect 22100 -7956 22152 -7924
rect 22217 -7936 22263 -7924
rect 23156 -7897 23800 -7866
rect 23156 -7931 23185 -7897
rect 23219 -7931 23277 -7897
rect 23311 -7900 23369 -7897
rect 23403 -7900 23461 -7897
rect 23495 -7900 23553 -7897
rect 23500 -7931 23553 -7900
rect 23587 -7931 23645 -7897
rect 23679 -7931 23737 -7897
rect 23771 -7931 23800 -7897
rect 21392 -7962 21506 -7956
rect 21392 -7996 21460 -7962
rect 21494 -7996 21506 -7962
rect 21042 -8060 21202 -8000
rect 21392 -8002 21506 -7996
rect 21566 -7962 21982 -7956
rect 21566 -7996 21578 -7962
rect 21612 -7996 21696 -7962
rect 21730 -7996 21814 -7962
rect 21848 -7996 21932 -7962
rect 21966 -7996 21982 -7962
rect 21566 -8002 21982 -7996
rect 22038 -7962 22152 -7956
rect 23156 -7962 23300 -7931
rect 22038 -7996 22050 -7962
rect 22084 -7996 22152 -7962
rect 22038 -8002 22152 -7996
rect 21042 -8628 21122 -8060
rect 21009 -8640 21122 -8628
rect 20944 -9028 21015 -8640
rect 20892 -9040 21015 -9028
rect 21049 -9040 21122 -8640
rect 18882 -9052 18995 -9040
rect 21009 -9052 21122 -9040
rect 18882 -9280 18962 -9052
rect 19119 -9078 20885 -9072
rect 19119 -9112 19131 -9078
rect 19499 -9112 19589 -9078
rect 19957 -9112 20047 -9078
rect 20415 -9112 20505 -9078
rect 20873 -9112 20885 -9078
rect 19119 -9118 20885 -9112
rect 18802 -9300 18962 -9280
rect 21042 -9280 21122 -9052
rect 21182 -9280 21202 -8060
rect 23200 -8100 23300 -7962
rect 23500 -7962 23800 -7931
rect 23500 -8100 23600 -7962
rect 21042 -9300 21202 -9280
rect 17380 -9380 17620 -9360
rect 16499 -9550 16539 -9384
rect 16499 -9584 16540 -9550
rect 16390 -9590 16470 -9584
rect 16500 -9650 16540 -9584
rect 16460 -9660 16540 -9650
rect 16460 -9720 16470 -9660
rect 16530 -9720 16540 -9660
rect 16460 -9730 16540 -9720
rect 16780 -10500 16876 -10494
rect 16700 -10510 16876 -10500
rect 16700 -10850 16710 -10510
rect 16800 -10523 16876 -10510
rect 16800 -10557 16811 -10523
rect 16845 -10557 16876 -10523
rect 16800 -10615 16876 -10557
rect 17324 -10500 17420 -10494
rect 17324 -10510 17520 -10500
rect 17324 -10523 17420 -10510
rect 17324 -10557 17355 -10523
rect 17389 -10557 17420 -10523
rect 17111 -10610 17169 -10603
rect 16800 -10649 16811 -10615
rect 16845 -10649 16876 -10615
rect 16800 -10707 16876 -10649
rect 16800 -10741 16811 -10707
rect 16845 -10741 16876 -10707
rect 16800 -10799 16876 -10741
rect 17020 -10618 17169 -10610
rect 17020 -10620 17120 -10618
rect 17020 -10740 17030 -10620
rect 17160 -10738 17169 -10618
rect 17130 -10740 17169 -10738
rect 17020 -10750 17169 -10740
rect 17111 -10753 17169 -10750
rect 17324 -10615 17420 -10557
rect 17324 -10649 17355 -10615
rect 17389 -10649 17420 -10615
rect 17324 -10707 17420 -10649
rect 17324 -10741 17355 -10707
rect 17389 -10741 17420 -10707
rect 16800 -10833 16811 -10799
rect 16845 -10833 16876 -10799
rect 16800 -10850 16876 -10833
rect 16700 -10860 16876 -10850
rect 16780 -10862 16876 -10860
rect 17324 -10799 17420 -10741
rect 17324 -10833 17355 -10799
rect 17389 -10833 17420 -10799
rect 17324 -10850 17420 -10833
rect 17510 -10850 17520 -10510
rect 17324 -10860 17520 -10850
rect 17324 -10862 17420 -10860
rect 6000 -11248 14000 -11000
rect 6000 -11300 6614 -11248
rect 6666 -11300 6934 -11248
rect 6986 -11300 7254 -11248
rect 7306 -11300 7574 -11248
rect 7626 -11300 7894 -11248
rect 7946 -11300 8214 -11248
rect 8266 -11300 8534 -11248
rect 8586 -11300 8854 -11248
rect 8906 -11300 9174 -11248
rect 9226 -11300 9494 -11248
rect 9546 -11300 9814 -11248
rect 9866 -11300 10134 -11248
rect 10186 -11300 10454 -11248
rect 10506 -11300 10774 -11248
rect 10826 -11300 11094 -11248
rect 11146 -11300 11414 -11248
rect 11466 -11300 11734 -11248
rect 11786 -11300 12054 -11248
rect 12106 -11300 12374 -11248
rect 12426 -11300 12694 -11248
rect 12746 -11300 13014 -11248
rect 13066 -11300 13334 -11248
rect 13386 -11300 14000 -11248
rect 6000 -11454 14000 -11300
rect 6000 -11506 6244 -11454
rect 6296 -11506 13710 -11454
rect 13762 -11506 14000 -11454
rect 6000 -11540 14000 -11506
rect 6000 -11774 6540 -11540
rect 6000 -11826 6244 -11774
rect 6296 -11826 6540 -11774
rect 6000 -12094 6540 -11826
rect 6000 -12146 6244 -12094
rect 6296 -12146 6540 -12094
rect 6000 -12414 6540 -12146
rect 6000 -12466 6244 -12414
rect 6296 -12466 6540 -12414
rect 6000 -12734 6540 -12466
rect 6000 -12786 6244 -12734
rect 6296 -12786 6540 -12734
rect 6000 -13054 6540 -12786
rect 6000 -13106 6244 -13054
rect 6296 -13106 6540 -13054
rect 6000 -13374 6540 -13106
rect 6000 -13426 6244 -13374
rect 6296 -13426 6540 -13374
rect 6000 -13694 6540 -13426
rect 6000 -13746 6244 -13694
rect 6296 -13746 6540 -13694
rect 6000 -14014 6540 -13746
rect 6000 -14066 6244 -14014
rect 6296 -14066 6540 -14014
rect 6000 -14334 6540 -14066
rect 6000 -14386 6244 -14334
rect 6296 -14386 6540 -14334
rect 6000 -14654 6540 -14386
rect 6000 -14706 6244 -14654
rect 6296 -14706 6540 -14654
rect 6000 -14974 6540 -14706
rect 6000 -15026 6244 -14974
rect 6296 -15026 6540 -14974
rect 6000 -15294 6540 -15026
rect 6000 -15346 6244 -15294
rect 6296 -15346 6540 -15294
rect 6000 -15614 6540 -15346
rect 6000 -15666 6244 -15614
rect 6296 -15666 6540 -15614
rect 6000 -15934 6540 -15666
rect 6000 -15986 6244 -15934
rect 6296 -15986 6540 -15934
rect 6000 -16254 6540 -15986
rect 6000 -16306 6244 -16254
rect 6296 -16306 6540 -16254
rect 6000 -16574 6540 -16306
rect 6000 -16626 6244 -16574
rect 6296 -16626 6540 -16574
rect 6000 -16894 6540 -16626
rect 6000 -16946 6244 -16894
rect 6296 -16946 6540 -16894
rect 6000 -17214 6540 -16946
rect 6000 -17266 6244 -17214
rect 6296 -17266 6540 -17214
rect 6000 -17534 6540 -17266
rect 6000 -17586 6244 -17534
rect 6296 -17586 6540 -17534
rect 6000 -17854 6540 -17586
rect 6000 -17906 6244 -17854
rect 6296 -17906 6540 -17854
rect 6000 -18174 6540 -17906
rect 6000 -18226 6244 -18174
rect 6296 -18226 6540 -18174
rect 6000 -18460 6540 -18226
rect 13460 -11774 14000 -11540
rect 13460 -11826 13710 -11774
rect 13762 -11826 14000 -11774
rect 13460 -12094 14000 -11826
rect 13460 -12146 13710 -12094
rect 13762 -12146 14000 -12094
rect 13460 -12414 14000 -12146
rect 13460 -12466 13710 -12414
rect 13762 -12466 14000 -12414
rect 13460 -12734 14000 -12466
rect 13460 -12786 13710 -12734
rect 13762 -12786 14000 -12734
rect 13460 -13054 14000 -12786
rect 13460 -13106 13710 -13054
rect 13762 -13106 14000 -13054
rect 13460 -13374 14000 -13106
rect 13460 -13426 13710 -13374
rect 13762 -13426 14000 -13374
rect 13460 -13694 14000 -13426
rect 13460 -13746 13710 -13694
rect 13762 -13746 14000 -13694
rect 13460 -14014 14000 -13746
rect 13460 -14066 13710 -14014
rect 13762 -14066 14000 -14014
rect 13460 -14334 14000 -14066
rect 13460 -14386 13710 -14334
rect 13762 -14386 14000 -14334
rect 13460 -14654 14000 -14386
rect 13460 -14706 13710 -14654
rect 13762 -14706 14000 -14654
rect 13460 -14974 14000 -14706
rect 13460 -15026 13710 -14974
rect 13762 -15026 14000 -14974
rect 13460 -15294 14000 -15026
rect 13460 -15346 13710 -15294
rect 13762 -15346 14000 -15294
rect 13460 -15614 14000 -15346
rect 13460 -15666 13710 -15614
rect 13762 -15666 14000 -15614
rect 13460 -15934 14000 -15666
rect 13460 -15986 13710 -15934
rect 13762 -15986 14000 -15934
rect 13460 -16254 14000 -15986
rect 13460 -16306 13710 -16254
rect 13762 -16306 14000 -16254
rect 13460 -16574 14000 -16306
rect 13460 -16626 13710 -16574
rect 13762 -16626 14000 -16574
rect 13460 -16894 14000 -16626
rect 13460 -16946 13710 -16894
rect 13762 -16946 14000 -16894
rect 13460 -17214 14000 -16946
rect 13460 -17266 13710 -17214
rect 13762 -17266 14000 -17214
rect 13460 -17534 14000 -17266
rect 13460 -17586 13710 -17534
rect 13762 -17586 14000 -17534
rect 13460 -17854 14000 -17586
rect 13460 -17906 13710 -17854
rect 13762 -17906 14000 -17854
rect 13460 -18174 14000 -17906
rect 13460 -18226 13710 -18174
rect 13762 -18226 14000 -18174
rect 13460 -18460 14000 -18226
rect 6000 -18494 14000 -18460
rect 6000 -18546 6244 -18494
rect 6296 -18546 13710 -18494
rect 13762 -18546 14000 -18494
rect 6000 -18704 14000 -18546
rect 6000 -18756 6614 -18704
rect 6666 -18756 6934 -18704
rect 6986 -18756 7254 -18704
rect 7306 -18756 7574 -18704
rect 7626 -18756 7894 -18704
rect 7946 -18756 8214 -18704
rect 8266 -18756 8534 -18704
rect 8586 -18756 8854 -18704
rect 8906 -18756 9174 -18704
rect 9226 -18756 9494 -18704
rect 9546 -18756 9814 -18704
rect 9866 -18756 10134 -18704
rect 10186 -18756 10454 -18704
rect 10506 -18756 10774 -18704
rect 10826 -18756 11094 -18704
rect 11146 -18756 11414 -18704
rect 11466 -18756 11734 -18704
rect 11786 -18756 12054 -18704
rect 12106 -18756 12374 -18704
rect 12426 -18756 12694 -18704
rect 12746 -18756 13014 -18704
rect 13066 -18756 13334 -18704
rect 13386 -18756 14000 -18704
rect 6000 -19000 14000 -18756
rect 18000 -11248 26000 -11000
rect 18000 -11300 18614 -11248
rect 18666 -11300 18934 -11248
rect 18986 -11300 19254 -11248
rect 19306 -11300 19574 -11248
rect 19626 -11300 19894 -11248
rect 19946 -11300 20214 -11248
rect 20266 -11300 20534 -11248
rect 20586 -11300 20854 -11248
rect 20906 -11300 21174 -11248
rect 21226 -11300 21494 -11248
rect 21546 -11300 21814 -11248
rect 21866 -11300 22134 -11248
rect 22186 -11300 22454 -11248
rect 22506 -11300 22774 -11248
rect 22826 -11300 23094 -11248
rect 23146 -11300 23414 -11248
rect 23466 -11300 23734 -11248
rect 23786 -11300 24054 -11248
rect 24106 -11300 24374 -11248
rect 24426 -11300 24694 -11248
rect 24746 -11300 25014 -11248
rect 25066 -11300 25334 -11248
rect 25386 -11300 26000 -11248
rect 18000 -11454 26000 -11300
rect 18000 -11506 18244 -11454
rect 18296 -11506 25710 -11454
rect 25762 -11506 26000 -11454
rect 18000 -11540 26000 -11506
rect 18000 -11774 18540 -11540
rect 18000 -11826 18244 -11774
rect 18296 -11826 18540 -11774
rect 18000 -12094 18540 -11826
rect 18000 -12146 18244 -12094
rect 18296 -12146 18540 -12094
rect 18000 -12414 18540 -12146
rect 18000 -12466 18244 -12414
rect 18296 -12466 18540 -12414
rect 18000 -12734 18540 -12466
rect 18000 -12786 18244 -12734
rect 18296 -12786 18540 -12734
rect 18000 -13054 18540 -12786
rect 18000 -13106 18244 -13054
rect 18296 -13106 18540 -13054
rect 18000 -13374 18540 -13106
rect 18000 -13426 18244 -13374
rect 18296 -13426 18540 -13374
rect 18000 -13694 18540 -13426
rect 18000 -13746 18244 -13694
rect 18296 -13746 18540 -13694
rect 18000 -14014 18540 -13746
rect 18000 -14066 18244 -14014
rect 18296 -14066 18540 -14014
rect 18000 -14334 18540 -14066
rect 18000 -14386 18244 -14334
rect 18296 -14386 18540 -14334
rect 18000 -14654 18540 -14386
rect 18000 -14706 18244 -14654
rect 18296 -14706 18540 -14654
rect 18000 -14974 18540 -14706
rect 18000 -15026 18244 -14974
rect 18296 -15026 18540 -14974
rect 18000 -15294 18540 -15026
rect 18000 -15346 18244 -15294
rect 18296 -15346 18540 -15294
rect 18000 -15614 18540 -15346
rect 18000 -15666 18244 -15614
rect 18296 -15666 18540 -15614
rect 18000 -15934 18540 -15666
rect 18000 -15986 18244 -15934
rect 18296 -15986 18540 -15934
rect 18000 -16254 18540 -15986
rect 18000 -16306 18244 -16254
rect 18296 -16306 18540 -16254
rect 18000 -16574 18540 -16306
rect 18000 -16626 18244 -16574
rect 18296 -16626 18540 -16574
rect 18000 -16894 18540 -16626
rect 18000 -16946 18244 -16894
rect 18296 -16946 18540 -16894
rect 18000 -17214 18540 -16946
rect 18000 -17266 18244 -17214
rect 18296 -17266 18540 -17214
rect 18000 -17534 18540 -17266
rect 18000 -17586 18244 -17534
rect 18296 -17586 18540 -17534
rect 18000 -17854 18540 -17586
rect 18000 -17906 18244 -17854
rect 18296 -17906 18540 -17854
rect 18000 -18174 18540 -17906
rect 18000 -18226 18244 -18174
rect 18296 -18226 18540 -18174
rect 18000 -18460 18540 -18226
rect 25460 -11774 26000 -11540
rect 25460 -11826 25710 -11774
rect 25762 -11826 26000 -11774
rect 25460 -12094 26000 -11826
rect 25460 -12146 25710 -12094
rect 25762 -12146 26000 -12094
rect 25460 -12414 26000 -12146
rect 25460 -12466 25710 -12414
rect 25762 -12466 26000 -12414
rect 25460 -12734 26000 -12466
rect 25460 -12786 25710 -12734
rect 25762 -12786 26000 -12734
rect 25460 -13054 26000 -12786
rect 25460 -13106 25710 -13054
rect 25762 -13106 26000 -13054
rect 25460 -13374 26000 -13106
rect 25460 -13426 25710 -13374
rect 25762 -13426 26000 -13374
rect 25460 -13694 26000 -13426
rect 25460 -13746 25710 -13694
rect 25762 -13746 26000 -13694
rect 25460 -14014 26000 -13746
rect 25460 -14066 25710 -14014
rect 25762 -14066 26000 -14014
rect 25460 -14334 26000 -14066
rect 25460 -14386 25710 -14334
rect 25762 -14386 26000 -14334
rect 25460 -14654 26000 -14386
rect 25460 -14706 25710 -14654
rect 25762 -14706 26000 -14654
rect 25460 -14974 26000 -14706
rect 25460 -15026 25710 -14974
rect 25762 -15026 26000 -14974
rect 25460 -15294 26000 -15026
rect 25460 -15346 25710 -15294
rect 25762 -15346 26000 -15294
rect 25460 -15614 26000 -15346
rect 25460 -15666 25710 -15614
rect 25762 -15666 26000 -15614
rect 25460 -15934 26000 -15666
rect 25460 -15986 25710 -15934
rect 25762 -15986 26000 -15934
rect 25460 -16254 26000 -15986
rect 25460 -16306 25710 -16254
rect 25762 -16306 26000 -16254
rect 25460 -16574 26000 -16306
rect 25460 -16626 25710 -16574
rect 25762 -16626 26000 -16574
rect 25460 -16894 26000 -16626
rect 25460 -16946 25710 -16894
rect 25762 -16946 26000 -16894
rect 25460 -17214 26000 -16946
rect 25460 -17266 25710 -17214
rect 25762 -17266 26000 -17214
rect 25460 -17534 26000 -17266
rect 25460 -17586 25710 -17534
rect 25762 -17586 26000 -17534
rect 25460 -17854 26000 -17586
rect 25460 -17906 25710 -17854
rect 25762 -17906 26000 -17854
rect 25460 -18174 26000 -17906
rect 25460 -18226 25710 -18174
rect 25762 -18226 26000 -18174
rect 25460 -18460 26000 -18226
rect 18000 -18494 26000 -18460
rect 18000 -18546 18244 -18494
rect 18296 -18546 25710 -18494
rect 25762 -18546 26000 -18494
rect 18000 -18704 26000 -18546
rect 18000 -18756 18614 -18704
rect 18666 -18756 18934 -18704
rect 18986 -18756 19254 -18704
rect 19306 -18756 19574 -18704
rect 19626 -18756 19894 -18704
rect 19946 -18756 20214 -18704
rect 20266 -18756 20534 -18704
rect 20586 -18756 20854 -18704
rect 20906 -18756 21174 -18704
rect 21226 -18756 21494 -18704
rect 21546 -18756 21814 -18704
rect 21866 -18756 22134 -18704
rect 22186 -18756 22454 -18704
rect 22506 -18756 22774 -18704
rect 22826 -18756 23094 -18704
rect 23146 -18756 23414 -18704
rect 23466 -18756 23734 -18704
rect 23786 -18756 24054 -18704
rect 24106 -18756 24374 -18704
rect 24426 -18756 24694 -18704
rect 24746 -18756 25014 -18704
rect 25066 -18756 25334 -18704
rect 25386 -18756 26000 -18704
rect 18000 -19000 26000 -18756
rect 30000 -11248 38000 -11000
rect 30000 -11300 30614 -11248
rect 30666 -11300 30934 -11248
rect 30986 -11300 31254 -11248
rect 31306 -11300 31574 -11248
rect 31626 -11300 31894 -11248
rect 31946 -11300 32214 -11248
rect 32266 -11300 32534 -11248
rect 32586 -11300 32854 -11248
rect 32906 -11300 33174 -11248
rect 33226 -11300 33494 -11248
rect 33546 -11300 33814 -11248
rect 33866 -11300 34134 -11248
rect 34186 -11300 34454 -11248
rect 34506 -11300 34774 -11248
rect 34826 -11300 35094 -11248
rect 35146 -11300 35414 -11248
rect 35466 -11300 35734 -11248
rect 35786 -11300 36054 -11248
rect 36106 -11300 36374 -11248
rect 36426 -11300 36694 -11248
rect 36746 -11300 37014 -11248
rect 37066 -11300 37334 -11248
rect 37386 -11300 38000 -11248
rect 30000 -11454 38000 -11300
rect 30000 -11506 30244 -11454
rect 30296 -11506 37710 -11454
rect 37762 -11506 38000 -11454
rect 30000 -11540 38000 -11506
rect 30000 -11774 30540 -11540
rect 30000 -11826 30244 -11774
rect 30296 -11826 30540 -11774
rect 30000 -12094 30540 -11826
rect 30000 -12146 30244 -12094
rect 30296 -12146 30540 -12094
rect 30000 -12414 30540 -12146
rect 30000 -12466 30244 -12414
rect 30296 -12466 30540 -12414
rect 30000 -12734 30540 -12466
rect 30000 -12786 30244 -12734
rect 30296 -12786 30540 -12734
rect 30000 -13054 30540 -12786
rect 30000 -13106 30244 -13054
rect 30296 -13106 30540 -13054
rect 30000 -13374 30540 -13106
rect 30000 -13426 30244 -13374
rect 30296 -13426 30540 -13374
rect 30000 -13694 30540 -13426
rect 30000 -13746 30244 -13694
rect 30296 -13746 30540 -13694
rect 30000 -14014 30540 -13746
rect 30000 -14066 30244 -14014
rect 30296 -14066 30540 -14014
rect 30000 -14334 30540 -14066
rect 30000 -14386 30244 -14334
rect 30296 -14386 30540 -14334
rect 30000 -14654 30540 -14386
rect 30000 -14706 30244 -14654
rect 30296 -14706 30540 -14654
rect 30000 -14974 30540 -14706
rect 30000 -15026 30244 -14974
rect 30296 -15026 30540 -14974
rect 30000 -15294 30540 -15026
rect 30000 -15346 30244 -15294
rect 30296 -15346 30540 -15294
rect 30000 -15614 30540 -15346
rect 30000 -15666 30244 -15614
rect 30296 -15666 30540 -15614
rect 30000 -15934 30540 -15666
rect 30000 -15986 30244 -15934
rect 30296 -15986 30540 -15934
rect 30000 -16254 30540 -15986
rect 30000 -16306 30244 -16254
rect 30296 -16306 30540 -16254
rect 30000 -16574 30540 -16306
rect 30000 -16626 30244 -16574
rect 30296 -16626 30540 -16574
rect 30000 -16894 30540 -16626
rect 30000 -16946 30244 -16894
rect 30296 -16946 30540 -16894
rect 30000 -17214 30540 -16946
rect 30000 -17266 30244 -17214
rect 30296 -17266 30540 -17214
rect 30000 -17534 30540 -17266
rect 30000 -17586 30244 -17534
rect 30296 -17586 30540 -17534
rect 30000 -17854 30540 -17586
rect 30000 -17906 30244 -17854
rect 30296 -17906 30540 -17854
rect 30000 -18174 30540 -17906
rect 30000 -18226 30244 -18174
rect 30296 -18226 30540 -18174
rect 30000 -18460 30540 -18226
rect 37460 -11774 38000 -11540
rect 37460 -11826 37710 -11774
rect 37762 -11826 38000 -11774
rect 37460 -12094 38000 -11826
rect 37460 -12146 37710 -12094
rect 37762 -12146 38000 -12094
rect 37460 -12414 38000 -12146
rect 37460 -12466 37710 -12414
rect 37762 -12466 38000 -12414
rect 37460 -12734 38000 -12466
rect 37460 -12786 37710 -12734
rect 37762 -12786 38000 -12734
rect 37460 -13054 38000 -12786
rect 37460 -13106 37710 -13054
rect 37762 -13106 38000 -13054
rect 37460 -13374 38000 -13106
rect 37460 -13426 37710 -13374
rect 37762 -13426 38000 -13374
rect 37460 -13694 38000 -13426
rect 37460 -13746 37710 -13694
rect 37762 -13746 38000 -13694
rect 37460 -14014 38000 -13746
rect 37460 -14066 37710 -14014
rect 37762 -14066 38000 -14014
rect 37460 -14334 38000 -14066
rect 37460 -14386 37710 -14334
rect 37762 -14386 38000 -14334
rect 37460 -14654 38000 -14386
rect 37460 -14706 37710 -14654
rect 37762 -14706 38000 -14654
rect 37460 -14974 38000 -14706
rect 37460 -15026 37710 -14974
rect 37762 -15026 38000 -14974
rect 37460 -15294 38000 -15026
rect 37460 -15346 37710 -15294
rect 37762 -15346 38000 -15294
rect 37460 -15614 38000 -15346
rect 37460 -15666 37710 -15614
rect 37762 -15666 38000 -15614
rect 37460 -15934 38000 -15666
rect 37460 -15986 37710 -15934
rect 37762 -15986 38000 -15934
rect 37460 -16254 38000 -15986
rect 37460 -16306 37710 -16254
rect 37762 -16306 38000 -16254
rect 37460 -16574 38000 -16306
rect 37460 -16626 37710 -16574
rect 37762 -16626 38000 -16574
rect 37460 -16894 38000 -16626
rect 37460 -16946 37710 -16894
rect 37762 -16946 38000 -16894
rect 37460 -17214 38000 -16946
rect 37460 -17266 37710 -17214
rect 37762 -17266 38000 -17214
rect 37460 -17534 38000 -17266
rect 37460 -17586 37710 -17534
rect 37762 -17586 38000 -17534
rect 37460 -17854 38000 -17586
rect 37460 -17906 37710 -17854
rect 37762 -17906 38000 -17854
rect 37460 -18174 38000 -17906
rect 37460 -18226 37710 -18174
rect 37762 -18226 38000 -18174
rect 37460 -18460 38000 -18226
rect 30000 -18494 38000 -18460
rect 30000 -18546 30244 -18494
rect 30296 -18546 37710 -18494
rect 37762 -18546 38000 -18494
rect 30000 -18704 38000 -18546
rect 30000 -18756 30614 -18704
rect 30666 -18756 30934 -18704
rect 30986 -18756 31254 -18704
rect 31306 -18756 31574 -18704
rect 31626 -18756 31894 -18704
rect 31946 -18756 32214 -18704
rect 32266 -18756 32534 -18704
rect 32586 -18756 32854 -18704
rect 32906 -18756 33174 -18704
rect 33226 -18756 33494 -18704
rect 33546 -18756 33814 -18704
rect 33866 -18756 34134 -18704
rect 34186 -18756 34454 -18704
rect 34506 -18756 34774 -18704
rect 34826 -18756 35094 -18704
rect 35146 -18756 35414 -18704
rect 35466 -18756 35734 -18704
rect 35786 -18756 36054 -18704
rect 36106 -18756 36374 -18704
rect 36426 -18756 36694 -18704
rect 36746 -18756 37014 -18704
rect 37066 -18756 37334 -18704
rect 37386 -18756 38000 -18704
rect 30000 -19000 38000 -18756
rect 42000 -11248 50000 -11000
rect 42000 -11300 42614 -11248
rect 42666 -11300 42934 -11248
rect 42986 -11300 43254 -11248
rect 43306 -11300 43574 -11248
rect 43626 -11300 43894 -11248
rect 43946 -11300 44214 -11248
rect 44266 -11300 44534 -11248
rect 44586 -11300 44854 -11248
rect 44906 -11300 45174 -11248
rect 45226 -11300 45494 -11248
rect 45546 -11300 45814 -11248
rect 45866 -11300 46134 -11248
rect 46186 -11300 46454 -11248
rect 46506 -11300 46774 -11248
rect 46826 -11300 47094 -11248
rect 47146 -11300 47414 -11248
rect 47466 -11300 47734 -11248
rect 47786 -11300 48054 -11248
rect 48106 -11300 48374 -11248
rect 48426 -11300 48694 -11248
rect 48746 -11300 49014 -11248
rect 49066 -11300 49334 -11248
rect 49386 -11300 50000 -11248
rect 42000 -11454 50000 -11300
rect 42000 -11506 42244 -11454
rect 42296 -11506 49710 -11454
rect 49762 -11506 50000 -11454
rect 42000 -11540 50000 -11506
rect 42000 -11774 42540 -11540
rect 42000 -11826 42244 -11774
rect 42296 -11826 42540 -11774
rect 42000 -12094 42540 -11826
rect 42000 -12146 42244 -12094
rect 42296 -12146 42540 -12094
rect 42000 -12414 42540 -12146
rect 42000 -12466 42244 -12414
rect 42296 -12466 42540 -12414
rect 42000 -12734 42540 -12466
rect 42000 -12786 42244 -12734
rect 42296 -12786 42540 -12734
rect 42000 -13054 42540 -12786
rect 42000 -13106 42244 -13054
rect 42296 -13106 42540 -13054
rect 42000 -13374 42540 -13106
rect 42000 -13426 42244 -13374
rect 42296 -13426 42540 -13374
rect 42000 -13694 42540 -13426
rect 42000 -13746 42244 -13694
rect 42296 -13746 42540 -13694
rect 42000 -14014 42540 -13746
rect 42000 -14066 42244 -14014
rect 42296 -14066 42540 -14014
rect 42000 -14334 42540 -14066
rect 42000 -14386 42244 -14334
rect 42296 -14386 42540 -14334
rect 42000 -14654 42540 -14386
rect 42000 -14706 42244 -14654
rect 42296 -14706 42540 -14654
rect 42000 -14974 42540 -14706
rect 42000 -15026 42244 -14974
rect 42296 -15026 42540 -14974
rect 42000 -15294 42540 -15026
rect 42000 -15346 42244 -15294
rect 42296 -15346 42540 -15294
rect 42000 -15614 42540 -15346
rect 42000 -15666 42244 -15614
rect 42296 -15666 42540 -15614
rect 42000 -15934 42540 -15666
rect 42000 -15986 42244 -15934
rect 42296 -15986 42540 -15934
rect 42000 -16254 42540 -15986
rect 42000 -16306 42244 -16254
rect 42296 -16306 42540 -16254
rect 42000 -16574 42540 -16306
rect 42000 -16626 42244 -16574
rect 42296 -16626 42540 -16574
rect 42000 -16894 42540 -16626
rect 42000 -16946 42244 -16894
rect 42296 -16946 42540 -16894
rect 42000 -17214 42540 -16946
rect 42000 -17266 42244 -17214
rect 42296 -17266 42540 -17214
rect 42000 -17534 42540 -17266
rect 42000 -17586 42244 -17534
rect 42296 -17586 42540 -17534
rect 42000 -17854 42540 -17586
rect 42000 -17906 42244 -17854
rect 42296 -17906 42540 -17854
rect 42000 -18174 42540 -17906
rect 42000 -18226 42244 -18174
rect 42296 -18226 42540 -18174
rect 42000 -18460 42540 -18226
rect 49460 -11774 50000 -11540
rect 49460 -11826 49710 -11774
rect 49762 -11826 50000 -11774
rect 49460 -12094 50000 -11826
rect 49460 -12146 49710 -12094
rect 49762 -12146 50000 -12094
rect 49460 -12414 50000 -12146
rect 49460 -12466 49710 -12414
rect 49762 -12466 50000 -12414
rect 49460 -12734 50000 -12466
rect 49460 -12786 49710 -12734
rect 49762 -12786 50000 -12734
rect 49460 -13054 50000 -12786
rect 49460 -13106 49710 -13054
rect 49762 -13106 50000 -13054
rect 49460 -13374 50000 -13106
rect 49460 -13426 49710 -13374
rect 49762 -13426 50000 -13374
rect 49460 -13694 50000 -13426
rect 49460 -13746 49710 -13694
rect 49762 -13746 50000 -13694
rect 49460 -14014 50000 -13746
rect 49460 -14066 49710 -14014
rect 49762 -14066 50000 -14014
rect 49460 -14334 50000 -14066
rect 49460 -14386 49710 -14334
rect 49762 -14386 50000 -14334
rect 49460 -14654 50000 -14386
rect 49460 -14706 49710 -14654
rect 49762 -14706 50000 -14654
rect 49460 -14974 50000 -14706
rect 49460 -15026 49710 -14974
rect 49762 -15026 50000 -14974
rect 49460 -15294 50000 -15026
rect 49460 -15346 49710 -15294
rect 49762 -15346 50000 -15294
rect 49460 -15614 50000 -15346
rect 49460 -15666 49710 -15614
rect 49762 -15666 50000 -15614
rect 49460 -15934 50000 -15666
rect 49460 -15986 49710 -15934
rect 49762 -15986 50000 -15934
rect 49460 -16254 50000 -15986
rect 49460 -16306 49710 -16254
rect 49762 -16306 50000 -16254
rect 49460 -16574 50000 -16306
rect 49460 -16626 49710 -16574
rect 49762 -16626 50000 -16574
rect 49460 -16894 50000 -16626
rect 49460 -16946 49710 -16894
rect 49762 -16946 50000 -16894
rect 49460 -17214 50000 -16946
rect 49460 -17266 49710 -17214
rect 49762 -17266 50000 -17214
rect 49460 -17534 50000 -17266
rect 49460 -17586 49710 -17534
rect 49762 -17586 50000 -17534
rect 49460 -17854 50000 -17586
rect 49460 -17906 49710 -17854
rect 49762 -17906 50000 -17854
rect 49460 -18174 50000 -17906
rect 49460 -18226 49710 -18174
rect 49762 -18226 50000 -18174
rect 49460 -18460 50000 -18226
rect 42000 -18494 50000 -18460
rect 42000 -18546 42244 -18494
rect 42296 -18546 49710 -18494
rect 49762 -18546 50000 -18494
rect 42000 -18704 50000 -18546
rect 42000 -18756 42614 -18704
rect 42666 -18756 42934 -18704
rect 42986 -18756 43254 -18704
rect 43306 -18756 43574 -18704
rect 43626 -18756 43894 -18704
rect 43946 -18756 44214 -18704
rect 44266 -18756 44534 -18704
rect 44586 -18756 44854 -18704
rect 44906 -18756 45174 -18704
rect 45226 -18756 45494 -18704
rect 45546 -18756 45814 -18704
rect 45866 -18756 46134 -18704
rect 46186 -18756 46454 -18704
rect 46506 -18756 46774 -18704
rect 46826 -18756 47094 -18704
rect 47146 -18756 47414 -18704
rect 47466 -18756 47734 -18704
rect 47786 -18756 48054 -18704
rect 48106 -18756 48374 -18704
rect 48426 -18756 48694 -18704
rect 48746 -18756 49014 -18704
rect 49066 -18756 49334 -18704
rect 49386 -18756 50000 -18704
rect 42000 -19000 50000 -18756
rect 6000 -23248 14000 -23000
rect 6000 -23300 6614 -23248
rect 6666 -23300 6934 -23248
rect 6986 -23300 7254 -23248
rect 7306 -23300 7574 -23248
rect 7626 -23300 7894 -23248
rect 7946 -23300 8214 -23248
rect 8266 -23300 8534 -23248
rect 8586 -23300 8854 -23248
rect 8906 -23300 9174 -23248
rect 9226 -23300 9494 -23248
rect 9546 -23300 9814 -23248
rect 9866 -23300 10134 -23248
rect 10186 -23300 10454 -23248
rect 10506 -23300 10774 -23248
rect 10826 -23300 11094 -23248
rect 11146 -23300 11414 -23248
rect 11466 -23300 11734 -23248
rect 11786 -23300 12054 -23248
rect 12106 -23300 12374 -23248
rect 12426 -23300 12694 -23248
rect 12746 -23300 13014 -23248
rect 13066 -23300 13334 -23248
rect 13386 -23300 14000 -23248
rect 6000 -23454 14000 -23300
rect 6000 -23506 6244 -23454
rect 6296 -23506 13710 -23454
rect 13762 -23506 14000 -23454
rect 6000 -23540 14000 -23506
rect 6000 -23774 6540 -23540
rect 6000 -23826 6244 -23774
rect 6296 -23826 6540 -23774
rect 6000 -24094 6540 -23826
rect 6000 -24146 6244 -24094
rect 6296 -24146 6540 -24094
rect 6000 -24414 6540 -24146
rect 6000 -24466 6244 -24414
rect 6296 -24466 6540 -24414
rect 6000 -24734 6540 -24466
rect 6000 -24786 6244 -24734
rect 6296 -24786 6540 -24734
rect 6000 -25054 6540 -24786
rect 6000 -25106 6244 -25054
rect 6296 -25106 6540 -25054
rect 6000 -25374 6540 -25106
rect 6000 -25426 6244 -25374
rect 6296 -25426 6540 -25374
rect 6000 -25694 6540 -25426
rect 6000 -25746 6244 -25694
rect 6296 -25746 6540 -25694
rect 6000 -26014 6540 -25746
rect 6000 -26066 6244 -26014
rect 6296 -26066 6540 -26014
rect 6000 -26334 6540 -26066
rect 6000 -26386 6244 -26334
rect 6296 -26386 6540 -26334
rect 6000 -26654 6540 -26386
rect 6000 -26706 6244 -26654
rect 6296 -26706 6540 -26654
rect 6000 -26974 6540 -26706
rect 6000 -27026 6244 -26974
rect 6296 -27026 6540 -26974
rect 6000 -27294 6540 -27026
rect 6000 -27346 6244 -27294
rect 6296 -27346 6540 -27294
rect 6000 -27614 6540 -27346
rect 6000 -27666 6244 -27614
rect 6296 -27666 6540 -27614
rect 6000 -27934 6540 -27666
rect 6000 -27986 6244 -27934
rect 6296 -27986 6540 -27934
rect 6000 -28254 6540 -27986
rect 6000 -28306 6244 -28254
rect 6296 -28306 6540 -28254
rect 6000 -28574 6540 -28306
rect 6000 -28626 6244 -28574
rect 6296 -28626 6540 -28574
rect 6000 -28894 6540 -28626
rect 6000 -28946 6244 -28894
rect 6296 -28946 6540 -28894
rect 6000 -29214 6540 -28946
rect 6000 -29266 6244 -29214
rect 6296 -29266 6540 -29214
rect 6000 -29534 6540 -29266
rect 6000 -29586 6244 -29534
rect 6296 -29586 6540 -29534
rect 6000 -29854 6540 -29586
rect 6000 -29906 6244 -29854
rect 6296 -29906 6540 -29854
rect 6000 -30174 6540 -29906
rect 6000 -30226 6244 -30174
rect 6296 -30226 6540 -30174
rect 6000 -30460 6540 -30226
rect 13460 -23774 14000 -23540
rect 13460 -23826 13710 -23774
rect 13762 -23826 14000 -23774
rect 13460 -24094 14000 -23826
rect 13460 -24146 13710 -24094
rect 13762 -24146 14000 -24094
rect 13460 -24414 14000 -24146
rect 13460 -24466 13710 -24414
rect 13762 -24466 14000 -24414
rect 13460 -24734 14000 -24466
rect 13460 -24786 13710 -24734
rect 13762 -24786 14000 -24734
rect 13460 -25054 14000 -24786
rect 13460 -25106 13710 -25054
rect 13762 -25106 14000 -25054
rect 13460 -25374 14000 -25106
rect 13460 -25426 13710 -25374
rect 13762 -25426 14000 -25374
rect 13460 -25694 14000 -25426
rect 13460 -25746 13710 -25694
rect 13762 -25746 14000 -25694
rect 13460 -26014 14000 -25746
rect 13460 -26066 13710 -26014
rect 13762 -26066 14000 -26014
rect 13460 -26334 14000 -26066
rect 13460 -26386 13710 -26334
rect 13762 -26386 14000 -26334
rect 13460 -26654 14000 -26386
rect 13460 -26706 13710 -26654
rect 13762 -26706 14000 -26654
rect 13460 -26974 14000 -26706
rect 13460 -27026 13710 -26974
rect 13762 -27026 14000 -26974
rect 13460 -27294 14000 -27026
rect 13460 -27346 13710 -27294
rect 13762 -27346 14000 -27294
rect 13460 -27614 14000 -27346
rect 13460 -27666 13710 -27614
rect 13762 -27666 14000 -27614
rect 13460 -27934 14000 -27666
rect 13460 -27986 13710 -27934
rect 13762 -27986 14000 -27934
rect 13460 -28254 14000 -27986
rect 13460 -28306 13710 -28254
rect 13762 -28306 14000 -28254
rect 13460 -28574 14000 -28306
rect 13460 -28626 13710 -28574
rect 13762 -28626 14000 -28574
rect 13460 -28894 14000 -28626
rect 13460 -28946 13710 -28894
rect 13762 -28946 14000 -28894
rect 13460 -29214 14000 -28946
rect 13460 -29266 13710 -29214
rect 13762 -29266 14000 -29214
rect 13460 -29534 14000 -29266
rect 13460 -29586 13710 -29534
rect 13762 -29586 14000 -29534
rect 13460 -29854 14000 -29586
rect 13460 -29906 13710 -29854
rect 13762 -29906 14000 -29854
rect 13460 -30174 14000 -29906
rect 13460 -30226 13710 -30174
rect 13762 -30226 14000 -30174
rect 13460 -30460 14000 -30226
rect 6000 -30494 14000 -30460
rect 6000 -30546 6244 -30494
rect 6296 -30546 13710 -30494
rect 13762 -30546 14000 -30494
rect 6000 -30704 14000 -30546
rect 6000 -30756 6614 -30704
rect 6666 -30756 6934 -30704
rect 6986 -30756 7254 -30704
rect 7306 -30756 7574 -30704
rect 7626 -30756 7894 -30704
rect 7946 -30756 8214 -30704
rect 8266 -30756 8534 -30704
rect 8586 -30756 8854 -30704
rect 8906 -30756 9174 -30704
rect 9226 -30756 9494 -30704
rect 9546 -30756 9814 -30704
rect 9866 -30756 10134 -30704
rect 10186 -30756 10454 -30704
rect 10506 -30756 10774 -30704
rect 10826 -30756 11094 -30704
rect 11146 -30756 11414 -30704
rect 11466 -30756 11734 -30704
rect 11786 -30756 12054 -30704
rect 12106 -30756 12374 -30704
rect 12426 -30756 12694 -30704
rect 12746 -30756 13014 -30704
rect 13066 -30756 13334 -30704
rect 13386 -30756 14000 -30704
rect 6000 -31000 14000 -30756
rect 18000 -23248 26000 -23000
rect 18000 -23300 18614 -23248
rect 18666 -23300 18934 -23248
rect 18986 -23300 19254 -23248
rect 19306 -23300 19574 -23248
rect 19626 -23300 19894 -23248
rect 19946 -23300 20214 -23248
rect 20266 -23300 20534 -23248
rect 20586 -23300 20854 -23248
rect 20906 -23300 21174 -23248
rect 21226 -23300 21494 -23248
rect 21546 -23300 21814 -23248
rect 21866 -23300 22134 -23248
rect 22186 -23300 22454 -23248
rect 22506 -23300 22774 -23248
rect 22826 -23300 23094 -23248
rect 23146 -23300 23414 -23248
rect 23466 -23300 23734 -23248
rect 23786 -23300 24054 -23248
rect 24106 -23300 24374 -23248
rect 24426 -23300 24694 -23248
rect 24746 -23300 25014 -23248
rect 25066 -23300 25334 -23248
rect 25386 -23300 26000 -23248
rect 18000 -23454 26000 -23300
rect 18000 -23506 18244 -23454
rect 18296 -23506 25710 -23454
rect 25762 -23506 26000 -23454
rect 18000 -23540 26000 -23506
rect 18000 -23774 18540 -23540
rect 18000 -23826 18244 -23774
rect 18296 -23826 18540 -23774
rect 18000 -24094 18540 -23826
rect 18000 -24146 18244 -24094
rect 18296 -24146 18540 -24094
rect 18000 -24414 18540 -24146
rect 18000 -24466 18244 -24414
rect 18296 -24466 18540 -24414
rect 18000 -24734 18540 -24466
rect 18000 -24786 18244 -24734
rect 18296 -24786 18540 -24734
rect 18000 -25054 18540 -24786
rect 18000 -25106 18244 -25054
rect 18296 -25106 18540 -25054
rect 18000 -25374 18540 -25106
rect 18000 -25426 18244 -25374
rect 18296 -25426 18540 -25374
rect 18000 -25694 18540 -25426
rect 18000 -25746 18244 -25694
rect 18296 -25746 18540 -25694
rect 18000 -26014 18540 -25746
rect 18000 -26066 18244 -26014
rect 18296 -26066 18540 -26014
rect 18000 -26334 18540 -26066
rect 18000 -26386 18244 -26334
rect 18296 -26386 18540 -26334
rect 18000 -26654 18540 -26386
rect 18000 -26706 18244 -26654
rect 18296 -26706 18540 -26654
rect 18000 -26974 18540 -26706
rect 18000 -27026 18244 -26974
rect 18296 -27026 18540 -26974
rect 18000 -27294 18540 -27026
rect 18000 -27346 18244 -27294
rect 18296 -27346 18540 -27294
rect 18000 -27614 18540 -27346
rect 18000 -27666 18244 -27614
rect 18296 -27666 18540 -27614
rect 18000 -27934 18540 -27666
rect 18000 -27986 18244 -27934
rect 18296 -27986 18540 -27934
rect 18000 -28254 18540 -27986
rect 18000 -28306 18244 -28254
rect 18296 -28306 18540 -28254
rect 18000 -28574 18540 -28306
rect 18000 -28626 18244 -28574
rect 18296 -28626 18540 -28574
rect 18000 -28894 18540 -28626
rect 18000 -28946 18244 -28894
rect 18296 -28946 18540 -28894
rect 18000 -29214 18540 -28946
rect 18000 -29266 18244 -29214
rect 18296 -29266 18540 -29214
rect 18000 -29534 18540 -29266
rect 18000 -29586 18244 -29534
rect 18296 -29586 18540 -29534
rect 18000 -29854 18540 -29586
rect 18000 -29906 18244 -29854
rect 18296 -29906 18540 -29854
rect 18000 -30174 18540 -29906
rect 18000 -30226 18244 -30174
rect 18296 -30226 18540 -30174
rect 18000 -30460 18540 -30226
rect 25460 -23774 26000 -23540
rect 25460 -23826 25710 -23774
rect 25762 -23826 26000 -23774
rect 25460 -24094 26000 -23826
rect 25460 -24146 25710 -24094
rect 25762 -24146 26000 -24094
rect 25460 -24414 26000 -24146
rect 25460 -24466 25710 -24414
rect 25762 -24466 26000 -24414
rect 25460 -24734 26000 -24466
rect 25460 -24786 25710 -24734
rect 25762 -24786 26000 -24734
rect 25460 -25054 26000 -24786
rect 25460 -25106 25710 -25054
rect 25762 -25106 26000 -25054
rect 25460 -25374 26000 -25106
rect 25460 -25426 25710 -25374
rect 25762 -25426 26000 -25374
rect 25460 -25694 26000 -25426
rect 25460 -25746 25710 -25694
rect 25762 -25746 26000 -25694
rect 25460 -26014 26000 -25746
rect 25460 -26066 25710 -26014
rect 25762 -26066 26000 -26014
rect 25460 -26334 26000 -26066
rect 25460 -26386 25710 -26334
rect 25762 -26386 26000 -26334
rect 25460 -26654 26000 -26386
rect 25460 -26706 25710 -26654
rect 25762 -26706 26000 -26654
rect 25460 -26974 26000 -26706
rect 25460 -27026 25710 -26974
rect 25762 -27026 26000 -26974
rect 25460 -27294 26000 -27026
rect 25460 -27346 25710 -27294
rect 25762 -27346 26000 -27294
rect 25460 -27614 26000 -27346
rect 25460 -27666 25710 -27614
rect 25762 -27666 26000 -27614
rect 25460 -27934 26000 -27666
rect 25460 -27986 25710 -27934
rect 25762 -27986 26000 -27934
rect 25460 -28254 26000 -27986
rect 25460 -28306 25710 -28254
rect 25762 -28306 26000 -28254
rect 25460 -28574 26000 -28306
rect 25460 -28626 25710 -28574
rect 25762 -28626 26000 -28574
rect 25460 -28894 26000 -28626
rect 25460 -28946 25710 -28894
rect 25762 -28946 26000 -28894
rect 25460 -29214 26000 -28946
rect 25460 -29266 25710 -29214
rect 25762 -29266 26000 -29214
rect 25460 -29534 26000 -29266
rect 25460 -29586 25710 -29534
rect 25762 -29586 26000 -29534
rect 25460 -29854 26000 -29586
rect 25460 -29906 25710 -29854
rect 25762 -29906 26000 -29854
rect 25460 -30174 26000 -29906
rect 25460 -30226 25710 -30174
rect 25762 -30226 26000 -30174
rect 25460 -30460 26000 -30226
rect 18000 -30494 26000 -30460
rect 18000 -30546 18244 -30494
rect 18296 -30546 25710 -30494
rect 25762 -30546 26000 -30494
rect 18000 -30704 26000 -30546
rect 18000 -30756 18614 -30704
rect 18666 -30756 18934 -30704
rect 18986 -30756 19254 -30704
rect 19306 -30756 19574 -30704
rect 19626 -30756 19894 -30704
rect 19946 -30756 20214 -30704
rect 20266 -30756 20534 -30704
rect 20586 -30756 20854 -30704
rect 20906 -30756 21174 -30704
rect 21226 -30756 21494 -30704
rect 21546 -30756 21814 -30704
rect 21866 -30756 22134 -30704
rect 22186 -30756 22454 -30704
rect 22506 -30756 22774 -30704
rect 22826 -30756 23094 -30704
rect 23146 -30756 23414 -30704
rect 23466 -30756 23734 -30704
rect 23786 -30756 24054 -30704
rect 24106 -30756 24374 -30704
rect 24426 -30756 24694 -30704
rect 24746 -30756 25014 -30704
rect 25066 -30756 25334 -30704
rect 25386 -30756 26000 -30704
rect 18000 -31000 26000 -30756
rect 30000 -23248 38000 -23000
rect 30000 -23300 30614 -23248
rect 30666 -23300 30934 -23248
rect 30986 -23300 31254 -23248
rect 31306 -23300 31574 -23248
rect 31626 -23300 31894 -23248
rect 31946 -23300 32214 -23248
rect 32266 -23300 32534 -23248
rect 32586 -23300 32854 -23248
rect 32906 -23300 33174 -23248
rect 33226 -23300 33494 -23248
rect 33546 -23300 33814 -23248
rect 33866 -23300 34134 -23248
rect 34186 -23300 34454 -23248
rect 34506 -23300 34774 -23248
rect 34826 -23300 35094 -23248
rect 35146 -23300 35414 -23248
rect 35466 -23300 35734 -23248
rect 35786 -23300 36054 -23248
rect 36106 -23300 36374 -23248
rect 36426 -23300 36694 -23248
rect 36746 -23300 37014 -23248
rect 37066 -23300 37334 -23248
rect 37386 -23300 38000 -23248
rect 30000 -23454 38000 -23300
rect 30000 -23506 30244 -23454
rect 30296 -23506 37710 -23454
rect 37762 -23506 38000 -23454
rect 30000 -23540 38000 -23506
rect 30000 -23774 30540 -23540
rect 30000 -23826 30244 -23774
rect 30296 -23826 30540 -23774
rect 30000 -24094 30540 -23826
rect 30000 -24146 30244 -24094
rect 30296 -24146 30540 -24094
rect 30000 -24414 30540 -24146
rect 30000 -24466 30244 -24414
rect 30296 -24466 30540 -24414
rect 30000 -24734 30540 -24466
rect 30000 -24786 30244 -24734
rect 30296 -24786 30540 -24734
rect 30000 -25054 30540 -24786
rect 30000 -25106 30244 -25054
rect 30296 -25106 30540 -25054
rect 30000 -25374 30540 -25106
rect 30000 -25426 30244 -25374
rect 30296 -25426 30540 -25374
rect 30000 -25694 30540 -25426
rect 30000 -25746 30244 -25694
rect 30296 -25746 30540 -25694
rect 30000 -26014 30540 -25746
rect 30000 -26066 30244 -26014
rect 30296 -26066 30540 -26014
rect 30000 -26334 30540 -26066
rect 30000 -26386 30244 -26334
rect 30296 -26386 30540 -26334
rect 30000 -26654 30540 -26386
rect 30000 -26706 30244 -26654
rect 30296 -26706 30540 -26654
rect 30000 -26974 30540 -26706
rect 30000 -27026 30244 -26974
rect 30296 -27026 30540 -26974
rect 30000 -27294 30540 -27026
rect 30000 -27346 30244 -27294
rect 30296 -27346 30540 -27294
rect 30000 -27614 30540 -27346
rect 30000 -27666 30244 -27614
rect 30296 -27666 30540 -27614
rect 30000 -27934 30540 -27666
rect 30000 -27986 30244 -27934
rect 30296 -27986 30540 -27934
rect 30000 -28254 30540 -27986
rect 30000 -28306 30244 -28254
rect 30296 -28306 30540 -28254
rect 30000 -28574 30540 -28306
rect 30000 -28626 30244 -28574
rect 30296 -28626 30540 -28574
rect 30000 -28894 30540 -28626
rect 30000 -28946 30244 -28894
rect 30296 -28946 30540 -28894
rect 30000 -29214 30540 -28946
rect 30000 -29266 30244 -29214
rect 30296 -29266 30540 -29214
rect 30000 -29534 30540 -29266
rect 30000 -29586 30244 -29534
rect 30296 -29586 30540 -29534
rect 30000 -29854 30540 -29586
rect 30000 -29906 30244 -29854
rect 30296 -29906 30540 -29854
rect 30000 -30174 30540 -29906
rect 30000 -30226 30244 -30174
rect 30296 -30226 30540 -30174
rect 30000 -30460 30540 -30226
rect 37460 -23774 38000 -23540
rect 37460 -23826 37710 -23774
rect 37762 -23826 38000 -23774
rect 37460 -24094 38000 -23826
rect 37460 -24146 37710 -24094
rect 37762 -24146 38000 -24094
rect 37460 -24414 38000 -24146
rect 37460 -24466 37710 -24414
rect 37762 -24466 38000 -24414
rect 37460 -24734 38000 -24466
rect 37460 -24786 37710 -24734
rect 37762 -24786 38000 -24734
rect 37460 -25054 38000 -24786
rect 37460 -25106 37710 -25054
rect 37762 -25106 38000 -25054
rect 37460 -25374 38000 -25106
rect 37460 -25426 37710 -25374
rect 37762 -25426 38000 -25374
rect 37460 -25694 38000 -25426
rect 37460 -25746 37710 -25694
rect 37762 -25746 38000 -25694
rect 37460 -26014 38000 -25746
rect 37460 -26066 37710 -26014
rect 37762 -26066 38000 -26014
rect 37460 -26334 38000 -26066
rect 37460 -26386 37710 -26334
rect 37762 -26386 38000 -26334
rect 37460 -26654 38000 -26386
rect 37460 -26706 37710 -26654
rect 37762 -26706 38000 -26654
rect 37460 -26974 38000 -26706
rect 37460 -27026 37710 -26974
rect 37762 -27026 38000 -26974
rect 37460 -27294 38000 -27026
rect 37460 -27346 37710 -27294
rect 37762 -27346 38000 -27294
rect 37460 -27614 38000 -27346
rect 37460 -27666 37710 -27614
rect 37762 -27666 38000 -27614
rect 37460 -27934 38000 -27666
rect 37460 -27986 37710 -27934
rect 37762 -27986 38000 -27934
rect 37460 -28254 38000 -27986
rect 37460 -28306 37710 -28254
rect 37762 -28306 38000 -28254
rect 37460 -28574 38000 -28306
rect 37460 -28626 37710 -28574
rect 37762 -28626 38000 -28574
rect 37460 -28894 38000 -28626
rect 37460 -28946 37710 -28894
rect 37762 -28946 38000 -28894
rect 37460 -29214 38000 -28946
rect 37460 -29266 37710 -29214
rect 37762 -29266 38000 -29214
rect 37460 -29534 38000 -29266
rect 37460 -29586 37710 -29534
rect 37762 -29586 38000 -29534
rect 37460 -29854 38000 -29586
rect 37460 -29906 37710 -29854
rect 37762 -29906 38000 -29854
rect 37460 -30174 38000 -29906
rect 37460 -30226 37710 -30174
rect 37762 -30226 38000 -30174
rect 37460 -30460 38000 -30226
rect 30000 -30494 38000 -30460
rect 30000 -30546 30244 -30494
rect 30296 -30546 37710 -30494
rect 37762 -30546 38000 -30494
rect 30000 -30704 38000 -30546
rect 30000 -30756 30614 -30704
rect 30666 -30756 30934 -30704
rect 30986 -30756 31254 -30704
rect 31306 -30756 31574 -30704
rect 31626 -30756 31894 -30704
rect 31946 -30756 32214 -30704
rect 32266 -30756 32534 -30704
rect 32586 -30756 32854 -30704
rect 32906 -30756 33174 -30704
rect 33226 -30756 33494 -30704
rect 33546 -30756 33814 -30704
rect 33866 -30756 34134 -30704
rect 34186 -30756 34454 -30704
rect 34506 -30756 34774 -30704
rect 34826 -30756 35094 -30704
rect 35146 -30756 35414 -30704
rect 35466 -30756 35734 -30704
rect 35786 -30756 36054 -30704
rect 36106 -30756 36374 -30704
rect 36426 -30756 36694 -30704
rect 36746 -30756 37014 -30704
rect 37066 -30756 37334 -30704
rect 37386 -30756 38000 -30704
rect 30000 -31000 38000 -30756
rect 42000 -23248 50000 -23000
rect 42000 -23300 42614 -23248
rect 42666 -23300 42934 -23248
rect 42986 -23300 43254 -23248
rect 43306 -23300 43574 -23248
rect 43626 -23300 43894 -23248
rect 43946 -23300 44214 -23248
rect 44266 -23300 44534 -23248
rect 44586 -23300 44854 -23248
rect 44906 -23300 45174 -23248
rect 45226 -23300 45494 -23248
rect 45546 -23300 45814 -23248
rect 45866 -23300 46134 -23248
rect 46186 -23300 46454 -23248
rect 46506 -23300 46774 -23248
rect 46826 -23300 47094 -23248
rect 47146 -23300 47414 -23248
rect 47466 -23300 47734 -23248
rect 47786 -23300 48054 -23248
rect 48106 -23300 48374 -23248
rect 48426 -23300 48694 -23248
rect 48746 -23300 49014 -23248
rect 49066 -23300 49334 -23248
rect 49386 -23300 50000 -23248
rect 42000 -23454 50000 -23300
rect 42000 -23506 42244 -23454
rect 42296 -23506 49710 -23454
rect 49762 -23506 50000 -23454
rect 42000 -23540 50000 -23506
rect 42000 -23774 42540 -23540
rect 42000 -23826 42244 -23774
rect 42296 -23826 42540 -23774
rect 42000 -24094 42540 -23826
rect 42000 -24146 42244 -24094
rect 42296 -24146 42540 -24094
rect 42000 -24414 42540 -24146
rect 42000 -24466 42244 -24414
rect 42296 -24466 42540 -24414
rect 42000 -24734 42540 -24466
rect 42000 -24786 42244 -24734
rect 42296 -24786 42540 -24734
rect 42000 -25054 42540 -24786
rect 42000 -25106 42244 -25054
rect 42296 -25106 42540 -25054
rect 42000 -25374 42540 -25106
rect 42000 -25426 42244 -25374
rect 42296 -25426 42540 -25374
rect 42000 -25694 42540 -25426
rect 42000 -25746 42244 -25694
rect 42296 -25746 42540 -25694
rect 42000 -26014 42540 -25746
rect 42000 -26066 42244 -26014
rect 42296 -26066 42540 -26014
rect 42000 -26334 42540 -26066
rect 42000 -26386 42244 -26334
rect 42296 -26386 42540 -26334
rect 42000 -26654 42540 -26386
rect 42000 -26706 42244 -26654
rect 42296 -26706 42540 -26654
rect 42000 -26974 42540 -26706
rect 42000 -27026 42244 -26974
rect 42296 -27026 42540 -26974
rect 42000 -27294 42540 -27026
rect 42000 -27346 42244 -27294
rect 42296 -27346 42540 -27294
rect 42000 -27614 42540 -27346
rect 42000 -27666 42244 -27614
rect 42296 -27666 42540 -27614
rect 42000 -27934 42540 -27666
rect 42000 -27986 42244 -27934
rect 42296 -27986 42540 -27934
rect 42000 -28254 42540 -27986
rect 42000 -28306 42244 -28254
rect 42296 -28306 42540 -28254
rect 42000 -28574 42540 -28306
rect 42000 -28626 42244 -28574
rect 42296 -28626 42540 -28574
rect 42000 -28894 42540 -28626
rect 42000 -28946 42244 -28894
rect 42296 -28946 42540 -28894
rect 42000 -29214 42540 -28946
rect 42000 -29266 42244 -29214
rect 42296 -29266 42540 -29214
rect 42000 -29534 42540 -29266
rect 42000 -29586 42244 -29534
rect 42296 -29586 42540 -29534
rect 42000 -29854 42540 -29586
rect 42000 -29906 42244 -29854
rect 42296 -29906 42540 -29854
rect 42000 -30174 42540 -29906
rect 42000 -30226 42244 -30174
rect 42296 -30226 42540 -30174
rect 42000 -30460 42540 -30226
rect 49460 -23774 50000 -23540
rect 49460 -23826 49710 -23774
rect 49762 -23826 50000 -23774
rect 49460 -24094 50000 -23826
rect 49460 -24146 49710 -24094
rect 49762 -24146 50000 -24094
rect 49460 -24414 50000 -24146
rect 49460 -24466 49710 -24414
rect 49762 -24466 50000 -24414
rect 49460 -24734 50000 -24466
rect 49460 -24786 49710 -24734
rect 49762 -24786 50000 -24734
rect 49460 -25054 50000 -24786
rect 49460 -25106 49710 -25054
rect 49762 -25106 50000 -25054
rect 49460 -25374 50000 -25106
rect 49460 -25426 49710 -25374
rect 49762 -25426 50000 -25374
rect 49460 -25694 50000 -25426
rect 49460 -25746 49710 -25694
rect 49762 -25746 50000 -25694
rect 49460 -26014 50000 -25746
rect 49460 -26066 49710 -26014
rect 49762 -26066 50000 -26014
rect 49460 -26334 50000 -26066
rect 49460 -26386 49710 -26334
rect 49762 -26386 50000 -26334
rect 49460 -26654 50000 -26386
rect 49460 -26706 49710 -26654
rect 49762 -26706 50000 -26654
rect 49460 -26974 50000 -26706
rect 49460 -27026 49710 -26974
rect 49762 -27026 50000 -26974
rect 49460 -27294 50000 -27026
rect 49460 -27346 49710 -27294
rect 49762 -27346 50000 -27294
rect 49460 -27614 50000 -27346
rect 49460 -27666 49710 -27614
rect 49762 -27666 50000 -27614
rect 49460 -27934 50000 -27666
rect 49460 -27986 49710 -27934
rect 49762 -27986 50000 -27934
rect 49460 -28254 50000 -27986
rect 49460 -28306 49710 -28254
rect 49762 -28306 50000 -28254
rect 49460 -28574 50000 -28306
rect 49460 -28626 49710 -28574
rect 49762 -28626 50000 -28574
rect 49460 -28894 50000 -28626
rect 49460 -28946 49710 -28894
rect 49762 -28946 50000 -28894
rect 49460 -29214 50000 -28946
rect 49460 -29266 49710 -29214
rect 49762 -29266 50000 -29214
rect 49460 -29534 50000 -29266
rect 49460 -29586 49710 -29534
rect 49762 -29586 50000 -29534
rect 49460 -29854 50000 -29586
rect 49460 -29906 49710 -29854
rect 49762 -29906 50000 -29854
rect 49460 -30174 50000 -29906
rect 49460 -30226 49710 -30174
rect 49762 -30226 50000 -30174
rect 49460 -30460 50000 -30226
rect 42000 -30494 50000 -30460
rect 42000 -30546 42244 -30494
rect 42296 -30546 49710 -30494
rect 49762 -30546 50000 -30494
rect 42000 -30704 50000 -30546
rect 42000 -30756 42614 -30704
rect 42666 -30756 42934 -30704
rect 42986 -30756 43254 -30704
rect 43306 -30756 43574 -30704
rect 43626 -30756 43894 -30704
rect 43946 -30756 44214 -30704
rect 44266 -30756 44534 -30704
rect 44586 -30756 44854 -30704
rect 44906 -30756 45174 -30704
rect 45226 -30756 45494 -30704
rect 45546 -30756 45814 -30704
rect 45866 -30756 46134 -30704
rect 46186 -30756 46454 -30704
rect 46506 -30756 46774 -30704
rect 46826 -30756 47094 -30704
rect 47146 -30756 47414 -30704
rect 47466 -30756 47734 -30704
rect 47786 -30756 48054 -30704
rect 48106 -30756 48374 -30704
rect 48426 -30756 48694 -30704
rect 48746 -30756 49014 -30704
rect 49066 -30756 49334 -30704
rect 49386 -30756 50000 -30704
rect 42000 -31000 50000 -30756
<< via1 >>
rect 18088 -5403 18097 -3427
rect 18097 -5403 18131 -3427
rect 18131 -5403 18140 -3427
rect 18206 -5403 18215 -3427
rect 18215 -5403 18249 -3427
rect 18249 -5403 18258 -3427
rect 18324 -5403 18333 -3427
rect 18333 -5403 18367 -3427
rect 18367 -5403 18376 -3427
rect 18442 -5403 18451 -3427
rect 18451 -5403 18485 -3427
rect 18485 -5403 18494 -3427
rect 18560 -5403 18569 -3427
rect 18569 -5403 18603 -3427
rect 18603 -5403 18612 -3427
rect 18678 -5403 18687 -3427
rect 18687 -5403 18721 -3427
rect 18721 -5403 18730 -3427
rect 18796 -5403 18805 -3427
rect 18805 -5403 18839 -3427
rect 18839 -5403 18848 -3427
rect 18914 -5403 18923 -3427
rect 18923 -5403 18957 -3427
rect 18957 -5403 18966 -3427
rect 19032 -5403 19041 -3427
rect 19041 -5403 19075 -3427
rect 19075 -5403 19084 -3427
rect 19150 -5403 19159 -3427
rect 19159 -5403 19193 -3427
rect 19193 -5403 19202 -3427
rect 19268 -5403 19277 -3427
rect 19277 -5403 19311 -3427
rect 19311 -5403 19320 -3427
rect 19386 -5403 19395 -3427
rect 19395 -5403 19429 -3427
rect 19429 -5403 19438 -3427
rect 19504 -5403 19513 -3427
rect 19513 -5403 19547 -3427
rect 19547 -5403 19556 -3427
rect 19622 -5403 19631 -3427
rect 19631 -5403 19665 -3427
rect 19665 -5403 19674 -3427
rect 19740 -5403 19749 -3427
rect 19749 -5403 19783 -3427
rect 19783 -5403 19792 -3427
rect 19858 -5403 19867 -3427
rect 19867 -5403 19901 -3427
rect 19901 -5403 19910 -3427
rect 19976 -5403 19985 -3427
rect 19985 -5403 20019 -3427
rect 20019 -5403 20028 -3427
rect 20094 -5403 20103 -3427
rect 20103 -5403 20137 -3427
rect 20137 -5403 20146 -3427
rect 20212 -5403 20221 -3427
rect 20221 -5403 20255 -3427
rect 20255 -5403 20264 -3427
rect 20330 -5403 20339 -3427
rect 20339 -5403 20373 -3427
rect 20373 -5403 20382 -3427
rect 20448 -5403 20457 -3427
rect 20457 -5403 20491 -3427
rect 20491 -5403 20500 -3427
rect 20566 -5403 20575 -3427
rect 20575 -5403 20609 -3427
rect 20609 -5403 20618 -3427
rect 20684 -5403 20693 -3427
rect 20693 -5403 20727 -3427
rect 20727 -5403 20736 -3427
rect 20802 -5403 20811 -3427
rect 20811 -5403 20845 -3427
rect 20845 -5403 20854 -3427
rect 20920 -5403 20929 -3427
rect 20929 -5403 20963 -3427
rect 20963 -5403 20972 -3427
rect 21038 -5403 21047 -3427
rect 21047 -5403 21081 -3427
rect 21081 -5403 21090 -3427
rect 21156 -5403 21165 -3427
rect 21165 -5403 21199 -3427
rect 21199 -5403 21208 -3427
rect 21274 -5403 21283 -3427
rect 21283 -5403 21317 -3427
rect 21317 -5403 21326 -3427
rect 21392 -5403 21401 -3427
rect 21401 -5403 21435 -3427
rect 21435 -5403 21444 -3427
rect 21510 -5403 21519 -3427
rect 21519 -5403 21553 -3427
rect 21553 -5403 21562 -3427
rect 21628 -5403 21637 -3427
rect 21637 -5403 21671 -3427
rect 21671 -5403 21680 -3427
rect 21746 -5403 21755 -3427
rect 21755 -5403 21789 -3427
rect 21789 -5403 21798 -3427
rect 21864 -5403 21873 -3427
rect 21873 -5403 21907 -3427
rect 21907 -5403 21916 -3427
rect 19918 -5462 19970 -5456
rect 19918 -5496 19926 -5462
rect 19926 -5496 19960 -5462
rect 19960 -5496 19970 -5462
rect 19918 -5508 19970 -5496
rect 20033 -5552 20085 -5500
rect 18205 -5794 18257 -5742
rect 21746 -5794 21798 -5742
rect 17851 -7912 17860 -5936
rect 17860 -7912 17894 -5936
rect 17894 -7912 17903 -5936
rect 17969 -7912 17978 -5936
rect 17978 -7912 18012 -5936
rect 18012 -7912 18021 -5936
rect 18087 -7912 18096 -5936
rect 18096 -7912 18130 -5936
rect 18130 -7912 18139 -5936
rect 18205 -7912 18214 -5936
rect 18214 -7912 18248 -5936
rect 18248 -7912 18257 -5936
rect 18323 -7912 18332 -5936
rect 18332 -7912 18366 -5936
rect 18366 -7912 18375 -5936
rect 18441 -7912 18450 -5936
rect 18450 -7912 18484 -5936
rect 18484 -7912 18493 -5936
rect 18559 -7912 18568 -5936
rect 18568 -7912 18602 -5936
rect 18602 -7912 18611 -5936
rect 19015 -6112 19069 -6100
rect 19015 -6588 19025 -6112
rect 19025 -6588 19059 -6112
rect 19059 -6588 19069 -6112
rect 19015 -6600 19069 -6588
rect 19111 -6112 19165 -6100
rect 19111 -6588 19121 -6112
rect 19121 -6588 19155 -6112
rect 19155 -6588 19165 -6112
rect 19111 -6600 19165 -6588
rect 19207 -6112 19261 -6100
rect 19207 -6588 19217 -6112
rect 19217 -6588 19251 -6112
rect 19251 -6588 19261 -6112
rect 19207 -6600 19261 -6588
rect 19303 -6112 19357 -6100
rect 19303 -6588 19313 -6112
rect 19313 -6588 19347 -6112
rect 19347 -6588 19357 -6112
rect 19303 -6600 19357 -6588
rect 19399 -6112 19453 -6100
rect 19399 -6588 19409 -6112
rect 19409 -6588 19443 -6112
rect 19443 -6588 19453 -6112
rect 19399 -6600 19453 -6588
rect 19495 -6112 19549 -6100
rect 19495 -6588 19505 -6112
rect 19505 -6588 19539 -6112
rect 19539 -6588 19549 -6112
rect 19495 -6600 19549 -6588
rect 19591 -6112 19645 -6100
rect 19591 -6588 19601 -6112
rect 19601 -6588 19635 -6112
rect 19635 -6588 19645 -6112
rect 19591 -6600 19645 -6588
rect 19687 -6112 19741 -6100
rect 19687 -6588 19697 -6112
rect 19697 -6588 19731 -6112
rect 19731 -6588 19741 -6112
rect 19687 -6600 19741 -6588
rect 19783 -6112 19837 -6100
rect 19783 -6588 19793 -6112
rect 19793 -6588 19827 -6112
rect 19827 -6588 19837 -6112
rect 19783 -6600 19837 -6588
rect 19879 -6112 19933 -6100
rect 19879 -6588 19889 -6112
rect 19889 -6588 19923 -6112
rect 19923 -6588 19933 -6112
rect 19879 -6600 19933 -6588
rect 19975 -6112 20029 -6100
rect 19975 -6588 19985 -6112
rect 19985 -6588 20019 -6112
rect 20019 -6588 20029 -6112
rect 19975 -6600 20029 -6588
rect 20071 -6112 20125 -6100
rect 20071 -6588 20081 -6112
rect 20081 -6588 20115 -6112
rect 20115 -6588 20125 -6112
rect 20071 -6600 20125 -6588
rect 20167 -6112 20221 -6100
rect 20167 -6588 20177 -6112
rect 20177 -6588 20211 -6112
rect 20211 -6588 20221 -6112
rect 20167 -6600 20221 -6588
rect 20263 -6112 20317 -6100
rect 20263 -6588 20273 -6112
rect 20273 -6588 20307 -6112
rect 20307 -6588 20317 -6112
rect 20263 -6600 20317 -6588
rect 20359 -6112 20413 -6100
rect 20359 -6588 20369 -6112
rect 20369 -6588 20403 -6112
rect 20403 -6588 20413 -6112
rect 20359 -6600 20413 -6588
rect 20455 -6112 20509 -6100
rect 20455 -6588 20465 -6112
rect 20465 -6588 20499 -6112
rect 20499 -6588 20509 -6112
rect 20455 -6600 20509 -6588
rect 20551 -6112 20605 -6100
rect 20551 -6588 20561 -6112
rect 20561 -6588 20595 -6112
rect 20595 -6588 20605 -6112
rect 20551 -6600 20605 -6588
rect 20647 -6112 20701 -6100
rect 20647 -6588 20657 -6112
rect 20657 -6588 20691 -6112
rect 20691 -6588 20701 -6112
rect 20647 -6600 20701 -6588
rect 20743 -6112 20797 -6100
rect 20743 -6588 20753 -6112
rect 20753 -6588 20787 -6112
rect 20787 -6588 20797 -6112
rect 20743 -6600 20797 -6588
rect 20839 -6112 20893 -6100
rect 20839 -6588 20849 -6112
rect 20849 -6588 20883 -6112
rect 20883 -6588 20893 -6112
rect 20839 -6600 20893 -6588
rect 20935 -6112 20989 -6100
rect 20935 -6588 20945 -6112
rect 20945 -6588 20979 -6112
rect 20979 -6588 20989 -6112
rect 20935 -6600 20989 -6588
rect 19297 -6650 19363 -6644
rect 19297 -6684 19313 -6650
rect 19313 -6684 19347 -6650
rect 19347 -6684 19363 -6650
rect 19297 -6700 19363 -6684
rect 19489 -6650 19555 -6644
rect 19489 -6684 19505 -6650
rect 19505 -6684 19539 -6650
rect 19539 -6684 19555 -6650
rect 19489 -6700 19555 -6684
rect 19681 -6650 19747 -6644
rect 19681 -6684 19697 -6650
rect 19697 -6684 19731 -6650
rect 19731 -6684 19747 -6650
rect 19681 -6700 19747 -6684
rect 19873 -6650 19939 -6644
rect 19873 -6684 19889 -6650
rect 19889 -6684 19923 -6650
rect 19923 -6684 19939 -6650
rect 19873 -6700 19939 -6684
rect 20065 -6650 20131 -6644
rect 20065 -6684 20081 -6650
rect 20081 -6684 20115 -6650
rect 20115 -6684 20131 -6650
rect 20065 -6700 20131 -6684
rect 20257 -6650 20323 -6644
rect 20257 -6684 20273 -6650
rect 20273 -6684 20307 -6650
rect 20307 -6684 20323 -6650
rect 20257 -6700 20323 -6684
rect 20449 -6650 20515 -6644
rect 20449 -6684 20465 -6650
rect 20465 -6684 20499 -6650
rect 20499 -6684 20515 -6650
rect 20449 -6700 20515 -6684
rect 20641 -6650 20707 -6644
rect 20641 -6684 20657 -6650
rect 20657 -6684 20691 -6650
rect 20691 -6684 20707 -6650
rect 20641 -6700 20707 -6684
rect 19058 -7002 19122 -6938
rect 16666 -8494 17135 -8485
rect 16666 -8528 17135 -8494
rect 16666 -8537 17135 -8528
rect 16400 -9580 16460 -9520
rect 16590 -9108 17019 -9100
rect 16590 -9161 17019 -9108
rect 16590 -9170 17019 -9161
rect 17400 -9360 17460 -8440
rect 17460 -9360 17600 -8440
rect 18822 -9280 18882 -8060
rect 19060 -9028 19069 -7052
rect 19069 -9028 19103 -7052
rect 19103 -9028 19112 -7052
rect 19518 -9028 19527 -7052
rect 19527 -9028 19561 -7052
rect 19561 -9028 19570 -7052
rect 19976 -9028 19985 -7052
rect 19985 -9028 20019 -7052
rect 20019 -9028 20028 -7052
rect 20434 -9028 20443 -7052
rect 20443 -9028 20477 -7052
rect 20477 -9028 20486 -7052
rect 20892 -9028 20901 -7052
rect 20901 -9028 20935 -7052
rect 20935 -9028 20944 -7052
rect 21392 -7912 21401 -5936
rect 21401 -7912 21435 -5936
rect 21435 -7912 21444 -5936
rect 21510 -7912 21519 -5936
rect 21519 -7912 21553 -5936
rect 21553 -7912 21562 -5936
rect 21628 -7912 21637 -5936
rect 21637 -7912 21671 -5936
rect 21671 -7912 21680 -5936
rect 21746 -7912 21755 -5936
rect 21755 -7912 21789 -5936
rect 21789 -7912 21798 -5936
rect 21864 -7912 21873 -5936
rect 21873 -7912 21907 -5936
rect 21907 -7912 21916 -5936
rect 21982 -7912 21991 -5936
rect 21991 -7912 22025 -5936
rect 22025 -7912 22034 -5936
rect 22100 -7912 22109 -5936
rect 22109 -7912 22143 -5936
rect 22143 -7912 22152 -5936
rect 22472 -6660 22582 -6270
rect 22702 -6660 22812 -6270
rect 23300 -7353 23500 -7200
rect 23300 -7387 23311 -7353
rect 23311 -7387 23369 -7353
rect 23369 -7387 23403 -7353
rect 23403 -7387 23461 -7353
rect 23461 -7387 23495 -7353
rect 23495 -7387 23500 -7353
rect 23300 -7400 23500 -7387
rect 23270 -7662 23410 -7640
rect 23270 -7702 23280 -7662
rect 23280 -7702 23400 -7662
rect 23400 -7702 23410 -7662
rect 23270 -7720 23410 -7702
rect 23550 -7662 23690 -7640
rect 23550 -7702 23556 -7662
rect 23556 -7702 23676 -7662
rect 23676 -7702 23690 -7662
rect 23550 -7720 23690 -7702
rect 23300 -7931 23311 -7900
rect 23311 -7931 23369 -7900
rect 23369 -7931 23403 -7900
rect 23403 -7931 23461 -7900
rect 23461 -7931 23495 -7900
rect 23495 -7931 23500 -7900
rect 21122 -9280 21182 -8060
rect 23300 -8100 23500 -7931
rect 16470 -9720 16530 -9660
rect 16710 -10850 16800 -10510
rect 17030 -10738 17120 -10620
rect 17120 -10738 17130 -10620
rect 17030 -10740 17130 -10738
rect 17420 -10850 17510 -10510
rect 6614 -11300 6666 -11248
rect 6934 -11300 6986 -11248
rect 7254 -11300 7306 -11248
rect 7574 -11300 7626 -11248
rect 7894 -11300 7946 -11248
rect 8214 -11300 8266 -11248
rect 8534 -11300 8586 -11248
rect 8854 -11300 8906 -11248
rect 9174 -11300 9226 -11248
rect 9494 -11300 9546 -11248
rect 9814 -11300 9866 -11248
rect 10134 -11300 10186 -11248
rect 10454 -11300 10506 -11248
rect 10774 -11300 10826 -11248
rect 11094 -11300 11146 -11248
rect 11414 -11300 11466 -11248
rect 11734 -11300 11786 -11248
rect 12054 -11300 12106 -11248
rect 12374 -11300 12426 -11248
rect 12694 -11300 12746 -11248
rect 13014 -11300 13066 -11248
rect 13334 -11300 13386 -11248
rect 6244 -11506 6296 -11454
rect 13710 -11506 13762 -11454
rect 6244 -11826 6296 -11774
rect 6244 -12146 6296 -12094
rect 6244 -12466 6296 -12414
rect 6244 -12786 6296 -12734
rect 6244 -13106 6296 -13054
rect 6244 -13426 6296 -13374
rect 6244 -13746 6296 -13694
rect 6244 -14066 6296 -14014
rect 6244 -14386 6296 -14334
rect 6244 -14706 6296 -14654
rect 6244 -15026 6296 -14974
rect 6244 -15346 6296 -15294
rect 6244 -15666 6296 -15614
rect 6244 -15986 6296 -15934
rect 6244 -16306 6296 -16254
rect 6244 -16626 6296 -16574
rect 6244 -16946 6296 -16894
rect 6244 -17266 6296 -17214
rect 6244 -17586 6296 -17534
rect 6244 -17906 6296 -17854
rect 6244 -18226 6296 -18174
rect 13710 -11826 13762 -11774
rect 13710 -12146 13762 -12094
rect 13710 -12466 13762 -12414
rect 13710 -12786 13762 -12734
rect 13710 -13106 13762 -13054
rect 13710 -13426 13762 -13374
rect 13710 -13746 13762 -13694
rect 13710 -14066 13762 -14014
rect 13710 -14386 13762 -14334
rect 13710 -14706 13762 -14654
rect 13710 -15026 13762 -14974
rect 13710 -15346 13762 -15294
rect 13710 -15666 13762 -15614
rect 13710 -15986 13762 -15934
rect 13710 -16306 13762 -16254
rect 13710 -16626 13762 -16574
rect 13710 -16946 13762 -16894
rect 13710 -17266 13762 -17214
rect 13710 -17586 13762 -17534
rect 13710 -17906 13762 -17854
rect 13710 -18226 13762 -18174
rect 6244 -18546 6296 -18494
rect 13710 -18546 13762 -18494
rect 6614 -18756 6666 -18704
rect 6934 -18756 6986 -18704
rect 7254 -18756 7306 -18704
rect 7574 -18756 7626 -18704
rect 7894 -18756 7946 -18704
rect 8214 -18756 8266 -18704
rect 8534 -18756 8586 -18704
rect 8854 -18756 8906 -18704
rect 9174 -18756 9226 -18704
rect 9494 -18756 9546 -18704
rect 9814 -18756 9866 -18704
rect 10134 -18756 10186 -18704
rect 10454 -18756 10506 -18704
rect 10774 -18756 10826 -18704
rect 11094 -18756 11146 -18704
rect 11414 -18756 11466 -18704
rect 11734 -18756 11786 -18704
rect 12054 -18756 12106 -18704
rect 12374 -18756 12426 -18704
rect 12694 -18756 12746 -18704
rect 13014 -18756 13066 -18704
rect 13334 -18756 13386 -18704
rect 18614 -11300 18666 -11248
rect 18934 -11300 18986 -11248
rect 19254 -11300 19306 -11248
rect 19574 -11300 19626 -11248
rect 19894 -11300 19946 -11248
rect 20214 -11300 20266 -11248
rect 20534 -11300 20586 -11248
rect 20854 -11300 20906 -11248
rect 21174 -11300 21226 -11248
rect 21494 -11300 21546 -11248
rect 21814 -11300 21866 -11248
rect 22134 -11300 22186 -11248
rect 22454 -11300 22506 -11248
rect 22774 -11300 22826 -11248
rect 23094 -11300 23146 -11248
rect 23414 -11300 23466 -11248
rect 23734 -11300 23786 -11248
rect 24054 -11300 24106 -11248
rect 24374 -11300 24426 -11248
rect 24694 -11300 24746 -11248
rect 25014 -11300 25066 -11248
rect 25334 -11300 25386 -11248
rect 18244 -11506 18296 -11454
rect 25710 -11506 25762 -11454
rect 18244 -11826 18296 -11774
rect 18244 -12146 18296 -12094
rect 18244 -12466 18296 -12414
rect 18244 -12786 18296 -12734
rect 18244 -13106 18296 -13054
rect 18244 -13426 18296 -13374
rect 18244 -13746 18296 -13694
rect 18244 -14066 18296 -14014
rect 18244 -14386 18296 -14334
rect 18244 -14706 18296 -14654
rect 18244 -15026 18296 -14974
rect 18244 -15346 18296 -15294
rect 18244 -15666 18296 -15614
rect 18244 -15986 18296 -15934
rect 18244 -16306 18296 -16254
rect 18244 -16626 18296 -16574
rect 18244 -16946 18296 -16894
rect 18244 -17266 18296 -17214
rect 18244 -17586 18296 -17534
rect 18244 -17906 18296 -17854
rect 18244 -18226 18296 -18174
rect 25710 -11826 25762 -11774
rect 25710 -12146 25762 -12094
rect 25710 -12466 25762 -12414
rect 25710 -12786 25762 -12734
rect 25710 -13106 25762 -13054
rect 25710 -13426 25762 -13374
rect 25710 -13746 25762 -13694
rect 25710 -14066 25762 -14014
rect 25710 -14386 25762 -14334
rect 25710 -14706 25762 -14654
rect 25710 -15026 25762 -14974
rect 25710 -15346 25762 -15294
rect 25710 -15666 25762 -15614
rect 25710 -15986 25762 -15934
rect 25710 -16306 25762 -16254
rect 25710 -16626 25762 -16574
rect 25710 -16946 25762 -16894
rect 25710 -17266 25762 -17214
rect 25710 -17586 25762 -17534
rect 25710 -17906 25762 -17854
rect 25710 -18226 25762 -18174
rect 18244 -18546 18296 -18494
rect 25710 -18546 25762 -18494
rect 18614 -18756 18666 -18704
rect 18934 -18756 18986 -18704
rect 19254 -18756 19306 -18704
rect 19574 -18756 19626 -18704
rect 19894 -18756 19946 -18704
rect 20214 -18756 20266 -18704
rect 20534 -18756 20586 -18704
rect 20854 -18756 20906 -18704
rect 21174 -18756 21226 -18704
rect 21494 -18756 21546 -18704
rect 21814 -18756 21866 -18704
rect 22134 -18756 22186 -18704
rect 22454 -18756 22506 -18704
rect 22774 -18756 22826 -18704
rect 23094 -18756 23146 -18704
rect 23414 -18756 23466 -18704
rect 23734 -18756 23786 -18704
rect 24054 -18756 24106 -18704
rect 24374 -18756 24426 -18704
rect 24694 -18756 24746 -18704
rect 25014 -18756 25066 -18704
rect 25334 -18756 25386 -18704
rect 30614 -11300 30666 -11248
rect 30934 -11300 30986 -11248
rect 31254 -11300 31306 -11248
rect 31574 -11300 31626 -11248
rect 31894 -11300 31946 -11248
rect 32214 -11300 32266 -11248
rect 32534 -11300 32586 -11248
rect 32854 -11300 32906 -11248
rect 33174 -11300 33226 -11248
rect 33494 -11300 33546 -11248
rect 33814 -11300 33866 -11248
rect 34134 -11300 34186 -11248
rect 34454 -11300 34506 -11248
rect 34774 -11300 34826 -11248
rect 35094 -11300 35146 -11248
rect 35414 -11300 35466 -11248
rect 35734 -11300 35786 -11248
rect 36054 -11300 36106 -11248
rect 36374 -11300 36426 -11248
rect 36694 -11300 36746 -11248
rect 37014 -11300 37066 -11248
rect 37334 -11300 37386 -11248
rect 30244 -11506 30296 -11454
rect 37710 -11506 37762 -11454
rect 30244 -11826 30296 -11774
rect 30244 -12146 30296 -12094
rect 30244 -12466 30296 -12414
rect 30244 -12786 30296 -12734
rect 30244 -13106 30296 -13054
rect 30244 -13426 30296 -13374
rect 30244 -13746 30296 -13694
rect 30244 -14066 30296 -14014
rect 30244 -14386 30296 -14334
rect 30244 -14706 30296 -14654
rect 30244 -15026 30296 -14974
rect 30244 -15346 30296 -15294
rect 30244 -15666 30296 -15614
rect 30244 -15986 30296 -15934
rect 30244 -16306 30296 -16254
rect 30244 -16626 30296 -16574
rect 30244 -16946 30296 -16894
rect 30244 -17266 30296 -17214
rect 30244 -17586 30296 -17534
rect 30244 -17906 30296 -17854
rect 30244 -18226 30296 -18174
rect 37710 -11826 37762 -11774
rect 37710 -12146 37762 -12094
rect 37710 -12466 37762 -12414
rect 37710 -12786 37762 -12734
rect 37710 -13106 37762 -13054
rect 37710 -13426 37762 -13374
rect 37710 -13746 37762 -13694
rect 37710 -14066 37762 -14014
rect 37710 -14386 37762 -14334
rect 37710 -14706 37762 -14654
rect 37710 -15026 37762 -14974
rect 37710 -15346 37762 -15294
rect 37710 -15666 37762 -15614
rect 37710 -15986 37762 -15934
rect 37710 -16306 37762 -16254
rect 37710 -16626 37762 -16574
rect 37710 -16946 37762 -16894
rect 37710 -17266 37762 -17214
rect 37710 -17586 37762 -17534
rect 37710 -17906 37762 -17854
rect 37710 -18226 37762 -18174
rect 30244 -18546 30296 -18494
rect 37710 -18546 37762 -18494
rect 30614 -18756 30666 -18704
rect 30934 -18756 30986 -18704
rect 31254 -18756 31306 -18704
rect 31574 -18756 31626 -18704
rect 31894 -18756 31946 -18704
rect 32214 -18756 32266 -18704
rect 32534 -18756 32586 -18704
rect 32854 -18756 32906 -18704
rect 33174 -18756 33226 -18704
rect 33494 -18756 33546 -18704
rect 33814 -18756 33866 -18704
rect 34134 -18756 34186 -18704
rect 34454 -18756 34506 -18704
rect 34774 -18756 34826 -18704
rect 35094 -18756 35146 -18704
rect 35414 -18756 35466 -18704
rect 35734 -18756 35786 -18704
rect 36054 -18756 36106 -18704
rect 36374 -18756 36426 -18704
rect 36694 -18756 36746 -18704
rect 37014 -18756 37066 -18704
rect 37334 -18756 37386 -18704
rect 42614 -11300 42666 -11248
rect 42934 -11300 42986 -11248
rect 43254 -11300 43306 -11248
rect 43574 -11300 43626 -11248
rect 43894 -11300 43946 -11248
rect 44214 -11300 44266 -11248
rect 44534 -11300 44586 -11248
rect 44854 -11300 44906 -11248
rect 45174 -11300 45226 -11248
rect 45494 -11300 45546 -11248
rect 45814 -11300 45866 -11248
rect 46134 -11300 46186 -11248
rect 46454 -11300 46506 -11248
rect 46774 -11300 46826 -11248
rect 47094 -11300 47146 -11248
rect 47414 -11300 47466 -11248
rect 47734 -11300 47786 -11248
rect 48054 -11300 48106 -11248
rect 48374 -11300 48426 -11248
rect 48694 -11300 48746 -11248
rect 49014 -11300 49066 -11248
rect 49334 -11300 49386 -11248
rect 42244 -11506 42296 -11454
rect 49710 -11506 49762 -11454
rect 42244 -11826 42296 -11774
rect 42244 -12146 42296 -12094
rect 42244 -12466 42296 -12414
rect 42244 -12786 42296 -12734
rect 42244 -13106 42296 -13054
rect 42244 -13426 42296 -13374
rect 42244 -13746 42296 -13694
rect 42244 -14066 42296 -14014
rect 42244 -14386 42296 -14334
rect 42244 -14706 42296 -14654
rect 42244 -15026 42296 -14974
rect 42244 -15346 42296 -15294
rect 42244 -15666 42296 -15614
rect 42244 -15986 42296 -15934
rect 42244 -16306 42296 -16254
rect 42244 -16626 42296 -16574
rect 42244 -16946 42296 -16894
rect 42244 -17266 42296 -17214
rect 42244 -17586 42296 -17534
rect 42244 -17906 42296 -17854
rect 42244 -18226 42296 -18174
rect 49710 -11826 49762 -11774
rect 49710 -12146 49762 -12094
rect 49710 -12466 49762 -12414
rect 49710 -12786 49762 -12734
rect 49710 -13106 49762 -13054
rect 49710 -13426 49762 -13374
rect 49710 -13746 49762 -13694
rect 49710 -14066 49762 -14014
rect 49710 -14386 49762 -14334
rect 49710 -14706 49762 -14654
rect 49710 -15026 49762 -14974
rect 49710 -15346 49762 -15294
rect 49710 -15666 49762 -15614
rect 49710 -15986 49762 -15934
rect 49710 -16306 49762 -16254
rect 49710 -16626 49762 -16574
rect 49710 -16946 49762 -16894
rect 49710 -17266 49762 -17214
rect 49710 -17586 49762 -17534
rect 49710 -17906 49762 -17854
rect 49710 -18226 49762 -18174
rect 42244 -18546 42296 -18494
rect 49710 -18546 49762 -18494
rect 42614 -18756 42666 -18704
rect 42934 -18756 42986 -18704
rect 43254 -18756 43306 -18704
rect 43574 -18756 43626 -18704
rect 43894 -18756 43946 -18704
rect 44214 -18756 44266 -18704
rect 44534 -18756 44586 -18704
rect 44854 -18756 44906 -18704
rect 45174 -18756 45226 -18704
rect 45494 -18756 45546 -18704
rect 45814 -18756 45866 -18704
rect 46134 -18756 46186 -18704
rect 46454 -18756 46506 -18704
rect 46774 -18756 46826 -18704
rect 47094 -18756 47146 -18704
rect 47414 -18756 47466 -18704
rect 47734 -18756 47786 -18704
rect 48054 -18756 48106 -18704
rect 48374 -18756 48426 -18704
rect 48694 -18756 48746 -18704
rect 49014 -18756 49066 -18704
rect 49334 -18756 49386 -18704
rect 6614 -23300 6666 -23248
rect 6934 -23300 6986 -23248
rect 7254 -23300 7306 -23248
rect 7574 -23300 7626 -23248
rect 7894 -23300 7946 -23248
rect 8214 -23300 8266 -23248
rect 8534 -23300 8586 -23248
rect 8854 -23300 8906 -23248
rect 9174 -23300 9226 -23248
rect 9494 -23300 9546 -23248
rect 9814 -23300 9866 -23248
rect 10134 -23300 10186 -23248
rect 10454 -23300 10506 -23248
rect 10774 -23300 10826 -23248
rect 11094 -23300 11146 -23248
rect 11414 -23300 11466 -23248
rect 11734 -23300 11786 -23248
rect 12054 -23300 12106 -23248
rect 12374 -23300 12426 -23248
rect 12694 -23300 12746 -23248
rect 13014 -23300 13066 -23248
rect 13334 -23300 13386 -23248
rect 6244 -23506 6296 -23454
rect 13710 -23506 13762 -23454
rect 6244 -23826 6296 -23774
rect 6244 -24146 6296 -24094
rect 6244 -24466 6296 -24414
rect 6244 -24786 6296 -24734
rect 6244 -25106 6296 -25054
rect 6244 -25426 6296 -25374
rect 6244 -25746 6296 -25694
rect 6244 -26066 6296 -26014
rect 6244 -26386 6296 -26334
rect 6244 -26706 6296 -26654
rect 6244 -27026 6296 -26974
rect 6244 -27346 6296 -27294
rect 6244 -27666 6296 -27614
rect 6244 -27986 6296 -27934
rect 6244 -28306 6296 -28254
rect 6244 -28626 6296 -28574
rect 6244 -28946 6296 -28894
rect 6244 -29266 6296 -29214
rect 6244 -29586 6296 -29534
rect 6244 -29906 6296 -29854
rect 6244 -30226 6296 -30174
rect 13710 -23826 13762 -23774
rect 13710 -24146 13762 -24094
rect 13710 -24466 13762 -24414
rect 13710 -24786 13762 -24734
rect 13710 -25106 13762 -25054
rect 13710 -25426 13762 -25374
rect 13710 -25746 13762 -25694
rect 13710 -26066 13762 -26014
rect 13710 -26386 13762 -26334
rect 13710 -26706 13762 -26654
rect 13710 -27026 13762 -26974
rect 13710 -27346 13762 -27294
rect 13710 -27666 13762 -27614
rect 13710 -27986 13762 -27934
rect 13710 -28306 13762 -28254
rect 13710 -28626 13762 -28574
rect 13710 -28946 13762 -28894
rect 13710 -29266 13762 -29214
rect 13710 -29586 13762 -29534
rect 13710 -29906 13762 -29854
rect 13710 -30226 13762 -30174
rect 6244 -30546 6296 -30494
rect 13710 -30546 13762 -30494
rect 6614 -30756 6666 -30704
rect 6934 -30756 6986 -30704
rect 7254 -30756 7306 -30704
rect 7574 -30756 7626 -30704
rect 7894 -30756 7946 -30704
rect 8214 -30756 8266 -30704
rect 8534 -30756 8586 -30704
rect 8854 -30756 8906 -30704
rect 9174 -30756 9226 -30704
rect 9494 -30756 9546 -30704
rect 9814 -30756 9866 -30704
rect 10134 -30756 10186 -30704
rect 10454 -30756 10506 -30704
rect 10774 -30756 10826 -30704
rect 11094 -30756 11146 -30704
rect 11414 -30756 11466 -30704
rect 11734 -30756 11786 -30704
rect 12054 -30756 12106 -30704
rect 12374 -30756 12426 -30704
rect 12694 -30756 12746 -30704
rect 13014 -30756 13066 -30704
rect 13334 -30756 13386 -30704
rect 18614 -23300 18666 -23248
rect 18934 -23300 18986 -23248
rect 19254 -23300 19306 -23248
rect 19574 -23300 19626 -23248
rect 19894 -23300 19946 -23248
rect 20214 -23300 20266 -23248
rect 20534 -23300 20586 -23248
rect 20854 -23300 20906 -23248
rect 21174 -23300 21226 -23248
rect 21494 -23300 21546 -23248
rect 21814 -23300 21866 -23248
rect 22134 -23300 22186 -23248
rect 22454 -23300 22506 -23248
rect 22774 -23300 22826 -23248
rect 23094 -23300 23146 -23248
rect 23414 -23300 23466 -23248
rect 23734 -23300 23786 -23248
rect 24054 -23300 24106 -23248
rect 24374 -23300 24426 -23248
rect 24694 -23300 24746 -23248
rect 25014 -23300 25066 -23248
rect 25334 -23300 25386 -23248
rect 18244 -23506 18296 -23454
rect 25710 -23506 25762 -23454
rect 18244 -23826 18296 -23774
rect 18244 -24146 18296 -24094
rect 18244 -24466 18296 -24414
rect 18244 -24786 18296 -24734
rect 18244 -25106 18296 -25054
rect 18244 -25426 18296 -25374
rect 18244 -25746 18296 -25694
rect 18244 -26066 18296 -26014
rect 18244 -26386 18296 -26334
rect 18244 -26706 18296 -26654
rect 18244 -27026 18296 -26974
rect 18244 -27346 18296 -27294
rect 18244 -27666 18296 -27614
rect 18244 -27986 18296 -27934
rect 18244 -28306 18296 -28254
rect 18244 -28626 18296 -28574
rect 18244 -28946 18296 -28894
rect 18244 -29266 18296 -29214
rect 18244 -29586 18296 -29534
rect 18244 -29906 18296 -29854
rect 18244 -30226 18296 -30174
rect 25710 -23826 25762 -23774
rect 25710 -24146 25762 -24094
rect 25710 -24466 25762 -24414
rect 25710 -24786 25762 -24734
rect 25710 -25106 25762 -25054
rect 25710 -25426 25762 -25374
rect 25710 -25746 25762 -25694
rect 25710 -26066 25762 -26014
rect 25710 -26386 25762 -26334
rect 25710 -26706 25762 -26654
rect 25710 -27026 25762 -26974
rect 25710 -27346 25762 -27294
rect 25710 -27666 25762 -27614
rect 25710 -27986 25762 -27934
rect 25710 -28306 25762 -28254
rect 25710 -28626 25762 -28574
rect 25710 -28946 25762 -28894
rect 25710 -29266 25762 -29214
rect 25710 -29586 25762 -29534
rect 25710 -29906 25762 -29854
rect 25710 -30226 25762 -30174
rect 18244 -30546 18296 -30494
rect 25710 -30546 25762 -30494
rect 18614 -30756 18666 -30704
rect 18934 -30756 18986 -30704
rect 19254 -30756 19306 -30704
rect 19574 -30756 19626 -30704
rect 19894 -30756 19946 -30704
rect 20214 -30756 20266 -30704
rect 20534 -30756 20586 -30704
rect 20854 -30756 20906 -30704
rect 21174 -30756 21226 -30704
rect 21494 -30756 21546 -30704
rect 21814 -30756 21866 -30704
rect 22134 -30756 22186 -30704
rect 22454 -30756 22506 -30704
rect 22774 -30756 22826 -30704
rect 23094 -30756 23146 -30704
rect 23414 -30756 23466 -30704
rect 23734 -30756 23786 -30704
rect 24054 -30756 24106 -30704
rect 24374 -30756 24426 -30704
rect 24694 -30756 24746 -30704
rect 25014 -30756 25066 -30704
rect 25334 -30756 25386 -30704
rect 30614 -23300 30666 -23248
rect 30934 -23300 30986 -23248
rect 31254 -23300 31306 -23248
rect 31574 -23300 31626 -23248
rect 31894 -23300 31946 -23248
rect 32214 -23300 32266 -23248
rect 32534 -23300 32586 -23248
rect 32854 -23300 32906 -23248
rect 33174 -23300 33226 -23248
rect 33494 -23300 33546 -23248
rect 33814 -23300 33866 -23248
rect 34134 -23300 34186 -23248
rect 34454 -23300 34506 -23248
rect 34774 -23300 34826 -23248
rect 35094 -23300 35146 -23248
rect 35414 -23300 35466 -23248
rect 35734 -23300 35786 -23248
rect 36054 -23300 36106 -23248
rect 36374 -23300 36426 -23248
rect 36694 -23300 36746 -23248
rect 37014 -23300 37066 -23248
rect 37334 -23300 37386 -23248
rect 30244 -23506 30296 -23454
rect 37710 -23506 37762 -23454
rect 30244 -23826 30296 -23774
rect 30244 -24146 30296 -24094
rect 30244 -24466 30296 -24414
rect 30244 -24786 30296 -24734
rect 30244 -25106 30296 -25054
rect 30244 -25426 30296 -25374
rect 30244 -25746 30296 -25694
rect 30244 -26066 30296 -26014
rect 30244 -26386 30296 -26334
rect 30244 -26706 30296 -26654
rect 30244 -27026 30296 -26974
rect 30244 -27346 30296 -27294
rect 30244 -27666 30296 -27614
rect 30244 -27986 30296 -27934
rect 30244 -28306 30296 -28254
rect 30244 -28626 30296 -28574
rect 30244 -28946 30296 -28894
rect 30244 -29266 30296 -29214
rect 30244 -29586 30296 -29534
rect 30244 -29906 30296 -29854
rect 30244 -30226 30296 -30174
rect 37710 -23826 37762 -23774
rect 37710 -24146 37762 -24094
rect 37710 -24466 37762 -24414
rect 37710 -24786 37762 -24734
rect 37710 -25106 37762 -25054
rect 37710 -25426 37762 -25374
rect 37710 -25746 37762 -25694
rect 37710 -26066 37762 -26014
rect 37710 -26386 37762 -26334
rect 37710 -26706 37762 -26654
rect 37710 -27026 37762 -26974
rect 37710 -27346 37762 -27294
rect 37710 -27666 37762 -27614
rect 37710 -27986 37762 -27934
rect 37710 -28306 37762 -28254
rect 37710 -28626 37762 -28574
rect 37710 -28946 37762 -28894
rect 37710 -29266 37762 -29214
rect 37710 -29586 37762 -29534
rect 37710 -29906 37762 -29854
rect 37710 -30226 37762 -30174
rect 30244 -30546 30296 -30494
rect 37710 -30546 37762 -30494
rect 30614 -30756 30666 -30704
rect 30934 -30756 30986 -30704
rect 31254 -30756 31306 -30704
rect 31574 -30756 31626 -30704
rect 31894 -30756 31946 -30704
rect 32214 -30756 32266 -30704
rect 32534 -30756 32586 -30704
rect 32854 -30756 32906 -30704
rect 33174 -30756 33226 -30704
rect 33494 -30756 33546 -30704
rect 33814 -30756 33866 -30704
rect 34134 -30756 34186 -30704
rect 34454 -30756 34506 -30704
rect 34774 -30756 34826 -30704
rect 35094 -30756 35146 -30704
rect 35414 -30756 35466 -30704
rect 35734 -30756 35786 -30704
rect 36054 -30756 36106 -30704
rect 36374 -30756 36426 -30704
rect 36694 -30756 36746 -30704
rect 37014 -30756 37066 -30704
rect 37334 -30756 37386 -30704
rect 42614 -23300 42666 -23248
rect 42934 -23300 42986 -23248
rect 43254 -23300 43306 -23248
rect 43574 -23300 43626 -23248
rect 43894 -23300 43946 -23248
rect 44214 -23300 44266 -23248
rect 44534 -23300 44586 -23248
rect 44854 -23300 44906 -23248
rect 45174 -23300 45226 -23248
rect 45494 -23300 45546 -23248
rect 45814 -23300 45866 -23248
rect 46134 -23300 46186 -23248
rect 46454 -23300 46506 -23248
rect 46774 -23300 46826 -23248
rect 47094 -23300 47146 -23248
rect 47414 -23300 47466 -23248
rect 47734 -23300 47786 -23248
rect 48054 -23300 48106 -23248
rect 48374 -23300 48426 -23248
rect 48694 -23300 48746 -23248
rect 49014 -23300 49066 -23248
rect 49334 -23300 49386 -23248
rect 42244 -23506 42296 -23454
rect 49710 -23506 49762 -23454
rect 42244 -23826 42296 -23774
rect 42244 -24146 42296 -24094
rect 42244 -24466 42296 -24414
rect 42244 -24786 42296 -24734
rect 42244 -25106 42296 -25054
rect 42244 -25426 42296 -25374
rect 42244 -25746 42296 -25694
rect 42244 -26066 42296 -26014
rect 42244 -26386 42296 -26334
rect 42244 -26706 42296 -26654
rect 42244 -27026 42296 -26974
rect 42244 -27346 42296 -27294
rect 42244 -27666 42296 -27614
rect 42244 -27986 42296 -27934
rect 42244 -28306 42296 -28254
rect 42244 -28626 42296 -28574
rect 42244 -28946 42296 -28894
rect 42244 -29266 42296 -29214
rect 42244 -29586 42296 -29534
rect 42244 -29906 42296 -29854
rect 42244 -30226 42296 -30174
rect 49710 -23826 49762 -23774
rect 49710 -24146 49762 -24094
rect 49710 -24466 49762 -24414
rect 49710 -24786 49762 -24734
rect 49710 -25106 49762 -25054
rect 49710 -25426 49762 -25374
rect 49710 -25746 49762 -25694
rect 49710 -26066 49762 -26014
rect 49710 -26386 49762 -26334
rect 49710 -26706 49762 -26654
rect 49710 -27026 49762 -26974
rect 49710 -27346 49762 -27294
rect 49710 -27666 49762 -27614
rect 49710 -27986 49762 -27934
rect 49710 -28306 49762 -28254
rect 49710 -28626 49762 -28574
rect 49710 -28946 49762 -28894
rect 49710 -29266 49762 -29214
rect 49710 -29586 49762 -29534
rect 49710 -29906 49762 -29854
rect 49710 -30226 49762 -30174
rect 42244 -30546 42296 -30494
rect 49710 -30546 49762 -30494
rect 42614 -30756 42666 -30704
rect 42934 -30756 42986 -30704
rect 43254 -30756 43306 -30704
rect 43574 -30756 43626 -30704
rect 43894 -30756 43946 -30704
rect 44214 -30756 44266 -30704
rect 44534 -30756 44586 -30704
rect 44854 -30756 44906 -30704
rect 45174 -30756 45226 -30704
rect 45494 -30756 45546 -30704
rect 45814 -30756 45866 -30704
rect 46134 -30756 46186 -30704
rect 46454 -30756 46506 -30704
rect 46774 -30756 46826 -30704
rect 47094 -30756 47146 -30704
rect 47414 -30756 47466 -30704
rect 47734 -30756 47786 -30704
rect 48054 -30756 48106 -30704
rect 48374 -30756 48426 -30704
rect 48694 -30756 48746 -30704
rect 49014 -30756 49066 -30704
rect 49334 -30756 49386 -30704
<< metal2 >>
rect 18200 -2500 21600 -2400
rect 18200 -2900 18300 -2500
rect 18110 -3000 18300 -2900
rect 21500 -2900 21600 -2500
rect 21800 -2900 23400 -2800
rect 21500 -3000 23400 -2900
rect 18110 -3100 21894 -3000
rect 18110 -3164 18210 -3100
rect 18602 -3164 18702 -3100
rect 19002 -3164 19102 -3100
rect 19402 -3164 19502 -3100
rect 19802 -3164 19902 -3100
rect 20102 -3164 20202 -3100
rect 20502 -3164 20602 -3100
rect 20902 -3164 21002 -3100
rect 21302 -3164 21402 -3100
rect 21794 -3164 21894 -3100
rect 18088 -3266 21916 -3164
rect 18088 -3427 18140 -3266
rect 18088 -5415 18140 -5403
rect 18206 -3427 18258 -3415
rect 18206 -5512 18258 -5403
rect 18324 -3427 18376 -3266
rect 18324 -5415 18376 -5403
rect 18442 -3427 18494 -3415
rect 18442 -5512 18494 -5403
rect 18560 -3427 18612 -3266
rect 18560 -5415 18612 -5403
rect 18678 -3427 18730 -3415
rect 18678 -5512 18730 -5403
rect 18796 -3427 18848 -3266
rect 18796 -5415 18848 -5403
rect 18914 -3427 18966 -3415
rect 18914 -5512 18966 -5403
rect 19032 -3427 19084 -3266
rect 19032 -5415 19084 -5403
rect 19150 -3427 19202 -3415
rect 18206 -5564 18966 -5512
rect 19150 -5512 19202 -5403
rect 19268 -3427 19320 -3266
rect 19268 -5415 19320 -5403
rect 19386 -3427 19438 -3415
rect 19386 -5512 19438 -5403
rect 19504 -3427 19556 -3266
rect 19504 -5415 19556 -5403
rect 19622 -3427 19674 -3415
rect 19622 -5415 19674 -5403
rect 19740 -3427 19792 -3266
rect 19740 -5415 19792 -5403
rect 19858 -3427 19910 -3415
rect 19858 -5422 19910 -5403
rect 19976 -3427 20028 -3266
rect 19976 -5416 20028 -5403
rect 20094 -3427 20146 -3415
rect 19858 -5512 19890 -5422
rect 20094 -5444 20146 -5403
rect 20212 -3427 20264 -3266
rect 20212 -5415 20264 -5403
rect 20330 -3427 20382 -3415
rect 20330 -5415 20382 -5403
rect 20448 -3427 20500 -3266
rect 20448 -5415 20500 -5403
rect 20566 -3427 20618 -3415
rect 19942 -5450 20148 -5444
rect 19150 -5542 19890 -5512
rect 19918 -5456 20148 -5450
rect 19970 -5472 20148 -5456
rect 19918 -5514 19970 -5508
rect 20027 -5542 20033 -5500
rect 19150 -5552 20033 -5542
rect 20085 -5552 20091 -5500
rect 19150 -5564 20091 -5552
rect 20119 -5512 20148 -5472
rect 20566 -5510 20618 -5403
rect 20684 -3427 20736 -3266
rect 20802 -3427 20854 -3415
rect 20684 -5415 20736 -5403
rect 20801 -5403 20802 -5335
rect 20801 -5415 20854 -5403
rect 20920 -3427 20972 -3266
rect 21038 -3427 21090 -3415
rect 20920 -5415 20972 -5403
rect 21037 -5403 21038 -5335
rect 21037 -5415 21090 -5403
rect 21156 -3427 21208 -3266
rect 21274 -3427 21326 -3415
rect 21156 -5415 21208 -5403
rect 21273 -5403 21274 -5335
rect 21273 -5415 21326 -5403
rect 21392 -3427 21444 -3266
rect 21510 -3427 21562 -3415
rect 21392 -5415 21444 -5403
rect 21509 -5403 21510 -5335
rect 21509 -5415 21562 -5403
rect 21628 -3427 21680 -3266
rect 21746 -3427 21798 -3415
rect 21628 -5415 21680 -5403
rect 21745 -5403 21746 -5335
rect 20382 -5511 20618 -5510
rect 20801 -5511 20853 -5415
rect 20382 -5512 20853 -5511
rect 20119 -5562 20853 -5512
rect 20119 -5564 20382 -5562
rect 20566 -5563 20853 -5562
rect 21037 -5512 21089 -5415
rect 21273 -5512 21325 -5415
rect 21509 -5512 21561 -5415
rect 21745 -5512 21798 -5403
rect 21864 -3427 21916 -3266
rect 21864 -5415 21916 -5403
rect 18442 -5634 18494 -5564
rect 18087 -5686 18494 -5634
rect 18087 -5731 18139 -5686
rect 18323 -5731 18375 -5686
rect 18087 -5740 18375 -5731
rect 18087 -5796 18203 -5740
rect 18259 -5796 18375 -5740
rect 18087 -5805 18375 -5796
rect 17851 -5936 17903 -5924
rect 17851 -8064 17903 -7912
rect 17969 -5936 18021 -5924
rect 17969 -8064 18021 -7912
rect 18087 -5936 18139 -5805
rect 18087 -7924 18139 -7912
rect 18205 -5936 18257 -5924
rect 18205 -8064 18257 -7912
rect 18323 -5936 18375 -5805
rect 19386 -5890 19438 -5564
rect 19858 -5570 20091 -5564
rect 20566 -5890 20618 -5563
rect 21037 -5564 21798 -5512
rect 21872 -5560 22002 -5550
rect 21509 -5634 21561 -5564
rect 21872 -5634 21882 -5560
rect 21509 -5650 21882 -5634
rect 21992 -5650 22002 -5560
rect 21509 -5686 22002 -5650
rect 18323 -7924 18375 -7912
rect 18441 -5936 18493 -5924
rect 18441 -8040 18493 -7912
rect 18559 -5936 18611 -5924
rect 19297 -6030 19939 -5890
rect 19297 -6100 19363 -6030
rect 19489 -6100 19555 -6030
rect 19681 -6100 19747 -6030
rect 19873 -6100 19939 -6030
rect 20065 -6030 20707 -5890
rect 20065 -6100 20131 -6030
rect 20257 -6100 20323 -6030
rect 20449 -6100 20515 -6030
rect 20641 -6100 20707 -6030
rect 21392 -5936 21444 -5924
rect 19009 -6600 19015 -6100
rect 19069 -6600 19075 -6100
rect 19105 -6600 19111 -6100
rect 19165 -6600 19171 -6100
rect 19201 -6600 19207 -6100
rect 19261 -6600 19267 -6100
rect 19297 -6600 19303 -6100
rect 19357 -6600 19363 -6100
rect 19393 -6600 19399 -6100
rect 19453 -6600 19459 -6100
rect 19489 -6600 19495 -6100
rect 19549 -6600 19555 -6100
rect 19585 -6600 19591 -6100
rect 19645 -6600 19651 -6100
rect 19681 -6600 19687 -6100
rect 19741 -6600 19747 -6100
rect 19777 -6600 19783 -6100
rect 19837 -6600 19843 -6100
rect 19873 -6600 19879 -6100
rect 19933 -6600 19939 -6100
rect 19969 -6600 19975 -6100
rect 20029 -6600 20035 -6100
rect 20065 -6600 20071 -6100
rect 20125 -6600 20131 -6100
rect 20161 -6600 20167 -6100
rect 20221 -6600 20227 -6100
rect 20257 -6600 20263 -6100
rect 20317 -6600 20323 -6100
rect 20353 -6600 20359 -6100
rect 20413 -6600 20419 -6100
rect 20449 -6600 20455 -6100
rect 20509 -6600 20515 -6100
rect 20545 -6600 20551 -6100
rect 20605 -6600 20611 -6100
rect 20641 -6600 20647 -6100
rect 20701 -6600 20707 -6100
rect 20737 -6600 20743 -6100
rect 20797 -6600 20803 -6100
rect 20833 -6600 20839 -6100
rect 20893 -6600 20899 -6100
rect 20929 -6600 20935 -6100
rect 20989 -6600 20995 -6100
rect 19207 -6760 19261 -6600
rect 19297 -6644 19363 -6638
rect 19297 -6720 19363 -6706
rect 19399 -6760 19453 -6600
rect 19489 -6644 19555 -6638
rect 19489 -6720 19555 -6706
rect 19591 -6760 19645 -6600
rect 19681 -6644 19747 -6638
rect 19681 -6720 19747 -6706
rect 19783 -6760 19837 -6600
rect 19873 -6644 19939 -6638
rect 19873 -6720 19939 -6706
rect 19975 -6760 20029 -6600
rect 20065 -6644 20131 -6638
rect 20065 -6720 20131 -6706
rect 20167 -6760 20221 -6600
rect 20257 -6644 20323 -6638
rect 20257 -6720 20323 -6706
rect 20359 -6760 20413 -6600
rect 20449 -6644 20515 -6638
rect 20449 -6720 20515 -6706
rect 20551 -6760 20605 -6600
rect 20641 -6644 20707 -6638
rect 20641 -6720 20707 -6706
rect 20743 -6760 20797 -6600
rect 19207 -6830 20797 -6760
rect 19207 -6916 19261 -6830
rect 19399 -6916 19453 -6830
rect 19591 -6916 19645 -6830
rect 19783 -6916 19837 -6830
rect 19975 -6916 20029 -6830
rect 20167 -6916 20221 -6830
rect 20359 -6916 20413 -6830
rect 20551 -6916 20605 -6830
rect 20743 -6916 20797 -6830
rect 18800 -6938 19122 -6930
rect 18800 -6940 19058 -6938
rect 18800 -7000 18810 -6940
rect 18970 -7000 19058 -6940
rect 18800 -7002 19058 -7000
rect 18800 -7010 19122 -7002
rect 19207 -7008 20797 -6916
rect 18559 -8040 18611 -7912
rect 19060 -7052 19112 -7040
rect 18441 -8060 18902 -8040
rect 18441 -8064 18822 -8060
rect 17802 -8134 18822 -8064
rect 16900 -8268 17150 -8249
rect 16900 -8485 16920 -8268
rect 17130 -8485 17150 -8268
rect 17802 -8300 17902 -8134
rect 18002 -8300 18102 -8134
rect 18202 -8300 18302 -8134
rect 18402 -8140 18822 -8134
rect 18402 -8300 18502 -8140
rect 18602 -8300 18702 -8140
rect 18802 -8300 18822 -8140
rect 16649 -8537 16666 -8485
rect 17135 -8537 17150 -8485
rect 17380 -8440 17620 -8420
rect 16567 -9170 16590 -9100
rect 17019 -9170 17038 -9100
rect 16600 -9348 16800 -9170
rect 16600 -9510 16680 -9348
rect 17380 -9360 17400 -8440
rect 17600 -9200 17620 -8440
rect 17760 -8500 18822 -8300
rect 17760 -8800 18702 -8500
rect 18802 -8800 18822 -8500
rect 17760 -8900 18822 -8800
rect 17760 -9200 18702 -8900
rect 18802 -9200 18822 -8900
rect 17600 -9280 18822 -9200
rect 18882 -9200 18902 -8060
rect 19060 -9180 19112 -9028
rect 19518 -7052 19570 -7008
rect 19518 -9040 19570 -9028
rect 19976 -7052 20028 -7040
rect 19976 -9180 20028 -9028
rect 20434 -7052 20486 -7008
rect 20434 -9040 20486 -9028
rect 20892 -7052 20944 -7040
rect 21392 -8040 21444 -7912
rect 21510 -5936 21562 -5924
rect 21510 -8040 21562 -7912
rect 21628 -5936 21680 -5686
rect 21741 -5740 21802 -5731
rect 21741 -5796 21744 -5740
rect 21800 -5796 21802 -5740
rect 21741 -5805 21802 -5796
rect 21628 -7924 21680 -7912
rect 21746 -5936 21798 -5924
rect 20892 -9180 20944 -9028
rect 19060 -9200 20944 -9180
rect 21102 -8060 21562 -8040
rect 21102 -9200 21122 -8060
rect 18882 -9280 21122 -9200
rect 21182 -8064 21562 -8060
rect 21746 -8064 21798 -7912
rect 21864 -5936 21916 -5686
rect 21864 -7924 21916 -7912
rect 21982 -5936 22034 -5924
rect 21982 -8064 22034 -7912
rect 22100 -5936 22152 -5924
rect 22452 -6270 22602 -6250
rect 22452 -6660 22472 -6270
rect 22582 -6660 22602 -6270
rect 22452 -6680 22602 -6660
rect 22682 -6270 22832 -6250
rect 22682 -6660 22702 -6270
rect 22812 -6660 22832 -6270
rect 22682 -6680 22832 -6660
rect 23200 -7200 23400 -3000
rect 23200 -7400 23300 -7200
rect 23500 -7400 23600 -7200
rect 23260 -7480 23420 -7470
rect 23260 -7540 23270 -7480
rect 23410 -7540 23420 -7480
rect 23260 -7640 23420 -7540
rect 23260 -7720 23270 -7640
rect 23410 -7720 23420 -7640
rect 23540 -7720 23550 -7640
rect 23690 -7720 23700 -7640
rect 23540 -7800 23700 -7720
rect 23540 -7860 23550 -7800
rect 23690 -7860 23700 -7800
rect 23540 -7870 23700 -7860
rect 22100 -8064 22152 -7912
rect 21182 -8134 22152 -8064
rect 23200 -8100 23300 -7900
rect 23500 -8100 23600 -7900
rect 21182 -8140 21602 -8134
rect 21182 -8400 21202 -8140
rect 21302 -8300 21402 -8140
rect 21502 -8300 21602 -8140
rect 21702 -8300 21802 -8134
rect 21902 -8300 22002 -8134
rect 23200 -8300 23400 -8100
rect 21302 -8400 23400 -8300
rect 21182 -8500 23400 -8400
rect 21182 -8800 21202 -8500
rect 21302 -8800 22200 -8500
rect 21182 -8900 22200 -8800
rect 21182 -9200 21202 -8900
rect 21302 -9200 22200 -8900
rect 21182 -9280 22200 -9200
rect 17600 -9360 22200 -9280
rect 17380 -9500 22200 -9360
rect 16390 -9520 16470 -9510
rect 16390 -9580 16400 -9520
rect 16460 -9580 16470 -9520
rect 16390 -9590 16470 -9580
rect 16600 -9570 16610 -9510
rect 16670 -9570 16680 -9510
rect 16600 -9584 16680 -9570
rect 16460 -9660 16540 -9650
rect 16460 -9720 16470 -9660
rect 16530 -9720 16540 -9660
rect 16460 -9730 16540 -9720
rect 15950 -10510 16810 -10500
rect 15950 -10850 16710 -10510
rect 16800 -10850 16810 -10510
rect 17410 -10510 17520 -9500
rect 17600 -9600 19000 -9500
rect 17600 -10200 17700 -9600
rect 18900 -10200 19000 -9600
rect 17600 -10300 19000 -10200
rect 20800 -9600 22200 -9500
rect 20800 -10200 20900 -9600
rect 22100 -10200 22200 -9600
rect 20800 -10300 22200 -10200
rect 17020 -10620 17140 -10610
rect 17020 -10740 17030 -10620
rect 17130 -10740 17140 -10620
rect 17020 -10750 17140 -10740
rect 15950 -10860 16810 -10850
rect 17410 -10850 17420 -10510
rect 17510 -10850 17520 -10510
rect 17410 -10860 17520 -10850
rect 6000 -11110 14000 -11000
rect 15950 -11110 16170 -10860
rect 6000 -11246 16170 -11110
rect 6000 -11302 6612 -11246
rect 6668 -11302 6932 -11246
rect 6988 -11302 7252 -11246
rect 7308 -11302 7572 -11246
rect 7628 -11302 7892 -11246
rect 7948 -11302 8212 -11246
rect 8268 -11302 8532 -11246
rect 8588 -11302 8852 -11246
rect 8908 -11302 9172 -11246
rect 9228 -11302 9492 -11246
rect 9548 -11302 9812 -11246
rect 9868 -11302 10132 -11246
rect 10188 -11302 10452 -11246
rect 10508 -11302 10772 -11246
rect 10828 -11302 11092 -11246
rect 11148 -11302 11412 -11246
rect 11468 -11302 11732 -11246
rect 11788 -11302 12052 -11246
rect 12108 -11302 12372 -11246
rect 12428 -11302 12692 -11246
rect 12748 -11302 13012 -11246
rect 13068 -11302 13332 -11246
rect 13388 -11302 16170 -11246
rect 6000 -11310 16170 -11302
rect 18000 -11246 26000 -11000
rect 18000 -11302 18612 -11246
rect 18668 -11302 18932 -11246
rect 18988 -11302 19252 -11246
rect 19308 -11302 19572 -11246
rect 19628 -11302 19892 -11246
rect 19948 -11302 20212 -11246
rect 20268 -11302 20532 -11246
rect 20588 -11302 20852 -11246
rect 20908 -11302 21172 -11246
rect 21228 -11302 21492 -11246
rect 21548 -11302 21812 -11246
rect 21868 -11302 22132 -11246
rect 22188 -11302 22452 -11246
rect 22508 -11302 22772 -11246
rect 22828 -11302 23092 -11246
rect 23148 -11302 23412 -11246
rect 23468 -11302 23732 -11246
rect 23788 -11302 24052 -11246
rect 24108 -11302 24372 -11246
rect 24428 -11302 24692 -11246
rect 24748 -11302 25012 -11246
rect 25068 -11302 25332 -11246
rect 25388 -11302 26000 -11246
rect 6000 -11452 14000 -11310
rect 6000 -11508 6242 -11452
rect 6298 -11508 13708 -11452
rect 13764 -11508 14000 -11452
rect 6000 -11540 14000 -11508
rect 6000 -11772 6540 -11540
rect 6000 -11828 6242 -11772
rect 6298 -11828 6540 -11772
rect 6000 -12092 6540 -11828
rect 6000 -12148 6242 -12092
rect 6298 -12148 6540 -12092
rect 6000 -12412 6540 -12148
rect 6000 -12468 6242 -12412
rect 6298 -12468 6540 -12412
rect 6000 -12732 6540 -12468
rect 6000 -12788 6242 -12732
rect 6298 -12788 6540 -12732
rect 6000 -13052 6540 -12788
rect 6000 -13108 6242 -13052
rect 6298 -13108 6540 -13052
rect 6000 -13372 6540 -13108
rect 6000 -13428 6242 -13372
rect 6298 -13428 6540 -13372
rect 6000 -13692 6540 -13428
rect 6000 -13748 6242 -13692
rect 6298 -13748 6540 -13692
rect 6000 -14012 6540 -13748
rect 6000 -14068 6242 -14012
rect 6298 -14068 6540 -14012
rect 6000 -14332 6540 -14068
rect 6000 -14388 6242 -14332
rect 6298 -14388 6540 -14332
rect 6000 -14652 6540 -14388
rect 6000 -14708 6242 -14652
rect 6298 -14708 6540 -14652
rect 6000 -14972 6540 -14708
rect 6000 -15028 6242 -14972
rect 6298 -15028 6540 -14972
rect 6000 -15292 6540 -15028
rect 6000 -15348 6242 -15292
rect 6298 -15348 6540 -15292
rect 6000 -15612 6540 -15348
rect 6000 -15668 6242 -15612
rect 6298 -15668 6540 -15612
rect 6000 -15932 6540 -15668
rect 6000 -15988 6242 -15932
rect 6298 -15988 6540 -15932
rect 6000 -16252 6540 -15988
rect 6000 -16308 6242 -16252
rect 6298 -16308 6540 -16252
rect 6000 -16572 6540 -16308
rect 6000 -16628 6242 -16572
rect 6298 -16628 6540 -16572
rect 6000 -16892 6540 -16628
rect 6000 -16948 6242 -16892
rect 6298 -16948 6540 -16892
rect 6000 -17212 6540 -16948
rect 6000 -17268 6242 -17212
rect 6298 -17268 6540 -17212
rect 6000 -17532 6540 -17268
rect 6000 -17588 6242 -17532
rect 6298 -17588 6540 -17532
rect 6000 -17852 6540 -17588
rect 6000 -17908 6242 -17852
rect 6298 -17908 6540 -17852
rect 6000 -18172 6540 -17908
rect 6000 -18228 6242 -18172
rect 6298 -18228 6540 -18172
rect 6000 -18460 6540 -18228
rect 13460 -11772 14000 -11540
rect 13460 -11828 13708 -11772
rect 13764 -11828 14000 -11772
rect 13460 -12092 14000 -11828
rect 13460 -12148 13708 -12092
rect 13764 -12148 14000 -12092
rect 13460 -12412 14000 -12148
rect 13460 -12468 13708 -12412
rect 13764 -12468 14000 -12412
rect 13460 -12732 14000 -12468
rect 13460 -12788 13708 -12732
rect 13764 -12788 14000 -12732
rect 13460 -13052 14000 -12788
rect 13460 -13108 13708 -13052
rect 13764 -13108 14000 -13052
rect 13460 -13372 14000 -13108
rect 13460 -13428 13708 -13372
rect 13764 -13428 14000 -13372
rect 13460 -13692 14000 -13428
rect 13460 -13748 13708 -13692
rect 13764 -13748 14000 -13692
rect 13460 -14012 14000 -13748
rect 13460 -14068 13708 -14012
rect 13764 -14068 14000 -14012
rect 13460 -14332 14000 -14068
rect 13460 -14388 13708 -14332
rect 13764 -14388 14000 -14332
rect 13460 -14652 14000 -14388
rect 13460 -14708 13708 -14652
rect 13764 -14708 14000 -14652
rect 13460 -14972 14000 -14708
rect 13460 -15028 13708 -14972
rect 13764 -15028 14000 -14972
rect 13460 -15292 14000 -15028
rect 13460 -15348 13708 -15292
rect 13764 -15348 14000 -15292
rect 13460 -15612 14000 -15348
rect 13460 -15668 13708 -15612
rect 13764 -15668 14000 -15612
rect 13460 -15932 14000 -15668
rect 13460 -15988 13708 -15932
rect 13764 -15988 14000 -15932
rect 13460 -16252 14000 -15988
rect 13460 -16308 13708 -16252
rect 13764 -16308 14000 -16252
rect 13460 -16572 14000 -16308
rect 13460 -16628 13708 -16572
rect 13764 -16628 14000 -16572
rect 13460 -16892 14000 -16628
rect 13460 -16948 13708 -16892
rect 13764 -16948 14000 -16892
rect 13460 -17212 14000 -16948
rect 13460 -17268 13708 -17212
rect 13764 -17268 14000 -17212
rect 13460 -17532 14000 -17268
rect 13460 -17588 13708 -17532
rect 13764 -17588 14000 -17532
rect 13460 -17852 14000 -17588
rect 13460 -17908 13708 -17852
rect 13764 -17908 14000 -17852
rect 13460 -18172 14000 -17908
rect 13460 -18228 13708 -18172
rect 13764 -18228 14000 -18172
rect 13460 -18460 14000 -18228
rect 6000 -18492 14000 -18460
rect 6000 -18548 6242 -18492
rect 6298 -18548 13708 -18492
rect 13764 -18548 14000 -18492
rect 6000 -18702 14000 -18548
rect 6000 -18758 6612 -18702
rect 6668 -18758 6932 -18702
rect 6988 -18758 7252 -18702
rect 7308 -18758 7572 -18702
rect 7628 -18758 7892 -18702
rect 7948 -18758 8212 -18702
rect 8268 -18758 8532 -18702
rect 8588 -18758 8852 -18702
rect 8908 -18758 9172 -18702
rect 9228 -18758 9492 -18702
rect 9548 -18758 9812 -18702
rect 9868 -18758 10132 -18702
rect 10188 -18758 10452 -18702
rect 10508 -18758 10772 -18702
rect 10828 -18758 11092 -18702
rect 11148 -18758 11412 -18702
rect 11468 -18758 11732 -18702
rect 11788 -18758 12052 -18702
rect 12108 -18758 12372 -18702
rect 12428 -18758 12692 -18702
rect 12748 -18758 13012 -18702
rect 13068 -18758 13332 -18702
rect 13388 -18758 14000 -18702
rect 6000 -19000 14000 -18758
rect 18000 -11452 26000 -11302
rect 18000 -11508 18242 -11452
rect 18298 -11508 25708 -11452
rect 25764 -11508 26000 -11452
rect 18000 -11540 26000 -11508
rect 18000 -11772 18540 -11540
rect 18000 -11828 18242 -11772
rect 18298 -11828 18540 -11772
rect 18000 -12092 18540 -11828
rect 18000 -12148 18242 -12092
rect 18298 -12148 18540 -12092
rect 18000 -12412 18540 -12148
rect 18000 -12468 18242 -12412
rect 18298 -12468 18540 -12412
rect 18000 -12732 18540 -12468
rect 18000 -12788 18242 -12732
rect 18298 -12788 18540 -12732
rect 18000 -13052 18540 -12788
rect 18000 -13108 18242 -13052
rect 18298 -13108 18540 -13052
rect 18000 -13372 18540 -13108
rect 18000 -13428 18242 -13372
rect 18298 -13428 18540 -13372
rect 18000 -13692 18540 -13428
rect 18000 -13748 18242 -13692
rect 18298 -13748 18540 -13692
rect 18000 -14012 18540 -13748
rect 18000 -14068 18242 -14012
rect 18298 -14068 18540 -14012
rect 18000 -14332 18540 -14068
rect 18000 -14388 18242 -14332
rect 18298 -14388 18540 -14332
rect 18000 -14652 18540 -14388
rect 18000 -14708 18242 -14652
rect 18298 -14708 18540 -14652
rect 18000 -14972 18540 -14708
rect 18000 -15028 18242 -14972
rect 18298 -15028 18540 -14972
rect 18000 -15292 18540 -15028
rect 18000 -15348 18242 -15292
rect 18298 -15348 18540 -15292
rect 18000 -15612 18540 -15348
rect 18000 -15668 18242 -15612
rect 18298 -15668 18540 -15612
rect 18000 -15932 18540 -15668
rect 18000 -15988 18242 -15932
rect 18298 -15988 18540 -15932
rect 18000 -16252 18540 -15988
rect 18000 -16308 18242 -16252
rect 18298 -16308 18540 -16252
rect 18000 -16572 18540 -16308
rect 18000 -16628 18242 -16572
rect 18298 -16628 18540 -16572
rect 18000 -16892 18540 -16628
rect 18000 -16948 18242 -16892
rect 18298 -16948 18540 -16892
rect 18000 -17212 18540 -16948
rect 18000 -17268 18242 -17212
rect 18298 -17268 18540 -17212
rect 18000 -17532 18540 -17268
rect 18000 -17588 18242 -17532
rect 18298 -17588 18540 -17532
rect 18000 -17852 18540 -17588
rect 18000 -17908 18242 -17852
rect 18298 -17908 18540 -17852
rect 18000 -18172 18540 -17908
rect 18000 -18228 18242 -18172
rect 18298 -18228 18540 -18172
rect 18000 -18460 18540 -18228
rect 25460 -11772 26000 -11540
rect 25460 -11828 25708 -11772
rect 25764 -11828 26000 -11772
rect 25460 -12092 26000 -11828
rect 25460 -12148 25708 -12092
rect 25764 -12148 26000 -12092
rect 25460 -12412 26000 -12148
rect 25460 -12468 25708 -12412
rect 25764 -12468 26000 -12412
rect 25460 -12732 26000 -12468
rect 25460 -12788 25708 -12732
rect 25764 -12788 26000 -12732
rect 25460 -13052 26000 -12788
rect 25460 -13108 25708 -13052
rect 25764 -13108 26000 -13052
rect 25460 -13372 26000 -13108
rect 25460 -13428 25708 -13372
rect 25764 -13428 26000 -13372
rect 25460 -13692 26000 -13428
rect 25460 -13748 25708 -13692
rect 25764 -13748 26000 -13692
rect 25460 -14012 26000 -13748
rect 25460 -14068 25708 -14012
rect 25764 -14068 26000 -14012
rect 25460 -14332 26000 -14068
rect 25460 -14388 25708 -14332
rect 25764 -14388 26000 -14332
rect 25460 -14652 26000 -14388
rect 25460 -14708 25708 -14652
rect 25764 -14708 26000 -14652
rect 25460 -14972 26000 -14708
rect 25460 -15028 25708 -14972
rect 25764 -15028 26000 -14972
rect 25460 -15292 26000 -15028
rect 25460 -15348 25708 -15292
rect 25764 -15348 26000 -15292
rect 25460 -15612 26000 -15348
rect 25460 -15668 25708 -15612
rect 25764 -15668 26000 -15612
rect 25460 -15932 26000 -15668
rect 25460 -15988 25708 -15932
rect 25764 -15988 26000 -15932
rect 25460 -16252 26000 -15988
rect 25460 -16308 25708 -16252
rect 25764 -16308 26000 -16252
rect 25460 -16572 26000 -16308
rect 25460 -16628 25708 -16572
rect 25764 -16628 26000 -16572
rect 25460 -16892 26000 -16628
rect 25460 -16948 25708 -16892
rect 25764 -16948 26000 -16892
rect 25460 -17212 26000 -16948
rect 25460 -17268 25708 -17212
rect 25764 -17268 26000 -17212
rect 25460 -17532 26000 -17268
rect 25460 -17588 25708 -17532
rect 25764 -17588 26000 -17532
rect 25460 -17852 26000 -17588
rect 25460 -17908 25708 -17852
rect 25764 -17908 26000 -17852
rect 25460 -18172 26000 -17908
rect 25460 -18228 25708 -18172
rect 25764 -18228 26000 -18172
rect 25460 -18460 26000 -18228
rect 18000 -18492 26000 -18460
rect 18000 -18548 18242 -18492
rect 18298 -18548 25708 -18492
rect 25764 -18548 26000 -18492
rect 18000 -18702 26000 -18548
rect 18000 -18758 18612 -18702
rect 18668 -18758 18932 -18702
rect 18988 -18758 19252 -18702
rect 19308 -18758 19572 -18702
rect 19628 -18758 19892 -18702
rect 19948 -18758 20212 -18702
rect 20268 -18758 20532 -18702
rect 20588 -18758 20852 -18702
rect 20908 -18758 21172 -18702
rect 21228 -18758 21492 -18702
rect 21548 -18758 21812 -18702
rect 21868 -18758 22132 -18702
rect 22188 -18758 22452 -18702
rect 22508 -18758 22772 -18702
rect 22828 -18758 23092 -18702
rect 23148 -18758 23412 -18702
rect 23468 -18758 23732 -18702
rect 23788 -18758 24052 -18702
rect 24108 -18758 24372 -18702
rect 24428 -18758 24692 -18702
rect 24748 -18758 25012 -18702
rect 25068 -18758 25332 -18702
rect 25388 -18758 26000 -18702
rect 18000 -19000 26000 -18758
rect 30000 -11246 38000 -11000
rect 30000 -11302 30612 -11246
rect 30668 -11302 30932 -11246
rect 30988 -11302 31252 -11246
rect 31308 -11302 31572 -11246
rect 31628 -11302 31892 -11246
rect 31948 -11302 32212 -11246
rect 32268 -11302 32532 -11246
rect 32588 -11302 32852 -11246
rect 32908 -11302 33172 -11246
rect 33228 -11302 33492 -11246
rect 33548 -11302 33812 -11246
rect 33868 -11302 34132 -11246
rect 34188 -11302 34452 -11246
rect 34508 -11302 34772 -11246
rect 34828 -11302 35092 -11246
rect 35148 -11302 35412 -11246
rect 35468 -11302 35732 -11246
rect 35788 -11302 36052 -11246
rect 36108 -11302 36372 -11246
rect 36428 -11302 36692 -11246
rect 36748 -11302 37012 -11246
rect 37068 -11302 37332 -11246
rect 37388 -11302 38000 -11246
rect 30000 -11452 38000 -11302
rect 30000 -11508 30242 -11452
rect 30298 -11508 37708 -11452
rect 37764 -11508 38000 -11452
rect 30000 -11540 38000 -11508
rect 30000 -11772 30540 -11540
rect 30000 -11828 30242 -11772
rect 30298 -11828 30540 -11772
rect 30000 -12092 30540 -11828
rect 30000 -12148 30242 -12092
rect 30298 -12148 30540 -12092
rect 30000 -12412 30540 -12148
rect 30000 -12468 30242 -12412
rect 30298 -12468 30540 -12412
rect 30000 -12732 30540 -12468
rect 30000 -12788 30242 -12732
rect 30298 -12788 30540 -12732
rect 30000 -13052 30540 -12788
rect 30000 -13108 30242 -13052
rect 30298 -13108 30540 -13052
rect 30000 -13372 30540 -13108
rect 30000 -13428 30242 -13372
rect 30298 -13428 30540 -13372
rect 30000 -13692 30540 -13428
rect 30000 -13748 30242 -13692
rect 30298 -13748 30540 -13692
rect 30000 -14012 30540 -13748
rect 30000 -14068 30242 -14012
rect 30298 -14068 30540 -14012
rect 30000 -14332 30540 -14068
rect 30000 -14388 30242 -14332
rect 30298 -14388 30540 -14332
rect 30000 -14652 30540 -14388
rect 30000 -14708 30242 -14652
rect 30298 -14708 30540 -14652
rect 30000 -14972 30540 -14708
rect 30000 -15028 30242 -14972
rect 30298 -15028 30540 -14972
rect 30000 -15292 30540 -15028
rect 30000 -15348 30242 -15292
rect 30298 -15348 30540 -15292
rect 30000 -15612 30540 -15348
rect 30000 -15668 30242 -15612
rect 30298 -15668 30540 -15612
rect 30000 -15932 30540 -15668
rect 30000 -15988 30242 -15932
rect 30298 -15988 30540 -15932
rect 30000 -16252 30540 -15988
rect 30000 -16308 30242 -16252
rect 30298 -16308 30540 -16252
rect 30000 -16572 30540 -16308
rect 30000 -16628 30242 -16572
rect 30298 -16628 30540 -16572
rect 30000 -16892 30540 -16628
rect 30000 -16948 30242 -16892
rect 30298 -16948 30540 -16892
rect 30000 -17212 30540 -16948
rect 30000 -17268 30242 -17212
rect 30298 -17268 30540 -17212
rect 30000 -17532 30540 -17268
rect 30000 -17588 30242 -17532
rect 30298 -17588 30540 -17532
rect 30000 -17852 30540 -17588
rect 30000 -17908 30242 -17852
rect 30298 -17908 30540 -17852
rect 30000 -18172 30540 -17908
rect 30000 -18228 30242 -18172
rect 30298 -18228 30540 -18172
rect 30000 -18460 30540 -18228
rect 37460 -11772 38000 -11540
rect 37460 -11828 37708 -11772
rect 37764 -11828 38000 -11772
rect 37460 -12092 38000 -11828
rect 37460 -12148 37708 -12092
rect 37764 -12148 38000 -12092
rect 37460 -12412 38000 -12148
rect 37460 -12468 37708 -12412
rect 37764 -12468 38000 -12412
rect 37460 -12732 38000 -12468
rect 37460 -12788 37708 -12732
rect 37764 -12788 38000 -12732
rect 37460 -13052 38000 -12788
rect 37460 -13108 37708 -13052
rect 37764 -13108 38000 -13052
rect 37460 -13372 38000 -13108
rect 37460 -13428 37708 -13372
rect 37764 -13428 38000 -13372
rect 37460 -13692 38000 -13428
rect 37460 -13748 37708 -13692
rect 37764 -13748 38000 -13692
rect 37460 -14012 38000 -13748
rect 37460 -14068 37708 -14012
rect 37764 -14068 38000 -14012
rect 37460 -14332 38000 -14068
rect 37460 -14388 37708 -14332
rect 37764 -14388 38000 -14332
rect 37460 -14652 38000 -14388
rect 37460 -14708 37708 -14652
rect 37764 -14708 38000 -14652
rect 37460 -14972 38000 -14708
rect 37460 -15028 37708 -14972
rect 37764 -15028 38000 -14972
rect 37460 -15292 38000 -15028
rect 37460 -15348 37708 -15292
rect 37764 -15348 38000 -15292
rect 37460 -15612 38000 -15348
rect 37460 -15668 37708 -15612
rect 37764 -15668 38000 -15612
rect 37460 -15932 38000 -15668
rect 37460 -15988 37708 -15932
rect 37764 -15988 38000 -15932
rect 37460 -16252 38000 -15988
rect 37460 -16308 37708 -16252
rect 37764 -16308 38000 -16252
rect 37460 -16572 38000 -16308
rect 37460 -16628 37708 -16572
rect 37764 -16628 38000 -16572
rect 37460 -16892 38000 -16628
rect 37460 -16948 37708 -16892
rect 37764 -16948 38000 -16892
rect 37460 -17212 38000 -16948
rect 37460 -17268 37708 -17212
rect 37764 -17268 38000 -17212
rect 37460 -17532 38000 -17268
rect 37460 -17588 37708 -17532
rect 37764 -17588 38000 -17532
rect 37460 -17852 38000 -17588
rect 37460 -17908 37708 -17852
rect 37764 -17908 38000 -17852
rect 37460 -18172 38000 -17908
rect 37460 -18228 37708 -18172
rect 37764 -18228 38000 -18172
rect 37460 -18460 38000 -18228
rect 30000 -18492 38000 -18460
rect 30000 -18548 30242 -18492
rect 30298 -18548 37708 -18492
rect 37764 -18548 38000 -18492
rect 30000 -18702 38000 -18548
rect 30000 -18758 30612 -18702
rect 30668 -18758 30932 -18702
rect 30988 -18758 31252 -18702
rect 31308 -18758 31572 -18702
rect 31628 -18758 31892 -18702
rect 31948 -18758 32212 -18702
rect 32268 -18758 32532 -18702
rect 32588 -18758 32852 -18702
rect 32908 -18758 33172 -18702
rect 33228 -18758 33492 -18702
rect 33548 -18758 33812 -18702
rect 33868 -18758 34132 -18702
rect 34188 -18758 34452 -18702
rect 34508 -18758 34772 -18702
rect 34828 -18758 35092 -18702
rect 35148 -18758 35412 -18702
rect 35468 -18758 35732 -18702
rect 35788 -18758 36052 -18702
rect 36108 -18758 36372 -18702
rect 36428 -18758 36692 -18702
rect 36748 -18758 37012 -18702
rect 37068 -18758 37332 -18702
rect 37388 -18758 38000 -18702
rect 30000 -19000 38000 -18758
rect 42000 -11246 50000 -11000
rect 42000 -11302 42612 -11246
rect 42668 -11302 42932 -11246
rect 42988 -11302 43252 -11246
rect 43308 -11302 43572 -11246
rect 43628 -11302 43892 -11246
rect 43948 -11302 44212 -11246
rect 44268 -11302 44532 -11246
rect 44588 -11302 44852 -11246
rect 44908 -11302 45172 -11246
rect 45228 -11302 45492 -11246
rect 45548 -11302 45812 -11246
rect 45868 -11302 46132 -11246
rect 46188 -11302 46452 -11246
rect 46508 -11302 46772 -11246
rect 46828 -11302 47092 -11246
rect 47148 -11302 47412 -11246
rect 47468 -11302 47732 -11246
rect 47788 -11302 48052 -11246
rect 48108 -11302 48372 -11246
rect 48428 -11302 48692 -11246
rect 48748 -11302 49012 -11246
rect 49068 -11302 49332 -11246
rect 49388 -11302 50000 -11246
rect 42000 -11452 50000 -11302
rect 42000 -11508 42242 -11452
rect 42298 -11508 49708 -11452
rect 49764 -11508 50000 -11452
rect 42000 -11540 50000 -11508
rect 42000 -11772 42540 -11540
rect 42000 -11828 42242 -11772
rect 42298 -11828 42540 -11772
rect 42000 -12092 42540 -11828
rect 42000 -12148 42242 -12092
rect 42298 -12148 42540 -12092
rect 42000 -12412 42540 -12148
rect 42000 -12468 42242 -12412
rect 42298 -12468 42540 -12412
rect 42000 -12732 42540 -12468
rect 42000 -12788 42242 -12732
rect 42298 -12788 42540 -12732
rect 42000 -13052 42540 -12788
rect 42000 -13108 42242 -13052
rect 42298 -13108 42540 -13052
rect 42000 -13372 42540 -13108
rect 42000 -13428 42242 -13372
rect 42298 -13428 42540 -13372
rect 42000 -13692 42540 -13428
rect 42000 -13748 42242 -13692
rect 42298 -13748 42540 -13692
rect 42000 -14012 42540 -13748
rect 42000 -14068 42242 -14012
rect 42298 -14068 42540 -14012
rect 42000 -14332 42540 -14068
rect 42000 -14388 42242 -14332
rect 42298 -14388 42540 -14332
rect 42000 -14652 42540 -14388
rect 42000 -14708 42242 -14652
rect 42298 -14708 42540 -14652
rect 42000 -14972 42540 -14708
rect 42000 -15028 42242 -14972
rect 42298 -15028 42540 -14972
rect 42000 -15292 42540 -15028
rect 42000 -15348 42242 -15292
rect 42298 -15348 42540 -15292
rect 42000 -15612 42540 -15348
rect 42000 -15668 42242 -15612
rect 42298 -15668 42540 -15612
rect 42000 -15932 42540 -15668
rect 42000 -15988 42242 -15932
rect 42298 -15988 42540 -15932
rect 42000 -16252 42540 -15988
rect 42000 -16308 42242 -16252
rect 42298 -16308 42540 -16252
rect 42000 -16572 42540 -16308
rect 42000 -16628 42242 -16572
rect 42298 -16628 42540 -16572
rect 42000 -16892 42540 -16628
rect 42000 -16948 42242 -16892
rect 42298 -16948 42540 -16892
rect 42000 -17212 42540 -16948
rect 42000 -17268 42242 -17212
rect 42298 -17268 42540 -17212
rect 42000 -17532 42540 -17268
rect 42000 -17588 42242 -17532
rect 42298 -17588 42540 -17532
rect 42000 -17852 42540 -17588
rect 42000 -17908 42242 -17852
rect 42298 -17908 42540 -17852
rect 42000 -18172 42540 -17908
rect 42000 -18228 42242 -18172
rect 42298 -18228 42540 -18172
rect 42000 -18460 42540 -18228
rect 49460 -11772 50000 -11540
rect 49460 -11828 49708 -11772
rect 49764 -11828 50000 -11772
rect 49460 -12092 50000 -11828
rect 49460 -12148 49708 -12092
rect 49764 -12148 50000 -12092
rect 49460 -12412 50000 -12148
rect 49460 -12468 49708 -12412
rect 49764 -12468 50000 -12412
rect 49460 -12732 50000 -12468
rect 49460 -12788 49708 -12732
rect 49764 -12788 50000 -12732
rect 49460 -13052 50000 -12788
rect 49460 -13108 49708 -13052
rect 49764 -13108 50000 -13052
rect 49460 -13372 50000 -13108
rect 49460 -13428 49708 -13372
rect 49764 -13428 50000 -13372
rect 49460 -13692 50000 -13428
rect 49460 -13748 49708 -13692
rect 49764 -13748 50000 -13692
rect 49460 -14012 50000 -13748
rect 49460 -14068 49708 -14012
rect 49764 -14068 50000 -14012
rect 49460 -14332 50000 -14068
rect 49460 -14388 49708 -14332
rect 49764 -14388 50000 -14332
rect 49460 -14652 50000 -14388
rect 49460 -14708 49708 -14652
rect 49764 -14708 50000 -14652
rect 49460 -14972 50000 -14708
rect 49460 -15028 49708 -14972
rect 49764 -15028 50000 -14972
rect 49460 -15292 50000 -15028
rect 49460 -15348 49708 -15292
rect 49764 -15348 50000 -15292
rect 49460 -15612 50000 -15348
rect 49460 -15668 49708 -15612
rect 49764 -15668 50000 -15612
rect 49460 -15932 50000 -15668
rect 49460 -15988 49708 -15932
rect 49764 -15988 50000 -15932
rect 49460 -16252 50000 -15988
rect 49460 -16308 49708 -16252
rect 49764 -16308 50000 -16252
rect 49460 -16572 50000 -16308
rect 49460 -16628 49708 -16572
rect 49764 -16628 50000 -16572
rect 49460 -16892 50000 -16628
rect 49460 -16948 49708 -16892
rect 49764 -16948 50000 -16892
rect 49460 -17212 50000 -16948
rect 49460 -17268 49708 -17212
rect 49764 -17268 50000 -17212
rect 49460 -17532 50000 -17268
rect 49460 -17588 49708 -17532
rect 49764 -17588 50000 -17532
rect 49460 -17852 50000 -17588
rect 49460 -17908 49708 -17852
rect 49764 -17908 50000 -17852
rect 49460 -18172 50000 -17908
rect 49460 -18228 49708 -18172
rect 49764 -18228 50000 -18172
rect 49460 -18460 50000 -18228
rect 42000 -18492 50000 -18460
rect 42000 -18548 42242 -18492
rect 42298 -18548 49708 -18492
rect 49764 -18548 50000 -18492
rect 42000 -18702 50000 -18548
rect 42000 -18758 42612 -18702
rect 42668 -18758 42932 -18702
rect 42988 -18758 43252 -18702
rect 43308 -18758 43572 -18702
rect 43628 -18758 43892 -18702
rect 43948 -18758 44212 -18702
rect 44268 -18758 44532 -18702
rect 44588 -18758 44852 -18702
rect 44908 -18758 45172 -18702
rect 45228 -18758 45492 -18702
rect 45548 -18758 45812 -18702
rect 45868 -18758 46132 -18702
rect 46188 -18758 46452 -18702
rect 46508 -18758 46772 -18702
rect 46828 -18758 47092 -18702
rect 47148 -18758 47412 -18702
rect 47468 -18758 47732 -18702
rect 47788 -18758 48052 -18702
rect 48108 -18758 48372 -18702
rect 48428 -18758 48692 -18702
rect 48748 -18758 49012 -18702
rect 49068 -18758 49332 -18702
rect 49388 -18758 50000 -18702
rect 42000 -19000 50000 -18758
rect 6000 -23246 14000 -23000
rect 6000 -23302 6612 -23246
rect 6668 -23302 6932 -23246
rect 6988 -23302 7252 -23246
rect 7308 -23302 7572 -23246
rect 7628 -23302 7892 -23246
rect 7948 -23302 8212 -23246
rect 8268 -23302 8532 -23246
rect 8588 -23302 8852 -23246
rect 8908 -23302 9172 -23246
rect 9228 -23302 9492 -23246
rect 9548 -23302 9812 -23246
rect 9868 -23302 10132 -23246
rect 10188 -23302 10452 -23246
rect 10508 -23302 10772 -23246
rect 10828 -23302 11092 -23246
rect 11148 -23302 11412 -23246
rect 11468 -23302 11732 -23246
rect 11788 -23302 12052 -23246
rect 12108 -23302 12372 -23246
rect 12428 -23302 12692 -23246
rect 12748 -23302 13012 -23246
rect 13068 -23302 13332 -23246
rect 13388 -23302 14000 -23246
rect 6000 -23452 14000 -23302
rect 6000 -23508 6242 -23452
rect 6298 -23508 13708 -23452
rect 13764 -23508 14000 -23452
rect 6000 -23540 14000 -23508
rect 6000 -23772 6540 -23540
rect 6000 -23828 6242 -23772
rect 6298 -23828 6540 -23772
rect 6000 -24092 6540 -23828
rect 6000 -24148 6242 -24092
rect 6298 -24148 6540 -24092
rect 6000 -24412 6540 -24148
rect 6000 -24468 6242 -24412
rect 6298 -24468 6540 -24412
rect 6000 -24732 6540 -24468
rect 6000 -24788 6242 -24732
rect 6298 -24788 6540 -24732
rect 6000 -25052 6540 -24788
rect 6000 -25108 6242 -25052
rect 6298 -25108 6540 -25052
rect 6000 -25372 6540 -25108
rect 6000 -25428 6242 -25372
rect 6298 -25428 6540 -25372
rect 6000 -25692 6540 -25428
rect 6000 -25748 6242 -25692
rect 6298 -25748 6540 -25692
rect 6000 -26012 6540 -25748
rect 6000 -26068 6242 -26012
rect 6298 -26068 6540 -26012
rect 6000 -26332 6540 -26068
rect 6000 -26388 6242 -26332
rect 6298 -26388 6540 -26332
rect 6000 -26652 6540 -26388
rect 6000 -26708 6242 -26652
rect 6298 -26708 6540 -26652
rect 6000 -26972 6540 -26708
rect 6000 -27028 6242 -26972
rect 6298 -27028 6540 -26972
rect 6000 -27292 6540 -27028
rect 6000 -27348 6242 -27292
rect 6298 -27348 6540 -27292
rect 6000 -27612 6540 -27348
rect 6000 -27668 6242 -27612
rect 6298 -27668 6540 -27612
rect 6000 -27932 6540 -27668
rect 6000 -27988 6242 -27932
rect 6298 -27988 6540 -27932
rect 6000 -28252 6540 -27988
rect 6000 -28308 6242 -28252
rect 6298 -28308 6540 -28252
rect 6000 -28572 6540 -28308
rect 6000 -28628 6242 -28572
rect 6298 -28628 6540 -28572
rect 6000 -28892 6540 -28628
rect 6000 -28948 6242 -28892
rect 6298 -28948 6540 -28892
rect 6000 -29212 6540 -28948
rect 6000 -29268 6242 -29212
rect 6298 -29268 6540 -29212
rect 6000 -29532 6540 -29268
rect 6000 -29588 6242 -29532
rect 6298 -29588 6540 -29532
rect 6000 -29852 6540 -29588
rect 6000 -29908 6242 -29852
rect 6298 -29908 6540 -29852
rect 6000 -30172 6540 -29908
rect 6000 -30228 6242 -30172
rect 6298 -30228 6540 -30172
rect 6000 -30460 6540 -30228
rect 13460 -23772 14000 -23540
rect 13460 -23828 13708 -23772
rect 13764 -23828 14000 -23772
rect 13460 -24092 14000 -23828
rect 13460 -24148 13708 -24092
rect 13764 -24148 14000 -24092
rect 13460 -24412 14000 -24148
rect 13460 -24468 13708 -24412
rect 13764 -24468 14000 -24412
rect 13460 -24732 14000 -24468
rect 13460 -24788 13708 -24732
rect 13764 -24788 14000 -24732
rect 13460 -25052 14000 -24788
rect 13460 -25108 13708 -25052
rect 13764 -25108 14000 -25052
rect 13460 -25372 14000 -25108
rect 13460 -25428 13708 -25372
rect 13764 -25428 14000 -25372
rect 13460 -25692 14000 -25428
rect 13460 -25748 13708 -25692
rect 13764 -25748 14000 -25692
rect 13460 -26012 14000 -25748
rect 13460 -26068 13708 -26012
rect 13764 -26068 14000 -26012
rect 13460 -26332 14000 -26068
rect 13460 -26388 13708 -26332
rect 13764 -26388 14000 -26332
rect 13460 -26652 14000 -26388
rect 13460 -26708 13708 -26652
rect 13764 -26708 14000 -26652
rect 13460 -26972 14000 -26708
rect 13460 -27028 13708 -26972
rect 13764 -27028 14000 -26972
rect 13460 -27292 14000 -27028
rect 13460 -27348 13708 -27292
rect 13764 -27348 14000 -27292
rect 13460 -27612 14000 -27348
rect 13460 -27668 13708 -27612
rect 13764 -27668 14000 -27612
rect 13460 -27932 14000 -27668
rect 13460 -27988 13708 -27932
rect 13764 -27988 14000 -27932
rect 13460 -28252 14000 -27988
rect 13460 -28308 13708 -28252
rect 13764 -28308 14000 -28252
rect 13460 -28572 14000 -28308
rect 13460 -28628 13708 -28572
rect 13764 -28628 14000 -28572
rect 13460 -28892 14000 -28628
rect 13460 -28948 13708 -28892
rect 13764 -28948 14000 -28892
rect 13460 -29212 14000 -28948
rect 13460 -29268 13708 -29212
rect 13764 -29268 14000 -29212
rect 13460 -29532 14000 -29268
rect 13460 -29588 13708 -29532
rect 13764 -29588 14000 -29532
rect 13460 -29852 14000 -29588
rect 13460 -29908 13708 -29852
rect 13764 -29908 14000 -29852
rect 13460 -30172 14000 -29908
rect 13460 -30228 13708 -30172
rect 13764 -30228 14000 -30172
rect 13460 -30460 14000 -30228
rect 6000 -30492 14000 -30460
rect 6000 -30548 6242 -30492
rect 6298 -30548 13708 -30492
rect 13764 -30548 14000 -30492
rect 6000 -30702 14000 -30548
rect 6000 -30758 6612 -30702
rect 6668 -30758 6932 -30702
rect 6988 -30758 7252 -30702
rect 7308 -30758 7572 -30702
rect 7628 -30758 7892 -30702
rect 7948 -30758 8212 -30702
rect 8268 -30758 8532 -30702
rect 8588 -30758 8852 -30702
rect 8908 -30758 9172 -30702
rect 9228 -30758 9492 -30702
rect 9548 -30758 9812 -30702
rect 9868 -30758 10132 -30702
rect 10188 -30758 10452 -30702
rect 10508 -30758 10772 -30702
rect 10828 -30758 11092 -30702
rect 11148 -30758 11412 -30702
rect 11468 -30758 11732 -30702
rect 11788 -30758 12052 -30702
rect 12108 -30758 12372 -30702
rect 12428 -30758 12692 -30702
rect 12748 -30758 13012 -30702
rect 13068 -30758 13332 -30702
rect 13388 -30758 14000 -30702
rect 6000 -31000 14000 -30758
rect 18000 -23246 26000 -23000
rect 18000 -23302 18612 -23246
rect 18668 -23302 18932 -23246
rect 18988 -23302 19252 -23246
rect 19308 -23302 19572 -23246
rect 19628 -23302 19892 -23246
rect 19948 -23302 20212 -23246
rect 20268 -23302 20532 -23246
rect 20588 -23302 20852 -23246
rect 20908 -23302 21172 -23246
rect 21228 -23302 21492 -23246
rect 21548 -23302 21812 -23246
rect 21868 -23302 22132 -23246
rect 22188 -23302 22452 -23246
rect 22508 -23302 22772 -23246
rect 22828 -23302 23092 -23246
rect 23148 -23302 23412 -23246
rect 23468 -23302 23732 -23246
rect 23788 -23302 24052 -23246
rect 24108 -23302 24372 -23246
rect 24428 -23302 24692 -23246
rect 24748 -23302 25012 -23246
rect 25068 -23302 25332 -23246
rect 25388 -23302 26000 -23246
rect 18000 -23452 26000 -23302
rect 18000 -23508 18242 -23452
rect 18298 -23508 25708 -23452
rect 25764 -23508 26000 -23452
rect 18000 -23540 26000 -23508
rect 18000 -23772 18540 -23540
rect 18000 -23828 18242 -23772
rect 18298 -23828 18540 -23772
rect 18000 -24092 18540 -23828
rect 18000 -24148 18242 -24092
rect 18298 -24148 18540 -24092
rect 18000 -24412 18540 -24148
rect 18000 -24468 18242 -24412
rect 18298 -24468 18540 -24412
rect 18000 -24732 18540 -24468
rect 18000 -24788 18242 -24732
rect 18298 -24788 18540 -24732
rect 18000 -25052 18540 -24788
rect 18000 -25108 18242 -25052
rect 18298 -25108 18540 -25052
rect 18000 -25372 18540 -25108
rect 18000 -25428 18242 -25372
rect 18298 -25428 18540 -25372
rect 18000 -25692 18540 -25428
rect 18000 -25748 18242 -25692
rect 18298 -25748 18540 -25692
rect 18000 -26012 18540 -25748
rect 18000 -26068 18242 -26012
rect 18298 -26068 18540 -26012
rect 18000 -26332 18540 -26068
rect 18000 -26388 18242 -26332
rect 18298 -26388 18540 -26332
rect 18000 -26652 18540 -26388
rect 18000 -26708 18242 -26652
rect 18298 -26708 18540 -26652
rect 18000 -26972 18540 -26708
rect 18000 -27028 18242 -26972
rect 18298 -27028 18540 -26972
rect 18000 -27292 18540 -27028
rect 18000 -27348 18242 -27292
rect 18298 -27348 18540 -27292
rect 18000 -27612 18540 -27348
rect 18000 -27668 18242 -27612
rect 18298 -27668 18540 -27612
rect 18000 -27932 18540 -27668
rect 18000 -27988 18242 -27932
rect 18298 -27988 18540 -27932
rect 18000 -28252 18540 -27988
rect 18000 -28308 18242 -28252
rect 18298 -28308 18540 -28252
rect 18000 -28572 18540 -28308
rect 18000 -28628 18242 -28572
rect 18298 -28628 18540 -28572
rect 18000 -28892 18540 -28628
rect 18000 -28948 18242 -28892
rect 18298 -28948 18540 -28892
rect 18000 -29212 18540 -28948
rect 18000 -29268 18242 -29212
rect 18298 -29268 18540 -29212
rect 18000 -29532 18540 -29268
rect 18000 -29588 18242 -29532
rect 18298 -29588 18540 -29532
rect 18000 -29852 18540 -29588
rect 18000 -29908 18242 -29852
rect 18298 -29908 18540 -29852
rect 18000 -30172 18540 -29908
rect 18000 -30228 18242 -30172
rect 18298 -30228 18540 -30172
rect 18000 -30460 18540 -30228
rect 25460 -23772 26000 -23540
rect 25460 -23828 25708 -23772
rect 25764 -23828 26000 -23772
rect 25460 -24092 26000 -23828
rect 25460 -24148 25708 -24092
rect 25764 -24148 26000 -24092
rect 25460 -24412 26000 -24148
rect 25460 -24468 25708 -24412
rect 25764 -24468 26000 -24412
rect 25460 -24732 26000 -24468
rect 25460 -24788 25708 -24732
rect 25764 -24788 26000 -24732
rect 25460 -25052 26000 -24788
rect 25460 -25108 25708 -25052
rect 25764 -25108 26000 -25052
rect 25460 -25372 26000 -25108
rect 25460 -25428 25708 -25372
rect 25764 -25428 26000 -25372
rect 25460 -25692 26000 -25428
rect 25460 -25748 25708 -25692
rect 25764 -25748 26000 -25692
rect 25460 -26012 26000 -25748
rect 25460 -26068 25708 -26012
rect 25764 -26068 26000 -26012
rect 25460 -26332 26000 -26068
rect 25460 -26388 25708 -26332
rect 25764 -26388 26000 -26332
rect 25460 -26652 26000 -26388
rect 25460 -26708 25708 -26652
rect 25764 -26708 26000 -26652
rect 25460 -26972 26000 -26708
rect 25460 -27028 25708 -26972
rect 25764 -27028 26000 -26972
rect 25460 -27292 26000 -27028
rect 25460 -27348 25708 -27292
rect 25764 -27348 26000 -27292
rect 25460 -27612 26000 -27348
rect 25460 -27668 25708 -27612
rect 25764 -27668 26000 -27612
rect 25460 -27932 26000 -27668
rect 25460 -27988 25708 -27932
rect 25764 -27988 26000 -27932
rect 25460 -28252 26000 -27988
rect 25460 -28308 25708 -28252
rect 25764 -28308 26000 -28252
rect 25460 -28572 26000 -28308
rect 25460 -28628 25708 -28572
rect 25764 -28628 26000 -28572
rect 25460 -28892 26000 -28628
rect 25460 -28948 25708 -28892
rect 25764 -28948 26000 -28892
rect 25460 -29212 26000 -28948
rect 25460 -29268 25708 -29212
rect 25764 -29268 26000 -29212
rect 25460 -29532 26000 -29268
rect 25460 -29588 25708 -29532
rect 25764 -29588 26000 -29532
rect 25460 -29852 26000 -29588
rect 25460 -29908 25708 -29852
rect 25764 -29908 26000 -29852
rect 25460 -30172 26000 -29908
rect 25460 -30228 25708 -30172
rect 25764 -30228 26000 -30172
rect 25460 -30460 26000 -30228
rect 18000 -30492 26000 -30460
rect 18000 -30548 18242 -30492
rect 18298 -30548 25708 -30492
rect 25764 -30548 26000 -30492
rect 18000 -30702 26000 -30548
rect 18000 -30758 18612 -30702
rect 18668 -30758 18932 -30702
rect 18988 -30758 19252 -30702
rect 19308 -30758 19572 -30702
rect 19628 -30758 19892 -30702
rect 19948 -30758 20212 -30702
rect 20268 -30758 20532 -30702
rect 20588 -30758 20852 -30702
rect 20908 -30758 21172 -30702
rect 21228 -30758 21492 -30702
rect 21548 -30758 21812 -30702
rect 21868 -30758 22132 -30702
rect 22188 -30758 22452 -30702
rect 22508 -30758 22772 -30702
rect 22828 -30758 23092 -30702
rect 23148 -30758 23412 -30702
rect 23468 -30758 23732 -30702
rect 23788 -30758 24052 -30702
rect 24108 -30758 24372 -30702
rect 24428 -30758 24692 -30702
rect 24748 -30758 25012 -30702
rect 25068 -30758 25332 -30702
rect 25388 -30758 26000 -30702
rect 18000 -31000 26000 -30758
rect 30000 -23246 38000 -23000
rect 30000 -23302 30612 -23246
rect 30668 -23302 30932 -23246
rect 30988 -23302 31252 -23246
rect 31308 -23302 31572 -23246
rect 31628 -23302 31892 -23246
rect 31948 -23302 32212 -23246
rect 32268 -23302 32532 -23246
rect 32588 -23302 32852 -23246
rect 32908 -23302 33172 -23246
rect 33228 -23302 33492 -23246
rect 33548 -23302 33812 -23246
rect 33868 -23302 34132 -23246
rect 34188 -23302 34452 -23246
rect 34508 -23302 34772 -23246
rect 34828 -23302 35092 -23246
rect 35148 -23302 35412 -23246
rect 35468 -23302 35732 -23246
rect 35788 -23302 36052 -23246
rect 36108 -23302 36372 -23246
rect 36428 -23302 36692 -23246
rect 36748 -23302 37012 -23246
rect 37068 -23302 37332 -23246
rect 37388 -23302 38000 -23246
rect 30000 -23452 38000 -23302
rect 30000 -23508 30242 -23452
rect 30298 -23508 37708 -23452
rect 37764 -23508 38000 -23452
rect 30000 -23540 38000 -23508
rect 30000 -23772 30540 -23540
rect 30000 -23828 30242 -23772
rect 30298 -23828 30540 -23772
rect 30000 -24092 30540 -23828
rect 30000 -24148 30242 -24092
rect 30298 -24148 30540 -24092
rect 30000 -24412 30540 -24148
rect 30000 -24468 30242 -24412
rect 30298 -24468 30540 -24412
rect 30000 -24732 30540 -24468
rect 30000 -24788 30242 -24732
rect 30298 -24788 30540 -24732
rect 30000 -25052 30540 -24788
rect 30000 -25108 30242 -25052
rect 30298 -25108 30540 -25052
rect 30000 -25372 30540 -25108
rect 30000 -25428 30242 -25372
rect 30298 -25428 30540 -25372
rect 30000 -25692 30540 -25428
rect 30000 -25748 30242 -25692
rect 30298 -25748 30540 -25692
rect 30000 -26012 30540 -25748
rect 30000 -26068 30242 -26012
rect 30298 -26068 30540 -26012
rect 30000 -26332 30540 -26068
rect 30000 -26388 30242 -26332
rect 30298 -26388 30540 -26332
rect 30000 -26652 30540 -26388
rect 30000 -26708 30242 -26652
rect 30298 -26708 30540 -26652
rect 30000 -26972 30540 -26708
rect 30000 -27028 30242 -26972
rect 30298 -27028 30540 -26972
rect 30000 -27292 30540 -27028
rect 30000 -27348 30242 -27292
rect 30298 -27348 30540 -27292
rect 30000 -27612 30540 -27348
rect 30000 -27668 30242 -27612
rect 30298 -27668 30540 -27612
rect 30000 -27932 30540 -27668
rect 30000 -27988 30242 -27932
rect 30298 -27988 30540 -27932
rect 30000 -28252 30540 -27988
rect 30000 -28308 30242 -28252
rect 30298 -28308 30540 -28252
rect 30000 -28572 30540 -28308
rect 30000 -28628 30242 -28572
rect 30298 -28628 30540 -28572
rect 30000 -28892 30540 -28628
rect 30000 -28948 30242 -28892
rect 30298 -28948 30540 -28892
rect 30000 -29212 30540 -28948
rect 30000 -29268 30242 -29212
rect 30298 -29268 30540 -29212
rect 30000 -29532 30540 -29268
rect 30000 -29588 30242 -29532
rect 30298 -29588 30540 -29532
rect 30000 -29852 30540 -29588
rect 30000 -29908 30242 -29852
rect 30298 -29908 30540 -29852
rect 30000 -30172 30540 -29908
rect 30000 -30228 30242 -30172
rect 30298 -30228 30540 -30172
rect 30000 -30460 30540 -30228
rect 37460 -23772 38000 -23540
rect 37460 -23828 37708 -23772
rect 37764 -23828 38000 -23772
rect 37460 -24092 38000 -23828
rect 37460 -24148 37708 -24092
rect 37764 -24148 38000 -24092
rect 37460 -24412 38000 -24148
rect 37460 -24468 37708 -24412
rect 37764 -24468 38000 -24412
rect 37460 -24732 38000 -24468
rect 37460 -24788 37708 -24732
rect 37764 -24788 38000 -24732
rect 37460 -25052 38000 -24788
rect 37460 -25108 37708 -25052
rect 37764 -25108 38000 -25052
rect 37460 -25372 38000 -25108
rect 37460 -25428 37708 -25372
rect 37764 -25428 38000 -25372
rect 37460 -25692 38000 -25428
rect 37460 -25748 37708 -25692
rect 37764 -25748 38000 -25692
rect 37460 -26012 38000 -25748
rect 37460 -26068 37708 -26012
rect 37764 -26068 38000 -26012
rect 37460 -26332 38000 -26068
rect 37460 -26388 37708 -26332
rect 37764 -26388 38000 -26332
rect 37460 -26652 38000 -26388
rect 37460 -26708 37708 -26652
rect 37764 -26708 38000 -26652
rect 37460 -26972 38000 -26708
rect 37460 -27028 37708 -26972
rect 37764 -27028 38000 -26972
rect 37460 -27292 38000 -27028
rect 37460 -27348 37708 -27292
rect 37764 -27348 38000 -27292
rect 37460 -27612 38000 -27348
rect 37460 -27668 37708 -27612
rect 37764 -27668 38000 -27612
rect 37460 -27932 38000 -27668
rect 37460 -27988 37708 -27932
rect 37764 -27988 38000 -27932
rect 37460 -28252 38000 -27988
rect 37460 -28308 37708 -28252
rect 37764 -28308 38000 -28252
rect 37460 -28572 38000 -28308
rect 37460 -28628 37708 -28572
rect 37764 -28628 38000 -28572
rect 37460 -28892 38000 -28628
rect 37460 -28948 37708 -28892
rect 37764 -28948 38000 -28892
rect 37460 -29212 38000 -28948
rect 37460 -29268 37708 -29212
rect 37764 -29268 38000 -29212
rect 37460 -29532 38000 -29268
rect 37460 -29588 37708 -29532
rect 37764 -29588 38000 -29532
rect 37460 -29852 38000 -29588
rect 37460 -29908 37708 -29852
rect 37764 -29908 38000 -29852
rect 37460 -30172 38000 -29908
rect 37460 -30228 37708 -30172
rect 37764 -30228 38000 -30172
rect 37460 -30460 38000 -30228
rect 30000 -30492 38000 -30460
rect 30000 -30548 30242 -30492
rect 30298 -30548 37708 -30492
rect 37764 -30548 38000 -30492
rect 30000 -30702 38000 -30548
rect 30000 -30758 30612 -30702
rect 30668 -30758 30932 -30702
rect 30988 -30758 31252 -30702
rect 31308 -30758 31572 -30702
rect 31628 -30758 31892 -30702
rect 31948 -30758 32212 -30702
rect 32268 -30758 32532 -30702
rect 32588 -30758 32852 -30702
rect 32908 -30758 33172 -30702
rect 33228 -30758 33492 -30702
rect 33548 -30758 33812 -30702
rect 33868 -30758 34132 -30702
rect 34188 -30758 34452 -30702
rect 34508 -30758 34772 -30702
rect 34828 -30758 35092 -30702
rect 35148 -30758 35412 -30702
rect 35468 -30758 35732 -30702
rect 35788 -30758 36052 -30702
rect 36108 -30758 36372 -30702
rect 36428 -30758 36692 -30702
rect 36748 -30758 37012 -30702
rect 37068 -30758 37332 -30702
rect 37388 -30758 38000 -30702
rect 30000 -31000 38000 -30758
rect 42000 -23246 50000 -23000
rect 42000 -23302 42612 -23246
rect 42668 -23302 42932 -23246
rect 42988 -23302 43252 -23246
rect 43308 -23302 43572 -23246
rect 43628 -23302 43892 -23246
rect 43948 -23302 44212 -23246
rect 44268 -23302 44532 -23246
rect 44588 -23302 44852 -23246
rect 44908 -23302 45172 -23246
rect 45228 -23302 45492 -23246
rect 45548 -23302 45812 -23246
rect 45868 -23302 46132 -23246
rect 46188 -23302 46452 -23246
rect 46508 -23302 46772 -23246
rect 46828 -23302 47092 -23246
rect 47148 -23302 47412 -23246
rect 47468 -23302 47732 -23246
rect 47788 -23302 48052 -23246
rect 48108 -23302 48372 -23246
rect 48428 -23302 48692 -23246
rect 48748 -23302 49012 -23246
rect 49068 -23302 49332 -23246
rect 49388 -23302 50000 -23246
rect 42000 -23452 50000 -23302
rect 42000 -23508 42242 -23452
rect 42298 -23508 49708 -23452
rect 49764 -23508 50000 -23452
rect 42000 -23540 50000 -23508
rect 42000 -23772 42540 -23540
rect 42000 -23828 42242 -23772
rect 42298 -23828 42540 -23772
rect 42000 -24092 42540 -23828
rect 42000 -24148 42242 -24092
rect 42298 -24148 42540 -24092
rect 42000 -24412 42540 -24148
rect 42000 -24468 42242 -24412
rect 42298 -24468 42540 -24412
rect 42000 -24732 42540 -24468
rect 42000 -24788 42242 -24732
rect 42298 -24788 42540 -24732
rect 42000 -25052 42540 -24788
rect 42000 -25108 42242 -25052
rect 42298 -25108 42540 -25052
rect 42000 -25372 42540 -25108
rect 42000 -25428 42242 -25372
rect 42298 -25428 42540 -25372
rect 42000 -25692 42540 -25428
rect 42000 -25748 42242 -25692
rect 42298 -25748 42540 -25692
rect 42000 -26012 42540 -25748
rect 42000 -26068 42242 -26012
rect 42298 -26068 42540 -26012
rect 42000 -26332 42540 -26068
rect 42000 -26388 42242 -26332
rect 42298 -26388 42540 -26332
rect 42000 -26652 42540 -26388
rect 42000 -26708 42242 -26652
rect 42298 -26708 42540 -26652
rect 42000 -26972 42540 -26708
rect 42000 -27028 42242 -26972
rect 42298 -27028 42540 -26972
rect 42000 -27292 42540 -27028
rect 42000 -27348 42242 -27292
rect 42298 -27348 42540 -27292
rect 42000 -27612 42540 -27348
rect 42000 -27668 42242 -27612
rect 42298 -27668 42540 -27612
rect 42000 -27932 42540 -27668
rect 42000 -27988 42242 -27932
rect 42298 -27988 42540 -27932
rect 42000 -28252 42540 -27988
rect 42000 -28308 42242 -28252
rect 42298 -28308 42540 -28252
rect 42000 -28572 42540 -28308
rect 42000 -28628 42242 -28572
rect 42298 -28628 42540 -28572
rect 42000 -28892 42540 -28628
rect 42000 -28948 42242 -28892
rect 42298 -28948 42540 -28892
rect 42000 -29212 42540 -28948
rect 42000 -29268 42242 -29212
rect 42298 -29268 42540 -29212
rect 42000 -29532 42540 -29268
rect 42000 -29588 42242 -29532
rect 42298 -29588 42540 -29532
rect 42000 -29852 42540 -29588
rect 42000 -29908 42242 -29852
rect 42298 -29908 42540 -29852
rect 42000 -30172 42540 -29908
rect 42000 -30228 42242 -30172
rect 42298 -30228 42540 -30172
rect 42000 -30460 42540 -30228
rect 49460 -23772 50000 -23540
rect 49460 -23828 49708 -23772
rect 49764 -23828 50000 -23772
rect 49460 -24092 50000 -23828
rect 49460 -24148 49708 -24092
rect 49764 -24148 50000 -24092
rect 49460 -24412 50000 -24148
rect 49460 -24468 49708 -24412
rect 49764 -24468 50000 -24412
rect 49460 -24732 50000 -24468
rect 49460 -24788 49708 -24732
rect 49764 -24788 50000 -24732
rect 49460 -25052 50000 -24788
rect 49460 -25108 49708 -25052
rect 49764 -25108 50000 -25052
rect 49460 -25372 50000 -25108
rect 49460 -25428 49708 -25372
rect 49764 -25428 50000 -25372
rect 49460 -25692 50000 -25428
rect 49460 -25748 49708 -25692
rect 49764 -25748 50000 -25692
rect 49460 -26012 50000 -25748
rect 49460 -26068 49708 -26012
rect 49764 -26068 50000 -26012
rect 49460 -26332 50000 -26068
rect 49460 -26388 49708 -26332
rect 49764 -26388 50000 -26332
rect 49460 -26652 50000 -26388
rect 49460 -26708 49708 -26652
rect 49764 -26708 50000 -26652
rect 49460 -26972 50000 -26708
rect 49460 -27028 49708 -26972
rect 49764 -27028 50000 -26972
rect 49460 -27292 50000 -27028
rect 49460 -27348 49708 -27292
rect 49764 -27348 50000 -27292
rect 49460 -27612 50000 -27348
rect 49460 -27668 49708 -27612
rect 49764 -27668 50000 -27612
rect 49460 -27932 50000 -27668
rect 49460 -27988 49708 -27932
rect 49764 -27988 50000 -27932
rect 49460 -28252 50000 -27988
rect 49460 -28308 49708 -28252
rect 49764 -28308 50000 -28252
rect 49460 -28572 50000 -28308
rect 49460 -28628 49708 -28572
rect 49764 -28628 50000 -28572
rect 49460 -28892 50000 -28628
rect 49460 -28948 49708 -28892
rect 49764 -28948 50000 -28892
rect 49460 -29212 50000 -28948
rect 49460 -29268 49708 -29212
rect 49764 -29268 50000 -29212
rect 49460 -29532 50000 -29268
rect 49460 -29588 49708 -29532
rect 49764 -29588 50000 -29532
rect 49460 -29852 50000 -29588
rect 49460 -29908 49708 -29852
rect 49764 -29908 50000 -29852
rect 49460 -30172 50000 -29908
rect 49460 -30228 49708 -30172
rect 49764 -30228 50000 -30172
rect 49460 -30460 50000 -30228
rect 42000 -30492 50000 -30460
rect 42000 -30548 42242 -30492
rect 42298 -30548 49708 -30492
rect 49764 -30548 50000 -30492
rect 42000 -30702 50000 -30548
rect 42000 -30758 42612 -30702
rect 42668 -30758 42932 -30702
rect 42988 -30758 43252 -30702
rect 43308 -30758 43572 -30702
rect 43628 -30758 43892 -30702
rect 43948 -30758 44212 -30702
rect 44268 -30758 44532 -30702
rect 44588 -30758 44852 -30702
rect 44908 -30758 45172 -30702
rect 45228 -30758 45492 -30702
rect 45548 -30758 45812 -30702
rect 45868 -30758 46132 -30702
rect 46188 -30758 46452 -30702
rect 46508 -30758 46772 -30702
rect 46828 -30758 47092 -30702
rect 47148 -30758 47412 -30702
rect 47468 -30758 47732 -30702
rect 47788 -30758 48052 -30702
rect 48108 -30758 48372 -30702
rect 48428 -30758 48692 -30702
rect 48748 -30758 49012 -30702
rect 49068 -30758 49332 -30702
rect 49388 -30758 50000 -30702
rect 42000 -31000 50000 -30758
<< via2 >>
rect 18300 -3000 21500 -2500
rect 18203 -5742 18259 -5740
rect 18203 -5794 18205 -5742
rect 18205 -5794 18257 -5742
rect 18257 -5794 18259 -5742
rect 18203 -5796 18259 -5794
rect 21882 -5650 21992 -5560
rect 19297 -6700 19363 -6650
rect 19297 -6706 19363 -6700
rect 19489 -6700 19555 -6650
rect 19489 -6706 19555 -6700
rect 19681 -6700 19747 -6650
rect 19681 -6706 19747 -6700
rect 19873 -6700 19939 -6650
rect 19873 -6706 19939 -6700
rect 20065 -6700 20131 -6650
rect 20065 -6706 20131 -6700
rect 20257 -6700 20323 -6650
rect 20257 -6706 20323 -6700
rect 20449 -6700 20515 -6650
rect 20449 -6706 20515 -6700
rect 20641 -6700 20707 -6650
rect 20641 -6706 20707 -6700
rect 18810 -7000 18970 -6940
rect 16920 -8485 17130 -8268
rect 16920 -8488 17130 -8485
rect 17400 -9360 17600 -8440
rect 21744 -5742 21800 -5740
rect 21744 -5794 21746 -5742
rect 21746 -5794 21798 -5742
rect 21798 -5794 21800 -5742
rect 21744 -5796 21800 -5794
rect 22472 -6660 22582 -6270
rect 22702 -6660 22812 -6270
rect 23270 -7540 23410 -7480
rect 23550 -7860 23690 -7800
rect 16400 -9580 16460 -9520
rect 16610 -9570 16670 -9510
rect 16470 -9720 16530 -9660
rect 17700 -10200 18900 -9600
rect 20900 -10200 22100 -9600
rect 17040 -10740 17120 -10620
rect 6612 -11248 6668 -11246
rect 6612 -11300 6614 -11248
rect 6614 -11300 6666 -11248
rect 6666 -11300 6668 -11248
rect 6612 -11302 6668 -11300
rect 6932 -11248 6988 -11246
rect 6932 -11300 6934 -11248
rect 6934 -11300 6986 -11248
rect 6986 -11300 6988 -11248
rect 6932 -11302 6988 -11300
rect 7252 -11248 7308 -11246
rect 7252 -11300 7254 -11248
rect 7254 -11300 7306 -11248
rect 7306 -11300 7308 -11248
rect 7252 -11302 7308 -11300
rect 7572 -11248 7628 -11246
rect 7572 -11300 7574 -11248
rect 7574 -11300 7626 -11248
rect 7626 -11300 7628 -11248
rect 7572 -11302 7628 -11300
rect 7892 -11248 7948 -11246
rect 7892 -11300 7894 -11248
rect 7894 -11300 7946 -11248
rect 7946 -11300 7948 -11248
rect 7892 -11302 7948 -11300
rect 8212 -11248 8268 -11246
rect 8212 -11300 8214 -11248
rect 8214 -11300 8266 -11248
rect 8266 -11300 8268 -11248
rect 8212 -11302 8268 -11300
rect 8532 -11248 8588 -11246
rect 8532 -11300 8534 -11248
rect 8534 -11300 8586 -11248
rect 8586 -11300 8588 -11248
rect 8532 -11302 8588 -11300
rect 8852 -11248 8908 -11246
rect 8852 -11300 8854 -11248
rect 8854 -11300 8906 -11248
rect 8906 -11300 8908 -11248
rect 8852 -11302 8908 -11300
rect 9172 -11248 9228 -11246
rect 9172 -11300 9174 -11248
rect 9174 -11300 9226 -11248
rect 9226 -11300 9228 -11248
rect 9172 -11302 9228 -11300
rect 9492 -11248 9548 -11246
rect 9492 -11300 9494 -11248
rect 9494 -11300 9546 -11248
rect 9546 -11300 9548 -11248
rect 9492 -11302 9548 -11300
rect 9812 -11248 9868 -11246
rect 9812 -11300 9814 -11248
rect 9814 -11300 9866 -11248
rect 9866 -11300 9868 -11248
rect 9812 -11302 9868 -11300
rect 10132 -11248 10188 -11246
rect 10132 -11300 10134 -11248
rect 10134 -11300 10186 -11248
rect 10186 -11300 10188 -11248
rect 10132 -11302 10188 -11300
rect 10452 -11248 10508 -11246
rect 10452 -11300 10454 -11248
rect 10454 -11300 10506 -11248
rect 10506 -11300 10508 -11248
rect 10452 -11302 10508 -11300
rect 10772 -11248 10828 -11246
rect 10772 -11300 10774 -11248
rect 10774 -11300 10826 -11248
rect 10826 -11300 10828 -11248
rect 10772 -11302 10828 -11300
rect 11092 -11248 11148 -11246
rect 11092 -11300 11094 -11248
rect 11094 -11300 11146 -11248
rect 11146 -11300 11148 -11248
rect 11092 -11302 11148 -11300
rect 11412 -11248 11468 -11246
rect 11412 -11300 11414 -11248
rect 11414 -11300 11466 -11248
rect 11466 -11300 11468 -11248
rect 11412 -11302 11468 -11300
rect 11732 -11248 11788 -11246
rect 11732 -11300 11734 -11248
rect 11734 -11300 11786 -11248
rect 11786 -11300 11788 -11248
rect 11732 -11302 11788 -11300
rect 12052 -11248 12108 -11246
rect 12052 -11300 12054 -11248
rect 12054 -11300 12106 -11248
rect 12106 -11300 12108 -11248
rect 12052 -11302 12108 -11300
rect 12372 -11248 12428 -11246
rect 12372 -11300 12374 -11248
rect 12374 -11300 12426 -11248
rect 12426 -11300 12428 -11248
rect 12372 -11302 12428 -11300
rect 12692 -11248 12748 -11246
rect 12692 -11300 12694 -11248
rect 12694 -11300 12746 -11248
rect 12746 -11300 12748 -11248
rect 12692 -11302 12748 -11300
rect 13012 -11248 13068 -11246
rect 13012 -11300 13014 -11248
rect 13014 -11300 13066 -11248
rect 13066 -11300 13068 -11248
rect 13012 -11302 13068 -11300
rect 13332 -11248 13388 -11246
rect 13332 -11300 13334 -11248
rect 13334 -11300 13386 -11248
rect 13386 -11300 13388 -11248
rect 13332 -11302 13388 -11300
rect 18612 -11248 18668 -11246
rect 18612 -11300 18614 -11248
rect 18614 -11300 18666 -11248
rect 18666 -11300 18668 -11248
rect 18612 -11302 18668 -11300
rect 18932 -11248 18988 -11246
rect 18932 -11300 18934 -11248
rect 18934 -11300 18986 -11248
rect 18986 -11300 18988 -11248
rect 18932 -11302 18988 -11300
rect 19252 -11248 19308 -11246
rect 19252 -11300 19254 -11248
rect 19254 -11300 19306 -11248
rect 19306 -11300 19308 -11248
rect 19252 -11302 19308 -11300
rect 19572 -11248 19628 -11246
rect 19572 -11300 19574 -11248
rect 19574 -11300 19626 -11248
rect 19626 -11300 19628 -11248
rect 19572 -11302 19628 -11300
rect 19892 -11248 19948 -11246
rect 19892 -11300 19894 -11248
rect 19894 -11300 19946 -11248
rect 19946 -11300 19948 -11248
rect 19892 -11302 19948 -11300
rect 20212 -11248 20268 -11246
rect 20212 -11300 20214 -11248
rect 20214 -11300 20266 -11248
rect 20266 -11300 20268 -11248
rect 20212 -11302 20268 -11300
rect 20532 -11248 20588 -11246
rect 20532 -11300 20534 -11248
rect 20534 -11300 20586 -11248
rect 20586 -11300 20588 -11248
rect 20532 -11302 20588 -11300
rect 20852 -11248 20908 -11246
rect 20852 -11300 20854 -11248
rect 20854 -11300 20906 -11248
rect 20906 -11300 20908 -11248
rect 20852 -11302 20908 -11300
rect 21172 -11248 21228 -11246
rect 21172 -11300 21174 -11248
rect 21174 -11300 21226 -11248
rect 21226 -11300 21228 -11248
rect 21172 -11302 21228 -11300
rect 21492 -11248 21548 -11246
rect 21492 -11300 21494 -11248
rect 21494 -11300 21546 -11248
rect 21546 -11300 21548 -11248
rect 21492 -11302 21548 -11300
rect 21812 -11248 21868 -11246
rect 21812 -11300 21814 -11248
rect 21814 -11300 21866 -11248
rect 21866 -11300 21868 -11248
rect 21812 -11302 21868 -11300
rect 22132 -11248 22188 -11246
rect 22132 -11300 22134 -11248
rect 22134 -11300 22186 -11248
rect 22186 -11300 22188 -11248
rect 22132 -11302 22188 -11300
rect 22452 -11248 22508 -11246
rect 22452 -11300 22454 -11248
rect 22454 -11300 22506 -11248
rect 22506 -11300 22508 -11248
rect 22452 -11302 22508 -11300
rect 22772 -11248 22828 -11246
rect 22772 -11300 22774 -11248
rect 22774 -11300 22826 -11248
rect 22826 -11300 22828 -11248
rect 22772 -11302 22828 -11300
rect 23092 -11248 23148 -11246
rect 23092 -11300 23094 -11248
rect 23094 -11300 23146 -11248
rect 23146 -11300 23148 -11248
rect 23092 -11302 23148 -11300
rect 23412 -11248 23468 -11246
rect 23412 -11300 23414 -11248
rect 23414 -11300 23466 -11248
rect 23466 -11300 23468 -11248
rect 23412 -11302 23468 -11300
rect 23732 -11248 23788 -11246
rect 23732 -11300 23734 -11248
rect 23734 -11300 23786 -11248
rect 23786 -11300 23788 -11248
rect 23732 -11302 23788 -11300
rect 24052 -11248 24108 -11246
rect 24052 -11300 24054 -11248
rect 24054 -11300 24106 -11248
rect 24106 -11300 24108 -11248
rect 24052 -11302 24108 -11300
rect 24372 -11248 24428 -11246
rect 24372 -11300 24374 -11248
rect 24374 -11300 24426 -11248
rect 24426 -11300 24428 -11248
rect 24372 -11302 24428 -11300
rect 24692 -11248 24748 -11246
rect 24692 -11300 24694 -11248
rect 24694 -11300 24746 -11248
rect 24746 -11300 24748 -11248
rect 24692 -11302 24748 -11300
rect 25012 -11248 25068 -11246
rect 25012 -11300 25014 -11248
rect 25014 -11300 25066 -11248
rect 25066 -11300 25068 -11248
rect 25012 -11302 25068 -11300
rect 25332 -11248 25388 -11246
rect 25332 -11300 25334 -11248
rect 25334 -11300 25386 -11248
rect 25386 -11300 25388 -11248
rect 25332 -11302 25388 -11300
rect 6242 -11454 6298 -11452
rect 6242 -11506 6244 -11454
rect 6244 -11506 6296 -11454
rect 6296 -11506 6298 -11454
rect 6242 -11508 6298 -11506
rect 13708 -11454 13764 -11452
rect 13708 -11506 13710 -11454
rect 13710 -11506 13762 -11454
rect 13762 -11506 13764 -11454
rect 13708 -11508 13764 -11506
rect 6242 -11774 6298 -11772
rect 6242 -11826 6244 -11774
rect 6244 -11826 6296 -11774
rect 6296 -11826 6298 -11774
rect 6242 -11828 6298 -11826
rect 6242 -12094 6298 -12092
rect 6242 -12146 6244 -12094
rect 6244 -12146 6296 -12094
rect 6296 -12146 6298 -12094
rect 6242 -12148 6298 -12146
rect 6242 -12414 6298 -12412
rect 6242 -12466 6244 -12414
rect 6244 -12466 6296 -12414
rect 6296 -12466 6298 -12414
rect 6242 -12468 6298 -12466
rect 6242 -12734 6298 -12732
rect 6242 -12786 6244 -12734
rect 6244 -12786 6296 -12734
rect 6296 -12786 6298 -12734
rect 6242 -12788 6298 -12786
rect 6242 -13054 6298 -13052
rect 6242 -13106 6244 -13054
rect 6244 -13106 6296 -13054
rect 6296 -13106 6298 -13054
rect 6242 -13108 6298 -13106
rect 6242 -13374 6298 -13372
rect 6242 -13426 6244 -13374
rect 6244 -13426 6296 -13374
rect 6296 -13426 6298 -13374
rect 6242 -13428 6298 -13426
rect 6242 -13694 6298 -13692
rect 6242 -13746 6244 -13694
rect 6244 -13746 6296 -13694
rect 6296 -13746 6298 -13694
rect 6242 -13748 6298 -13746
rect 6242 -14014 6298 -14012
rect 6242 -14066 6244 -14014
rect 6244 -14066 6296 -14014
rect 6296 -14066 6298 -14014
rect 6242 -14068 6298 -14066
rect 6242 -14334 6298 -14332
rect 6242 -14386 6244 -14334
rect 6244 -14386 6296 -14334
rect 6296 -14386 6298 -14334
rect 6242 -14388 6298 -14386
rect 6242 -14654 6298 -14652
rect 6242 -14706 6244 -14654
rect 6244 -14706 6296 -14654
rect 6296 -14706 6298 -14654
rect 6242 -14708 6298 -14706
rect 6242 -14974 6298 -14972
rect 6242 -15026 6244 -14974
rect 6244 -15026 6296 -14974
rect 6296 -15026 6298 -14974
rect 6242 -15028 6298 -15026
rect 6242 -15294 6298 -15292
rect 6242 -15346 6244 -15294
rect 6244 -15346 6296 -15294
rect 6296 -15346 6298 -15294
rect 6242 -15348 6298 -15346
rect 6242 -15614 6298 -15612
rect 6242 -15666 6244 -15614
rect 6244 -15666 6296 -15614
rect 6296 -15666 6298 -15614
rect 6242 -15668 6298 -15666
rect 6242 -15934 6298 -15932
rect 6242 -15986 6244 -15934
rect 6244 -15986 6296 -15934
rect 6296 -15986 6298 -15934
rect 6242 -15988 6298 -15986
rect 6242 -16254 6298 -16252
rect 6242 -16306 6244 -16254
rect 6244 -16306 6296 -16254
rect 6296 -16306 6298 -16254
rect 6242 -16308 6298 -16306
rect 6242 -16574 6298 -16572
rect 6242 -16626 6244 -16574
rect 6244 -16626 6296 -16574
rect 6296 -16626 6298 -16574
rect 6242 -16628 6298 -16626
rect 6242 -16894 6298 -16892
rect 6242 -16946 6244 -16894
rect 6244 -16946 6296 -16894
rect 6296 -16946 6298 -16894
rect 6242 -16948 6298 -16946
rect 6242 -17214 6298 -17212
rect 6242 -17266 6244 -17214
rect 6244 -17266 6296 -17214
rect 6296 -17266 6298 -17214
rect 6242 -17268 6298 -17266
rect 6242 -17534 6298 -17532
rect 6242 -17586 6244 -17534
rect 6244 -17586 6296 -17534
rect 6296 -17586 6298 -17534
rect 6242 -17588 6298 -17586
rect 6242 -17854 6298 -17852
rect 6242 -17906 6244 -17854
rect 6244 -17906 6296 -17854
rect 6296 -17906 6298 -17854
rect 6242 -17908 6298 -17906
rect 6242 -18174 6298 -18172
rect 6242 -18226 6244 -18174
rect 6244 -18226 6296 -18174
rect 6296 -18226 6298 -18174
rect 6242 -18228 6298 -18226
rect 13708 -11774 13764 -11772
rect 13708 -11826 13710 -11774
rect 13710 -11826 13762 -11774
rect 13762 -11826 13764 -11774
rect 13708 -11828 13764 -11826
rect 13708 -12094 13764 -12092
rect 13708 -12146 13710 -12094
rect 13710 -12146 13762 -12094
rect 13762 -12146 13764 -12094
rect 13708 -12148 13764 -12146
rect 13708 -12414 13764 -12412
rect 13708 -12466 13710 -12414
rect 13710 -12466 13762 -12414
rect 13762 -12466 13764 -12414
rect 13708 -12468 13764 -12466
rect 13708 -12734 13764 -12732
rect 13708 -12786 13710 -12734
rect 13710 -12786 13762 -12734
rect 13762 -12786 13764 -12734
rect 13708 -12788 13764 -12786
rect 13708 -13054 13764 -13052
rect 13708 -13106 13710 -13054
rect 13710 -13106 13762 -13054
rect 13762 -13106 13764 -13054
rect 13708 -13108 13764 -13106
rect 13708 -13374 13764 -13372
rect 13708 -13426 13710 -13374
rect 13710 -13426 13762 -13374
rect 13762 -13426 13764 -13374
rect 13708 -13428 13764 -13426
rect 13708 -13694 13764 -13692
rect 13708 -13746 13710 -13694
rect 13710 -13746 13762 -13694
rect 13762 -13746 13764 -13694
rect 13708 -13748 13764 -13746
rect 13708 -14014 13764 -14012
rect 13708 -14066 13710 -14014
rect 13710 -14066 13762 -14014
rect 13762 -14066 13764 -14014
rect 13708 -14068 13764 -14066
rect 13708 -14334 13764 -14332
rect 13708 -14386 13710 -14334
rect 13710 -14386 13762 -14334
rect 13762 -14386 13764 -14334
rect 13708 -14388 13764 -14386
rect 13708 -14654 13764 -14652
rect 13708 -14706 13710 -14654
rect 13710 -14706 13762 -14654
rect 13762 -14706 13764 -14654
rect 13708 -14708 13764 -14706
rect 13708 -14974 13764 -14972
rect 13708 -15026 13710 -14974
rect 13710 -15026 13762 -14974
rect 13762 -15026 13764 -14974
rect 13708 -15028 13764 -15026
rect 13708 -15294 13764 -15292
rect 13708 -15346 13710 -15294
rect 13710 -15346 13762 -15294
rect 13762 -15346 13764 -15294
rect 13708 -15348 13764 -15346
rect 13708 -15614 13764 -15612
rect 13708 -15666 13710 -15614
rect 13710 -15666 13762 -15614
rect 13762 -15666 13764 -15614
rect 13708 -15668 13764 -15666
rect 13708 -15934 13764 -15932
rect 13708 -15986 13710 -15934
rect 13710 -15986 13762 -15934
rect 13762 -15986 13764 -15934
rect 13708 -15988 13764 -15986
rect 13708 -16254 13764 -16252
rect 13708 -16306 13710 -16254
rect 13710 -16306 13762 -16254
rect 13762 -16306 13764 -16254
rect 13708 -16308 13764 -16306
rect 13708 -16574 13764 -16572
rect 13708 -16626 13710 -16574
rect 13710 -16626 13762 -16574
rect 13762 -16626 13764 -16574
rect 13708 -16628 13764 -16626
rect 13708 -16894 13764 -16892
rect 13708 -16946 13710 -16894
rect 13710 -16946 13762 -16894
rect 13762 -16946 13764 -16894
rect 13708 -16948 13764 -16946
rect 13708 -17214 13764 -17212
rect 13708 -17266 13710 -17214
rect 13710 -17266 13762 -17214
rect 13762 -17266 13764 -17214
rect 13708 -17268 13764 -17266
rect 13708 -17534 13764 -17532
rect 13708 -17586 13710 -17534
rect 13710 -17586 13762 -17534
rect 13762 -17586 13764 -17534
rect 13708 -17588 13764 -17586
rect 13708 -17854 13764 -17852
rect 13708 -17906 13710 -17854
rect 13710 -17906 13762 -17854
rect 13762 -17906 13764 -17854
rect 13708 -17908 13764 -17906
rect 13708 -18174 13764 -18172
rect 13708 -18226 13710 -18174
rect 13710 -18226 13762 -18174
rect 13762 -18226 13764 -18174
rect 13708 -18228 13764 -18226
rect 6242 -18494 6298 -18492
rect 6242 -18546 6244 -18494
rect 6244 -18546 6296 -18494
rect 6296 -18546 6298 -18494
rect 6242 -18548 6298 -18546
rect 13708 -18494 13764 -18492
rect 13708 -18546 13710 -18494
rect 13710 -18546 13762 -18494
rect 13762 -18546 13764 -18494
rect 13708 -18548 13764 -18546
rect 6612 -18704 6668 -18702
rect 6612 -18756 6614 -18704
rect 6614 -18756 6666 -18704
rect 6666 -18756 6668 -18704
rect 6612 -18758 6668 -18756
rect 6932 -18704 6988 -18702
rect 6932 -18756 6934 -18704
rect 6934 -18756 6986 -18704
rect 6986 -18756 6988 -18704
rect 6932 -18758 6988 -18756
rect 7252 -18704 7308 -18702
rect 7252 -18756 7254 -18704
rect 7254 -18756 7306 -18704
rect 7306 -18756 7308 -18704
rect 7252 -18758 7308 -18756
rect 7572 -18704 7628 -18702
rect 7572 -18756 7574 -18704
rect 7574 -18756 7626 -18704
rect 7626 -18756 7628 -18704
rect 7572 -18758 7628 -18756
rect 7892 -18704 7948 -18702
rect 7892 -18756 7894 -18704
rect 7894 -18756 7946 -18704
rect 7946 -18756 7948 -18704
rect 7892 -18758 7948 -18756
rect 8212 -18704 8268 -18702
rect 8212 -18756 8214 -18704
rect 8214 -18756 8266 -18704
rect 8266 -18756 8268 -18704
rect 8212 -18758 8268 -18756
rect 8532 -18704 8588 -18702
rect 8532 -18756 8534 -18704
rect 8534 -18756 8586 -18704
rect 8586 -18756 8588 -18704
rect 8532 -18758 8588 -18756
rect 8852 -18704 8908 -18702
rect 8852 -18756 8854 -18704
rect 8854 -18756 8906 -18704
rect 8906 -18756 8908 -18704
rect 8852 -18758 8908 -18756
rect 9172 -18704 9228 -18702
rect 9172 -18756 9174 -18704
rect 9174 -18756 9226 -18704
rect 9226 -18756 9228 -18704
rect 9172 -18758 9228 -18756
rect 9492 -18704 9548 -18702
rect 9492 -18756 9494 -18704
rect 9494 -18756 9546 -18704
rect 9546 -18756 9548 -18704
rect 9492 -18758 9548 -18756
rect 9812 -18704 9868 -18702
rect 9812 -18756 9814 -18704
rect 9814 -18756 9866 -18704
rect 9866 -18756 9868 -18704
rect 9812 -18758 9868 -18756
rect 10132 -18704 10188 -18702
rect 10132 -18756 10134 -18704
rect 10134 -18756 10186 -18704
rect 10186 -18756 10188 -18704
rect 10132 -18758 10188 -18756
rect 10452 -18704 10508 -18702
rect 10452 -18756 10454 -18704
rect 10454 -18756 10506 -18704
rect 10506 -18756 10508 -18704
rect 10452 -18758 10508 -18756
rect 10772 -18704 10828 -18702
rect 10772 -18756 10774 -18704
rect 10774 -18756 10826 -18704
rect 10826 -18756 10828 -18704
rect 10772 -18758 10828 -18756
rect 11092 -18704 11148 -18702
rect 11092 -18756 11094 -18704
rect 11094 -18756 11146 -18704
rect 11146 -18756 11148 -18704
rect 11092 -18758 11148 -18756
rect 11412 -18704 11468 -18702
rect 11412 -18756 11414 -18704
rect 11414 -18756 11466 -18704
rect 11466 -18756 11468 -18704
rect 11412 -18758 11468 -18756
rect 11732 -18704 11788 -18702
rect 11732 -18756 11734 -18704
rect 11734 -18756 11786 -18704
rect 11786 -18756 11788 -18704
rect 11732 -18758 11788 -18756
rect 12052 -18704 12108 -18702
rect 12052 -18756 12054 -18704
rect 12054 -18756 12106 -18704
rect 12106 -18756 12108 -18704
rect 12052 -18758 12108 -18756
rect 12372 -18704 12428 -18702
rect 12372 -18756 12374 -18704
rect 12374 -18756 12426 -18704
rect 12426 -18756 12428 -18704
rect 12372 -18758 12428 -18756
rect 12692 -18704 12748 -18702
rect 12692 -18756 12694 -18704
rect 12694 -18756 12746 -18704
rect 12746 -18756 12748 -18704
rect 12692 -18758 12748 -18756
rect 13012 -18704 13068 -18702
rect 13012 -18756 13014 -18704
rect 13014 -18756 13066 -18704
rect 13066 -18756 13068 -18704
rect 13012 -18758 13068 -18756
rect 13332 -18704 13388 -18702
rect 13332 -18756 13334 -18704
rect 13334 -18756 13386 -18704
rect 13386 -18756 13388 -18704
rect 13332 -18758 13388 -18756
rect 18242 -11454 18298 -11452
rect 18242 -11506 18244 -11454
rect 18244 -11506 18296 -11454
rect 18296 -11506 18298 -11454
rect 18242 -11508 18298 -11506
rect 25708 -11454 25764 -11452
rect 25708 -11506 25710 -11454
rect 25710 -11506 25762 -11454
rect 25762 -11506 25764 -11454
rect 25708 -11508 25764 -11506
rect 18242 -11774 18298 -11772
rect 18242 -11826 18244 -11774
rect 18244 -11826 18296 -11774
rect 18296 -11826 18298 -11774
rect 18242 -11828 18298 -11826
rect 18242 -12094 18298 -12092
rect 18242 -12146 18244 -12094
rect 18244 -12146 18296 -12094
rect 18296 -12146 18298 -12094
rect 18242 -12148 18298 -12146
rect 18242 -12414 18298 -12412
rect 18242 -12466 18244 -12414
rect 18244 -12466 18296 -12414
rect 18296 -12466 18298 -12414
rect 18242 -12468 18298 -12466
rect 18242 -12734 18298 -12732
rect 18242 -12786 18244 -12734
rect 18244 -12786 18296 -12734
rect 18296 -12786 18298 -12734
rect 18242 -12788 18298 -12786
rect 18242 -13054 18298 -13052
rect 18242 -13106 18244 -13054
rect 18244 -13106 18296 -13054
rect 18296 -13106 18298 -13054
rect 18242 -13108 18298 -13106
rect 18242 -13374 18298 -13372
rect 18242 -13426 18244 -13374
rect 18244 -13426 18296 -13374
rect 18296 -13426 18298 -13374
rect 18242 -13428 18298 -13426
rect 18242 -13694 18298 -13692
rect 18242 -13746 18244 -13694
rect 18244 -13746 18296 -13694
rect 18296 -13746 18298 -13694
rect 18242 -13748 18298 -13746
rect 18242 -14014 18298 -14012
rect 18242 -14066 18244 -14014
rect 18244 -14066 18296 -14014
rect 18296 -14066 18298 -14014
rect 18242 -14068 18298 -14066
rect 18242 -14334 18298 -14332
rect 18242 -14386 18244 -14334
rect 18244 -14386 18296 -14334
rect 18296 -14386 18298 -14334
rect 18242 -14388 18298 -14386
rect 18242 -14654 18298 -14652
rect 18242 -14706 18244 -14654
rect 18244 -14706 18296 -14654
rect 18296 -14706 18298 -14654
rect 18242 -14708 18298 -14706
rect 18242 -14974 18298 -14972
rect 18242 -15026 18244 -14974
rect 18244 -15026 18296 -14974
rect 18296 -15026 18298 -14974
rect 18242 -15028 18298 -15026
rect 18242 -15294 18298 -15292
rect 18242 -15346 18244 -15294
rect 18244 -15346 18296 -15294
rect 18296 -15346 18298 -15294
rect 18242 -15348 18298 -15346
rect 18242 -15614 18298 -15612
rect 18242 -15666 18244 -15614
rect 18244 -15666 18296 -15614
rect 18296 -15666 18298 -15614
rect 18242 -15668 18298 -15666
rect 18242 -15934 18298 -15932
rect 18242 -15986 18244 -15934
rect 18244 -15986 18296 -15934
rect 18296 -15986 18298 -15934
rect 18242 -15988 18298 -15986
rect 18242 -16254 18298 -16252
rect 18242 -16306 18244 -16254
rect 18244 -16306 18296 -16254
rect 18296 -16306 18298 -16254
rect 18242 -16308 18298 -16306
rect 18242 -16574 18298 -16572
rect 18242 -16626 18244 -16574
rect 18244 -16626 18296 -16574
rect 18296 -16626 18298 -16574
rect 18242 -16628 18298 -16626
rect 18242 -16894 18298 -16892
rect 18242 -16946 18244 -16894
rect 18244 -16946 18296 -16894
rect 18296 -16946 18298 -16894
rect 18242 -16948 18298 -16946
rect 18242 -17214 18298 -17212
rect 18242 -17266 18244 -17214
rect 18244 -17266 18296 -17214
rect 18296 -17266 18298 -17214
rect 18242 -17268 18298 -17266
rect 18242 -17534 18298 -17532
rect 18242 -17586 18244 -17534
rect 18244 -17586 18296 -17534
rect 18296 -17586 18298 -17534
rect 18242 -17588 18298 -17586
rect 18242 -17854 18298 -17852
rect 18242 -17906 18244 -17854
rect 18244 -17906 18296 -17854
rect 18296 -17906 18298 -17854
rect 18242 -17908 18298 -17906
rect 18242 -18174 18298 -18172
rect 18242 -18226 18244 -18174
rect 18244 -18226 18296 -18174
rect 18296 -18226 18298 -18174
rect 18242 -18228 18298 -18226
rect 25708 -11774 25764 -11772
rect 25708 -11826 25710 -11774
rect 25710 -11826 25762 -11774
rect 25762 -11826 25764 -11774
rect 25708 -11828 25764 -11826
rect 25708 -12094 25764 -12092
rect 25708 -12146 25710 -12094
rect 25710 -12146 25762 -12094
rect 25762 -12146 25764 -12094
rect 25708 -12148 25764 -12146
rect 25708 -12414 25764 -12412
rect 25708 -12466 25710 -12414
rect 25710 -12466 25762 -12414
rect 25762 -12466 25764 -12414
rect 25708 -12468 25764 -12466
rect 25708 -12734 25764 -12732
rect 25708 -12786 25710 -12734
rect 25710 -12786 25762 -12734
rect 25762 -12786 25764 -12734
rect 25708 -12788 25764 -12786
rect 25708 -13054 25764 -13052
rect 25708 -13106 25710 -13054
rect 25710 -13106 25762 -13054
rect 25762 -13106 25764 -13054
rect 25708 -13108 25764 -13106
rect 25708 -13374 25764 -13372
rect 25708 -13426 25710 -13374
rect 25710 -13426 25762 -13374
rect 25762 -13426 25764 -13374
rect 25708 -13428 25764 -13426
rect 25708 -13694 25764 -13692
rect 25708 -13746 25710 -13694
rect 25710 -13746 25762 -13694
rect 25762 -13746 25764 -13694
rect 25708 -13748 25764 -13746
rect 25708 -14014 25764 -14012
rect 25708 -14066 25710 -14014
rect 25710 -14066 25762 -14014
rect 25762 -14066 25764 -14014
rect 25708 -14068 25764 -14066
rect 25708 -14334 25764 -14332
rect 25708 -14386 25710 -14334
rect 25710 -14386 25762 -14334
rect 25762 -14386 25764 -14334
rect 25708 -14388 25764 -14386
rect 25708 -14654 25764 -14652
rect 25708 -14706 25710 -14654
rect 25710 -14706 25762 -14654
rect 25762 -14706 25764 -14654
rect 25708 -14708 25764 -14706
rect 25708 -14974 25764 -14972
rect 25708 -15026 25710 -14974
rect 25710 -15026 25762 -14974
rect 25762 -15026 25764 -14974
rect 25708 -15028 25764 -15026
rect 25708 -15294 25764 -15292
rect 25708 -15346 25710 -15294
rect 25710 -15346 25762 -15294
rect 25762 -15346 25764 -15294
rect 25708 -15348 25764 -15346
rect 25708 -15614 25764 -15612
rect 25708 -15666 25710 -15614
rect 25710 -15666 25762 -15614
rect 25762 -15666 25764 -15614
rect 25708 -15668 25764 -15666
rect 25708 -15934 25764 -15932
rect 25708 -15986 25710 -15934
rect 25710 -15986 25762 -15934
rect 25762 -15986 25764 -15934
rect 25708 -15988 25764 -15986
rect 25708 -16254 25764 -16252
rect 25708 -16306 25710 -16254
rect 25710 -16306 25762 -16254
rect 25762 -16306 25764 -16254
rect 25708 -16308 25764 -16306
rect 25708 -16574 25764 -16572
rect 25708 -16626 25710 -16574
rect 25710 -16626 25762 -16574
rect 25762 -16626 25764 -16574
rect 25708 -16628 25764 -16626
rect 25708 -16894 25764 -16892
rect 25708 -16946 25710 -16894
rect 25710 -16946 25762 -16894
rect 25762 -16946 25764 -16894
rect 25708 -16948 25764 -16946
rect 25708 -17214 25764 -17212
rect 25708 -17266 25710 -17214
rect 25710 -17266 25762 -17214
rect 25762 -17266 25764 -17214
rect 25708 -17268 25764 -17266
rect 25708 -17534 25764 -17532
rect 25708 -17586 25710 -17534
rect 25710 -17586 25762 -17534
rect 25762 -17586 25764 -17534
rect 25708 -17588 25764 -17586
rect 25708 -17854 25764 -17852
rect 25708 -17906 25710 -17854
rect 25710 -17906 25762 -17854
rect 25762 -17906 25764 -17854
rect 25708 -17908 25764 -17906
rect 25708 -18174 25764 -18172
rect 25708 -18226 25710 -18174
rect 25710 -18226 25762 -18174
rect 25762 -18226 25764 -18174
rect 25708 -18228 25764 -18226
rect 18242 -18494 18298 -18492
rect 18242 -18546 18244 -18494
rect 18244 -18546 18296 -18494
rect 18296 -18546 18298 -18494
rect 18242 -18548 18298 -18546
rect 25708 -18494 25764 -18492
rect 25708 -18546 25710 -18494
rect 25710 -18546 25762 -18494
rect 25762 -18546 25764 -18494
rect 25708 -18548 25764 -18546
rect 18612 -18704 18668 -18702
rect 18612 -18756 18614 -18704
rect 18614 -18756 18666 -18704
rect 18666 -18756 18668 -18704
rect 18612 -18758 18668 -18756
rect 18932 -18704 18988 -18702
rect 18932 -18756 18934 -18704
rect 18934 -18756 18986 -18704
rect 18986 -18756 18988 -18704
rect 18932 -18758 18988 -18756
rect 19252 -18704 19308 -18702
rect 19252 -18756 19254 -18704
rect 19254 -18756 19306 -18704
rect 19306 -18756 19308 -18704
rect 19252 -18758 19308 -18756
rect 19572 -18704 19628 -18702
rect 19572 -18756 19574 -18704
rect 19574 -18756 19626 -18704
rect 19626 -18756 19628 -18704
rect 19572 -18758 19628 -18756
rect 19892 -18704 19948 -18702
rect 19892 -18756 19894 -18704
rect 19894 -18756 19946 -18704
rect 19946 -18756 19948 -18704
rect 19892 -18758 19948 -18756
rect 20212 -18704 20268 -18702
rect 20212 -18756 20214 -18704
rect 20214 -18756 20266 -18704
rect 20266 -18756 20268 -18704
rect 20212 -18758 20268 -18756
rect 20532 -18704 20588 -18702
rect 20532 -18756 20534 -18704
rect 20534 -18756 20586 -18704
rect 20586 -18756 20588 -18704
rect 20532 -18758 20588 -18756
rect 20852 -18704 20908 -18702
rect 20852 -18756 20854 -18704
rect 20854 -18756 20906 -18704
rect 20906 -18756 20908 -18704
rect 20852 -18758 20908 -18756
rect 21172 -18704 21228 -18702
rect 21172 -18756 21174 -18704
rect 21174 -18756 21226 -18704
rect 21226 -18756 21228 -18704
rect 21172 -18758 21228 -18756
rect 21492 -18704 21548 -18702
rect 21492 -18756 21494 -18704
rect 21494 -18756 21546 -18704
rect 21546 -18756 21548 -18704
rect 21492 -18758 21548 -18756
rect 21812 -18704 21868 -18702
rect 21812 -18756 21814 -18704
rect 21814 -18756 21866 -18704
rect 21866 -18756 21868 -18704
rect 21812 -18758 21868 -18756
rect 22132 -18704 22188 -18702
rect 22132 -18756 22134 -18704
rect 22134 -18756 22186 -18704
rect 22186 -18756 22188 -18704
rect 22132 -18758 22188 -18756
rect 22452 -18704 22508 -18702
rect 22452 -18756 22454 -18704
rect 22454 -18756 22506 -18704
rect 22506 -18756 22508 -18704
rect 22452 -18758 22508 -18756
rect 22772 -18704 22828 -18702
rect 22772 -18756 22774 -18704
rect 22774 -18756 22826 -18704
rect 22826 -18756 22828 -18704
rect 22772 -18758 22828 -18756
rect 23092 -18704 23148 -18702
rect 23092 -18756 23094 -18704
rect 23094 -18756 23146 -18704
rect 23146 -18756 23148 -18704
rect 23092 -18758 23148 -18756
rect 23412 -18704 23468 -18702
rect 23412 -18756 23414 -18704
rect 23414 -18756 23466 -18704
rect 23466 -18756 23468 -18704
rect 23412 -18758 23468 -18756
rect 23732 -18704 23788 -18702
rect 23732 -18756 23734 -18704
rect 23734 -18756 23786 -18704
rect 23786 -18756 23788 -18704
rect 23732 -18758 23788 -18756
rect 24052 -18704 24108 -18702
rect 24052 -18756 24054 -18704
rect 24054 -18756 24106 -18704
rect 24106 -18756 24108 -18704
rect 24052 -18758 24108 -18756
rect 24372 -18704 24428 -18702
rect 24372 -18756 24374 -18704
rect 24374 -18756 24426 -18704
rect 24426 -18756 24428 -18704
rect 24372 -18758 24428 -18756
rect 24692 -18704 24748 -18702
rect 24692 -18756 24694 -18704
rect 24694 -18756 24746 -18704
rect 24746 -18756 24748 -18704
rect 24692 -18758 24748 -18756
rect 25012 -18704 25068 -18702
rect 25012 -18756 25014 -18704
rect 25014 -18756 25066 -18704
rect 25066 -18756 25068 -18704
rect 25012 -18758 25068 -18756
rect 25332 -18704 25388 -18702
rect 25332 -18756 25334 -18704
rect 25334 -18756 25386 -18704
rect 25386 -18756 25388 -18704
rect 25332 -18758 25388 -18756
rect 30612 -11248 30668 -11246
rect 30612 -11300 30614 -11248
rect 30614 -11300 30666 -11248
rect 30666 -11300 30668 -11248
rect 30612 -11302 30668 -11300
rect 30932 -11248 30988 -11246
rect 30932 -11300 30934 -11248
rect 30934 -11300 30986 -11248
rect 30986 -11300 30988 -11248
rect 30932 -11302 30988 -11300
rect 31252 -11248 31308 -11246
rect 31252 -11300 31254 -11248
rect 31254 -11300 31306 -11248
rect 31306 -11300 31308 -11248
rect 31252 -11302 31308 -11300
rect 31572 -11248 31628 -11246
rect 31572 -11300 31574 -11248
rect 31574 -11300 31626 -11248
rect 31626 -11300 31628 -11248
rect 31572 -11302 31628 -11300
rect 31892 -11248 31948 -11246
rect 31892 -11300 31894 -11248
rect 31894 -11300 31946 -11248
rect 31946 -11300 31948 -11248
rect 31892 -11302 31948 -11300
rect 32212 -11248 32268 -11246
rect 32212 -11300 32214 -11248
rect 32214 -11300 32266 -11248
rect 32266 -11300 32268 -11248
rect 32212 -11302 32268 -11300
rect 32532 -11248 32588 -11246
rect 32532 -11300 32534 -11248
rect 32534 -11300 32586 -11248
rect 32586 -11300 32588 -11248
rect 32532 -11302 32588 -11300
rect 32852 -11248 32908 -11246
rect 32852 -11300 32854 -11248
rect 32854 -11300 32906 -11248
rect 32906 -11300 32908 -11248
rect 32852 -11302 32908 -11300
rect 33172 -11248 33228 -11246
rect 33172 -11300 33174 -11248
rect 33174 -11300 33226 -11248
rect 33226 -11300 33228 -11248
rect 33172 -11302 33228 -11300
rect 33492 -11248 33548 -11246
rect 33492 -11300 33494 -11248
rect 33494 -11300 33546 -11248
rect 33546 -11300 33548 -11248
rect 33492 -11302 33548 -11300
rect 33812 -11248 33868 -11246
rect 33812 -11300 33814 -11248
rect 33814 -11300 33866 -11248
rect 33866 -11300 33868 -11248
rect 33812 -11302 33868 -11300
rect 34132 -11248 34188 -11246
rect 34132 -11300 34134 -11248
rect 34134 -11300 34186 -11248
rect 34186 -11300 34188 -11248
rect 34132 -11302 34188 -11300
rect 34452 -11248 34508 -11246
rect 34452 -11300 34454 -11248
rect 34454 -11300 34506 -11248
rect 34506 -11300 34508 -11248
rect 34452 -11302 34508 -11300
rect 34772 -11248 34828 -11246
rect 34772 -11300 34774 -11248
rect 34774 -11300 34826 -11248
rect 34826 -11300 34828 -11248
rect 34772 -11302 34828 -11300
rect 35092 -11248 35148 -11246
rect 35092 -11300 35094 -11248
rect 35094 -11300 35146 -11248
rect 35146 -11300 35148 -11248
rect 35092 -11302 35148 -11300
rect 35412 -11248 35468 -11246
rect 35412 -11300 35414 -11248
rect 35414 -11300 35466 -11248
rect 35466 -11300 35468 -11248
rect 35412 -11302 35468 -11300
rect 35732 -11248 35788 -11246
rect 35732 -11300 35734 -11248
rect 35734 -11300 35786 -11248
rect 35786 -11300 35788 -11248
rect 35732 -11302 35788 -11300
rect 36052 -11248 36108 -11246
rect 36052 -11300 36054 -11248
rect 36054 -11300 36106 -11248
rect 36106 -11300 36108 -11248
rect 36052 -11302 36108 -11300
rect 36372 -11248 36428 -11246
rect 36372 -11300 36374 -11248
rect 36374 -11300 36426 -11248
rect 36426 -11300 36428 -11248
rect 36372 -11302 36428 -11300
rect 36692 -11248 36748 -11246
rect 36692 -11300 36694 -11248
rect 36694 -11300 36746 -11248
rect 36746 -11300 36748 -11248
rect 36692 -11302 36748 -11300
rect 37012 -11248 37068 -11246
rect 37012 -11300 37014 -11248
rect 37014 -11300 37066 -11248
rect 37066 -11300 37068 -11248
rect 37012 -11302 37068 -11300
rect 37332 -11248 37388 -11246
rect 37332 -11300 37334 -11248
rect 37334 -11300 37386 -11248
rect 37386 -11300 37388 -11248
rect 37332 -11302 37388 -11300
rect 30242 -11454 30298 -11452
rect 30242 -11506 30244 -11454
rect 30244 -11506 30296 -11454
rect 30296 -11506 30298 -11454
rect 30242 -11508 30298 -11506
rect 37708 -11454 37764 -11452
rect 37708 -11506 37710 -11454
rect 37710 -11506 37762 -11454
rect 37762 -11506 37764 -11454
rect 37708 -11508 37764 -11506
rect 30242 -11774 30298 -11772
rect 30242 -11826 30244 -11774
rect 30244 -11826 30296 -11774
rect 30296 -11826 30298 -11774
rect 30242 -11828 30298 -11826
rect 30242 -12094 30298 -12092
rect 30242 -12146 30244 -12094
rect 30244 -12146 30296 -12094
rect 30296 -12146 30298 -12094
rect 30242 -12148 30298 -12146
rect 30242 -12414 30298 -12412
rect 30242 -12466 30244 -12414
rect 30244 -12466 30296 -12414
rect 30296 -12466 30298 -12414
rect 30242 -12468 30298 -12466
rect 30242 -12734 30298 -12732
rect 30242 -12786 30244 -12734
rect 30244 -12786 30296 -12734
rect 30296 -12786 30298 -12734
rect 30242 -12788 30298 -12786
rect 30242 -13054 30298 -13052
rect 30242 -13106 30244 -13054
rect 30244 -13106 30296 -13054
rect 30296 -13106 30298 -13054
rect 30242 -13108 30298 -13106
rect 30242 -13374 30298 -13372
rect 30242 -13426 30244 -13374
rect 30244 -13426 30296 -13374
rect 30296 -13426 30298 -13374
rect 30242 -13428 30298 -13426
rect 30242 -13694 30298 -13692
rect 30242 -13746 30244 -13694
rect 30244 -13746 30296 -13694
rect 30296 -13746 30298 -13694
rect 30242 -13748 30298 -13746
rect 30242 -14014 30298 -14012
rect 30242 -14066 30244 -14014
rect 30244 -14066 30296 -14014
rect 30296 -14066 30298 -14014
rect 30242 -14068 30298 -14066
rect 30242 -14334 30298 -14332
rect 30242 -14386 30244 -14334
rect 30244 -14386 30296 -14334
rect 30296 -14386 30298 -14334
rect 30242 -14388 30298 -14386
rect 30242 -14654 30298 -14652
rect 30242 -14706 30244 -14654
rect 30244 -14706 30296 -14654
rect 30296 -14706 30298 -14654
rect 30242 -14708 30298 -14706
rect 30242 -14974 30298 -14972
rect 30242 -15026 30244 -14974
rect 30244 -15026 30296 -14974
rect 30296 -15026 30298 -14974
rect 30242 -15028 30298 -15026
rect 30242 -15294 30298 -15292
rect 30242 -15346 30244 -15294
rect 30244 -15346 30296 -15294
rect 30296 -15346 30298 -15294
rect 30242 -15348 30298 -15346
rect 30242 -15614 30298 -15612
rect 30242 -15666 30244 -15614
rect 30244 -15666 30296 -15614
rect 30296 -15666 30298 -15614
rect 30242 -15668 30298 -15666
rect 30242 -15934 30298 -15932
rect 30242 -15986 30244 -15934
rect 30244 -15986 30296 -15934
rect 30296 -15986 30298 -15934
rect 30242 -15988 30298 -15986
rect 30242 -16254 30298 -16252
rect 30242 -16306 30244 -16254
rect 30244 -16306 30296 -16254
rect 30296 -16306 30298 -16254
rect 30242 -16308 30298 -16306
rect 30242 -16574 30298 -16572
rect 30242 -16626 30244 -16574
rect 30244 -16626 30296 -16574
rect 30296 -16626 30298 -16574
rect 30242 -16628 30298 -16626
rect 30242 -16894 30298 -16892
rect 30242 -16946 30244 -16894
rect 30244 -16946 30296 -16894
rect 30296 -16946 30298 -16894
rect 30242 -16948 30298 -16946
rect 30242 -17214 30298 -17212
rect 30242 -17266 30244 -17214
rect 30244 -17266 30296 -17214
rect 30296 -17266 30298 -17214
rect 30242 -17268 30298 -17266
rect 30242 -17534 30298 -17532
rect 30242 -17586 30244 -17534
rect 30244 -17586 30296 -17534
rect 30296 -17586 30298 -17534
rect 30242 -17588 30298 -17586
rect 30242 -17854 30298 -17852
rect 30242 -17906 30244 -17854
rect 30244 -17906 30296 -17854
rect 30296 -17906 30298 -17854
rect 30242 -17908 30298 -17906
rect 30242 -18174 30298 -18172
rect 30242 -18226 30244 -18174
rect 30244 -18226 30296 -18174
rect 30296 -18226 30298 -18174
rect 30242 -18228 30298 -18226
rect 37708 -11774 37764 -11772
rect 37708 -11826 37710 -11774
rect 37710 -11826 37762 -11774
rect 37762 -11826 37764 -11774
rect 37708 -11828 37764 -11826
rect 37708 -12094 37764 -12092
rect 37708 -12146 37710 -12094
rect 37710 -12146 37762 -12094
rect 37762 -12146 37764 -12094
rect 37708 -12148 37764 -12146
rect 37708 -12414 37764 -12412
rect 37708 -12466 37710 -12414
rect 37710 -12466 37762 -12414
rect 37762 -12466 37764 -12414
rect 37708 -12468 37764 -12466
rect 37708 -12734 37764 -12732
rect 37708 -12786 37710 -12734
rect 37710 -12786 37762 -12734
rect 37762 -12786 37764 -12734
rect 37708 -12788 37764 -12786
rect 37708 -13054 37764 -13052
rect 37708 -13106 37710 -13054
rect 37710 -13106 37762 -13054
rect 37762 -13106 37764 -13054
rect 37708 -13108 37764 -13106
rect 37708 -13374 37764 -13372
rect 37708 -13426 37710 -13374
rect 37710 -13426 37762 -13374
rect 37762 -13426 37764 -13374
rect 37708 -13428 37764 -13426
rect 37708 -13694 37764 -13692
rect 37708 -13746 37710 -13694
rect 37710 -13746 37762 -13694
rect 37762 -13746 37764 -13694
rect 37708 -13748 37764 -13746
rect 37708 -14014 37764 -14012
rect 37708 -14066 37710 -14014
rect 37710 -14066 37762 -14014
rect 37762 -14066 37764 -14014
rect 37708 -14068 37764 -14066
rect 37708 -14334 37764 -14332
rect 37708 -14386 37710 -14334
rect 37710 -14386 37762 -14334
rect 37762 -14386 37764 -14334
rect 37708 -14388 37764 -14386
rect 37708 -14654 37764 -14652
rect 37708 -14706 37710 -14654
rect 37710 -14706 37762 -14654
rect 37762 -14706 37764 -14654
rect 37708 -14708 37764 -14706
rect 37708 -14974 37764 -14972
rect 37708 -15026 37710 -14974
rect 37710 -15026 37762 -14974
rect 37762 -15026 37764 -14974
rect 37708 -15028 37764 -15026
rect 37708 -15294 37764 -15292
rect 37708 -15346 37710 -15294
rect 37710 -15346 37762 -15294
rect 37762 -15346 37764 -15294
rect 37708 -15348 37764 -15346
rect 37708 -15614 37764 -15612
rect 37708 -15666 37710 -15614
rect 37710 -15666 37762 -15614
rect 37762 -15666 37764 -15614
rect 37708 -15668 37764 -15666
rect 37708 -15934 37764 -15932
rect 37708 -15986 37710 -15934
rect 37710 -15986 37762 -15934
rect 37762 -15986 37764 -15934
rect 37708 -15988 37764 -15986
rect 37708 -16254 37764 -16252
rect 37708 -16306 37710 -16254
rect 37710 -16306 37762 -16254
rect 37762 -16306 37764 -16254
rect 37708 -16308 37764 -16306
rect 37708 -16574 37764 -16572
rect 37708 -16626 37710 -16574
rect 37710 -16626 37762 -16574
rect 37762 -16626 37764 -16574
rect 37708 -16628 37764 -16626
rect 37708 -16894 37764 -16892
rect 37708 -16946 37710 -16894
rect 37710 -16946 37762 -16894
rect 37762 -16946 37764 -16894
rect 37708 -16948 37764 -16946
rect 37708 -17214 37764 -17212
rect 37708 -17266 37710 -17214
rect 37710 -17266 37762 -17214
rect 37762 -17266 37764 -17214
rect 37708 -17268 37764 -17266
rect 37708 -17534 37764 -17532
rect 37708 -17586 37710 -17534
rect 37710 -17586 37762 -17534
rect 37762 -17586 37764 -17534
rect 37708 -17588 37764 -17586
rect 37708 -17854 37764 -17852
rect 37708 -17906 37710 -17854
rect 37710 -17906 37762 -17854
rect 37762 -17906 37764 -17854
rect 37708 -17908 37764 -17906
rect 37708 -18174 37764 -18172
rect 37708 -18226 37710 -18174
rect 37710 -18226 37762 -18174
rect 37762 -18226 37764 -18174
rect 37708 -18228 37764 -18226
rect 30242 -18494 30298 -18492
rect 30242 -18546 30244 -18494
rect 30244 -18546 30296 -18494
rect 30296 -18546 30298 -18494
rect 30242 -18548 30298 -18546
rect 37708 -18494 37764 -18492
rect 37708 -18546 37710 -18494
rect 37710 -18546 37762 -18494
rect 37762 -18546 37764 -18494
rect 37708 -18548 37764 -18546
rect 30612 -18704 30668 -18702
rect 30612 -18756 30614 -18704
rect 30614 -18756 30666 -18704
rect 30666 -18756 30668 -18704
rect 30612 -18758 30668 -18756
rect 30932 -18704 30988 -18702
rect 30932 -18756 30934 -18704
rect 30934 -18756 30986 -18704
rect 30986 -18756 30988 -18704
rect 30932 -18758 30988 -18756
rect 31252 -18704 31308 -18702
rect 31252 -18756 31254 -18704
rect 31254 -18756 31306 -18704
rect 31306 -18756 31308 -18704
rect 31252 -18758 31308 -18756
rect 31572 -18704 31628 -18702
rect 31572 -18756 31574 -18704
rect 31574 -18756 31626 -18704
rect 31626 -18756 31628 -18704
rect 31572 -18758 31628 -18756
rect 31892 -18704 31948 -18702
rect 31892 -18756 31894 -18704
rect 31894 -18756 31946 -18704
rect 31946 -18756 31948 -18704
rect 31892 -18758 31948 -18756
rect 32212 -18704 32268 -18702
rect 32212 -18756 32214 -18704
rect 32214 -18756 32266 -18704
rect 32266 -18756 32268 -18704
rect 32212 -18758 32268 -18756
rect 32532 -18704 32588 -18702
rect 32532 -18756 32534 -18704
rect 32534 -18756 32586 -18704
rect 32586 -18756 32588 -18704
rect 32532 -18758 32588 -18756
rect 32852 -18704 32908 -18702
rect 32852 -18756 32854 -18704
rect 32854 -18756 32906 -18704
rect 32906 -18756 32908 -18704
rect 32852 -18758 32908 -18756
rect 33172 -18704 33228 -18702
rect 33172 -18756 33174 -18704
rect 33174 -18756 33226 -18704
rect 33226 -18756 33228 -18704
rect 33172 -18758 33228 -18756
rect 33492 -18704 33548 -18702
rect 33492 -18756 33494 -18704
rect 33494 -18756 33546 -18704
rect 33546 -18756 33548 -18704
rect 33492 -18758 33548 -18756
rect 33812 -18704 33868 -18702
rect 33812 -18756 33814 -18704
rect 33814 -18756 33866 -18704
rect 33866 -18756 33868 -18704
rect 33812 -18758 33868 -18756
rect 34132 -18704 34188 -18702
rect 34132 -18756 34134 -18704
rect 34134 -18756 34186 -18704
rect 34186 -18756 34188 -18704
rect 34132 -18758 34188 -18756
rect 34452 -18704 34508 -18702
rect 34452 -18756 34454 -18704
rect 34454 -18756 34506 -18704
rect 34506 -18756 34508 -18704
rect 34452 -18758 34508 -18756
rect 34772 -18704 34828 -18702
rect 34772 -18756 34774 -18704
rect 34774 -18756 34826 -18704
rect 34826 -18756 34828 -18704
rect 34772 -18758 34828 -18756
rect 35092 -18704 35148 -18702
rect 35092 -18756 35094 -18704
rect 35094 -18756 35146 -18704
rect 35146 -18756 35148 -18704
rect 35092 -18758 35148 -18756
rect 35412 -18704 35468 -18702
rect 35412 -18756 35414 -18704
rect 35414 -18756 35466 -18704
rect 35466 -18756 35468 -18704
rect 35412 -18758 35468 -18756
rect 35732 -18704 35788 -18702
rect 35732 -18756 35734 -18704
rect 35734 -18756 35786 -18704
rect 35786 -18756 35788 -18704
rect 35732 -18758 35788 -18756
rect 36052 -18704 36108 -18702
rect 36052 -18756 36054 -18704
rect 36054 -18756 36106 -18704
rect 36106 -18756 36108 -18704
rect 36052 -18758 36108 -18756
rect 36372 -18704 36428 -18702
rect 36372 -18756 36374 -18704
rect 36374 -18756 36426 -18704
rect 36426 -18756 36428 -18704
rect 36372 -18758 36428 -18756
rect 36692 -18704 36748 -18702
rect 36692 -18756 36694 -18704
rect 36694 -18756 36746 -18704
rect 36746 -18756 36748 -18704
rect 36692 -18758 36748 -18756
rect 37012 -18704 37068 -18702
rect 37012 -18756 37014 -18704
rect 37014 -18756 37066 -18704
rect 37066 -18756 37068 -18704
rect 37012 -18758 37068 -18756
rect 37332 -18704 37388 -18702
rect 37332 -18756 37334 -18704
rect 37334 -18756 37386 -18704
rect 37386 -18756 37388 -18704
rect 37332 -18758 37388 -18756
rect 42612 -11248 42668 -11246
rect 42612 -11300 42614 -11248
rect 42614 -11300 42666 -11248
rect 42666 -11300 42668 -11248
rect 42612 -11302 42668 -11300
rect 42932 -11248 42988 -11246
rect 42932 -11300 42934 -11248
rect 42934 -11300 42986 -11248
rect 42986 -11300 42988 -11248
rect 42932 -11302 42988 -11300
rect 43252 -11248 43308 -11246
rect 43252 -11300 43254 -11248
rect 43254 -11300 43306 -11248
rect 43306 -11300 43308 -11248
rect 43252 -11302 43308 -11300
rect 43572 -11248 43628 -11246
rect 43572 -11300 43574 -11248
rect 43574 -11300 43626 -11248
rect 43626 -11300 43628 -11248
rect 43572 -11302 43628 -11300
rect 43892 -11248 43948 -11246
rect 43892 -11300 43894 -11248
rect 43894 -11300 43946 -11248
rect 43946 -11300 43948 -11248
rect 43892 -11302 43948 -11300
rect 44212 -11248 44268 -11246
rect 44212 -11300 44214 -11248
rect 44214 -11300 44266 -11248
rect 44266 -11300 44268 -11248
rect 44212 -11302 44268 -11300
rect 44532 -11248 44588 -11246
rect 44532 -11300 44534 -11248
rect 44534 -11300 44586 -11248
rect 44586 -11300 44588 -11248
rect 44532 -11302 44588 -11300
rect 44852 -11248 44908 -11246
rect 44852 -11300 44854 -11248
rect 44854 -11300 44906 -11248
rect 44906 -11300 44908 -11248
rect 44852 -11302 44908 -11300
rect 45172 -11248 45228 -11246
rect 45172 -11300 45174 -11248
rect 45174 -11300 45226 -11248
rect 45226 -11300 45228 -11248
rect 45172 -11302 45228 -11300
rect 45492 -11248 45548 -11246
rect 45492 -11300 45494 -11248
rect 45494 -11300 45546 -11248
rect 45546 -11300 45548 -11248
rect 45492 -11302 45548 -11300
rect 45812 -11248 45868 -11246
rect 45812 -11300 45814 -11248
rect 45814 -11300 45866 -11248
rect 45866 -11300 45868 -11248
rect 45812 -11302 45868 -11300
rect 46132 -11248 46188 -11246
rect 46132 -11300 46134 -11248
rect 46134 -11300 46186 -11248
rect 46186 -11300 46188 -11248
rect 46132 -11302 46188 -11300
rect 46452 -11248 46508 -11246
rect 46452 -11300 46454 -11248
rect 46454 -11300 46506 -11248
rect 46506 -11300 46508 -11248
rect 46452 -11302 46508 -11300
rect 46772 -11248 46828 -11246
rect 46772 -11300 46774 -11248
rect 46774 -11300 46826 -11248
rect 46826 -11300 46828 -11248
rect 46772 -11302 46828 -11300
rect 47092 -11248 47148 -11246
rect 47092 -11300 47094 -11248
rect 47094 -11300 47146 -11248
rect 47146 -11300 47148 -11248
rect 47092 -11302 47148 -11300
rect 47412 -11248 47468 -11246
rect 47412 -11300 47414 -11248
rect 47414 -11300 47466 -11248
rect 47466 -11300 47468 -11248
rect 47412 -11302 47468 -11300
rect 47732 -11248 47788 -11246
rect 47732 -11300 47734 -11248
rect 47734 -11300 47786 -11248
rect 47786 -11300 47788 -11248
rect 47732 -11302 47788 -11300
rect 48052 -11248 48108 -11246
rect 48052 -11300 48054 -11248
rect 48054 -11300 48106 -11248
rect 48106 -11300 48108 -11248
rect 48052 -11302 48108 -11300
rect 48372 -11248 48428 -11246
rect 48372 -11300 48374 -11248
rect 48374 -11300 48426 -11248
rect 48426 -11300 48428 -11248
rect 48372 -11302 48428 -11300
rect 48692 -11248 48748 -11246
rect 48692 -11300 48694 -11248
rect 48694 -11300 48746 -11248
rect 48746 -11300 48748 -11248
rect 48692 -11302 48748 -11300
rect 49012 -11248 49068 -11246
rect 49012 -11300 49014 -11248
rect 49014 -11300 49066 -11248
rect 49066 -11300 49068 -11248
rect 49012 -11302 49068 -11300
rect 49332 -11248 49388 -11246
rect 49332 -11300 49334 -11248
rect 49334 -11300 49386 -11248
rect 49386 -11300 49388 -11248
rect 49332 -11302 49388 -11300
rect 42242 -11454 42298 -11452
rect 42242 -11506 42244 -11454
rect 42244 -11506 42296 -11454
rect 42296 -11506 42298 -11454
rect 42242 -11508 42298 -11506
rect 49708 -11454 49764 -11452
rect 49708 -11506 49710 -11454
rect 49710 -11506 49762 -11454
rect 49762 -11506 49764 -11454
rect 49708 -11508 49764 -11506
rect 42242 -11774 42298 -11772
rect 42242 -11826 42244 -11774
rect 42244 -11826 42296 -11774
rect 42296 -11826 42298 -11774
rect 42242 -11828 42298 -11826
rect 42242 -12094 42298 -12092
rect 42242 -12146 42244 -12094
rect 42244 -12146 42296 -12094
rect 42296 -12146 42298 -12094
rect 42242 -12148 42298 -12146
rect 42242 -12414 42298 -12412
rect 42242 -12466 42244 -12414
rect 42244 -12466 42296 -12414
rect 42296 -12466 42298 -12414
rect 42242 -12468 42298 -12466
rect 42242 -12734 42298 -12732
rect 42242 -12786 42244 -12734
rect 42244 -12786 42296 -12734
rect 42296 -12786 42298 -12734
rect 42242 -12788 42298 -12786
rect 42242 -13054 42298 -13052
rect 42242 -13106 42244 -13054
rect 42244 -13106 42296 -13054
rect 42296 -13106 42298 -13054
rect 42242 -13108 42298 -13106
rect 42242 -13374 42298 -13372
rect 42242 -13426 42244 -13374
rect 42244 -13426 42296 -13374
rect 42296 -13426 42298 -13374
rect 42242 -13428 42298 -13426
rect 42242 -13694 42298 -13692
rect 42242 -13746 42244 -13694
rect 42244 -13746 42296 -13694
rect 42296 -13746 42298 -13694
rect 42242 -13748 42298 -13746
rect 42242 -14014 42298 -14012
rect 42242 -14066 42244 -14014
rect 42244 -14066 42296 -14014
rect 42296 -14066 42298 -14014
rect 42242 -14068 42298 -14066
rect 42242 -14334 42298 -14332
rect 42242 -14386 42244 -14334
rect 42244 -14386 42296 -14334
rect 42296 -14386 42298 -14334
rect 42242 -14388 42298 -14386
rect 42242 -14654 42298 -14652
rect 42242 -14706 42244 -14654
rect 42244 -14706 42296 -14654
rect 42296 -14706 42298 -14654
rect 42242 -14708 42298 -14706
rect 42242 -14974 42298 -14972
rect 42242 -15026 42244 -14974
rect 42244 -15026 42296 -14974
rect 42296 -15026 42298 -14974
rect 42242 -15028 42298 -15026
rect 42242 -15294 42298 -15292
rect 42242 -15346 42244 -15294
rect 42244 -15346 42296 -15294
rect 42296 -15346 42298 -15294
rect 42242 -15348 42298 -15346
rect 42242 -15614 42298 -15612
rect 42242 -15666 42244 -15614
rect 42244 -15666 42296 -15614
rect 42296 -15666 42298 -15614
rect 42242 -15668 42298 -15666
rect 42242 -15934 42298 -15932
rect 42242 -15986 42244 -15934
rect 42244 -15986 42296 -15934
rect 42296 -15986 42298 -15934
rect 42242 -15988 42298 -15986
rect 42242 -16254 42298 -16252
rect 42242 -16306 42244 -16254
rect 42244 -16306 42296 -16254
rect 42296 -16306 42298 -16254
rect 42242 -16308 42298 -16306
rect 42242 -16574 42298 -16572
rect 42242 -16626 42244 -16574
rect 42244 -16626 42296 -16574
rect 42296 -16626 42298 -16574
rect 42242 -16628 42298 -16626
rect 42242 -16894 42298 -16892
rect 42242 -16946 42244 -16894
rect 42244 -16946 42296 -16894
rect 42296 -16946 42298 -16894
rect 42242 -16948 42298 -16946
rect 42242 -17214 42298 -17212
rect 42242 -17266 42244 -17214
rect 42244 -17266 42296 -17214
rect 42296 -17266 42298 -17214
rect 42242 -17268 42298 -17266
rect 42242 -17534 42298 -17532
rect 42242 -17586 42244 -17534
rect 42244 -17586 42296 -17534
rect 42296 -17586 42298 -17534
rect 42242 -17588 42298 -17586
rect 42242 -17854 42298 -17852
rect 42242 -17906 42244 -17854
rect 42244 -17906 42296 -17854
rect 42296 -17906 42298 -17854
rect 42242 -17908 42298 -17906
rect 42242 -18174 42298 -18172
rect 42242 -18226 42244 -18174
rect 42244 -18226 42296 -18174
rect 42296 -18226 42298 -18174
rect 42242 -18228 42298 -18226
rect 49708 -11774 49764 -11772
rect 49708 -11826 49710 -11774
rect 49710 -11826 49762 -11774
rect 49762 -11826 49764 -11774
rect 49708 -11828 49764 -11826
rect 49708 -12094 49764 -12092
rect 49708 -12146 49710 -12094
rect 49710 -12146 49762 -12094
rect 49762 -12146 49764 -12094
rect 49708 -12148 49764 -12146
rect 49708 -12414 49764 -12412
rect 49708 -12466 49710 -12414
rect 49710 -12466 49762 -12414
rect 49762 -12466 49764 -12414
rect 49708 -12468 49764 -12466
rect 49708 -12734 49764 -12732
rect 49708 -12786 49710 -12734
rect 49710 -12786 49762 -12734
rect 49762 -12786 49764 -12734
rect 49708 -12788 49764 -12786
rect 49708 -13054 49764 -13052
rect 49708 -13106 49710 -13054
rect 49710 -13106 49762 -13054
rect 49762 -13106 49764 -13054
rect 49708 -13108 49764 -13106
rect 49708 -13374 49764 -13372
rect 49708 -13426 49710 -13374
rect 49710 -13426 49762 -13374
rect 49762 -13426 49764 -13374
rect 49708 -13428 49764 -13426
rect 49708 -13694 49764 -13692
rect 49708 -13746 49710 -13694
rect 49710 -13746 49762 -13694
rect 49762 -13746 49764 -13694
rect 49708 -13748 49764 -13746
rect 49708 -14014 49764 -14012
rect 49708 -14066 49710 -14014
rect 49710 -14066 49762 -14014
rect 49762 -14066 49764 -14014
rect 49708 -14068 49764 -14066
rect 49708 -14334 49764 -14332
rect 49708 -14386 49710 -14334
rect 49710 -14386 49762 -14334
rect 49762 -14386 49764 -14334
rect 49708 -14388 49764 -14386
rect 49708 -14654 49764 -14652
rect 49708 -14706 49710 -14654
rect 49710 -14706 49762 -14654
rect 49762 -14706 49764 -14654
rect 49708 -14708 49764 -14706
rect 49708 -14974 49764 -14972
rect 49708 -15026 49710 -14974
rect 49710 -15026 49762 -14974
rect 49762 -15026 49764 -14974
rect 49708 -15028 49764 -15026
rect 49708 -15294 49764 -15292
rect 49708 -15346 49710 -15294
rect 49710 -15346 49762 -15294
rect 49762 -15346 49764 -15294
rect 49708 -15348 49764 -15346
rect 49708 -15614 49764 -15612
rect 49708 -15666 49710 -15614
rect 49710 -15666 49762 -15614
rect 49762 -15666 49764 -15614
rect 49708 -15668 49764 -15666
rect 49708 -15934 49764 -15932
rect 49708 -15986 49710 -15934
rect 49710 -15986 49762 -15934
rect 49762 -15986 49764 -15934
rect 49708 -15988 49764 -15986
rect 49708 -16254 49764 -16252
rect 49708 -16306 49710 -16254
rect 49710 -16306 49762 -16254
rect 49762 -16306 49764 -16254
rect 49708 -16308 49764 -16306
rect 49708 -16574 49764 -16572
rect 49708 -16626 49710 -16574
rect 49710 -16626 49762 -16574
rect 49762 -16626 49764 -16574
rect 49708 -16628 49764 -16626
rect 49708 -16894 49764 -16892
rect 49708 -16946 49710 -16894
rect 49710 -16946 49762 -16894
rect 49762 -16946 49764 -16894
rect 49708 -16948 49764 -16946
rect 49708 -17214 49764 -17212
rect 49708 -17266 49710 -17214
rect 49710 -17266 49762 -17214
rect 49762 -17266 49764 -17214
rect 49708 -17268 49764 -17266
rect 49708 -17534 49764 -17532
rect 49708 -17586 49710 -17534
rect 49710 -17586 49762 -17534
rect 49762 -17586 49764 -17534
rect 49708 -17588 49764 -17586
rect 49708 -17854 49764 -17852
rect 49708 -17906 49710 -17854
rect 49710 -17906 49762 -17854
rect 49762 -17906 49764 -17854
rect 49708 -17908 49764 -17906
rect 49708 -18174 49764 -18172
rect 49708 -18226 49710 -18174
rect 49710 -18226 49762 -18174
rect 49762 -18226 49764 -18174
rect 49708 -18228 49764 -18226
rect 42242 -18494 42298 -18492
rect 42242 -18546 42244 -18494
rect 42244 -18546 42296 -18494
rect 42296 -18546 42298 -18494
rect 42242 -18548 42298 -18546
rect 49708 -18494 49764 -18492
rect 49708 -18546 49710 -18494
rect 49710 -18546 49762 -18494
rect 49762 -18546 49764 -18494
rect 49708 -18548 49764 -18546
rect 42612 -18704 42668 -18702
rect 42612 -18756 42614 -18704
rect 42614 -18756 42666 -18704
rect 42666 -18756 42668 -18704
rect 42612 -18758 42668 -18756
rect 42932 -18704 42988 -18702
rect 42932 -18756 42934 -18704
rect 42934 -18756 42986 -18704
rect 42986 -18756 42988 -18704
rect 42932 -18758 42988 -18756
rect 43252 -18704 43308 -18702
rect 43252 -18756 43254 -18704
rect 43254 -18756 43306 -18704
rect 43306 -18756 43308 -18704
rect 43252 -18758 43308 -18756
rect 43572 -18704 43628 -18702
rect 43572 -18756 43574 -18704
rect 43574 -18756 43626 -18704
rect 43626 -18756 43628 -18704
rect 43572 -18758 43628 -18756
rect 43892 -18704 43948 -18702
rect 43892 -18756 43894 -18704
rect 43894 -18756 43946 -18704
rect 43946 -18756 43948 -18704
rect 43892 -18758 43948 -18756
rect 44212 -18704 44268 -18702
rect 44212 -18756 44214 -18704
rect 44214 -18756 44266 -18704
rect 44266 -18756 44268 -18704
rect 44212 -18758 44268 -18756
rect 44532 -18704 44588 -18702
rect 44532 -18756 44534 -18704
rect 44534 -18756 44586 -18704
rect 44586 -18756 44588 -18704
rect 44532 -18758 44588 -18756
rect 44852 -18704 44908 -18702
rect 44852 -18756 44854 -18704
rect 44854 -18756 44906 -18704
rect 44906 -18756 44908 -18704
rect 44852 -18758 44908 -18756
rect 45172 -18704 45228 -18702
rect 45172 -18756 45174 -18704
rect 45174 -18756 45226 -18704
rect 45226 -18756 45228 -18704
rect 45172 -18758 45228 -18756
rect 45492 -18704 45548 -18702
rect 45492 -18756 45494 -18704
rect 45494 -18756 45546 -18704
rect 45546 -18756 45548 -18704
rect 45492 -18758 45548 -18756
rect 45812 -18704 45868 -18702
rect 45812 -18756 45814 -18704
rect 45814 -18756 45866 -18704
rect 45866 -18756 45868 -18704
rect 45812 -18758 45868 -18756
rect 46132 -18704 46188 -18702
rect 46132 -18756 46134 -18704
rect 46134 -18756 46186 -18704
rect 46186 -18756 46188 -18704
rect 46132 -18758 46188 -18756
rect 46452 -18704 46508 -18702
rect 46452 -18756 46454 -18704
rect 46454 -18756 46506 -18704
rect 46506 -18756 46508 -18704
rect 46452 -18758 46508 -18756
rect 46772 -18704 46828 -18702
rect 46772 -18756 46774 -18704
rect 46774 -18756 46826 -18704
rect 46826 -18756 46828 -18704
rect 46772 -18758 46828 -18756
rect 47092 -18704 47148 -18702
rect 47092 -18756 47094 -18704
rect 47094 -18756 47146 -18704
rect 47146 -18756 47148 -18704
rect 47092 -18758 47148 -18756
rect 47412 -18704 47468 -18702
rect 47412 -18756 47414 -18704
rect 47414 -18756 47466 -18704
rect 47466 -18756 47468 -18704
rect 47412 -18758 47468 -18756
rect 47732 -18704 47788 -18702
rect 47732 -18756 47734 -18704
rect 47734 -18756 47786 -18704
rect 47786 -18756 47788 -18704
rect 47732 -18758 47788 -18756
rect 48052 -18704 48108 -18702
rect 48052 -18756 48054 -18704
rect 48054 -18756 48106 -18704
rect 48106 -18756 48108 -18704
rect 48052 -18758 48108 -18756
rect 48372 -18704 48428 -18702
rect 48372 -18756 48374 -18704
rect 48374 -18756 48426 -18704
rect 48426 -18756 48428 -18704
rect 48372 -18758 48428 -18756
rect 48692 -18704 48748 -18702
rect 48692 -18756 48694 -18704
rect 48694 -18756 48746 -18704
rect 48746 -18756 48748 -18704
rect 48692 -18758 48748 -18756
rect 49012 -18704 49068 -18702
rect 49012 -18756 49014 -18704
rect 49014 -18756 49066 -18704
rect 49066 -18756 49068 -18704
rect 49012 -18758 49068 -18756
rect 49332 -18704 49388 -18702
rect 49332 -18756 49334 -18704
rect 49334 -18756 49386 -18704
rect 49386 -18756 49388 -18704
rect 49332 -18758 49388 -18756
rect 6612 -23248 6668 -23246
rect 6612 -23300 6614 -23248
rect 6614 -23300 6666 -23248
rect 6666 -23300 6668 -23248
rect 6612 -23302 6668 -23300
rect 6932 -23248 6988 -23246
rect 6932 -23300 6934 -23248
rect 6934 -23300 6986 -23248
rect 6986 -23300 6988 -23248
rect 6932 -23302 6988 -23300
rect 7252 -23248 7308 -23246
rect 7252 -23300 7254 -23248
rect 7254 -23300 7306 -23248
rect 7306 -23300 7308 -23248
rect 7252 -23302 7308 -23300
rect 7572 -23248 7628 -23246
rect 7572 -23300 7574 -23248
rect 7574 -23300 7626 -23248
rect 7626 -23300 7628 -23248
rect 7572 -23302 7628 -23300
rect 7892 -23248 7948 -23246
rect 7892 -23300 7894 -23248
rect 7894 -23300 7946 -23248
rect 7946 -23300 7948 -23248
rect 7892 -23302 7948 -23300
rect 8212 -23248 8268 -23246
rect 8212 -23300 8214 -23248
rect 8214 -23300 8266 -23248
rect 8266 -23300 8268 -23248
rect 8212 -23302 8268 -23300
rect 8532 -23248 8588 -23246
rect 8532 -23300 8534 -23248
rect 8534 -23300 8586 -23248
rect 8586 -23300 8588 -23248
rect 8532 -23302 8588 -23300
rect 8852 -23248 8908 -23246
rect 8852 -23300 8854 -23248
rect 8854 -23300 8906 -23248
rect 8906 -23300 8908 -23248
rect 8852 -23302 8908 -23300
rect 9172 -23248 9228 -23246
rect 9172 -23300 9174 -23248
rect 9174 -23300 9226 -23248
rect 9226 -23300 9228 -23248
rect 9172 -23302 9228 -23300
rect 9492 -23248 9548 -23246
rect 9492 -23300 9494 -23248
rect 9494 -23300 9546 -23248
rect 9546 -23300 9548 -23248
rect 9492 -23302 9548 -23300
rect 9812 -23248 9868 -23246
rect 9812 -23300 9814 -23248
rect 9814 -23300 9866 -23248
rect 9866 -23300 9868 -23248
rect 9812 -23302 9868 -23300
rect 10132 -23248 10188 -23246
rect 10132 -23300 10134 -23248
rect 10134 -23300 10186 -23248
rect 10186 -23300 10188 -23248
rect 10132 -23302 10188 -23300
rect 10452 -23248 10508 -23246
rect 10452 -23300 10454 -23248
rect 10454 -23300 10506 -23248
rect 10506 -23300 10508 -23248
rect 10452 -23302 10508 -23300
rect 10772 -23248 10828 -23246
rect 10772 -23300 10774 -23248
rect 10774 -23300 10826 -23248
rect 10826 -23300 10828 -23248
rect 10772 -23302 10828 -23300
rect 11092 -23248 11148 -23246
rect 11092 -23300 11094 -23248
rect 11094 -23300 11146 -23248
rect 11146 -23300 11148 -23248
rect 11092 -23302 11148 -23300
rect 11412 -23248 11468 -23246
rect 11412 -23300 11414 -23248
rect 11414 -23300 11466 -23248
rect 11466 -23300 11468 -23248
rect 11412 -23302 11468 -23300
rect 11732 -23248 11788 -23246
rect 11732 -23300 11734 -23248
rect 11734 -23300 11786 -23248
rect 11786 -23300 11788 -23248
rect 11732 -23302 11788 -23300
rect 12052 -23248 12108 -23246
rect 12052 -23300 12054 -23248
rect 12054 -23300 12106 -23248
rect 12106 -23300 12108 -23248
rect 12052 -23302 12108 -23300
rect 12372 -23248 12428 -23246
rect 12372 -23300 12374 -23248
rect 12374 -23300 12426 -23248
rect 12426 -23300 12428 -23248
rect 12372 -23302 12428 -23300
rect 12692 -23248 12748 -23246
rect 12692 -23300 12694 -23248
rect 12694 -23300 12746 -23248
rect 12746 -23300 12748 -23248
rect 12692 -23302 12748 -23300
rect 13012 -23248 13068 -23246
rect 13012 -23300 13014 -23248
rect 13014 -23300 13066 -23248
rect 13066 -23300 13068 -23248
rect 13012 -23302 13068 -23300
rect 13332 -23248 13388 -23246
rect 13332 -23300 13334 -23248
rect 13334 -23300 13386 -23248
rect 13386 -23300 13388 -23248
rect 13332 -23302 13388 -23300
rect 6242 -23454 6298 -23452
rect 6242 -23506 6244 -23454
rect 6244 -23506 6296 -23454
rect 6296 -23506 6298 -23454
rect 6242 -23508 6298 -23506
rect 13708 -23454 13764 -23452
rect 13708 -23506 13710 -23454
rect 13710 -23506 13762 -23454
rect 13762 -23506 13764 -23454
rect 13708 -23508 13764 -23506
rect 6242 -23774 6298 -23772
rect 6242 -23826 6244 -23774
rect 6244 -23826 6296 -23774
rect 6296 -23826 6298 -23774
rect 6242 -23828 6298 -23826
rect 6242 -24094 6298 -24092
rect 6242 -24146 6244 -24094
rect 6244 -24146 6296 -24094
rect 6296 -24146 6298 -24094
rect 6242 -24148 6298 -24146
rect 6242 -24414 6298 -24412
rect 6242 -24466 6244 -24414
rect 6244 -24466 6296 -24414
rect 6296 -24466 6298 -24414
rect 6242 -24468 6298 -24466
rect 6242 -24734 6298 -24732
rect 6242 -24786 6244 -24734
rect 6244 -24786 6296 -24734
rect 6296 -24786 6298 -24734
rect 6242 -24788 6298 -24786
rect 6242 -25054 6298 -25052
rect 6242 -25106 6244 -25054
rect 6244 -25106 6296 -25054
rect 6296 -25106 6298 -25054
rect 6242 -25108 6298 -25106
rect 6242 -25374 6298 -25372
rect 6242 -25426 6244 -25374
rect 6244 -25426 6296 -25374
rect 6296 -25426 6298 -25374
rect 6242 -25428 6298 -25426
rect 6242 -25694 6298 -25692
rect 6242 -25746 6244 -25694
rect 6244 -25746 6296 -25694
rect 6296 -25746 6298 -25694
rect 6242 -25748 6298 -25746
rect 6242 -26014 6298 -26012
rect 6242 -26066 6244 -26014
rect 6244 -26066 6296 -26014
rect 6296 -26066 6298 -26014
rect 6242 -26068 6298 -26066
rect 6242 -26334 6298 -26332
rect 6242 -26386 6244 -26334
rect 6244 -26386 6296 -26334
rect 6296 -26386 6298 -26334
rect 6242 -26388 6298 -26386
rect 6242 -26654 6298 -26652
rect 6242 -26706 6244 -26654
rect 6244 -26706 6296 -26654
rect 6296 -26706 6298 -26654
rect 6242 -26708 6298 -26706
rect 6242 -26974 6298 -26972
rect 6242 -27026 6244 -26974
rect 6244 -27026 6296 -26974
rect 6296 -27026 6298 -26974
rect 6242 -27028 6298 -27026
rect 6242 -27294 6298 -27292
rect 6242 -27346 6244 -27294
rect 6244 -27346 6296 -27294
rect 6296 -27346 6298 -27294
rect 6242 -27348 6298 -27346
rect 6242 -27614 6298 -27612
rect 6242 -27666 6244 -27614
rect 6244 -27666 6296 -27614
rect 6296 -27666 6298 -27614
rect 6242 -27668 6298 -27666
rect 6242 -27934 6298 -27932
rect 6242 -27986 6244 -27934
rect 6244 -27986 6296 -27934
rect 6296 -27986 6298 -27934
rect 6242 -27988 6298 -27986
rect 6242 -28254 6298 -28252
rect 6242 -28306 6244 -28254
rect 6244 -28306 6296 -28254
rect 6296 -28306 6298 -28254
rect 6242 -28308 6298 -28306
rect 6242 -28574 6298 -28572
rect 6242 -28626 6244 -28574
rect 6244 -28626 6296 -28574
rect 6296 -28626 6298 -28574
rect 6242 -28628 6298 -28626
rect 6242 -28894 6298 -28892
rect 6242 -28946 6244 -28894
rect 6244 -28946 6296 -28894
rect 6296 -28946 6298 -28894
rect 6242 -28948 6298 -28946
rect 6242 -29214 6298 -29212
rect 6242 -29266 6244 -29214
rect 6244 -29266 6296 -29214
rect 6296 -29266 6298 -29214
rect 6242 -29268 6298 -29266
rect 6242 -29534 6298 -29532
rect 6242 -29586 6244 -29534
rect 6244 -29586 6296 -29534
rect 6296 -29586 6298 -29534
rect 6242 -29588 6298 -29586
rect 6242 -29854 6298 -29852
rect 6242 -29906 6244 -29854
rect 6244 -29906 6296 -29854
rect 6296 -29906 6298 -29854
rect 6242 -29908 6298 -29906
rect 6242 -30174 6298 -30172
rect 6242 -30226 6244 -30174
rect 6244 -30226 6296 -30174
rect 6296 -30226 6298 -30174
rect 6242 -30228 6298 -30226
rect 13708 -23774 13764 -23772
rect 13708 -23826 13710 -23774
rect 13710 -23826 13762 -23774
rect 13762 -23826 13764 -23774
rect 13708 -23828 13764 -23826
rect 13708 -24094 13764 -24092
rect 13708 -24146 13710 -24094
rect 13710 -24146 13762 -24094
rect 13762 -24146 13764 -24094
rect 13708 -24148 13764 -24146
rect 13708 -24414 13764 -24412
rect 13708 -24466 13710 -24414
rect 13710 -24466 13762 -24414
rect 13762 -24466 13764 -24414
rect 13708 -24468 13764 -24466
rect 13708 -24734 13764 -24732
rect 13708 -24786 13710 -24734
rect 13710 -24786 13762 -24734
rect 13762 -24786 13764 -24734
rect 13708 -24788 13764 -24786
rect 13708 -25054 13764 -25052
rect 13708 -25106 13710 -25054
rect 13710 -25106 13762 -25054
rect 13762 -25106 13764 -25054
rect 13708 -25108 13764 -25106
rect 13708 -25374 13764 -25372
rect 13708 -25426 13710 -25374
rect 13710 -25426 13762 -25374
rect 13762 -25426 13764 -25374
rect 13708 -25428 13764 -25426
rect 13708 -25694 13764 -25692
rect 13708 -25746 13710 -25694
rect 13710 -25746 13762 -25694
rect 13762 -25746 13764 -25694
rect 13708 -25748 13764 -25746
rect 13708 -26014 13764 -26012
rect 13708 -26066 13710 -26014
rect 13710 -26066 13762 -26014
rect 13762 -26066 13764 -26014
rect 13708 -26068 13764 -26066
rect 13708 -26334 13764 -26332
rect 13708 -26386 13710 -26334
rect 13710 -26386 13762 -26334
rect 13762 -26386 13764 -26334
rect 13708 -26388 13764 -26386
rect 13708 -26654 13764 -26652
rect 13708 -26706 13710 -26654
rect 13710 -26706 13762 -26654
rect 13762 -26706 13764 -26654
rect 13708 -26708 13764 -26706
rect 13708 -26974 13764 -26972
rect 13708 -27026 13710 -26974
rect 13710 -27026 13762 -26974
rect 13762 -27026 13764 -26974
rect 13708 -27028 13764 -27026
rect 13708 -27294 13764 -27292
rect 13708 -27346 13710 -27294
rect 13710 -27346 13762 -27294
rect 13762 -27346 13764 -27294
rect 13708 -27348 13764 -27346
rect 13708 -27614 13764 -27612
rect 13708 -27666 13710 -27614
rect 13710 -27666 13762 -27614
rect 13762 -27666 13764 -27614
rect 13708 -27668 13764 -27666
rect 13708 -27934 13764 -27932
rect 13708 -27986 13710 -27934
rect 13710 -27986 13762 -27934
rect 13762 -27986 13764 -27934
rect 13708 -27988 13764 -27986
rect 13708 -28254 13764 -28252
rect 13708 -28306 13710 -28254
rect 13710 -28306 13762 -28254
rect 13762 -28306 13764 -28254
rect 13708 -28308 13764 -28306
rect 13708 -28574 13764 -28572
rect 13708 -28626 13710 -28574
rect 13710 -28626 13762 -28574
rect 13762 -28626 13764 -28574
rect 13708 -28628 13764 -28626
rect 13708 -28894 13764 -28892
rect 13708 -28946 13710 -28894
rect 13710 -28946 13762 -28894
rect 13762 -28946 13764 -28894
rect 13708 -28948 13764 -28946
rect 13708 -29214 13764 -29212
rect 13708 -29266 13710 -29214
rect 13710 -29266 13762 -29214
rect 13762 -29266 13764 -29214
rect 13708 -29268 13764 -29266
rect 13708 -29534 13764 -29532
rect 13708 -29586 13710 -29534
rect 13710 -29586 13762 -29534
rect 13762 -29586 13764 -29534
rect 13708 -29588 13764 -29586
rect 13708 -29854 13764 -29852
rect 13708 -29906 13710 -29854
rect 13710 -29906 13762 -29854
rect 13762 -29906 13764 -29854
rect 13708 -29908 13764 -29906
rect 13708 -30174 13764 -30172
rect 13708 -30226 13710 -30174
rect 13710 -30226 13762 -30174
rect 13762 -30226 13764 -30174
rect 13708 -30228 13764 -30226
rect 6242 -30494 6298 -30492
rect 6242 -30546 6244 -30494
rect 6244 -30546 6296 -30494
rect 6296 -30546 6298 -30494
rect 6242 -30548 6298 -30546
rect 13708 -30494 13764 -30492
rect 13708 -30546 13710 -30494
rect 13710 -30546 13762 -30494
rect 13762 -30546 13764 -30494
rect 13708 -30548 13764 -30546
rect 6612 -30704 6668 -30702
rect 6612 -30756 6614 -30704
rect 6614 -30756 6666 -30704
rect 6666 -30756 6668 -30704
rect 6612 -30758 6668 -30756
rect 6932 -30704 6988 -30702
rect 6932 -30756 6934 -30704
rect 6934 -30756 6986 -30704
rect 6986 -30756 6988 -30704
rect 6932 -30758 6988 -30756
rect 7252 -30704 7308 -30702
rect 7252 -30756 7254 -30704
rect 7254 -30756 7306 -30704
rect 7306 -30756 7308 -30704
rect 7252 -30758 7308 -30756
rect 7572 -30704 7628 -30702
rect 7572 -30756 7574 -30704
rect 7574 -30756 7626 -30704
rect 7626 -30756 7628 -30704
rect 7572 -30758 7628 -30756
rect 7892 -30704 7948 -30702
rect 7892 -30756 7894 -30704
rect 7894 -30756 7946 -30704
rect 7946 -30756 7948 -30704
rect 7892 -30758 7948 -30756
rect 8212 -30704 8268 -30702
rect 8212 -30756 8214 -30704
rect 8214 -30756 8266 -30704
rect 8266 -30756 8268 -30704
rect 8212 -30758 8268 -30756
rect 8532 -30704 8588 -30702
rect 8532 -30756 8534 -30704
rect 8534 -30756 8586 -30704
rect 8586 -30756 8588 -30704
rect 8532 -30758 8588 -30756
rect 8852 -30704 8908 -30702
rect 8852 -30756 8854 -30704
rect 8854 -30756 8906 -30704
rect 8906 -30756 8908 -30704
rect 8852 -30758 8908 -30756
rect 9172 -30704 9228 -30702
rect 9172 -30756 9174 -30704
rect 9174 -30756 9226 -30704
rect 9226 -30756 9228 -30704
rect 9172 -30758 9228 -30756
rect 9492 -30704 9548 -30702
rect 9492 -30756 9494 -30704
rect 9494 -30756 9546 -30704
rect 9546 -30756 9548 -30704
rect 9492 -30758 9548 -30756
rect 9812 -30704 9868 -30702
rect 9812 -30756 9814 -30704
rect 9814 -30756 9866 -30704
rect 9866 -30756 9868 -30704
rect 9812 -30758 9868 -30756
rect 10132 -30704 10188 -30702
rect 10132 -30756 10134 -30704
rect 10134 -30756 10186 -30704
rect 10186 -30756 10188 -30704
rect 10132 -30758 10188 -30756
rect 10452 -30704 10508 -30702
rect 10452 -30756 10454 -30704
rect 10454 -30756 10506 -30704
rect 10506 -30756 10508 -30704
rect 10452 -30758 10508 -30756
rect 10772 -30704 10828 -30702
rect 10772 -30756 10774 -30704
rect 10774 -30756 10826 -30704
rect 10826 -30756 10828 -30704
rect 10772 -30758 10828 -30756
rect 11092 -30704 11148 -30702
rect 11092 -30756 11094 -30704
rect 11094 -30756 11146 -30704
rect 11146 -30756 11148 -30704
rect 11092 -30758 11148 -30756
rect 11412 -30704 11468 -30702
rect 11412 -30756 11414 -30704
rect 11414 -30756 11466 -30704
rect 11466 -30756 11468 -30704
rect 11412 -30758 11468 -30756
rect 11732 -30704 11788 -30702
rect 11732 -30756 11734 -30704
rect 11734 -30756 11786 -30704
rect 11786 -30756 11788 -30704
rect 11732 -30758 11788 -30756
rect 12052 -30704 12108 -30702
rect 12052 -30756 12054 -30704
rect 12054 -30756 12106 -30704
rect 12106 -30756 12108 -30704
rect 12052 -30758 12108 -30756
rect 12372 -30704 12428 -30702
rect 12372 -30756 12374 -30704
rect 12374 -30756 12426 -30704
rect 12426 -30756 12428 -30704
rect 12372 -30758 12428 -30756
rect 12692 -30704 12748 -30702
rect 12692 -30756 12694 -30704
rect 12694 -30756 12746 -30704
rect 12746 -30756 12748 -30704
rect 12692 -30758 12748 -30756
rect 13012 -30704 13068 -30702
rect 13012 -30756 13014 -30704
rect 13014 -30756 13066 -30704
rect 13066 -30756 13068 -30704
rect 13012 -30758 13068 -30756
rect 13332 -30704 13388 -30702
rect 13332 -30756 13334 -30704
rect 13334 -30756 13386 -30704
rect 13386 -30756 13388 -30704
rect 13332 -30758 13388 -30756
rect 18612 -23248 18668 -23246
rect 18612 -23300 18614 -23248
rect 18614 -23300 18666 -23248
rect 18666 -23300 18668 -23248
rect 18612 -23302 18668 -23300
rect 18932 -23248 18988 -23246
rect 18932 -23300 18934 -23248
rect 18934 -23300 18986 -23248
rect 18986 -23300 18988 -23248
rect 18932 -23302 18988 -23300
rect 19252 -23248 19308 -23246
rect 19252 -23300 19254 -23248
rect 19254 -23300 19306 -23248
rect 19306 -23300 19308 -23248
rect 19252 -23302 19308 -23300
rect 19572 -23248 19628 -23246
rect 19572 -23300 19574 -23248
rect 19574 -23300 19626 -23248
rect 19626 -23300 19628 -23248
rect 19572 -23302 19628 -23300
rect 19892 -23248 19948 -23246
rect 19892 -23300 19894 -23248
rect 19894 -23300 19946 -23248
rect 19946 -23300 19948 -23248
rect 19892 -23302 19948 -23300
rect 20212 -23248 20268 -23246
rect 20212 -23300 20214 -23248
rect 20214 -23300 20266 -23248
rect 20266 -23300 20268 -23248
rect 20212 -23302 20268 -23300
rect 20532 -23248 20588 -23246
rect 20532 -23300 20534 -23248
rect 20534 -23300 20586 -23248
rect 20586 -23300 20588 -23248
rect 20532 -23302 20588 -23300
rect 20852 -23248 20908 -23246
rect 20852 -23300 20854 -23248
rect 20854 -23300 20906 -23248
rect 20906 -23300 20908 -23248
rect 20852 -23302 20908 -23300
rect 21172 -23248 21228 -23246
rect 21172 -23300 21174 -23248
rect 21174 -23300 21226 -23248
rect 21226 -23300 21228 -23248
rect 21172 -23302 21228 -23300
rect 21492 -23248 21548 -23246
rect 21492 -23300 21494 -23248
rect 21494 -23300 21546 -23248
rect 21546 -23300 21548 -23248
rect 21492 -23302 21548 -23300
rect 21812 -23248 21868 -23246
rect 21812 -23300 21814 -23248
rect 21814 -23300 21866 -23248
rect 21866 -23300 21868 -23248
rect 21812 -23302 21868 -23300
rect 22132 -23248 22188 -23246
rect 22132 -23300 22134 -23248
rect 22134 -23300 22186 -23248
rect 22186 -23300 22188 -23248
rect 22132 -23302 22188 -23300
rect 22452 -23248 22508 -23246
rect 22452 -23300 22454 -23248
rect 22454 -23300 22506 -23248
rect 22506 -23300 22508 -23248
rect 22452 -23302 22508 -23300
rect 22772 -23248 22828 -23246
rect 22772 -23300 22774 -23248
rect 22774 -23300 22826 -23248
rect 22826 -23300 22828 -23248
rect 22772 -23302 22828 -23300
rect 23092 -23248 23148 -23246
rect 23092 -23300 23094 -23248
rect 23094 -23300 23146 -23248
rect 23146 -23300 23148 -23248
rect 23092 -23302 23148 -23300
rect 23412 -23248 23468 -23246
rect 23412 -23300 23414 -23248
rect 23414 -23300 23466 -23248
rect 23466 -23300 23468 -23248
rect 23412 -23302 23468 -23300
rect 23732 -23248 23788 -23246
rect 23732 -23300 23734 -23248
rect 23734 -23300 23786 -23248
rect 23786 -23300 23788 -23248
rect 23732 -23302 23788 -23300
rect 24052 -23248 24108 -23246
rect 24052 -23300 24054 -23248
rect 24054 -23300 24106 -23248
rect 24106 -23300 24108 -23248
rect 24052 -23302 24108 -23300
rect 24372 -23248 24428 -23246
rect 24372 -23300 24374 -23248
rect 24374 -23300 24426 -23248
rect 24426 -23300 24428 -23248
rect 24372 -23302 24428 -23300
rect 24692 -23248 24748 -23246
rect 24692 -23300 24694 -23248
rect 24694 -23300 24746 -23248
rect 24746 -23300 24748 -23248
rect 24692 -23302 24748 -23300
rect 25012 -23248 25068 -23246
rect 25012 -23300 25014 -23248
rect 25014 -23300 25066 -23248
rect 25066 -23300 25068 -23248
rect 25012 -23302 25068 -23300
rect 25332 -23248 25388 -23246
rect 25332 -23300 25334 -23248
rect 25334 -23300 25386 -23248
rect 25386 -23300 25388 -23248
rect 25332 -23302 25388 -23300
rect 18242 -23454 18298 -23452
rect 18242 -23506 18244 -23454
rect 18244 -23506 18296 -23454
rect 18296 -23506 18298 -23454
rect 18242 -23508 18298 -23506
rect 25708 -23454 25764 -23452
rect 25708 -23506 25710 -23454
rect 25710 -23506 25762 -23454
rect 25762 -23506 25764 -23454
rect 25708 -23508 25764 -23506
rect 18242 -23774 18298 -23772
rect 18242 -23826 18244 -23774
rect 18244 -23826 18296 -23774
rect 18296 -23826 18298 -23774
rect 18242 -23828 18298 -23826
rect 18242 -24094 18298 -24092
rect 18242 -24146 18244 -24094
rect 18244 -24146 18296 -24094
rect 18296 -24146 18298 -24094
rect 18242 -24148 18298 -24146
rect 18242 -24414 18298 -24412
rect 18242 -24466 18244 -24414
rect 18244 -24466 18296 -24414
rect 18296 -24466 18298 -24414
rect 18242 -24468 18298 -24466
rect 18242 -24734 18298 -24732
rect 18242 -24786 18244 -24734
rect 18244 -24786 18296 -24734
rect 18296 -24786 18298 -24734
rect 18242 -24788 18298 -24786
rect 18242 -25054 18298 -25052
rect 18242 -25106 18244 -25054
rect 18244 -25106 18296 -25054
rect 18296 -25106 18298 -25054
rect 18242 -25108 18298 -25106
rect 18242 -25374 18298 -25372
rect 18242 -25426 18244 -25374
rect 18244 -25426 18296 -25374
rect 18296 -25426 18298 -25374
rect 18242 -25428 18298 -25426
rect 18242 -25694 18298 -25692
rect 18242 -25746 18244 -25694
rect 18244 -25746 18296 -25694
rect 18296 -25746 18298 -25694
rect 18242 -25748 18298 -25746
rect 18242 -26014 18298 -26012
rect 18242 -26066 18244 -26014
rect 18244 -26066 18296 -26014
rect 18296 -26066 18298 -26014
rect 18242 -26068 18298 -26066
rect 18242 -26334 18298 -26332
rect 18242 -26386 18244 -26334
rect 18244 -26386 18296 -26334
rect 18296 -26386 18298 -26334
rect 18242 -26388 18298 -26386
rect 18242 -26654 18298 -26652
rect 18242 -26706 18244 -26654
rect 18244 -26706 18296 -26654
rect 18296 -26706 18298 -26654
rect 18242 -26708 18298 -26706
rect 18242 -26974 18298 -26972
rect 18242 -27026 18244 -26974
rect 18244 -27026 18296 -26974
rect 18296 -27026 18298 -26974
rect 18242 -27028 18298 -27026
rect 18242 -27294 18298 -27292
rect 18242 -27346 18244 -27294
rect 18244 -27346 18296 -27294
rect 18296 -27346 18298 -27294
rect 18242 -27348 18298 -27346
rect 18242 -27614 18298 -27612
rect 18242 -27666 18244 -27614
rect 18244 -27666 18296 -27614
rect 18296 -27666 18298 -27614
rect 18242 -27668 18298 -27666
rect 18242 -27934 18298 -27932
rect 18242 -27986 18244 -27934
rect 18244 -27986 18296 -27934
rect 18296 -27986 18298 -27934
rect 18242 -27988 18298 -27986
rect 18242 -28254 18298 -28252
rect 18242 -28306 18244 -28254
rect 18244 -28306 18296 -28254
rect 18296 -28306 18298 -28254
rect 18242 -28308 18298 -28306
rect 18242 -28574 18298 -28572
rect 18242 -28626 18244 -28574
rect 18244 -28626 18296 -28574
rect 18296 -28626 18298 -28574
rect 18242 -28628 18298 -28626
rect 18242 -28894 18298 -28892
rect 18242 -28946 18244 -28894
rect 18244 -28946 18296 -28894
rect 18296 -28946 18298 -28894
rect 18242 -28948 18298 -28946
rect 18242 -29214 18298 -29212
rect 18242 -29266 18244 -29214
rect 18244 -29266 18296 -29214
rect 18296 -29266 18298 -29214
rect 18242 -29268 18298 -29266
rect 18242 -29534 18298 -29532
rect 18242 -29586 18244 -29534
rect 18244 -29586 18296 -29534
rect 18296 -29586 18298 -29534
rect 18242 -29588 18298 -29586
rect 18242 -29854 18298 -29852
rect 18242 -29906 18244 -29854
rect 18244 -29906 18296 -29854
rect 18296 -29906 18298 -29854
rect 18242 -29908 18298 -29906
rect 18242 -30174 18298 -30172
rect 18242 -30226 18244 -30174
rect 18244 -30226 18296 -30174
rect 18296 -30226 18298 -30174
rect 18242 -30228 18298 -30226
rect 25708 -23774 25764 -23772
rect 25708 -23826 25710 -23774
rect 25710 -23826 25762 -23774
rect 25762 -23826 25764 -23774
rect 25708 -23828 25764 -23826
rect 25708 -24094 25764 -24092
rect 25708 -24146 25710 -24094
rect 25710 -24146 25762 -24094
rect 25762 -24146 25764 -24094
rect 25708 -24148 25764 -24146
rect 25708 -24414 25764 -24412
rect 25708 -24466 25710 -24414
rect 25710 -24466 25762 -24414
rect 25762 -24466 25764 -24414
rect 25708 -24468 25764 -24466
rect 25708 -24734 25764 -24732
rect 25708 -24786 25710 -24734
rect 25710 -24786 25762 -24734
rect 25762 -24786 25764 -24734
rect 25708 -24788 25764 -24786
rect 25708 -25054 25764 -25052
rect 25708 -25106 25710 -25054
rect 25710 -25106 25762 -25054
rect 25762 -25106 25764 -25054
rect 25708 -25108 25764 -25106
rect 25708 -25374 25764 -25372
rect 25708 -25426 25710 -25374
rect 25710 -25426 25762 -25374
rect 25762 -25426 25764 -25374
rect 25708 -25428 25764 -25426
rect 25708 -25694 25764 -25692
rect 25708 -25746 25710 -25694
rect 25710 -25746 25762 -25694
rect 25762 -25746 25764 -25694
rect 25708 -25748 25764 -25746
rect 25708 -26014 25764 -26012
rect 25708 -26066 25710 -26014
rect 25710 -26066 25762 -26014
rect 25762 -26066 25764 -26014
rect 25708 -26068 25764 -26066
rect 25708 -26334 25764 -26332
rect 25708 -26386 25710 -26334
rect 25710 -26386 25762 -26334
rect 25762 -26386 25764 -26334
rect 25708 -26388 25764 -26386
rect 25708 -26654 25764 -26652
rect 25708 -26706 25710 -26654
rect 25710 -26706 25762 -26654
rect 25762 -26706 25764 -26654
rect 25708 -26708 25764 -26706
rect 25708 -26974 25764 -26972
rect 25708 -27026 25710 -26974
rect 25710 -27026 25762 -26974
rect 25762 -27026 25764 -26974
rect 25708 -27028 25764 -27026
rect 25708 -27294 25764 -27292
rect 25708 -27346 25710 -27294
rect 25710 -27346 25762 -27294
rect 25762 -27346 25764 -27294
rect 25708 -27348 25764 -27346
rect 25708 -27614 25764 -27612
rect 25708 -27666 25710 -27614
rect 25710 -27666 25762 -27614
rect 25762 -27666 25764 -27614
rect 25708 -27668 25764 -27666
rect 25708 -27934 25764 -27932
rect 25708 -27986 25710 -27934
rect 25710 -27986 25762 -27934
rect 25762 -27986 25764 -27934
rect 25708 -27988 25764 -27986
rect 25708 -28254 25764 -28252
rect 25708 -28306 25710 -28254
rect 25710 -28306 25762 -28254
rect 25762 -28306 25764 -28254
rect 25708 -28308 25764 -28306
rect 25708 -28574 25764 -28572
rect 25708 -28626 25710 -28574
rect 25710 -28626 25762 -28574
rect 25762 -28626 25764 -28574
rect 25708 -28628 25764 -28626
rect 25708 -28894 25764 -28892
rect 25708 -28946 25710 -28894
rect 25710 -28946 25762 -28894
rect 25762 -28946 25764 -28894
rect 25708 -28948 25764 -28946
rect 25708 -29214 25764 -29212
rect 25708 -29266 25710 -29214
rect 25710 -29266 25762 -29214
rect 25762 -29266 25764 -29214
rect 25708 -29268 25764 -29266
rect 25708 -29534 25764 -29532
rect 25708 -29586 25710 -29534
rect 25710 -29586 25762 -29534
rect 25762 -29586 25764 -29534
rect 25708 -29588 25764 -29586
rect 25708 -29854 25764 -29852
rect 25708 -29906 25710 -29854
rect 25710 -29906 25762 -29854
rect 25762 -29906 25764 -29854
rect 25708 -29908 25764 -29906
rect 25708 -30174 25764 -30172
rect 25708 -30226 25710 -30174
rect 25710 -30226 25762 -30174
rect 25762 -30226 25764 -30174
rect 25708 -30228 25764 -30226
rect 18242 -30494 18298 -30492
rect 18242 -30546 18244 -30494
rect 18244 -30546 18296 -30494
rect 18296 -30546 18298 -30494
rect 18242 -30548 18298 -30546
rect 25708 -30494 25764 -30492
rect 25708 -30546 25710 -30494
rect 25710 -30546 25762 -30494
rect 25762 -30546 25764 -30494
rect 25708 -30548 25764 -30546
rect 18612 -30704 18668 -30702
rect 18612 -30756 18614 -30704
rect 18614 -30756 18666 -30704
rect 18666 -30756 18668 -30704
rect 18612 -30758 18668 -30756
rect 18932 -30704 18988 -30702
rect 18932 -30756 18934 -30704
rect 18934 -30756 18986 -30704
rect 18986 -30756 18988 -30704
rect 18932 -30758 18988 -30756
rect 19252 -30704 19308 -30702
rect 19252 -30756 19254 -30704
rect 19254 -30756 19306 -30704
rect 19306 -30756 19308 -30704
rect 19252 -30758 19308 -30756
rect 19572 -30704 19628 -30702
rect 19572 -30756 19574 -30704
rect 19574 -30756 19626 -30704
rect 19626 -30756 19628 -30704
rect 19572 -30758 19628 -30756
rect 19892 -30704 19948 -30702
rect 19892 -30756 19894 -30704
rect 19894 -30756 19946 -30704
rect 19946 -30756 19948 -30704
rect 19892 -30758 19948 -30756
rect 20212 -30704 20268 -30702
rect 20212 -30756 20214 -30704
rect 20214 -30756 20266 -30704
rect 20266 -30756 20268 -30704
rect 20212 -30758 20268 -30756
rect 20532 -30704 20588 -30702
rect 20532 -30756 20534 -30704
rect 20534 -30756 20586 -30704
rect 20586 -30756 20588 -30704
rect 20532 -30758 20588 -30756
rect 20852 -30704 20908 -30702
rect 20852 -30756 20854 -30704
rect 20854 -30756 20906 -30704
rect 20906 -30756 20908 -30704
rect 20852 -30758 20908 -30756
rect 21172 -30704 21228 -30702
rect 21172 -30756 21174 -30704
rect 21174 -30756 21226 -30704
rect 21226 -30756 21228 -30704
rect 21172 -30758 21228 -30756
rect 21492 -30704 21548 -30702
rect 21492 -30756 21494 -30704
rect 21494 -30756 21546 -30704
rect 21546 -30756 21548 -30704
rect 21492 -30758 21548 -30756
rect 21812 -30704 21868 -30702
rect 21812 -30756 21814 -30704
rect 21814 -30756 21866 -30704
rect 21866 -30756 21868 -30704
rect 21812 -30758 21868 -30756
rect 22132 -30704 22188 -30702
rect 22132 -30756 22134 -30704
rect 22134 -30756 22186 -30704
rect 22186 -30756 22188 -30704
rect 22132 -30758 22188 -30756
rect 22452 -30704 22508 -30702
rect 22452 -30756 22454 -30704
rect 22454 -30756 22506 -30704
rect 22506 -30756 22508 -30704
rect 22452 -30758 22508 -30756
rect 22772 -30704 22828 -30702
rect 22772 -30756 22774 -30704
rect 22774 -30756 22826 -30704
rect 22826 -30756 22828 -30704
rect 22772 -30758 22828 -30756
rect 23092 -30704 23148 -30702
rect 23092 -30756 23094 -30704
rect 23094 -30756 23146 -30704
rect 23146 -30756 23148 -30704
rect 23092 -30758 23148 -30756
rect 23412 -30704 23468 -30702
rect 23412 -30756 23414 -30704
rect 23414 -30756 23466 -30704
rect 23466 -30756 23468 -30704
rect 23412 -30758 23468 -30756
rect 23732 -30704 23788 -30702
rect 23732 -30756 23734 -30704
rect 23734 -30756 23786 -30704
rect 23786 -30756 23788 -30704
rect 23732 -30758 23788 -30756
rect 24052 -30704 24108 -30702
rect 24052 -30756 24054 -30704
rect 24054 -30756 24106 -30704
rect 24106 -30756 24108 -30704
rect 24052 -30758 24108 -30756
rect 24372 -30704 24428 -30702
rect 24372 -30756 24374 -30704
rect 24374 -30756 24426 -30704
rect 24426 -30756 24428 -30704
rect 24372 -30758 24428 -30756
rect 24692 -30704 24748 -30702
rect 24692 -30756 24694 -30704
rect 24694 -30756 24746 -30704
rect 24746 -30756 24748 -30704
rect 24692 -30758 24748 -30756
rect 25012 -30704 25068 -30702
rect 25012 -30756 25014 -30704
rect 25014 -30756 25066 -30704
rect 25066 -30756 25068 -30704
rect 25012 -30758 25068 -30756
rect 25332 -30704 25388 -30702
rect 25332 -30756 25334 -30704
rect 25334 -30756 25386 -30704
rect 25386 -30756 25388 -30704
rect 25332 -30758 25388 -30756
rect 30612 -23248 30668 -23246
rect 30612 -23300 30614 -23248
rect 30614 -23300 30666 -23248
rect 30666 -23300 30668 -23248
rect 30612 -23302 30668 -23300
rect 30932 -23248 30988 -23246
rect 30932 -23300 30934 -23248
rect 30934 -23300 30986 -23248
rect 30986 -23300 30988 -23248
rect 30932 -23302 30988 -23300
rect 31252 -23248 31308 -23246
rect 31252 -23300 31254 -23248
rect 31254 -23300 31306 -23248
rect 31306 -23300 31308 -23248
rect 31252 -23302 31308 -23300
rect 31572 -23248 31628 -23246
rect 31572 -23300 31574 -23248
rect 31574 -23300 31626 -23248
rect 31626 -23300 31628 -23248
rect 31572 -23302 31628 -23300
rect 31892 -23248 31948 -23246
rect 31892 -23300 31894 -23248
rect 31894 -23300 31946 -23248
rect 31946 -23300 31948 -23248
rect 31892 -23302 31948 -23300
rect 32212 -23248 32268 -23246
rect 32212 -23300 32214 -23248
rect 32214 -23300 32266 -23248
rect 32266 -23300 32268 -23248
rect 32212 -23302 32268 -23300
rect 32532 -23248 32588 -23246
rect 32532 -23300 32534 -23248
rect 32534 -23300 32586 -23248
rect 32586 -23300 32588 -23248
rect 32532 -23302 32588 -23300
rect 32852 -23248 32908 -23246
rect 32852 -23300 32854 -23248
rect 32854 -23300 32906 -23248
rect 32906 -23300 32908 -23248
rect 32852 -23302 32908 -23300
rect 33172 -23248 33228 -23246
rect 33172 -23300 33174 -23248
rect 33174 -23300 33226 -23248
rect 33226 -23300 33228 -23248
rect 33172 -23302 33228 -23300
rect 33492 -23248 33548 -23246
rect 33492 -23300 33494 -23248
rect 33494 -23300 33546 -23248
rect 33546 -23300 33548 -23248
rect 33492 -23302 33548 -23300
rect 33812 -23248 33868 -23246
rect 33812 -23300 33814 -23248
rect 33814 -23300 33866 -23248
rect 33866 -23300 33868 -23248
rect 33812 -23302 33868 -23300
rect 34132 -23248 34188 -23246
rect 34132 -23300 34134 -23248
rect 34134 -23300 34186 -23248
rect 34186 -23300 34188 -23248
rect 34132 -23302 34188 -23300
rect 34452 -23248 34508 -23246
rect 34452 -23300 34454 -23248
rect 34454 -23300 34506 -23248
rect 34506 -23300 34508 -23248
rect 34452 -23302 34508 -23300
rect 34772 -23248 34828 -23246
rect 34772 -23300 34774 -23248
rect 34774 -23300 34826 -23248
rect 34826 -23300 34828 -23248
rect 34772 -23302 34828 -23300
rect 35092 -23248 35148 -23246
rect 35092 -23300 35094 -23248
rect 35094 -23300 35146 -23248
rect 35146 -23300 35148 -23248
rect 35092 -23302 35148 -23300
rect 35412 -23248 35468 -23246
rect 35412 -23300 35414 -23248
rect 35414 -23300 35466 -23248
rect 35466 -23300 35468 -23248
rect 35412 -23302 35468 -23300
rect 35732 -23248 35788 -23246
rect 35732 -23300 35734 -23248
rect 35734 -23300 35786 -23248
rect 35786 -23300 35788 -23248
rect 35732 -23302 35788 -23300
rect 36052 -23248 36108 -23246
rect 36052 -23300 36054 -23248
rect 36054 -23300 36106 -23248
rect 36106 -23300 36108 -23248
rect 36052 -23302 36108 -23300
rect 36372 -23248 36428 -23246
rect 36372 -23300 36374 -23248
rect 36374 -23300 36426 -23248
rect 36426 -23300 36428 -23248
rect 36372 -23302 36428 -23300
rect 36692 -23248 36748 -23246
rect 36692 -23300 36694 -23248
rect 36694 -23300 36746 -23248
rect 36746 -23300 36748 -23248
rect 36692 -23302 36748 -23300
rect 37012 -23248 37068 -23246
rect 37012 -23300 37014 -23248
rect 37014 -23300 37066 -23248
rect 37066 -23300 37068 -23248
rect 37012 -23302 37068 -23300
rect 37332 -23248 37388 -23246
rect 37332 -23300 37334 -23248
rect 37334 -23300 37386 -23248
rect 37386 -23300 37388 -23248
rect 37332 -23302 37388 -23300
rect 30242 -23454 30298 -23452
rect 30242 -23506 30244 -23454
rect 30244 -23506 30296 -23454
rect 30296 -23506 30298 -23454
rect 30242 -23508 30298 -23506
rect 37708 -23454 37764 -23452
rect 37708 -23506 37710 -23454
rect 37710 -23506 37762 -23454
rect 37762 -23506 37764 -23454
rect 37708 -23508 37764 -23506
rect 30242 -23774 30298 -23772
rect 30242 -23826 30244 -23774
rect 30244 -23826 30296 -23774
rect 30296 -23826 30298 -23774
rect 30242 -23828 30298 -23826
rect 30242 -24094 30298 -24092
rect 30242 -24146 30244 -24094
rect 30244 -24146 30296 -24094
rect 30296 -24146 30298 -24094
rect 30242 -24148 30298 -24146
rect 30242 -24414 30298 -24412
rect 30242 -24466 30244 -24414
rect 30244 -24466 30296 -24414
rect 30296 -24466 30298 -24414
rect 30242 -24468 30298 -24466
rect 30242 -24734 30298 -24732
rect 30242 -24786 30244 -24734
rect 30244 -24786 30296 -24734
rect 30296 -24786 30298 -24734
rect 30242 -24788 30298 -24786
rect 30242 -25054 30298 -25052
rect 30242 -25106 30244 -25054
rect 30244 -25106 30296 -25054
rect 30296 -25106 30298 -25054
rect 30242 -25108 30298 -25106
rect 30242 -25374 30298 -25372
rect 30242 -25426 30244 -25374
rect 30244 -25426 30296 -25374
rect 30296 -25426 30298 -25374
rect 30242 -25428 30298 -25426
rect 30242 -25694 30298 -25692
rect 30242 -25746 30244 -25694
rect 30244 -25746 30296 -25694
rect 30296 -25746 30298 -25694
rect 30242 -25748 30298 -25746
rect 30242 -26014 30298 -26012
rect 30242 -26066 30244 -26014
rect 30244 -26066 30296 -26014
rect 30296 -26066 30298 -26014
rect 30242 -26068 30298 -26066
rect 30242 -26334 30298 -26332
rect 30242 -26386 30244 -26334
rect 30244 -26386 30296 -26334
rect 30296 -26386 30298 -26334
rect 30242 -26388 30298 -26386
rect 30242 -26654 30298 -26652
rect 30242 -26706 30244 -26654
rect 30244 -26706 30296 -26654
rect 30296 -26706 30298 -26654
rect 30242 -26708 30298 -26706
rect 30242 -26974 30298 -26972
rect 30242 -27026 30244 -26974
rect 30244 -27026 30296 -26974
rect 30296 -27026 30298 -26974
rect 30242 -27028 30298 -27026
rect 30242 -27294 30298 -27292
rect 30242 -27346 30244 -27294
rect 30244 -27346 30296 -27294
rect 30296 -27346 30298 -27294
rect 30242 -27348 30298 -27346
rect 30242 -27614 30298 -27612
rect 30242 -27666 30244 -27614
rect 30244 -27666 30296 -27614
rect 30296 -27666 30298 -27614
rect 30242 -27668 30298 -27666
rect 30242 -27934 30298 -27932
rect 30242 -27986 30244 -27934
rect 30244 -27986 30296 -27934
rect 30296 -27986 30298 -27934
rect 30242 -27988 30298 -27986
rect 30242 -28254 30298 -28252
rect 30242 -28306 30244 -28254
rect 30244 -28306 30296 -28254
rect 30296 -28306 30298 -28254
rect 30242 -28308 30298 -28306
rect 30242 -28574 30298 -28572
rect 30242 -28626 30244 -28574
rect 30244 -28626 30296 -28574
rect 30296 -28626 30298 -28574
rect 30242 -28628 30298 -28626
rect 30242 -28894 30298 -28892
rect 30242 -28946 30244 -28894
rect 30244 -28946 30296 -28894
rect 30296 -28946 30298 -28894
rect 30242 -28948 30298 -28946
rect 30242 -29214 30298 -29212
rect 30242 -29266 30244 -29214
rect 30244 -29266 30296 -29214
rect 30296 -29266 30298 -29214
rect 30242 -29268 30298 -29266
rect 30242 -29534 30298 -29532
rect 30242 -29586 30244 -29534
rect 30244 -29586 30296 -29534
rect 30296 -29586 30298 -29534
rect 30242 -29588 30298 -29586
rect 30242 -29854 30298 -29852
rect 30242 -29906 30244 -29854
rect 30244 -29906 30296 -29854
rect 30296 -29906 30298 -29854
rect 30242 -29908 30298 -29906
rect 30242 -30174 30298 -30172
rect 30242 -30226 30244 -30174
rect 30244 -30226 30296 -30174
rect 30296 -30226 30298 -30174
rect 30242 -30228 30298 -30226
rect 37708 -23774 37764 -23772
rect 37708 -23826 37710 -23774
rect 37710 -23826 37762 -23774
rect 37762 -23826 37764 -23774
rect 37708 -23828 37764 -23826
rect 37708 -24094 37764 -24092
rect 37708 -24146 37710 -24094
rect 37710 -24146 37762 -24094
rect 37762 -24146 37764 -24094
rect 37708 -24148 37764 -24146
rect 37708 -24414 37764 -24412
rect 37708 -24466 37710 -24414
rect 37710 -24466 37762 -24414
rect 37762 -24466 37764 -24414
rect 37708 -24468 37764 -24466
rect 37708 -24734 37764 -24732
rect 37708 -24786 37710 -24734
rect 37710 -24786 37762 -24734
rect 37762 -24786 37764 -24734
rect 37708 -24788 37764 -24786
rect 37708 -25054 37764 -25052
rect 37708 -25106 37710 -25054
rect 37710 -25106 37762 -25054
rect 37762 -25106 37764 -25054
rect 37708 -25108 37764 -25106
rect 37708 -25374 37764 -25372
rect 37708 -25426 37710 -25374
rect 37710 -25426 37762 -25374
rect 37762 -25426 37764 -25374
rect 37708 -25428 37764 -25426
rect 37708 -25694 37764 -25692
rect 37708 -25746 37710 -25694
rect 37710 -25746 37762 -25694
rect 37762 -25746 37764 -25694
rect 37708 -25748 37764 -25746
rect 37708 -26014 37764 -26012
rect 37708 -26066 37710 -26014
rect 37710 -26066 37762 -26014
rect 37762 -26066 37764 -26014
rect 37708 -26068 37764 -26066
rect 37708 -26334 37764 -26332
rect 37708 -26386 37710 -26334
rect 37710 -26386 37762 -26334
rect 37762 -26386 37764 -26334
rect 37708 -26388 37764 -26386
rect 37708 -26654 37764 -26652
rect 37708 -26706 37710 -26654
rect 37710 -26706 37762 -26654
rect 37762 -26706 37764 -26654
rect 37708 -26708 37764 -26706
rect 37708 -26974 37764 -26972
rect 37708 -27026 37710 -26974
rect 37710 -27026 37762 -26974
rect 37762 -27026 37764 -26974
rect 37708 -27028 37764 -27026
rect 37708 -27294 37764 -27292
rect 37708 -27346 37710 -27294
rect 37710 -27346 37762 -27294
rect 37762 -27346 37764 -27294
rect 37708 -27348 37764 -27346
rect 37708 -27614 37764 -27612
rect 37708 -27666 37710 -27614
rect 37710 -27666 37762 -27614
rect 37762 -27666 37764 -27614
rect 37708 -27668 37764 -27666
rect 37708 -27934 37764 -27932
rect 37708 -27986 37710 -27934
rect 37710 -27986 37762 -27934
rect 37762 -27986 37764 -27934
rect 37708 -27988 37764 -27986
rect 37708 -28254 37764 -28252
rect 37708 -28306 37710 -28254
rect 37710 -28306 37762 -28254
rect 37762 -28306 37764 -28254
rect 37708 -28308 37764 -28306
rect 37708 -28574 37764 -28572
rect 37708 -28626 37710 -28574
rect 37710 -28626 37762 -28574
rect 37762 -28626 37764 -28574
rect 37708 -28628 37764 -28626
rect 37708 -28894 37764 -28892
rect 37708 -28946 37710 -28894
rect 37710 -28946 37762 -28894
rect 37762 -28946 37764 -28894
rect 37708 -28948 37764 -28946
rect 37708 -29214 37764 -29212
rect 37708 -29266 37710 -29214
rect 37710 -29266 37762 -29214
rect 37762 -29266 37764 -29214
rect 37708 -29268 37764 -29266
rect 37708 -29534 37764 -29532
rect 37708 -29586 37710 -29534
rect 37710 -29586 37762 -29534
rect 37762 -29586 37764 -29534
rect 37708 -29588 37764 -29586
rect 37708 -29854 37764 -29852
rect 37708 -29906 37710 -29854
rect 37710 -29906 37762 -29854
rect 37762 -29906 37764 -29854
rect 37708 -29908 37764 -29906
rect 37708 -30174 37764 -30172
rect 37708 -30226 37710 -30174
rect 37710 -30226 37762 -30174
rect 37762 -30226 37764 -30174
rect 37708 -30228 37764 -30226
rect 30242 -30494 30298 -30492
rect 30242 -30546 30244 -30494
rect 30244 -30546 30296 -30494
rect 30296 -30546 30298 -30494
rect 30242 -30548 30298 -30546
rect 37708 -30494 37764 -30492
rect 37708 -30546 37710 -30494
rect 37710 -30546 37762 -30494
rect 37762 -30546 37764 -30494
rect 37708 -30548 37764 -30546
rect 30612 -30704 30668 -30702
rect 30612 -30756 30614 -30704
rect 30614 -30756 30666 -30704
rect 30666 -30756 30668 -30704
rect 30612 -30758 30668 -30756
rect 30932 -30704 30988 -30702
rect 30932 -30756 30934 -30704
rect 30934 -30756 30986 -30704
rect 30986 -30756 30988 -30704
rect 30932 -30758 30988 -30756
rect 31252 -30704 31308 -30702
rect 31252 -30756 31254 -30704
rect 31254 -30756 31306 -30704
rect 31306 -30756 31308 -30704
rect 31252 -30758 31308 -30756
rect 31572 -30704 31628 -30702
rect 31572 -30756 31574 -30704
rect 31574 -30756 31626 -30704
rect 31626 -30756 31628 -30704
rect 31572 -30758 31628 -30756
rect 31892 -30704 31948 -30702
rect 31892 -30756 31894 -30704
rect 31894 -30756 31946 -30704
rect 31946 -30756 31948 -30704
rect 31892 -30758 31948 -30756
rect 32212 -30704 32268 -30702
rect 32212 -30756 32214 -30704
rect 32214 -30756 32266 -30704
rect 32266 -30756 32268 -30704
rect 32212 -30758 32268 -30756
rect 32532 -30704 32588 -30702
rect 32532 -30756 32534 -30704
rect 32534 -30756 32586 -30704
rect 32586 -30756 32588 -30704
rect 32532 -30758 32588 -30756
rect 32852 -30704 32908 -30702
rect 32852 -30756 32854 -30704
rect 32854 -30756 32906 -30704
rect 32906 -30756 32908 -30704
rect 32852 -30758 32908 -30756
rect 33172 -30704 33228 -30702
rect 33172 -30756 33174 -30704
rect 33174 -30756 33226 -30704
rect 33226 -30756 33228 -30704
rect 33172 -30758 33228 -30756
rect 33492 -30704 33548 -30702
rect 33492 -30756 33494 -30704
rect 33494 -30756 33546 -30704
rect 33546 -30756 33548 -30704
rect 33492 -30758 33548 -30756
rect 33812 -30704 33868 -30702
rect 33812 -30756 33814 -30704
rect 33814 -30756 33866 -30704
rect 33866 -30756 33868 -30704
rect 33812 -30758 33868 -30756
rect 34132 -30704 34188 -30702
rect 34132 -30756 34134 -30704
rect 34134 -30756 34186 -30704
rect 34186 -30756 34188 -30704
rect 34132 -30758 34188 -30756
rect 34452 -30704 34508 -30702
rect 34452 -30756 34454 -30704
rect 34454 -30756 34506 -30704
rect 34506 -30756 34508 -30704
rect 34452 -30758 34508 -30756
rect 34772 -30704 34828 -30702
rect 34772 -30756 34774 -30704
rect 34774 -30756 34826 -30704
rect 34826 -30756 34828 -30704
rect 34772 -30758 34828 -30756
rect 35092 -30704 35148 -30702
rect 35092 -30756 35094 -30704
rect 35094 -30756 35146 -30704
rect 35146 -30756 35148 -30704
rect 35092 -30758 35148 -30756
rect 35412 -30704 35468 -30702
rect 35412 -30756 35414 -30704
rect 35414 -30756 35466 -30704
rect 35466 -30756 35468 -30704
rect 35412 -30758 35468 -30756
rect 35732 -30704 35788 -30702
rect 35732 -30756 35734 -30704
rect 35734 -30756 35786 -30704
rect 35786 -30756 35788 -30704
rect 35732 -30758 35788 -30756
rect 36052 -30704 36108 -30702
rect 36052 -30756 36054 -30704
rect 36054 -30756 36106 -30704
rect 36106 -30756 36108 -30704
rect 36052 -30758 36108 -30756
rect 36372 -30704 36428 -30702
rect 36372 -30756 36374 -30704
rect 36374 -30756 36426 -30704
rect 36426 -30756 36428 -30704
rect 36372 -30758 36428 -30756
rect 36692 -30704 36748 -30702
rect 36692 -30756 36694 -30704
rect 36694 -30756 36746 -30704
rect 36746 -30756 36748 -30704
rect 36692 -30758 36748 -30756
rect 37012 -30704 37068 -30702
rect 37012 -30756 37014 -30704
rect 37014 -30756 37066 -30704
rect 37066 -30756 37068 -30704
rect 37012 -30758 37068 -30756
rect 37332 -30704 37388 -30702
rect 37332 -30756 37334 -30704
rect 37334 -30756 37386 -30704
rect 37386 -30756 37388 -30704
rect 37332 -30758 37388 -30756
rect 42612 -23248 42668 -23246
rect 42612 -23300 42614 -23248
rect 42614 -23300 42666 -23248
rect 42666 -23300 42668 -23248
rect 42612 -23302 42668 -23300
rect 42932 -23248 42988 -23246
rect 42932 -23300 42934 -23248
rect 42934 -23300 42986 -23248
rect 42986 -23300 42988 -23248
rect 42932 -23302 42988 -23300
rect 43252 -23248 43308 -23246
rect 43252 -23300 43254 -23248
rect 43254 -23300 43306 -23248
rect 43306 -23300 43308 -23248
rect 43252 -23302 43308 -23300
rect 43572 -23248 43628 -23246
rect 43572 -23300 43574 -23248
rect 43574 -23300 43626 -23248
rect 43626 -23300 43628 -23248
rect 43572 -23302 43628 -23300
rect 43892 -23248 43948 -23246
rect 43892 -23300 43894 -23248
rect 43894 -23300 43946 -23248
rect 43946 -23300 43948 -23248
rect 43892 -23302 43948 -23300
rect 44212 -23248 44268 -23246
rect 44212 -23300 44214 -23248
rect 44214 -23300 44266 -23248
rect 44266 -23300 44268 -23248
rect 44212 -23302 44268 -23300
rect 44532 -23248 44588 -23246
rect 44532 -23300 44534 -23248
rect 44534 -23300 44586 -23248
rect 44586 -23300 44588 -23248
rect 44532 -23302 44588 -23300
rect 44852 -23248 44908 -23246
rect 44852 -23300 44854 -23248
rect 44854 -23300 44906 -23248
rect 44906 -23300 44908 -23248
rect 44852 -23302 44908 -23300
rect 45172 -23248 45228 -23246
rect 45172 -23300 45174 -23248
rect 45174 -23300 45226 -23248
rect 45226 -23300 45228 -23248
rect 45172 -23302 45228 -23300
rect 45492 -23248 45548 -23246
rect 45492 -23300 45494 -23248
rect 45494 -23300 45546 -23248
rect 45546 -23300 45548 -23248
rect 45492 -23302 45548 -23300
rect 45812 -23248 45868 -23246
rect 45812 -23300 45814 -23248
rect 45814 -23300 45866 -23248
rect 45866 -23300 45868 -23248
rect 45812 -23302 45868 -23300
rect 46132 -23248 46188 -23246
rect 46132 -23300 46134 -23248
rect 46134 -23300 46186 -23248
rect 46186 -23300 46188 -23248
rect 46132 -23302 46188 -23300
rect 46452 -23248 46508 -23246
rect 46452 -23300 46454 -23248
rect 46454 -23300 46506 -23248
rect 46506 -23300 46508 -23248
rect 46452 -23302 46508 -23300
rect 46772 -23248 46828 -23246
rect 46772 -23300 46774 -23248
rect 46774 -23300 46826 -23248
rect 46826 -23300 46828 -23248
rect 46772 -23302 46828 -23300
rect 47092 -23248 47148 -23246
rect 47092 -23300 47094 -23248
rect 47094 -23300 47146 -23248
rect 47146 -23300 47148 -23248
rect 47092 -23302 47148 -23300
rect 47412 -23248 47468 -23246
rect 47412 -23300 47414 -23248
rect 47414 -23300 47466 -23248
rect 47466 -23300 47468 -23248
rect 47412 -23302 47468 -23300
rect 47732 -23248 47788 -23246
rect 47732 -23300 47734 -23248
rect 47734 -23300 47786 -23248
rect 47786 -23300 47788 -23248
rect 47732 -23302 47788 -23300
rect 48052 -23248 48108 -23246
rect 48052 -23300 48054 -23248
rect 48054 -23300 48106 -23248
rect 48106 -23300 48108 -23248
rect 48052 -23302 48108 -23300
rect 48372 -23248 48428 -23246
rect 48372 -23300 48374 -23248
rect 48374 -23300 48426 -23248
rect 48426 -23300 48428 -23248
rect 48372 -23302 48428 -23300
rect 48692 -23248 48748 -23246
rect 48692 -23300 48694 -23248
rect 48694 -23300 48746 -23248
rect 48746 -23300 48748 -23248
rect 48692 -23302 48748 -23300
rect 49012 -23248 49068 -23246
rect 49012 -23300 49014 -23248
rect 49014 -23300 49066 -23248
rect 49066 -23300 49068 -23248
rect 49012 -23302 49068 -23300
rect 49332 -23248 49388 -23246
rect 49332 -23300 49334 -23248
rect 49334 -23300 49386 -23248
rect 49386 -23300 49388 -23248
rect 49332 -23302 49388 -23300
rect 42242 -23454 42298 -23452
rect 42242 -23506 42244 -23454
rect 42244 -23506 42296 -23454
rect 42296 -23506 42298 -23454
rect 42242 -23508 42298 -23506
rect 49708 -23454 49764 -23452
rect 49708 -23506 49710 -23454
rect 49710 -23506 49762 -23454
rect 49762 -23506 49764 -23454
rect 49708 -23508 49764 -23506
rect 42242 -23774 42298 -23772
rect 42242 -23826 42244 -23774
rect 42244 -23826 42296 -23774
rect 42296 -23826 42298 -23774
rect 42242 -23828 42298 -23826
rect 42242 -24094 42298 -24092
rect 42242 -24146 42244 -24094
rect 42244 -24146 42296 -24094
rect 42296 -24146 42298 -24094
rect 42242 -24148 42298 -24146
rect 42242 -24414 42298 -24412
rect 42242 -24466 42244 -24414
rect 42244 -24466 42296 -24414
rect 42296 -24466 42298 -24414
rect 42242 -24468 42298 -24466
rect 42242 -24734 42298 -24732
rect 42242 -24786 42244 -24734
rect 42244 -24786 42296 -24734
rect 42296 -24786 42298 -24734
rect 42242 -24788 42298 -24786
rect 42242 -25054 42298 -25052
rect 42242 -25106 42244 -25054
rect 42244 -25106 42296 -25054
rect 42296 -25106 42298 -25054
rect 42242 -25108 42298 -25106
rect 42242 -25374 42298 -25372
rect 42242 -25426 42244 -25374
rect 42244 -25426 42296 -25374
rect 42296 -25426 42298 -25374
rect 42242 -25428 42298 -25426
rect 42242 -25694 42298 -25692
rect 42242 -25746 42244 -25694
rect 42244 -25746 42296 -25694
rect 42296 -25746 42298 -25694
rect 42242 -25748 42298 -25746
rect 42242 -26014 42298 -26012
rect 42242 -26066 42244 -26014
rect 42244 -26066 42296 -26014
rect 42296 -26066 42298 -26014
rect 42242 -26068 42298 -26066
rect 42242 -26334 42298 -26332
rect 42242 -26386 42244 -26334
rect 42244 -26386 42296 -26334
rect 42296 -26386 42298 -26334
rect 42242 -26388 42298 -26386
rect 42242 -26654 42298 -26652
rect 42242 -26706 42244 -26654
rect 42244 -26706 42296 -26654
rect 42296 -26706 42298 -26654
rect 42242 -26708 42298 -26706
rect 42242 -26974 42298 -26972
rect 42242 -27026 42244 -26974
rect 42244 -27026 42296 -26974
rect 42296 -27026 42298 -26974
rect 42242 -27028 42298 -27026
rect 42242 -27294 42298 -27292
rect 42242 -27346 42244 -27294
rect 42244 -27346 42296 -27294
rect 42296 -27346 42298 -27294
rect 42242 -27348 42298 -27346
rect 42242 -27614 42298 -27612
rect 42242 -27666 42244 -27614
rect 42244 -27666 42296 -27614
rect 42296 -27666 42298 -27614
rect 42242 -27668 42298 -27666
rect 42242 -27934 42298 -27932
rect 42242 -27986 42244 -27934
rect 42244 -27986 42296 -27934
rect 42296 -27986 42298 -27934
rect 42242 -27988 42298 -27986
rect 42242 -28254 42298 -28252
rect 42242 -28306 42244 -28254
rect 42244 -28306 42296 -28254
rect 42296 -28306 42298 -28254
rect 42242 -28308 42298 -28306
rect 42242 -28574 42298 -28572
rect 42242 -28626 42244 -28574
rect 42244 -28626 42296 -28574
rect 42296 -28626 42298 -28574
rect 42242 -28628 42298 -28626
rect 42242 -28894 42298 -28892
rect 42242 -28946 42244 -28894
rect 42244 -28946 42296 -28894
rect 42296 -28946 42298 -28894
rect 42242 -28948 42298 -28946
rect 42242 -29214 42298 -29212
rect 42242 -29266 42244 -29214
rect 42244 -29266 42296 -29214
rect 42296 -29266 42298 -29214
rect 42242 -29268 42298 -29266
rect 42242 -29534 42298 -29532
rect 42242 -29586 42244 -29534
rect 42244 -29586 42296 -29534
rect 42296 -29586 42298 -29534
rect 42242 -29588 42298 -29586
rect 42242 -29854 42298 -29852
rect 42242 -29906 42244 -29854
rect 42244 -29906 42296 -29854
rect 42296 -29906 42298 -29854
rect 42242 -29908 42298 -29906
rect 42242 -30174 42298 -30172
rect 42242 -30226 42244 -30174
rect 42244 -30226 42296 -30174
rect 42296 -30226 42298 -30174
rect 42242 -30228 42298 -30226
rect 49708 -23774 49764 -23772
rect 49708 -23826 49710 -23774
rect 49710 -23826 49762 -23774
rect 49762 -23826 49764 -23774
rect 49708 -23828 49764 -23826
rect 49708 -24094 49764 -24092
rect 49708 -24146 49710 -24094
rect 49710 -24146 49762 -24094
rect 49762 -24146 49764 -24094
rect 49708 -24148 49764 -24146
rect 49708 -24414 49764 -24412
rect 49708 -24466 49710 -24414
rect 49710 -24466 49762 -24414
rect 49762 -24466 49764 -24414
rect 49708 -24468 49764 -24466
rect 49708 -24734 49764 -24732
rect 49708 -24786 49710 -24734
rect 49710 -24786 49762 -24734
rect 49762 -24786 49764 -24734
rect 49708 -24788 49764 -24786
rect 49708 -25054 49764 -25052
rect 49708 -25106 49710 -25054
rect 49710 -25106 49762 -25054
rect 49762 -25106 49764 -25054
rect 49708 -25108 49764 -25106
rect 49708 -25374 49764 -25372
rect 49708 -25426 49710 -25374
rect 49710 -25426 49762 -25374
rect 49762 -25426 49764 -25374
rect 49708 -25428 49764 -25426
rect 49708 -25694 49764 -25692
rect 49708 -25746 49710 -25694
rect 49710 -25746 49762 -25694
rect 49762 -25746 49764 -25694
rect 49708 -25748 49764 -25746
rect 49708 -26014 49764 -26012
rect 49708 -26066 49710 -26014
rect 49710 -26066 49762 -26014
rect 49762 -26066 49764 -26014
rect 49708 -26068 49764 -26066
rect 49708 -26334 49764 -26332
rect 49708 -26386 49710 -26334
rect 49710 -26386 49762 -26334
rect 49762 -26386 49764 -26334
rect 49708 -26388 49764 -26386
rect 49708 -26654 49764 -26652
rect 49708 -26706 49710 -26654
rect 49710 -26706 49762 -26654
rect 49762 -26706 49764 -26654
rect 49708 -26708 49764 -26706
rect 49708 -26974 49764 -26972
rect 49708 -27026 49710 -26974
rect 49710 -27026 49762 -26974
rect 49762 -27026 49764 -26974
rect 49708 -27028 49764 -27026
rect 49708 -27294 49764 -27292
rect 49708 -27346 49710 -27294
rect 49710 -27346 49762 -27294
rect 49762 -27346 49764 -27294
rect 49708 -27348 49764 -27346
rect 49708 -27614 49764 -27612
rect 49708 -27666 49710 -27614
rect 49710 -27666 49762 -27614
rect 49762 -27666 49764 -27614
rect 49708 -27668 49764 -27666
rect 49708 -27934 49764 -27932
rect 49708 -27986 49710 -27934
rect 49710 -27986 49762 -27934
rect 49762 -27986 49764 -27934
rect 49708 -27988 49764 -27986
rect 49708 -28254 49764 -28252
rect 49708 -28306 49710 -28254
rect 49710 -28306 49762 -28254
rect 49762 -28306 49764 -28254
rect 49708 -28308 49764 -28306
rect 49708 -28574 49764 -28572
rect 49708 -28626 49710 -28574
rect 49710 -28626 49762 -28574
rect 49762 -28626 49764 -28574
rect 49708 -28628 49764 -28626
rect 49708 -28894 49764 -28892
rect 49708 -28946 49710 -28894
rect 49710 -28946 49762 -28894
rect 49762 -28946 49764 -28894
rect 49708 -28948 49764 -28946
rect 49708 -29214 49764 -29212
rect 49708 -29266 49710 -29214
rect 49710 -29266 49762 -29214
rect 49762 -29266 49764 -29214
rect 49708 -29268 49764 -29266
rect 49708 -29534 49764 -29532
rect 49708 -29586 49710 -29534
rect 49710 -29586 49762 -29534
rect 49762 -29586 49764 -29534
rect 49708 -29588 49764 -29586
rect 49708 -29854 49764 -29852
rect 49708 -29906 49710 -29854
rect 49710 -29906 49762 -29854
rect 49762 -29906 49764 -29854
rect 49708 -29908 49764 -29906
rect 49708 -30174 49764 -30172
rect 49708 -30226 49710 -30174
rect 49710 -30226 49762 -30174
rect 49762 -30226 49764 -30174
rect 49708 -30228 49764 -30226
rect 42242 -30494 42298 -30492
rect 42242 -30546 42244 -30494
rect 42244 -30546 42296 -30494
rect 42296 -30546 42298 -30494
rect 42242 -30548 42298 -30546
rect 49708 -30494 49764 -30492
rect 49708 -30546 49710 -30494
rect 49710 -30546 49762 -30494
rect 49762 -30546 49764 -30494
rect 49708 -30548 49764 -30546
rect 42612 -30704 42668 -30702
rect 42612 -30756 42614 -30704
rect 42614 -30756 42666 -30704
rect 42666 -30756 42668 -30704
rect 42612 -30758 42668 -30756
rect 42932 -30704 42988 -30702
rect 42932 -30756 42934 -30704
rect 42934 -30756 42986 -30704
rect 42986 -30756 42988 -30704
rect 42932 -30758 42988 -30756
rect 43252 -30704 43308 -30702
rect 43252 -30756 43254 -30704
rect 43254 -30756 43306 -30704
rect 43306 -30756 43308 -30704
rect 43252 -30758 43308 -30756
rect 43572 -30704 43628 -30702
rect 43572 -30756 43574 -30704
rect 43574 -30756 43626 -30704
rect 43626 -30756 43628 -30704
rect 43572 -30758 43628 -30756
rect 43892 -30704 43948 -30702
rect 43892 -30756 43894 -30704
rect 43894 -30756 43946 -30704
rect 43946 -30756 43948 -30704
rect 43892 -30758 43948 -30756
rect 44212 -30704 44268 -30702
rect 44212 -30756 44214 -30704
rect 44214 -30756 44266 -30704
rect 44266 -30756 44268 -30704
rect 44212 -30758 44268 -30756
rect 44532 -30704 44588 -30702
rect 44532 -30756 44534 -30704
rect 44534 -30756 44586 -30704
rect 44586 -30756 44588 -30704
rect 44532 -30758 44588 -30756
rect 44852 -30704 44908 -30702
rect 44852 -30756 44854 -30704
rect 44854 -30756 44906 -30704
rect 44906 -30756 44908 -30704
rect 44852 -30758 44908 -30756
rect 45172 -30704 45228 -30702
rect 45172 -30756 45174 -30704
rect 45174 -30756 45226 -30704
rect 45226 -30756 45228 -30704
rect 45172 -30758 45228 -30756
rect 45492 -30704 45548 -30702
rect 45492 -30756 45494 -30704
rect 45494 -30756 45546 -30704
rect 45546 -30756 45548 -30704
rect 45492 -30758 45548 -30756
rect 45812 -30704 45868 -30702
rect 45812 -30756 45814 -30704
rect 45814 -30756 45866 -30704
rect 45866 -30756 45868 -30704
rect 45812 -30758 45868 -30756
rect 46132 -30704 46188 -30702
rect 46132 -30756 46134 -30704
rect 46134 -30756 46186 -30704
rect 46186 -30756 46188 -30704
rect 46132 -30758 46188 -30756
rect 46452 -30704 46508 -30702
rect 46452 -30756 46454 -30704
rect 46454 -30756 46506 -30704
rect 46506 -30756 46508 -30704
rect 46452 -30758 46508 -30756
rect 46772 -30704 46828 -30702
rect 46772 -30756 46774 -30704
rect 46774 -30756 46826 -30704
rect 46826 -30756 46828 -30704
rect 46772 -30758 46828 -30756
rect 47092 -30704 47148 -30702
rect 47092 -30756 47094 -30704
rect 47094 -30756 47146 -30704
rect 47146 -30756 47148 -30704
rect 47092 -30758 47148 -30756
rect 47412 -30704 47468 -30702
rect 47412 -30756 47414 -30704
rect 47414 -30756 47466 -30704
rect 47466 -30756 47468 -30704
rect 47412 -30758 47468 -30756
rect 47732 -30704 47788 -30702
rect 47732 -30756 47734 -30704
rect 47734 -30756 47786 -30704
rect 47786 -30756 47788 -30704
rect 47732 -30758 47788 -30756
rect 48052 -30704 48108 -30702
rect 48052 -30756 48054 -30704
rect 48054 -30756 48106 -30704
rect 48106 -30756 48108 -30704
rect 48052 -30758 48108 -30756
rect 48372 -30704 48428 -30702
rect 48372 -30756 48374 -30704
rect 48374 -30756 48426 -30704
rect 48426 -30756 48428 -30704
rect 48372 -30758 48428 -30756
rect 48692 -30704 48748 -30702
rect 48692 -30756 48694 -30704
rect 48694 -30756 48746 -30704
rect 48746 -30756 48748 -30704
rect 48692 -30758 48748 -30756
rect 49012 -30704 49068 -30702
rect 49012 -30756 49014 -30704
rect 49014 -30756 49066 -30704
rect 49066 -30756 49068 -30704
rect 49012 -30758 49068 -30756
rect 49332 -30704 49388 -30702
rect 49332 -30756 49334 -30704
rect 49334 -30756 49386 -30704
rect 49386 -30756 49388 -30704
rect 49332 -30758 49388 -30756
<< metal3 >>
rect 18200 -2500 21600 -2400
rect 13200 -9600 16000 -2700
rect 16400 -8000 17700 -2648
rect 18200 -3000 18300 -2500
rect 21500 -3000 21600 -2500
rect 18200 -3100 21600 -3000
rect 21872 -5560 22002 -5550
rect 21872 -5650 21882 -5560
rect 21992 -5650 22002 -5560
rect 22202 -5600 23002 -2900
rect 21872 -5660 22002 -5650
rect 22402 -5720 23002 -5600
rect 18195 -5740 22342 -5731
rect 18195 -5796 18203 -5740
rect 18259 -5796 21744 -5740
rect 21800 -5796 22342 -5740
rect 18195 -5805 22342 -5796
rect 18262 -5836 21741 -5805
rect 22268 -6251 22342 -5805
rect 22402 -5880 22422 -5720
rect 22982 -5880 23002 -5720
rect 22402 -5960 22432 -5880
rect 22972 -5960 23002 -5880
rect 22402 -5990 23002 -5960
rect 22712 -6250 22782 -5990
rect 22452 -6251 22602 -6250
rect 22268 -6270 22602 -6251
rect 22268 -6325 22472 -6270
rect 19291 -6650 19945 -6638
rect 19291 -6706 19297 -6650
rect 19363 -6706 19489 -6650
rect 19555 -6706 19681 -6650
rect 19747 -6706 19873 -6650
rect 19939 -6706 19945 -6650
rect 19291 -6720 19945 -6706
rect 20059 -6650 20713 -6638
rect 20059 -6706 20065 -6650
rect 20131 -6706 20257 -6650
rect 20323 -6706 20449 -6650
rect 20515 -6706 20641 -6650
rect 20707 -6706 20713 -6650
rect 22452 -6660 22472 -6325
rect 22582 -6660 22602 -6270
rect 22452 -6680 22602 -6660
rect 22682 -6270 22832 -6250
rect 22682 -6660 22702 -6270
rect 22812 -6660 22832 -6270
rect 22682 -6680 22832 -6660
rect 20059 -6720 20713 -6706
rect 19860 -6930 19940 -6720
rect 20060 -6780 20140 -6720
rect 20060 -6860 21200 -6780
rect 18800 -6940 18980 -6930
rect 18800 -7000 18810 -6940
rect 18970 -7000 18980 -6940
rect 16400 -8200 18100 -8000
rect 18800 -8200 18980 -7000
rect 19860 -7010 21040 -6930
rect 16400 -8248 17700 -8200
rect 16400 -8268 17300 -8248
rect 16400 -8488 16920 -8268
rect 17130 -8488 17300 -8268
rect 16400 -8748 17300 -8488
rect 16400 -9148 16500 -8748
rect 17200 -9148 17300 -8748
rect 16400 -9248 17300 -9148
rect 17380 -8440 17700 -8420
rect 17380 -9360 17400 -8440
rect 17680 -9360 17700 -8440
rect 17800 -8500 18980 -8200
rect 20960 -8260 21040 -7010
rect 21120 -8100 21200 -6860
rect 23080 -7480 24410 -7470
rect 23080 -7540 23270 -7480
rect 23410 -7540 24410 -7480
rect 23080 -7550 24410 -7540
rect 23080 -8100 23160 -7550
rect 21120 -8180 23160 -8100
rect 23290 -7800 24200 -7790
rect 23290 -7860 23550 -7800
rect 23690 -7860 24200 -7800
rect 23290 -7870 24200 -7860
rect 23290 -8260 23370 -7870
rect 20960 -8340 23370 -8260
rect 17380 -9380 17700 -9360
rect 16600 -9510 16680 -9500
rect 13200 -10200 13300 -9600
rect 15900 -10200 16000 -9600
rect 13200 -10300 16000 -10200
rect 16330 -9520 16470 -9510
rect 16330 -9580 16400 -9520
rect 16460 -9580 16470 -9520
rect 16330 -9590 16470 -9580
rect 16600 -9570 16610 -9510
rect 16670 -9570 16680 -9510
rect 16600 -9580 16680 -9570
rect 6000 -11242 14000 -11000
rect 6000 -11306 6608 -11242
rect 6672 -11306 6928 -11242
rect 6992 -11306 7248 -11242
rect 7312 -11306 7568 -11242
rect 7632 -11306 7888 -11242
rect 7952 -11306 8208 -11242
rect 8272 -11306 8528 -11242
rect 8592 -11306 8848 -11242
rect 8912 -11306 9168 -11242
rect 9232 -11306 9488 -11242
rect 9552 -11306 9808 -11242
rect 9872 -11306 10128 -11242
rect 10192 -11306 10448 -11242
rect 10512 -11306 10768 -11242
rect 10832 -11306 11088 -11242
rect 11152 -11306 11408 -11242
rect 11472 -11306 11728 -11242
rect 11792 -11306 12048 -11242
rect 12112 -11306 12368 -11242
rect 12432 -11306 12688 -11242
rect 12752 -11306 13008 -11242
rect 13072 -11306 13328 -11242
rect 13392 -11306 14000 -11242
rect 6000 -11448 14000 -11306
rect 6000 -11512 6238 -11448
rect 6302 -11512 13704 -11448
rect 13768 -11512 14000 -11448
rect 6000 -11540 14000 -11512
rect 6000 -11768 6540 -11540
rect 6000 -11832 6238 -11768
rect 6302 -11832 6540 -11768
rect 6000 -12088 6540 -11832
rect 6000 -12152 6238 -12088
rect 6302 -12152 6540 -12088
rect 6000 -12408 6540 -12152
rect 6000 -12472 6238 -12408
rect 6302 -12472 6540 -12408
rect 6000 -12728 6540 -12472
rect 6000 -12792 6238 -12728
rect 6302 -12792 6540 -12728
rect 6000 -13048 6540 -12792
rect 6000 -13112 6238 -13048
rect 6302 -13112 6540 -13048
rect 6000 -13368 6540 -13112
rect 6000 -13432 6238 -13368
rect 6302 -13432 6540 -13368
rect 6000 -13688 6540 -13432
rect 6000 -13752 6238 -13688
rect 6302 -13752 6540 -13688
rect 6000 -14008 6540 -13752
rect 6000 -14072 6238 -14008
rect 6302 -14072 6540 -14008
rect 6000 -14328 6540 -14072
rect 6000 -14392 6238 -14328
rect 6302 -14392 6540 -14328
rect 6000 -14648 6540 -14392
rect 6000 -14712 6238 -14648
rect 6302 -14712 6540 -14648
rect 6000 -14968 6540 -14712
rect 6000 -15032 6238 -14968
rect 6302 -15032 6540 -14968
rect 6000 -15288 6540 -15032
rect 6000 -15352 6238 -15288
rect 6302 -15352 6540 -15288
rect 6000 -15608 6540 -15352
rect 6000 -15672 6238 -15608
rect 6302 -15672 6540 -15608
rect 6000 -15928 6540 -15672
rect 6000 -15992 6238 -15928
rect 6302 -15992 6540 -15928
rect 6000 -16248 6540 -15992
rect 6000 -16312 6238 -16248
rect 6302 -16312 6540 -16248
rect 6000 -16568 6540 -16312
rect 6000 -16632 6238 -16568
rect 6302 -16632 6540 -16568
rect 6000 -16888 6540 -16632
rect 6000 -16952 6238 -16888
rect 6302 -16952 6540 -16888
rect 6000 -17208 6540 -16952
rect 6000 -17272 6238 -17208
rect 6302 -17272 6540 -17208
rect 6000 -17528 6540 -17272
rect 6000 -17592 6238 -17528
rect 6302 -17592 6540 -17528
rect 6000 -17848 6540 -17592
rect 6000 -17912 6238 -17848
rect 6302 -17912 6540 -17848
rect 6000 -18168 6540 -17912
rect 6000 -18232 6238 -18168
rect 6302 -18232 6540 -18168
rect 6000 -18460 6540 -18232
rect 13460 -11768 14000 -11540
rect 13460 -11832 13704 -11768
rect 13768 -11832 14000 -11768
rect 13460 -12088 14000 -11832
rect 13460 -12152 13704 -12088
rect 13768 -12152 14000 -12088
rect 13460 -12408 14000 -12152
rect 13460 -12472 13704 -12408
rect 13768 -12472 14000 -12408
rect 13460 -12728 14000 -12472
rect 13460 -12792 13704 -12728
rect 13768 -12792 14000 -12728
rect 13460 -13048 14000 -12792
rect 13460 -13112 13704 -13048
rect 13768 -13112 14000 -13048
rect 13460 -13368 14000 -13112
rect 13460 -13432 13704 -13368
rect 13768 -13432 14000 -13368
rect 13460 -13688 14000 -13432
rect 13460 -13752 13704 -13688
rect 13768 -13752 14000 -13688
rect 13460 -14008 14000 -13752
rect 13460 -14072 13704 -14008
rect 13768 -14072 14000 -14008
rect 13460 -14328 14000 -14072
rect 13460 -14392 13704 -14328
rect 13768 -14392 14000 -14328
rect 13460 -14648 14000 -14392
rect 13460 -14712 13704 -14648
rect 13768 -14712 14000 -14648
rect 13460 -14968 14000 -14712
rect 13460 -15032 13704 -14968
rect 13768 -15032 14000 -14968
rect 13460 -15288 14000 -15032
rect 13460 -15352 13704 -15288
rect 13768 -15352 14000 -15288
rect 13460 -15608 14000 -15352
rect 13460 -15672 13704 -15608
rect 13768 -15672 14000 -15608
rect 13460 -15928 14000 -15672
rect 13460 -15992 13704 -15928
rect 13768 -15992 14000 -15928
rect 13460 -16248 14000 -15992
rect 13460 -16312 13704 -16248
rect 13768 -16312 14000 -16248
rect 13460 -16568 14000 -16312
rect 13460 -16632 13704 -16568
rect 13768 -16632 14000 -16568
rect 13460 -16888 14000 -16632
rect 13460 -16952 13704 -16888
rect 13768 -16952 14000 -16888
rect 13460 -17208 14000 -16952
rect 13460 -17272 13704 -17208
rect 13768 -17272 14000 -17208
rect 13460 -17528 14000 -17272
rect 13460 -17592 13704 -17528
rect 13768 -17592 14000 -17528
rect 13460 -17848 14000 -17592
rect 13460 -17912 13704 -17848
rect 13768 -17912 14000 -17848
rect 13460 -18168 14000 -17912
rect 13460 -18232 13704 -18168
rect 13768 -18232 14000 -18168
rect 13460 -18460 14000 -18232
rect 6000 -18488 14000 -18460
rect 6000 -18552 6238 -18488
rect 6302 -18552 13704 -18488
rect 13768 -18552 14000 -18488
rect 6000 -18698 14000 -18552
rect 6000 -18762 6608 -18698
rect 6672 -18762 6928 -18698
rect 6992 -18762 7248 -18698
rect 7312 -18762 7568 -18698
rect 7632 -18762 7888 -18698
rect 7952 -18762 8208 -18698
rect 8272 -18762 8528 -18698
rect 8592 -18762 8848 -18698
rect 8912 -18762 9168 -18698
rect 9232 -18762 9488 -18698
rect 9552 -18762 9808 -18698
rect 9872 -18762 10128 -18698
rect 10192 -18762 10448 -18698
rect 10512 -18762 10768 -18698
rect 10832 -18762 11088 -18698
rect 11152 -18762 11408 -18698
rect 11472 -18762 11728 -18698
rect 11792 -18762 12048 -18698
rect 12112 -18762 12368 -18698
rect 12432 -18762 12688 -18698
rect 12752 -18762 13008 -18698
rect 13072 -18762 13328 -18698
rect 13392 -18762 14000 -18698
rect 6000 -19000 14000 -18762
rect 6000 -23242 14000 -23000
rect 6000 -23306 6608 -23242
rect 6672 -23306 6928 -23242
rect 6992 -23306 7248 -23242
rect 7312 -23306 7568 -23242
rect 7632 -23306 7888 -23242
rect 7952 -23306 8208 -23242
rect 8272 -23306 8528 -23242
rect 8592 -23306 8848 -23242
rect 8912 -23306 9168 -23242
rect 9232 -23306 9488 -23242
rect 9552 -23306 9808 -23242
rect 9872 -23306 10128 -23242
rect 10192 -23306 10448 -23242
rect 10512 -23306 10768 -23242
rect 10832 -23306 11088 -23242
rect 11152 -23306 11408 -23242
rect 11472 -23306 11728 -23242
rect 11792 -23306 12048 -23242
rect 12112 -23306 12368 -23242
rect 12432 -23306 12688 -23242
rect 12752 -23306 13008 -23242
rect 13072 -23306 13328 -23242
rect 13392 -23306 14000 -23242
rect 6000 -23448 14000 -23306
rect 6000 -23512 6238 -23448
rect 6302 -23512 13704 -23448
rect 13768 -23512 14000 -23448
rect 6000 -23540 14000 -23512
rect 6000 -23768 6540 -23540
rect 6000 -23832 6238 -23768
rect 6302 -23832 6540 -23768
rect 6000 -24088 6540 -23832
rect 6000 -24152 6238 -24088
rect 6302 -24152 6540 -24088
rect 6000 -24408 6540 -24152
rect 6000 -24472 6238 -24408
rect 6302 -24472 6540 -24408
rect 6000 -24728 6540 -24472
rect 6000 -24792 6238 -24728
rect 6302 -24792 6540 -24728
rect 6000 -25048 6540 -24792
rect 6000 -25112 6238 -25048
rect 6302 -25112 6540 -25048
rect 6000 -25368 6540 -25112
rect 6000 -25432 6238 -25368
rect 6302 -25432 6540 -25368
rect 6000 -25688 6540 -25432
rect 6000 -25752 6238 -25688
rect 6302 -25752 6540 -25688
rect 6000 -26008 6540 -25752
rect 6000 -26072 6238 -26008
rect 6302 -26072 6540 -26008
rect 6000 -26328 6540 -26072
rect 6000 -26392 6238 -26328
rect 6302 -26392 6540 -26328
rect 6000 -26648 6540 -26392
rect 6000 -26712 6238 -26648
rect 6302 -26712 6540 -26648
rect 6000 -26968 6540 -26712
rect 6000 -27032 6238 -26968
rect 6302 -27032 6540 -26968
rect 6000 -27288 6540 -27032
rect 6000 -27352 6238 -27288
rect 6302 -27352 6540 -27288
rect 6000 -27608 6540 -27352
rect 6000 -27672 6238 -27608
rect 6302 -27672 6540 -27608
rect 6000 -27928 6540 -27672
rect 6000 -27992 6238 -27928
rect 6302 -27992 6540 -27928
rect 6000 -28248 6540 -27992
rect 6000 -28312 6238 -28248
rect 6302 -28312 6540 -28248
rect 6000 -28568 6540 -28312
rect 6000 -28632 6238 -28568
rect 6302 -28632 6540 -28568
rect 6000 -28888 6540 -28632
rect 6000 -28952 6238 -28888
rect 6302 -28952 6540 -28888
rect 6000 -29208 6540 -28952
rect 6000 -29272 6238 -29208
rect 6302 -29272 6540 -29208
rect 6000 -29528 6540 -29272
rect 6000 -29592 6238 -29528
rect 6302 -29592 6540 -29528
rect 6000 -29848 6540 -29592
rect 6000 -29912 6238 -29848
rect 6302 -29912 6540 -29848
rect 6000 -30168 6540 -29912
rect 6000 -30232 6238 -30168
rect 6302 -30232 6540 -30168
rect 6000 -30460 6540 -30232
rect 13460 -23768 14000 -23540
rect 13460 -23832 13704 -23768
rect 13768 -23832 14000 -23768
rect 13460 -24088 14000 -23832
rect 13460 -24152 13704 -24088
rect 13768 -24152 14000 -24088
rect 13460 -24408 14000 -24152
rect 13460 -24472 13704 -24408
rect 13768 -24472 14000 -24408
rect 13460 -24728 14000 -24472
rect 13460 -24792 13704 -24728
rect 13768 -24792 14000 -24728
rect 13460 -25048 14000 -24792
rect 13460 -25112 13704 -25048
rect 13768 -25112 14000 -25048
rect 13460 -25368 14000 -25112
rect 13460 -25432 13704 -25368
rect 13768 -25432 14000 -25368
rect 13460 -25688 14000 -25432
rect 13460 -25752 13704 -25688
rect 13768 -25740 14000 -25688
rect 16330 -25740 16390 -9590
rect 13768 -25752 16390 -25740
rect 13460 -25800 16390 -25752
rect 16460 -9660 16540 -9650
rect 16460 -9720 16470 -9660
rect 16530 -9720 16540 -9660
rect 16460 -9730 16540 -9720
rect 16460 -25750 16520 -9730
rect 16600 -10610 16660 -9580
rect 17600 -9600 19000 -9500
rect 17600 -10200 17700 -9600
rect 18900 -10200 19000 -9600
rect 17600 -10300 19000 -10200
rect 20800 -9600 22200 -9500
rect 20800 -10200 20900 -9600
rect 22100 -10200 22200 -9600
rect 20800 -10300 22200 -10200
rect 16600 -10620 17140 -10610
rect 16600 -10740 17040 -10620
rect 17120 -10740 17140 -10620
rect 16600 -10750 17140 -10740
rect 16600 -22660 16660 -10750
rect 24120 -10800 24200 -7870
rect 24330 -10600 24410 -7550
rect 24330 -10680 26680 -10600
rect 24120 -10880 26480 -10800
rect 18000 -11242 26000 -11000
rect 18000 -11306 18608 -11242
rect 18672 -11306 18928 -11242
rect 18992 -11306 19248 -11242
rect 19312 -11306 19568 -11242
rect 19632 -11306 19888 -11242
rect 19952 -11306 20208 -11242
rect 20272 -11306 20528 -11242
rect 20592 -11306 20848 -11242
rect 20912 -11306 21168 -11242
rect 21232 -11306 21488 -11242
rect 21552 -11306 21808 -11242
rect 21872 -11306 22128 -11242
rect 22192 -11306 22448 -11242
rect 22512 -11306 22768 -11242
rect 22832 -11306 23088 -11242
rect 23152 -11306 23408 -11242
rect 23472 -11306 23728 -11242
rect 23792 -11306 24048 -11242
rect 24112 -11306 24368 -11242
rect 24432 -11306 24688 -11242
rect 24752 -11306 25008 -11242
rect 25072 -11306 25328 -11242
rect 25392 -11306 26000 -11242
rect 18000 -11448 26000 -11306
rect 18000 -11512 18238 -11448
rect 18302 -11512 25704 -11448
rect 25768 -11512 26000 -11448
rect 18000 -11540 26000 -11512
rect 18000 -11768 18540 -11540
rect 18000 -11832 18238 -11768
rect 18302 -11832 18540 -11768
rect 18000 -12088 18540 -11832
rect 18000 -12152 18238 -12088
rect 18302 -12152 18540 -12088
rect 18000 -12408 18540 -12152
rect 18000 -12472 18238 -12408
rect 18302 -12472 18540 -12408
rect 18000 -12728 18540 -12472
rect 18000 -12792 18238 -12728
rect 18302 -12792 18540 -12728
rect 18000 -13048 18540 -12792
rect 18000 -13112 18238 -13048
rect 18302 -13112 18540 -13048
rect 18000 -13368 18540 -13112
rect 18000 -13432 18238 -13368
rect 18302 -13432 18540 -13368
rect 18000 -13688 18540 -13432
rect 18000 -13752 18238 -13688
rect 18302 -13752 18540 -13688
rect 18000 -14008 18540 -13752
rect 18000 -14072 18238 -14008
rect 18302 -14072 18540 -14008
rect 18000 -14328 18540 -14072
rect 18000 -14392 18238 -14328
rect 18302 -14392 18540 -14328
rect 18000 -14648 18540 -14392
rect 18000 -14712 18238 -14648
rect 18302 -14712 18540 -14648
rect 18000 -14968 18540 -14712
rect 18000 -15032 18238 -14968
rect 18302 -15032 18540 -14968
rect 18000 -15288 18540 -15032
rect 18000 -15352 18238 -15288
rect 18302 -15352 18540 -15288
rect 18000 -15608 18540 -15352
rect 18000 -15672 18238 -15608
rect 18302 -15672 18540 -15608
rect 18000 -15928 18540 -15672
rect 18000 -15992 18238 -15928
rect 18302 -15992 18540 -15928
rect 18000 -16248 18540 -15992
rect 18000 -16312 18238 -16248
rect 18302 -16312 18540 -16248
rect 18000 -16568 18540 -16312
rect 18000 -16632 18238 -16568
rect 18302 -16632 18540 -16568
rect 18000 -16888 18540 -16632
rect 18000 -16952 18238 -16888
rect 18302 -16952 18540 -16888
rect 18000 -17208 18540 -16952
rect 18000 -17272 18238 -17208
rect 18302 -17272 18540 -17208
rect 18000 -17528 18540 -17272
rect 18000 -17592 18238 -17528
rect 18302 -17592 18540 -17528
rect 18000 -17848 18540 -17592
rect 18000 -17912 18238 -17848
rect 18302 -17912 18540 -17848
rect 18000 -18168 18540 -17912
rect 18000 -18232 18238 -18168
rect 18302 -18232 18540 -18168
rect 18000 -18460 18540 -18232
rect 25460 -11768 26000 -11540
rect 25460 -11832 25704 -11768
rect 25768 -11832 26000 -11768
rect 25460 -12088 26000 -11832
rect 25460 -12152 25704 -12088
rect 25768 -12152 26000 -12088
rect 25460 -12408 26000 -12152
rect 25460 -12472 25704 -12408
rect 25768 -12472 26000 -12408
rect 25460 -12728 26000 -12472
rect 25460 -12792 25704 -12728
rect 25768 -12792 26000 -12728
rect 25460 -13048 26000 -12792
rect 25460 -13112 25704 -13048
rect 25768 -13112 26000 -13048
rect 25460 -13368 26000 -13112
rect 25460 -13432 25704 -13368
rect 25768 -13432 26000 -13368
rect 25460 -13688 26000 -13432
rect 25460 -13752 25704 -13688
rect 25768 -13752 26000 -13688
rect 25460 -14008 26000 -13752
rect 25460 -14072 25704 -14008
rect 25768 -14072 26000 -14008
rect 25460 -14328 26000 -14072
rect 25460 -14392 25704 -14328
rect 25768 -14392 26000 -14328
rect 25460 -14648 26000 -14392
rect 25460 -14712 25704 -14648
rect 25768 -14712 26000 -14648
rect 25460 -14968 26000 -14712
rect 25460 -15032 25704 -14968
rect 25768 -15032 26000 -14968
rect 25460 -15288 26000 -15032
rect 25460 -15352 25704 -15288
rect 25768 -15352 26000 -15288
rect 25460 -15608 26000 -15352
rect 25460 -15672 25704 -15608
rect 25768 -15672 26000 -15608
rect 26400 -15590 26480 -10880
rect 26600 -15350 26680 -10680
rect 30000 -11242 38000 -11000
rect 30000 -11306 30608 -11242
rect 30672 -11306 30928 -11242
rect 30992 -11306 31248 -11242
rect 31312 -11306 31568 -11242
rect 31632 -11306 31888 -11242
rect 31952 -11306 32208 -11242
rect 32272 -11306 32528 -11242
rect 32592 -11306 32848 -11242
rect 32912 -11306 33168 -11242
rect 33232 -11306 33488 -11242
rect 33552 -11306 33808 -11242
rect 33872 -11306 34128 -11242
rect 34192 -11306 34448 -11242
rect 34512 -11306 34768 -11242
rect 34832 -11306 35088 -11242
rect 35152 -11306 35408 -11242
rect 35472 -11306 35728 -11242
rect 35792 -11306 36048 -11242
rect 36112 -11306 36368 -11242
rect 36432 -11306 36688 -11242
rect 36752 -11306 37008 -11242
rect 37072 -11306 37328 -11242
rect 37392 -11306 38000 -11242
rect 30000 -11448 38000 -11306
rect 30000 -11512 30238 -11448
rect 30302 -11512 37704 -11448
rect 37768 -11512 38000 -11448
rect 30000 -11540 38000 -11512
rect 30000 -11768 30540 -11540
rect 30000 -11832 30238 -11768
rect 30302 -11832 30540 -11768
rect 30000 -12088 30540 -11832
rect 30000 -12152 30238 -12088
rect 30302 -12152 30540 -12088
rect 30000 -12408 30540 -12152
rect 30000 -12472 30238 -12408
rect 30302 -12472 30540 -12408
rect 30000 -12728 30540 -12472
rect 30000 -12792 30238 -12728
rect 30302 -12792 30540 -12728
rect 30000 -13048 30540 -12792
rect 30000 -13112 30238 -13048
rect 30302 -13112 30540 -13048
rect 30000 -13368 30540 -13112
rect 30000 -13432 30238 -13368
rect 30302 -13432 30540 -13368
rect 30000 -13688 30540 -13432
rect 30000 -13752 30238 -13688
rect 30302 -13752 30540 -13688
rect 30000 -14008 30540 -13752
rect 30000 -14072 30238 -14008
rect 30302 -14072 30540 -14008
rect 30000 -14328 30540 -14072
rect 30000 -14392 30238 -14328
rect 30302 -14392 30540 -14328
rect 30000 -14648 30540 -14392
rect 30000 -14712 30238 -14648
rect 30302 -14712 30540 -14648
rect 30000 -14968 30540 -14712
rect 30000 -15032 30238 -14968
rect 30302 -15032 30540 -14968
rect 30000 -15288 30540 -15032
rect 30000 -15350 30238 -15288
rect 26600 -15352 30238 -15350
rect 30302 -15352 30540 -15288
rect 26600 -15430 30540 -15352
rect 26400 -15670 29170 -15590
rect 25460 -15928 26000 -15672
rect 25460 -15992 25704 -15928
rect 25768 -15992 26000 -15928
rect 25460 -16248 26000 -15992
rect 25460 -16312 25704 -16248
rect 25768 -16312 26000 -16248
rect 25460 -16568 26000 -16312
rect 25460 -16632 25704 -16568
rect 25768 -16632 26000 -16568
rect 25460 -16888 26000 -16632
rect 25460 -16952 25704 -16888
rect 25768 -16952 26000 -16888
rect 25460 -17208 26000 -16952
rect 25460 -17272 25704 -17208
rect 25768 -17272 26000 -17208
rect 25460 -17528 26000 -17272
rect 25460 -17592 25704 -17528
rect 25768 -17592 26000 -17528
rect 25460 -17848 26000 -17592
rect 25460 -17912 25704 -17848
rect 25768 -17912 26000 -17848
rect 25460 -18168 26000 -17912
rect 25460 -18232 25704 -18168
rect 25768 -18232 26000 -18168
rect 25460 -18460 26000 -18232
rect 18000 -18488 26000 -18460
rect 18000 -18552 18238 -18488
rect 18302 -18552 25704 -18488
rect 25768 -18552 26000 -18488
rect 18000 -18698 26000 -18552
rect 18000 -18762 18608 -18698
rect 18672 -18762 18928 -18698
rect 18992 -18762 19248 -18698
rect 19312 -18762 19568 -18698
rect 19632 -18762 19888 -18698
rect 19952 -18762 20208 -18698
rect 20272 -18762 20528 -18698
rect 20592 -18762 20848 -18698
rect 20912 -18762 21168 -18698
rect 21232 -18762 21488 -18698
rect 21552 -18762 21808 -18698
rect 21872 -18762 22128 -18698
rect 22192 -18762 22448 -18698
rect 22512 -18762 22768 -18698
rect 22832 -18762 23088 -18698
rect 23152 -18762 23408 -18698
rect 23472 -18762 23728 -18698
rect 23792 -18762 24048 -18698
rect 24112 -18762 24368 -18698
rect 24432 -18762 24688 -18698
rect 24752 -18762 25008 -18698
rect 25072 -18762 25328 -18698
rect 25392 -18762 26000 -18698
rect 18000 -19000 26000 -18762
rect 29090 -22240 29170 -15670
rect 30000 -15608 30540 -15430
rect 30000 -15672 30238 -15608
rect 30302 -15672 30540 -15608
rect 30000 -15928 30540 -15672
rect 30000 -15992 30238 -15928
rect 30302 -15992 30540 -15928
rect 30000 -16248 30540 -15992
rect 30000 -16312 30238 -16248
rect 30302 -16312 30540 -16248
rect 30000 -16568 30540 -16312
rect 30000 -16632 30238 -16568
rect 30302 -16632 30540 -16568
rect 30000 -16888 30540 -16632
rect 30000 -16952 30238 -16888
rect 30302 -16952 30540 -16888
rect 30000 -17208 30540 -16952
rect 30000 -17272 30238 -17208
rect 30302 -17272 30540 -17208
rect 30000 -17528 30540 -17272
rect 30000 -17592 30238 -17528
rect 30302 -17592 30540 -17528
rect 30000 -17848 30540 -17592
rect 30000 -17912 30238 -17848
rect 30302 -17912 30540 -17848
rect 30000 -18168 30540 -17912
rect 30000 -18232 30238 -18168
rect 30302 -18232 30540 -18168
rect 30000 -18460 30540 -18232
rect 37460 -11768 38000 -11540
rect 37460 -11832 37704 -11768
rect 37768 -11832 38000 -11768
rect 37460 -12088 38000 -11832
rect 37460 -12152 37704 -12088
rect 37768 -12152 38000 -12088
rect 37460 -12408 38000 -12152
rect 37460 -12472 37704 -12408
rect 37768 -12472 38000 -12408
rect 37460 -12728 38000 -12472
rect 37460 -12792 37704 -12728
rect 37768 -12792 38000 -12728
rect 37460 -13048 38000 -12792
rect 37460 -13112 37704 -13048
rect 37768 -13112 38000 -13048
rect 37460 -13368 38000 -13112
rect 37460 -13432 37704 -13368
rect 37768 -13432 38000 -13368
rect 37460 -13688 38000 -13432
rect 37460 -13752 37704 -13688
rect 37768 -13752 38000 -13688
rect 37460 -14008 38000 -13752
rect 37460 -14072 37704 -14008
rect 37768 -14072 38000 -14008
rect 37460 -14328 38000 -14072
rect 37460 -14392 37704 -14328
rect 37768 -14392 38000 -14328
rect 37460 -14648 38000 -14392
rect 37460 -14712 37704 -14648
rect 37768 -14712 38000 -14648
rect 37460 -14968 38000 -14712
rect 37460 -15032 37704 -14968
rect 37768 -15032 38000 -14968
rect 37460 -15288 38000 -15032
rect 37460 -15352 37704 -15288
rect 37768 -15352 38000 -15288
rect 37460 -15608 38000 -15352
rect 37460 -15672 37704 -15608
rect 37768 -15672 38000 -15608
rect 37460 -15928 38000 -15672
rect 37460 -15992 37704 -15928
rect 37768 -15992 38000 -15928
rect 37460 -16248 38000 -15992
rect 37460 -16312 37704 -16248
rect 37768 -16312 38000 -16248
rect 37460 -16568 38000 -16312
rect 37460 -16632 37704 -16568
rect 37768 -16632 38000 -16568
rect 37460 -16888 38000 -16632
rect 37460 -16952 37704 -16888
rect 37768 -16952 38000 -16888
rect 37460 -17208 38000 -16952
rect 37460 -17272 37704 -17208
rect 37768 -17272 38000 -17208
rect 37460 -17528 38000 -17272
rect 37460 -17592 37704 -17528
rect 37768 -17592 38000 -17528
rect 37460 -17848 38000 -17592
rect 37460 -17912 37704 -17848
rect 37768 -17912 38000 -17848
rect 37460 -18168 38000 -17912
rect 37460 -18232 37704 -18168
rect 37768 -18232 38000 -18168
rect 37460 -18460 38000 -18232
rect 30000 -18488 38000 -18460
rect 30000 -18552 30238 -18488
rect 30302 -18552 37704 -18488
rect 37768 -18552 38000 -18488
rect 30000 -18698 38000 -18552
rect 30000 -18762 30608 -18698
rect 30672 -18762 30928 -18698
rect 30992 -18762 31248 -18698
rect 31312 -18762 31568 -18698
rect 31632 -18762 31888 -18698
rect 31952 -18762 32208 -18698
rect 32272 -18762 32528 -18698
rect 32592 -18762 32848 -18698
rect 32912 -18762 33168 -18698
rect 33232 -18762 33488 -18698
rect 33552 -18762 33808 -18698
rect 33872 -18762 34128 -18698
rect 34192 -18762 34448 -18698
rect 34512 -18762 34768 -18698
rect 34832 -18762 35088 -18698
rect 35152 -18762 35408 -18698
rect 35472 -18762 35728 -18698
rect 35792 -18762 36048 -18698
rect 36112 -18762 36368 -18698
rect 36432 -18762 36688 -18698
rect 36752 -18762 37008 -18698
rect 37072 -18762 37328 -18698
rect 37392 -18762 38000 -18698
rect 30000 -19000 38000 -18762
rect 42000 -11242 50000 -11000
rect 42000 -11306 42608 -11242
rect 42672 -11306 42928 -11242
rect 42992 -11306 43248 -11242
rect 43312 -11306 43568 -11242
rect 43632 -11306 43888 -11242
rect 43952 -11306 44208 -11242
rect 44272 -11306 44528 -11242
rect 44592 -11306 44848 -11242
rect 44912 -11306 45168 -11242
rect 45232 -11306 45488 -11242
rect 45552 -11306 45808 -11242
rect 45872 -11306 46128 -11242
rect 46192 -11306 46448 -11242
rect 46512 -11306 46768 -11242
rect 46832 -11306 47088 -11242
rect 47152 -11306 47408 -11242
rect 47472 -11306 47728 -11242
rect 47792 -11306 48048 -11242
rect 48112 -11306 48368 -11242
rect 48432 -11306 48688 -11242
rect 48752 -11306 49008 -11242
rect 49072 -11306 49328 -11242
rect 49392 -11306 50000 -11242
rect 42000 -11448 50000 -11306
rect 42000 -11512 42238 -11448
rect 42302 -11512 49704 -11448
rect 49768 -11512 50000 -11448
rect 42000 -11540 50000 -11512
rect 42000 -11768 42540 -11540
rect 42000 -11832 42238 -11768
rect 42302 -11832 42540 -11768
rect 42000 -12088 42540 -11832
rect 42000 -12152 42238 -12088
rect 42302 -12152 42540 -12088
rect 42000 -12408 42540 -12152
rect 42000 -12472 42238 -12408
rect 42302 -12472 42540 -12408
rect 42000 -12728 42540 -12472
rect 42000 -12792 42238 -12728
rect 42302 -12792 42540 -12728
rect 42000 -13048 42540 -12792
rect 42000 -13112 42238 -13048
rect 42302 -13112 42540 -13048
rect 42000 -13368 42540 -13112
rect 42000 -13432 42238 -13368
rect 42302 -13432 42540 -13368
rect 42000 -13688 42540 -13432
rect 42000 -13752 42238 -13688
rect 42302 -13752 42540 -13688
rect 42000 -14008 42540 -13752
rect 42000 -14072 42238 -14008
rect 42302 -14072 42540 -14008
rect 42000 -14328 42540 -14072
rect 42000 -14392 42238 -14328
rect 42302 -14392 42540 -14328
rect 42000 -14648 42540 -14392
rect 42000 -14712 42238 -14648
rect 42302 -14712 42540 -14648
rect 42000 -14968 42540 -14712
rect 42000 -15032 42238 -14968
rect 42302 -15032 42540 -14968
rect 42000 -15288 42540 -15032
rect 42000 -15352 42238 -15288
rect 42302 -15352 42540 -15288
rect 42000 -15608 42540 -15352
rect 42000 -15672 42238 -15608
rect 42302 -15672 42540 -15608
rect 42000 -15928 42540 -15672
rect 42000 -15992 42238 -15928
rect 42302 -15992 42540 -15928
rect 42000 -16248 42540 -15992
rect 42000 -16312 42238 -16248
rect 42302 -16312 42540 -16248
rect 42000 -16568 42540 -16312
rect 42000 -16632 42238 -16568
rect 42302 -16632 42540 -16568
rect 42000 -16888 42540 -16632
rect 42000 -16952 42238 -16888
rect 42302 -16952 42540 -16888
rect 42000 -17208 42540 -16952
rect 42000 -17272 42238 -17208
rect 42302 -17272 42540 -17208
rect 42000 -17528 42540 -17272
rect 42000 -17592 42238 -17528
rect 42302 -17592 42540 -17528
rect 42000 -17848 42540 -17592
rect 42000 -17912 42238 -17848
rect 42302 -17912 42540 -17848
rect 42000 -18168 42540 -17912
rect 42000 -18232 42238 -18168
rect 42302 -18232 42540 -18168
rect 42000 -18460 42540 -18232
rect 49460 -11768 50000 -11540
rect 49460 -11832 49704 -11768
rect 49768 -11832 50000 -11768
rect 49460 -12088 50000 -11832
rect 49460 -12152 49704 -12088
rect 49768 -12152 50000 -12088
rect 49460 -12408 50000 -12152
rect 49460 -12472 49704 -12408
rect 49768 -12472 50000 -12408
rect 49460 -12728 50000 -12472
rect 49460 -12792 49704 -12728
rect 49768 -12792 50000 -12728
rect 49460 -13048 50000 -12792
rect 49460 -13112 49704 -13048
rect 49768 -13112 50000 -13048
rect 49460 -13368 50000 -13112
rect 49460 -13432 49704 -13368
rect 49768 -13432 50000 -13368
rect 49460 -13688 50000 -13432
rect 49460 -13752 49704 -13688
rect 49768 -13752 50000 -13688
rect 49460 -14008 50000 -13752
rect 49460 -14072 49704 -14008
rect 49768 -14072 50000 -14008
rect 49460 -14328 50000 -14072
rect 49460 -14392 49704 -14328
rect 49768 -14392 50000 -14328
rect 49460 -14648 50000 -14392
rect 49460 -14712 49704 -14648
rect 49768 -14712 50000 -14648
rect 49460 -14968 50000 -14712
rect 49460 -15032 49704 -14968
rect 49768 -15032 50000 -14968
rect 49460 -15288 50000 -15032
rect 49460 -15352 49704 -15288
rect 49768 -15352 50000 -15288
rect 49460 -15608 50000 -15352
rect 49460 -15672 49704 -15608
rect 49768 -15672 50000 -15608
rect 49460 -15928 50000 -15672
rect 49460 -15992 49704 -15928
rect 49768 -15992 50000 -15928
rect 49460 -16248 50000 -15992
rect 49460 -16312 49704 -16248
rect 49768 -16312 50000 -16248
rect 49460 -16568 50000 -16312
rect 49460 -16632 49704 -16568
rect 49768 -16632 50000 -16568
rect 49460 -16888 50000 -16632
rect 49460 -16952 49704 -16888
rect 49768 -16952 50000 -16888
rect 49460 -17208 50000 -16952
rect 49460 -17272 49704 -17208
rect 49768 -17272 50000 -17208
rect 49460 -17528 50000 -17272
rect 49460 -17592 49704 -17528
rect 49768 -17592 50000 -17528
rect 49460 -17848 50000 -17592
rect 49460 -17912 49704 -17848
rect 49768 -17912 50000 -17848
rect 49460 -18168 50000 -17912
rect 49460 -18232 49704 -18168
rect 49768 -18232 50000 -18168
rect 49460 -18460 50000 -18232
rect 42000 -18488 50000 -18460
rect 42000 -18552 42238 -18488
rect 42302 -18552 49704 -18488
rect 49768 -18552 50000 -18488
rect 42000 -18698 50000 -18552
rect 42000 -18762 42608 -18698
rect 42672 -18762 42928 -18698
rect 42992 -18762 43248 -18698
rect 43312 -18762 43568 -18698
rect 43632 -18762 43888 -18698
rect 43952 -18762 44208 -18698
rect 44272 -18762 44528 -18698
rect 44592 -18762 44848 -18698
rect 44912 -18762 45168 -18698
rect 45232 -18762 45488 -18698
rect 45552 -18762 45808 -18698
rect 45872 -18762 46128 -18698
rect 46192 -18762 46448 -18698
rect 46512 -18762 46768 -18698
rect 46832 -18762 47088 -18698
rect 47152 -18762 47408 -18698
rect 47472 -18762 47728 -18698
rect 47792 -18762 48048 -18698
rect 48112 -18762 48368 -18698
rect 48432 -18762 48688 -18698
rect 48752 -18762 49008 -18698
rect 49072 -18762 49328 -18698
rect 49392 -18762 50000 -18698
rect 42000 -19000 50000 -18762
rect 29090 -22320 42750 -22240
rect 16600 -22720 28300 -22660
rect 18000 -23242 26000 -23000
rect 18000 -23306 18608 -23242
rect 18672 -23306 18928 -23242
rect 18992 -23306 19248 -23242
rect 19312 -23306 19568 -23242
rect 19632 -23306 19888 -23242
rect 19952 -23306 20208 -23242
rect 20272 -23306 20528 -23242
rect 20592 -23306 20848 -23242
rect 20912 -23306 21168 -23242
rect 21232 -23306 21488 -23242
rect 21552 -23306 21808 -23242
rect 21872 -23306 22128 -23242
rect 22192 -23306 22448 -23242
rect 22512 -23306 22768 -23242
rect 22832 -23306 23088 -23242
rect 23152 -23306 23408 -23242
rect 23472 -23306 23728 -23242
rect 23792 -23306 24048 -23242
rect 24112 -23306 24368 -23242
rect 24432 -23306 24688 -23242
rect 24752 -23306 25008 -23242
rect 25072 -23306 25328 -23242
rect 25392 -23306 26000 -23242
rect 18000 -23448 26000 -23306
rect 18000 -23512 18238 -23448
rect 18302 -23512 25704 -23448
rect 25768 -23512 26000 -23448
rect 18000 -23540 26000 -23512
rect 18000 -23768 18540 -23540
rect 18000 -23832 18238 -23768
rect 18302 -23832 18540 -23768
rect 18000 -24088 18540 -23832
rect 18000 -24152 18238 -24088
rect 18302 -24152 18540 -24088
rect 18000 -24408 18540 -24152
rect 18000 -24472 18238 -24408
rect 18302 -24472 18540 -24408
rect 18000 -24728 18540 -24472
rect 18000 -24792 18238 -24728
rect 18302 -24792 18540 -24728
rect 18000 -25048 18540 -24792
rect 18000 -25112 18238 -25048
rect 18302 -25112 18540 -25048
rect 18000 -25368 18540 -25112
rect 18000 -25432 18238 -25368
rect 18302 -25432 18540 -25368
rect 18000 -25688 18540 -25432
rect 18000 -25750 18238 -25688
rect 16460 -25752 18238 -25750
rect 18302 -25752 18540 -25688
rect 13460 -26008 14000 -25800
rect 16460 -25810 18540 -25752
rect 13460 -26072 13704 -26008
rect 13768 -26072 14000 -26008
rect 13460 -26328 14000 -26072
rect 13460 -26392 13704 -26328
rect 13768 -26392 14000 -26328
rect 13460 -26648 14000 -26392
rect 13460 -26712 13704 -26648
rect 13768 -26712 14000 -26648
rect 13460 -26968 14000 -26712
rect 13460 -27032 13704 -26968
rect 13768 -27032 14000 -26968
rect 13460 -27288 14000 -27032
rect 13460 -27352 13704 -27288
rect 13768 -27352 14000 -27288
rect 13460 -27608 14000 -27352
rect 13460 -27672 13704 -27608
rect 13768 -27672 14000 -27608
rect 13460 -27928 14000 -27672
rect 13460 -27992 13704 -27928
rect 13768 -27992 14000 -27928
rect 13460 -28248 14000 -27992
rect 13460 -28312 13704 -28248
rect 13768 -28312 14000 -28248
rect 13460 -28568 14000 -28312
rect 13460 -28632 13704 -28568
rect 13768 -28632 14000 -28568
rect 13460 -28888 14000 -28632
rect 13460 -28952 13704 -28888
rect 13768 -28952 14000 -28888
rect 13460 -29208 14000 -28952
rect 13460 -29272 13704 -29208
rect 13768 -29272 14000 -29208
rect 13460 -29528 14000 -29272
rect 13460 -29592 13704 -29528
rect 13768 -29592 14000 -29528
rect 13460 -29848 14000 -29592
rect 13460 -29912 13704 -29848
rect 13768 -29912 14000 -29848
rect 13460 -30168 14000 -29912
rect 13460 -30232 13704 -30168
rect 13768 -30232 14000 -30168
rect 13460 -30460 14000 -30232
rect 6000 -30488 14000 -30460
rect 6000 -30552 6238 -30488
rect 6302 -30552 13704 -30488
rect 13768 -30552 14000 -30488
rect 6000 -30698 14000 -30552
rect 6000 -30762 6608 -30698
rect 6672 -30762 6928 -30698
rect 6992 -30762 7248 -30698
rect 7312 -30762 7568 -30698
rect 7632 -30762 7888 -30698
rect 7952 -30762 8208 -30698
rect 8272 -30762 8528 -30698
rect 8592 -30762 8848 -30698
rect 8912 -30762 9168 -30698
rect 9232 -30762 9488 -30698
rect 9552 -30762 9808 -30698
rect 9872 -30762 10128 -30698
rect 10192 -30762 10448 -30698
rect 10512 -30762 10768 -30698
rect 10832 -30762 11088 -30698
rect 11152 -30762 11408 -30698
rect 11472 -30762 11728 -30698
rect 11792 -30762 12048 -30698
rect 12112 -30762 12368 -30698
rect 12432 -30762 12688 -30698
rect 12752 -30762 13008 -30698
rect 13072 -30762 13328 -30698
rect 13392 -30762 14000 -30698
rect 6000 -31000 14000 -30762
rect 18000 -26008 18540 -25810
rect 18000 -26072 18238 -26008
rect 18302 -26072 18540 -26008
rect 18000 -26328 18540 -26072
rect 18000 -26392 18238 -26328
rect 18302 -26392 18540 -26328
rect 18000 -26648 18540 -26392
rect 18000 -26712 18238 -26648
rect 18302 -26712 18540 -26648
rect 18000 -26968 18540 -26712
rect 18000 -27032 18238 -26968
rect 18302 -27032 18540 -26968
rect 18000 -27288 18540 -27032
rect 18000 -27352 18238 -27288
rect 18302 -27352 18540 -27288
rect 18000 -27608 18540 -27352
rect 18000 -27672 18238 -27608
rect 18302 -27672 18540 -27608
rect 18000 -27928 18540 -27672
rect 18000 -27992 18238 -27928
rect 18302 -27992 18540 -27928
rect 18000 -28248 18540 -27992
rect 18000 -28312 18238 -28248
rect 18302 -28312 18540 -28248
rect 18000 -28568 18540 -28312
rect 18000 -28632 18238 -28568
rect 18302 -28632 18540 -28568
rect 18000 -28888 18540 -28632
rect 18000 -28952 18238 -28888
rect 18302 -28952 18540 -28888
rect 18000 -29208 18540 -28952
rect 18000 -29272 18238 -29208
rect 18302 -29272 18540 -29208
rect 18000 -29528 18540 -29272
rect 18000 -29592 18238 -29528
rect 18302 -29592 18540 -29528
rect 18000 -29848 18540 -29592
rect 18000 -29912 18238 -29848
rect 18302 -29912 18540 -29848
rect 18000 -30168 18540 -29912
rect 18000 -30232 18238 -30168
rect 18302 -30232 18540 -30168
rect 18000 -30460 18540 -30232
rect 25460 -23768 26000 -23540
rect 25460 -23832 25704 -23768
rect 25768 -23832 26000 -23768
rect 25460 -24088 26000 -23832
rect 25460 -24152 25704 -24088
rect 25768 -24152 26000 -24088
rect 25460 -24408 26000 -24152
rect 25460 -24472 25704 -24408
rect 25768 -24472 26000 -24408
rect 25460 -24728 26000 -24472
rect 25460 -24792 25704 -24728
rect 25768 -24792 26000 -24728
rect 25460 -25048 26000 -24792
rect 25460 -25112 25704 -25048
rect 25768 -25112 26000 -25048
rect 25460 -25368 26000 -25112
rect 25460 -25432 25704 -25368
rect 25768 -25432 26000 -25368
rect 25460 -25688 26000 -25432
rect 25460 -25752 25704 -25688
rect 25768 -25752 26000 -25688
rect 25460 -26008 26000 -25752
rect 28240 -25740 28300 -22720
rect 42670 -23000 42750 -22320
rect 30000 -23242 38000 -23000
rect 30000 -23306 30608 -23242
rect 30672 -23306 30928 -23242
rect 30992 -23306 31248 -23242
rect 31312 -23306 31568 -23242
rect 31632 -23306 31888 -23242
rect 31952 -23306 32208 -23242
rect 32272 -23306 32528 -23242
rect 32592 -23306 32848 -23242
rect 32912 -23306 33168 -23242
rect 33232 -23306 33488 -23242
rect 33552 -23306 33808 -23242
rect 33872 -23306 34128 -23242
rect 34192 -23306 34448 -23242
rect 34512 -23306 34768 -23242
rect 34832 -23306 35088 -23242
rect 35152 -23306 35408 -23242
rect 35472 -23306 35728 -23242
rect 35792 -23306 36048 -23242
rect 36112 -23306 36368 -23242
rect 36432 -23306 36688 -23242
rect 36752 -23306 37008 -23242
rect 37072 -23306 37328 -23242
rect 37392 -23306 38000 -23242
rect 30000 -23448 38000 -23306
rect 30000 -23512 30238 -23448
rect 30302 -23512 37704 -23448
rect 37768 -23512 38000 -23448
rect 30000 -23540 38000 -23512
rect 30000 -23768 30540 -23540
rect 30000 -23832 30238 -23768
rect 30302 -23832 30540 -23768
rect 30000 -24088 30540 -23832
rect 30000 -24152 30238 -24088
rect 30302 -24152 30540 -24088
rect 30000 -24408 30540 -24152
rect 30000 -24472 30238 -24408
rect 30302 -24472 30540 -24408
rect 30000 -24728 30540 -24472
rect 30000 -24792 30238 -24728
rect 30302 -24792 30540 -24728
rect 30000 -25048 30540 -24792
rect 30000 -25112 30238 -25048
rect 30302 -25112 30540 -25048
rect 30000 -25368 30540 -25112
rect 30000 -25432 30238 -25368
rect 30302 -25432 30540 -25368
rect 30000 -25688 30540 -25432
rect 30000 -25740 30238 -25688
rect 28240 -25752 30238 -25740
rect 30302 -25752 30540 -25688
rect 28240 -25800 30540 -25752
rect 25460 -26072 25704 -26008
rect 25768 -26072 26000 -26008
rect 25460 -26328 26000 -26072
rect 25460 -26392 25704 -26328
rect 25768 -26392 26000 -26328
rect 25460 -26648 26000 -26392
rect 25460 -26712 25704 -26648
rect 25768 -26712 26000 -26648
rect 25460 -26968 26000 -26712
rect 25460 -27032 25704 -26968
rect 25768 -27032 26000 -26968
rect 25460 -27288 26000 -27032
rect 25460 -27352 25704 -27288
rect 25768 -27352 26000 -27288
rect 25460 -27608 26000 -27352
rect 25460 -27672 25704 -27608
rect 25768 -27672 26000 -27608
rect 25460 -27928 26000 -27672
rect 25460 -27992 25704 -27928
rect 25768 -27992 26000 -27928
rect 25460 -28248 26000 -27992
rect 25460 -28312 25704 -28248
rect 25768 -28312 26000 -28248
rect 25460 -28568 26000 -28312
rect 25460 -28632 25704 -28568
rect 25768 -28632 26000 -28568
rect 25460 -28888 26000 -28632
rect 25460 -28952 25704 -28888
rect 25768 -28952 26000 -28888
rect 25460 -29208 26000 -28952
rect 25460 -29272 25704 -29208
rect 25768 -29272 26000 -29208
rect 25460 -29528 26000 -29272
rect 25460 -29592 25704 -29528
rect 25768 -29592 26000 -29528
rect 25460 -29848 26000 -29592
rect 25460 -29912 25704 -29848
rect 25768 -29912 26000 -29848
rect 25460 -30168 26000 -29912
rect 25460 -30232 25704 -30168
rect 25768 -30232 26000 -30168
rect 25460 -30460 26000 -30232
rect 18000 -30488 26000 -30460
rect 18000 -30552 18238 -30488
rect 18302 -30552 25704 -30488
rect 25768 -30552 26000 -30488
rect 18000 -30698 26000 -30552
rect 18000 -30762 18608 -30698
rect 18672 -30762 18928 -30698
rect 18992 -30762 19248 -30698
rect 19312 -30762 19568 -30698
rect 19632 -30762 19888 -30698
rect 19952 -30762 20208 -30698
rect 20272 -30762 20528 -30698
rect 20592 -30762 20848 -30698
rect 20912 -30762 21168 -30698
rect 21232 -30762 21488 -30698
rect 21552 -30762 21808 -30698
rect 21872 -30762 22128 -30698
rect 22192 -30762 22448 -30698
rect 22512 -30762 22768 -30698
rect 22832 -30762 23088 -30698
rect 23152 -30762 23408 -30698
rect 23472 -30762 23728 -30698
rect 23792 -30762 24048 -30698
rect 24112 -30762 24368 -30698
rect 24432 -30762 24688 -30698
rect 24752 -30762 25008 -30698
rect 25072 -30762 25328 -30698
rect 25392 -30762 26000 -30698
rect 18000 -31000 26000 -30762
rect 30000 -26008 30540 -25800
rect 30000 -26072 30238 -26008
rect 30302 -26072 30540 -26008
rect 30000 -26328 30540 -26072
rect 30000 -26392 30238 -26328
rect 30302 -26392 30540 -26328
rect 30000 -26648 30540 -26392
rect 30000 -26712 30238 -26648
rect 30302 -26712 30540 -26648
rect 30000 -26968 30540 -26712
rect 30000 -27032 30238 -26968
rect 30302 -27032 30540 -26968
rect 30000 -27288 30540 -27032
rect 30000 -27352 30238 -27288
rect 30302 -27352 30540 -27288
rect 30000 -27608 30540 -27352
rect 30000 -27672 30238 -27608
rect 30302 -27672 30540 -27608
rect 30000 -27928 30540 -27672
rect 30000 -27992 30238 -27928
rect 30302 -27992 30540 -27928
rect 30000 -28248 30540 -27992
rect 30000 -28312 30238 -28248
rect 30302 -28312 30540 -28248
rect 30000 -28568 30540 -28312
rect 30000 -28632 30238 -28568
rect 30302 -28632 30540 -28568
rect 30000 -28888 30540 -28632
rect 30000 -28952 30238 -28888
rect 30302 -28952 30540 -28888
rect 30000 -29208 30540 -28952
rect 30000 -29272 30238 -29208
rect 30302 -29272 30540 -29208
rect 30000 -29528 30540 -29272
rect 30000 -29592 30238 -29528
rect 30302 -29592 30540 -29528
rect 30000 -29848 30540 -29592
rect 30000 -29912 30238 -29848
rect 30302 -29912 30540 -29848
rect 30000 -30168 30540 -29912
rect 30000 -30232 30238 -30168
rect 30302 -30232 30540 -30168
rect 30000 -30460 30540 -30232
rect 37460 -23768 38000 -23540
rect 37460 -23832 37704 -23768
rect 37768 -23832 38000 -23768
rect 37460 -24088 38000 -23832
rect 37460 -24152 37704 -24088
rect 37768 -24152 38000 -24088
rect 37460 -24408 38000 -24152
rect 37460 -24472 37704 -24408
rect 37768 -24472 38000 -24408
rect 37460 -24728 38000 -24472
rect 37460 -24792 37704 -24728
rect 37768 -24792 38000 -24728
rect 37460 -25048 38000 -24792
rect 37460 -25112 37704 -25048
rect 37768 -25112 38000 -25048
rect 37460 -25368 38000 -25112
rect 37460 -25432 37704 -25368
rect 37768 -25432 38000 -25368
rect 37460 -25688 38000 -25432
rect 37460 -25752 37704 -25688
rect 37768 -25752 38000 -25688
rect 37460 -26008 38000 -25752
rect 37460 -26072 37704 -26008
rect 37768 -26072 38000 -26008
rect 37460 -26328 38000 -26072
rect 37460 -26392 37704 -26328
rect 37768 -26392 38000 -26328
rect 37460 -26648 38000 -26392
rect 37460 -26712 37704 -26648
rect 37768 -26712 38000 -26648
rect 37460 -26968 38000 -26712
rect 37460 -27032 37704 -26968
rect 37768 -27032 38000 -26968
rect 37460 -27288 38000 -27032
rect 37460 -27352 37704 -27288
rect 37768 -27352 38000 -27288
rect 37460 -27608 38000 -27352
rect 37460 -27672 37704 -27608
rect 37768 -27672 38000 -27608
rect 37460 -27928 38000 -27672
rect 37460 -27992 37704 -27928
rect 37768 -27992 38000 -27928
rect 37460 -28248 38000 -27992
rect 37460 -28312 37704 -28248
rect 37768 -28312 38000 -28248
rect 37460 -28568 38000 -28312
rect 37460 -28632 37704 -28568
rect 37768 -28632 38000 -28568
rect 37460 -28888 38000 -28632
rect 37460 -28952 37704 -28888
rect 37768 -28952 38000 -28888
rect 37460 -29208 38000 -28952
rect 37460 -29272 37704 -29208
rect 37768 -29272 38000 -29208
rect 37460 -29528 38000 -29272
rect 37460 -29592 37704 -29528
rect 37768 -29592 38000 -29528
rect 37460 -29848 38000 -29592
rect 37460 -29912 37704 -29848
rect 37768 -29912 38000 -29848
rect 37460 -30168 38000 -29912
rect 37460 -30232 37704 -30168
rect 37768 -30232 38000 -30168
rect 37460 -30460 38000 -30232
rect 30000 -30488 38000 -30460
rect 30000 -30552 30238 -30488
rect 30302 -30552 37704 -30488
rect 37768 -30552 38000 -30488
rect 30000 -30698 38000 -30552
rect 30000 -30762 30608 -30698
rect 30672 -30762 30928 -30698
rect 30992 -30762 31248 -30698
rect 31312 -30762 31568 -30698
rect 31632 -30762 31888 -30698
rect 31952 -30762 32208 -30698
rect 32272 -30762 32528 -30698
rect 32592 -30762 32848 -30698
rect 32912 -30762 33168 -30698
rect 33232 -30762 33488 -30698
rect 33552 -30762 33808 -30698
rect 33872 -30762 34128 -30698
rect 34192 -30762 34448 -30698
rect 34512 -30762 34768 -30698
rect 34832 -30762 35088 -30698
rect 35152 -30762 35408 -30698
rect 35472 -30762 35728 -30698
rect 35792 -30762 36048 -30698
rect 36112 -30762 36368 -30698
rect 36432 -30762 36688 -30698
rect 36752 -30762 37008 -30698
rect 37072 -30762 37328 -30698
rect 37392 -30762 38000 -30698
rect 30000 -31000 38000 -30762
rect 42000 -23242 50000 -23000
rect 42000 -23306 42608 -23242
rect 42672 -23306 42928 -23242
rect 42992 -23306 43248 -23242
rect 43312 -23306 43568 -23242
rect 43632 -23306 43888 -23242
rect 43952 -23306 44208 -23242
rect 44272 -23306 44528 -23242
rect 44592 -23306 44848 -23242
rect 44912 -23306 45168 -23242
rect 45232 -23306 45488 -23242
rect 45552 -23306 45808 -23242
rect 45872 -23306 46128 -23242
rect 46192 -23306 46448 -23242
rect 46512 -23306 46768 -23242
rect 46832 -23306 47088 -23242
rect 47152 -23306 47408 -23242
rect 47472 -23306 47728 -23242
rect 47792 -23306 48048 -23242
rect 48112 -23306 48368 -23242
rect 48432 -23306 48688 -23242
rect 48752 -23306 49008 -23242
rect 49072 -23306 49328 -23242
rect 49392 -23306 50000 -23242
rect 42000 -23448 50000 -23306
rect 42000 -23512 42238 -23448
rect 42302 -23512 49704 -23448
rect 49768 -23512 50000 -23448
rect 42000 -23540 50000 -23512
rect 42000 -23768 42540 -23540
rect 42000 -23832 42238 -23768
rect 42302 -23832 42540 -23768
rect 42000 -24088 42540 -23832
rect 42000 -24152 42238 -24088
rect 42302 -24152 42540 -24088
rect 42000 -24408 42540 -24152
rect 42000 -24472 42238 -24408
rect 42302 -24472 42540 -24408
rect 42000 -24728 42540 -24472
rect 42000 -24792 42238 -24728
rect 42302 -24792 42540 -24728
rect 42000 -25048 42540 -24792
rect 42000 -25112 42238 -25048
rect 42302 -25112 42540 -25048
rect 42000 -25368 42540 -25112
rect 42000 -25432 42238 -25368
rect 42302 -25432 42540 -25368
rect 42000 -25688 42540 -25432
rect 42000 -25752 42238 -25688
rect 42302 -25752 42540 -25688
rect 42000 -26008 42540 -25752
rect 42000 -26072 42238 -26008
rect 42302 -26072 42540 -26008
rect 42000 -26328 42540 -26072
rect 42000 -26392 42238 -26328
rect 42302 -26392 42540 -26328
rect 42000 -26648 42540 -26392
rect 42000 -26712 42238 -26648
rect 42302 -26712 42540 -26648
rect 42000 -26968 42540 -26712
rect 42000 -27032 42238 -26968
rect 42302 -27032 42540 -26968
rect 42000 -27288 42540 -27032
rect 42000 -27352 42238 -27288
rect 42302 -27352 42540 -27288
rect 42000 -27608 42540 -27352
rect 42000 -27672 42238 -27608
rect 42302 -27672 42540 -27608
rect 42000 -27928 42540 -27672
rect 42000 -27992 42238 -27928
rect 42302 -27992 42540 -27928
rect 42000 -28248 42540 -27992
rect 42000 -28312 42238 -28248
rect 42302 -28312 42540 -28248
rect 42000 -28568 42540 -28312
rect 42000 -28632 42238 -28568
rect 42302 -28632 42540 -28568
rect 42000 -28888 42540 -28632
rect 42000 -28952 42238 -28888
rect 42302 -28952 42540 -28888
rect 42000 -29208 42540 -28952
rect 42000 -29272 42238 -29208
rect 42302 -29272 42540 -29208
rect 42000 -29528 42540 -29272
rect 42000 -29592 42238 -29528
rect 42302 -29592 42540 -29528
rect 42000 -29848 42540 -29592
rect 42000 -29912 42238 -29848
rect 42302 -29912 42540 -29848
rect 42000 -30168 42540 -29912
rect 42000 -30232 42238 -30168
rect 42302 -30232 42540 -30168
rect 42000 -30460 42540 -30232
rect 49460 -23768 50000 -23540
rect 49460 -23832 49704 -23768
rect 49768 -23832 50000 -23768
rect 49460 -24088 50000 -23832
rect 49460 -24152 49704 -24088
rect 49768 -24152 50000 -24088
rect 49460 -24408 50000 -24152
rect 49460 -24472 49704 -24408
rect 49768 -24472 50000 -24408
rect 49460 -24728 50000 -24472
rect 49460 -24792 49704 -24728
rect 49768 -24792 50000 -24728
rect 49460 -25048 50000 -24792
rect 49460 -25112 49704 -25048
rect 49768 -25112 50000 -25048
rect 49460 -25368 50000 -25112
rect 49460 -25432 49704 -25368
rect 49768 -25432 50000 -25368
rect 49460 -25688 50000 -25432
rect 49460 -25752 49704 -25688
rect 49768 -25752 50000 -25688
rect 49460 -26008 50000 -25752
rect 49460 -26072 49704 -26008
rect 49768 -26072 50000 -26008
rect 49460 -26328 50000 -26072
rect 49460 -26392 49704 -26328
rect 49768 -26392 50000 -26328
rect 49460 -26648 50000 -26392
rect 49460 -26712 49704 -26648
rect 49768 -26712 50000 -26648
rect 49460 -26968 50000 -26712
rect 49460 -27032 49704 -26968
rect 49768 -27032 50000 -26968
rect 49460 -27288 50000 -27032
rect 49460 -27352 49704 -27288
rect 49768 -27352 50000 -27288
rect 49460 -27608 50000 -27352
rect 49460 -27672 49704 -27608
rect 49768 -27672 50000 -27608
rect 49460 -27928 50000 -27672
rect 49460 -27992 49704 -27928
rect 49768 -27992 50000 -27928
rect 49460 -28248 50000 -27992
rect 49460 -28312 49704 -28248
rect 49768 -28312 50000 -28248
rect 49460 -28568 50000 -28312
rect 49460 -28632 49704 -28568
rect 49768 -28632 50000 -28568
rect 49460 -28888 50000 -28632
rect 49460 -28952 49704 -28888
rect 49768 -28952 50000 -28888
rect 49460 -29208 50000 -28952
rect 49460 -29272 49704 -29208
rect 49768 -29272 50000 -29208
rect 49460 -29528 50000 -29272
rect 49460 -29592 49704 -29528
rect 49768 -29592 50000 -29528
rect 49460 -29848 50000 -29592
rect 49460 -29912 49704 -29848
rect 49768 -29912 50000 -29848
rect 49460 -30168 50000 -29912
rect 49460 -30232 49704 -30168
rect 49768 -30232 50000 -30168
rect 49460 -30460 50000 -30232
rect 42000 -30488 50000 -30460
rect 42000 -30552 42238 -30488
rect 42302 -30552 49704 -30488
rect 49768 -30552 50000 -30488
rect 42000 -30698 50000 -30552
rect 42000 -30762 42608 -30698
rect 42672 -30762 42928 -30698
rect 42992 -30762 43248 -30698
rect 43312 -30762 43568 -30698
rect 43632 -30762 43888 -30698
rect 43952 -30762 44208 -30698
rect 44272 -30762 44528 -30698
rect 44592 -30762 44848 -30698
rect 44912 -30762 45168 -30698
rect 45232 -30762 45488 -30698
rect 45552 -30762 45808 -30698
rect 45872 -30762 46128 -30698
rect 46192 -30762 46448 -30698
rect 46512 -30762 46768 -30698
rect 46832 -30762 47088 -30698
rect 47152 -30762 47408 -30698
rect 47472 -30762 47728 -30698
rect 47792 -30762 48048 -30698
rect 48112 -30762 48368 -30698
rect 48432 -30762 48688 -30698
rect 48752 -30762 49008 -30698
rect 49072 -30762 49328 -30698
rect 49392 -30762 50000 -30698
rect 42000 -31000 50000 -30762
<< via3 >>
rect 18300 -3000 21500 -2500
rect 21882 -5650 21992 -5560
rect 22422 -5880 22982 -5720
rect 22432 -5960 22972 -5880
rect 16500 -9148 17200 -8748
rect 17480 -9360 17600 -8440
rect 17600 -9360 17680 -8440
rect 13300 -10200 15900 -9600
rect 6608 -11246 6672 -11242
rect 6608 -11302 6612 -11246
rect 6612 -11302 6668 -11246
rect 6668 -11302 6672 -11246
rect 6608 -11306 6672 -11302
rect 6928 -11246 6992 -11242
rect 6928 -11302 6932 -11246
rect 6932 -11302 6988 -11246
rect 6988 -11302 6992 -11246
rect 6928 -11306 6992 -11302
rect 7248 -11246 7312 -11242
rect 7248 -11302 7252 -11246
rect 7252 -11302 7308 -11246
rect 7308 -11302 7312 -11246
rect 7248 -11306 7312 -11302
rect 7568 -11246 7632 -11242
rect 7568 -11302 7572 -11246
rect 7572 -11302 7628 -11246
rect 7628 -11302 7632 -11246
rect 7568 -11306 7632 -11302
rect 7888 -11246 7952 -11242
rect 7888 -11302 7892 -11246
rect 7892 -11302 7948 -11246
rect 7948 -11302 7952 -11246
rect 7888 -11306 7952 -11302
rect 8208 -11246 8272 -11242
rect 8208 -11302 8212 -11246
rect 8212 -11302 8268 -11246
rect 8268 -11302 8272 -11246
rect 8208 -11306 8272 -11302
rect 8528 -11246 8592 -11242
rect 8528 -11302 8532 -11246
rect 8532 -11302 8588 -11246
rect 8588 -11302 8592 -11246
rect 8528 -11306 8592 -11302
rect 8848 -11246 8912 -11242
rect 8848 -11302 8852 -11246
rect 8852 -11302 8908 -11246
rect 8908 -11302 8912 -11246
rect 8848 -11306 8912 -11302
rect 9168 -11246 9232 -11242
rect 9168 -11302 9172 -11246
rect 9172 -11302 9228 -11246
rect 9228 -11302 9232 -11246
rect 9168 -11306 9232 -11302
rect 9488 -11246 9552 -11242
rect 9488 -11302 9492 -11246
rect 9492 -11302 9548 -11246
rect 9548 -11302 9552 -11246
rect 9488 -11306 9552 -11302
rect 9808 -11246 9872 -11242
rect 9808 -11302 9812 -11246
rect 9812 -11302 9868 -11246
rect 9868 -11302 9872 -11246
rect 9808 -11306 9872 -11302
rect 10128 -11246 10192 -11242
rect 10128 -11302 10132 -11246
rect 10132 -11302 10188 -11246
rect 10188 -11302 10192 -11246
rect 10128 -11306 10192 -11302
rect 10448 -11246 10512 -11242
rect 10448 -11302 10452 -11246
rect 10452 -11302 10508 -11246
rect 10508 -11302 10512 -11246
rect 10448 -11306 10512 -11302
rect 10768 -11246 10832 -11242
rect 10768 -11302 10772 -11246
rect 10772 -11302 10828 -11246
rect 10828 -11302 10832 -11246
rect 10768 -11306 10832 -11302
rect 11088 -11246 11152 -11242
rect 11088 -11302 11092 -11246
rect 11092 -11302 11148 -11246
rect 11148 -11302 11152 -11246
rect 11088 -11306 11152 -11302
rect 11408 -11246 11472 -11242
rect 11408 -11302 11412 -11246
rect 11412 -11302 11468 -11246
rect 11468 -11302 11472 -11246
rect 11408 -11306 11472 -11302
rect 11728 -11246 11792 -11242
rect 11728 -11302 11732 -11246
rect 11732 -11302 11788 -11246
rect 11788 -11302 11792 -11246
rect 11728 -11306 11792 -11302
rect 12048 -11246 12112 -11242
rect 12048 -11302 12052 -11246
rect 12052 -11302 12108 -11246
rect 12108 -11302 12112 -11246
rect 12048 -11306 12112 -11302
rect 12368 -11246 12432 -11242
rect 12368 -11302 12372 -11246
rect 12372 -11302 12428 -11246
rect 12428 -11302 12432 -11246
rect 12368 -11306 12432 -11302
rect 12688 -11246 12752 -11242
rect 12688 -11302 12692 -11246
rect 12692 -11302 12748 -11246
rect 12748 -11302 12752 -11246
rect 12688 -11306 12752 -11302
rect 13008 -11246 13072 -11242
rect 13008 -11302 13012 -11246
rect 13012 -11302 13068 -11246
rect 13068 -11302 13072 -11246
rect 13008 -11306 13072 -11302
rect 13328 -11246 13392 -11242
rect 13328 -11302 13332 -11246
rect 13332 -11302 13388 -11246
rect 13388 -11302 13392 -11246
rect 13328 -11306 13392 -11302
rect 6238 -11452 6302 -11448
rect 6238 -11508 6242 -11452
rect 6242 -11508 6298 -11452
rect 6298 -11508 6302 -11452
rect 6238 -11512 6302 -11508
rect 13704 -11452 13768 -11448
rect 13704 -11508 13708 -11452
rect 13708 -11508 13764 -11452
rect 13764 -11508 13768 -11452
rect 13704 -11512 13768 -11508
rect 6238 -11772 6302 -11768
rect 6238 -11828 6242 -11772
rect 6242 -11828 6298 -11772
rect 6298 -11828 6302 -11772
rect 6238 -11832 6302 -11828
rect 6238 -12092 6302 -12088
rect 6238 -12148 6242 -12092
rect 6242 -12148 6298 -12092
rect 6298 -12148 6302 -12092
rect 6238 -12152 6302 -12148
rect 6238 -12412 6302 -12408
rect 6238 -12468 6242 -12412
rect 6242 -12468 6298 -12412
rect 6298 -12468 6302 -12412
rect 6238 -12472 6302 -12468
rect 6238 -12732 6302 -12728
rect 6238 -12788 6242 -12732
rect 6242 -12788 6298 -12732
rect 6298 -12788 6302 -12732
rect 6238 -12792 6302 -12788
rect 6238 -13052 6302 -13048
rect 6238 -13108 6242 -13052
rect 6242 -13108 6298 -13052
rect 6298 -13108 6302 -13052
rect 6238 -13112 6302 -13108
rect 6238 -13372 6302 -13368
rect 6238 -13428 6242 -13372
rect 6242 -13428 6298 -13372
rect 6298 -13428 6302 -13372
rect 6238 -13432 6302 -13428
rect 6238 -13692 6302 -13688
rect 6238 -13748 6242 -13692
rect 6242 -13748 6298 -13692
rect 6298 -13748 6302 -13692
rect 6238 -13752 6302 -13748
rect 6238 -14012 6302 -14008
rect 6238 -14068 6242 -14012
rect 6242 -14068 6298 -14012
rect 6298 -14068 6302 -14012
rect 6238 -14072 6302 -14068
rect 6238 -14332 6302 -14328
rect 6238 -14388 6242 -14332
rect 6242 -14388 6298 -14332
rect 6298 -14388 6302 -14332
rect 6238 -14392 6302 -14388
rect 6238 -14652 6302 -14648
rect 6238 -14708 6242 -14652
rect 6242 -14708 6298 -14652
rect 6298 -14708 6302 -14652
rect 6238 -14712 6302 -14708
rect 6238 -14972 6302 -14968
rect 6238 -15028 6242 -14972
rect 6242 -15028 6298 -14972
rect 6298 -15028 6302 -14972
rect 6238 -15032 6302 -15028
rect 6238 -15292 6302 -15288
rect 6238 -15348 6242 -15292
rect 6242 -15348 6298 -15292
rect 6298 -15348 6302 -15292
rect 6238 -15352 6302 -15348
rect 6238 -15612 6302 -15608
rect 6238 -15668 6242 -15612
rect 6242 -15668 6298 -15612
rect 6298 -15668 6302 -15612
rect 6238 -15672 6302 -15668
rect 6238 -15932 6302 -15928
rect 6238 -15988 6242 -15932
rect 6242 -15988 6298 -15932
rect 6298 -15988 6302 -15932
rect 6238 -15992 6302 -15988
rect 6238 -16252 6302 -16248
rect 6238 -16308 6242 -16252
rect 6242 -16308 6298 -16252
rect 6298 -16308 6302 -16252
rect 6238 -16312 6302 -16308
rect 6238 -16572 6302 -16568
rect 6238 -16628 6242 -16572
rect 6242 -16628 6298 -16572
rect 6298 -16628 6302 -16572
rect 6238 -16632 6302 -16628
rect 6238 -16892 6302 -16888
rect 6238 -16948 6242 -16892
rect 6242 -16948 6298 -16892
rect 6298 -16948 6302 -16892
rect 6238 -16952 6302 -16948
rect 6238 -17212 6302 -17208
rect 6238 -17268 6242 -17212
rect 6242 -17268 6298 -17212
rect 6298 -17268 6302 -17212
rect 6238 -17272 6302 -17268
rect 6238 -17532 6302 -17528
rect 6238 -17588 6242 -17532
rect 6242 -17588 6298 -17532
rect 6298 -17588 6302 -17532
rect 6238 -17592 6302 -17588
rect 6238 -17852 6302 -17848
rect 6238 -17908 6242 -17852
rect 6242 -17908 6298 -17852
rect 6298 -17908 6302 -17852
rect 6238 -17912 6302 -17908
rect 6238 -18172 6302 -18168
rect 6238 -18228 6242 -18172
rect 6242 -18228 6298 -18172
rect 6298 -18228 6302 -18172
rect 6238 -18232 6302 -18228
rect 13704 -11772 13768 -11768
rect 13704 -11828 13708 -11772
rect 13708 -11828 13764 -11772
rect 13764 -11828 13768 -11772
rect 13704 -11832 13768 -11828
rect 13704 -12092 13768 -12088
rect 13704 -12148 13708 -12092
rect 13708 -12148 13764 -12092
rect 13764 -12148 13768 -12092
rect 13704 -12152 13768 -12148
rect 13704 -12412 13768 -12408
rect 13704 -12468 13708 -12412
rect 13708 -12468 13764 -12412
rect 13764 -12468 13768 -12412
rect 13704 -12472 13768 -12468
rect 13704 -12732 13768 -12728
rect 13704 -12788 13708 -12732
rect 13708 -12788 13764 -12732
rect 13764 -12788 13768 -12732
rect 13704 -12792 13768 -12788
rect 13704 -13052 13768 -13048
rect 13704 -13108 13708 -13052
rect 13708 -13108 13764 -13052
rect 13764 -13108 13768 -13052
rect 13704 -13112 13768 -13108
rect 13704 -13372 13768 -13368
rect 13704 -13428 13708 -13372
rect 13708 -13428 13764 -13372
rect 13764 -13428 13768 -13372
rect 13704 -13432 13768 -13428
rect 13704 -13692 13768 -13688
rect 13704 -13748 13708 -13692
rect 13708 -13748 13764 -13692
rect 13764 -13748 13768 -13692
rect 13704 -13752 13768 -13748
rect 13704 -14012 13768 -14008
rect 13704 -14068 13708 -14012
rect 13708 -14068 13764 -14012
rect 13764 -14068 13768 -14012
rect 13704 -14072 13768 -14068
rect 13704 -14332 13768 -14328
rect 13704 -14388 13708 -14332
rect 13708 -14388 13764 -14332
rect 13764 -14388 13768 -14332
rect 13704 -14392 13768 -14388
rect 13704 -14652 13768 -14648
rect 13704 -14708 13708 -14652
rect 13708 -14708 13764 -14652
rect 13764 -14708 13768 -14652
rect 13704 -14712 13768 -14708
rect 13704 -14972 13768 -14968
rect 13704 -15028 13708 -14972
rect 13708 -15028 13764 -14972
rect 13764 -15028 13768 -14972
rect 13704 -15032 13768 -15028
rect 13704 -15292 13768 -15288
rect 13704 -15348 13708 -15292
rect 13708 -15348 13764 -15292
rect 13764 -15348 13768 -15292
rect 13704 -15352 13768 -15348
rect 13704 -15612 13768 -15608
rect 13704 -15668 13708 -15612
rect 13708 -15668 13764 -15612
rect 13764 -15668 13768 -15612
rect 13704 -15672 13768 -15668
rect 13704 -15932 13768 -15928
rect 13704 -15988 13708 -15932
rect 13708 -15988 13764 -15932
rect 13764 -15988 13768 -15932
rect 13704 -15992 13768 -15988
rect 13704 -16252 13768 -16248
rect 13704 -16308 13708 -16252
rect 13708 -16308 13764 -16252
rect 13764 -16308 13768 -16252
rect 13704 -16312 13768 -16308
rect 13704 -16572 13768 -16568
rect 13704 -16628 13708 -16572
rect 13708 -16628 13764 -16572
rect 13764 -16628 13768 -16572
rect 13704 -16632 13768 -16628
rect 13704 -16892 13768 -16888
rect 13704 -16948 13708 -16892
rect 13708 -16948 13764 -16892
rect 13764 -16948 13768 -16892
rect 13704 -16952 13768 -16948
rect 13704 -17212 13768 -17208
rect 13704 -17268 13708 -17212
rect 13708 -17268 13764 -17212
rect 13764 -17268 13768 -17212
rect 13704 -17272 13768 -17268
rect 13704 -17532 13768 -17528
rect 13704 -17588 13708 -17532
rect 13708 -17588 13764 -17532
rect 13764 -17588 13768 -17532
rect 13704 -17592 13768 -17588
rect 13704 -17852 13768 -17848
rect 13704 -17908 13708 -17852
rect 13708 -17908 13764 -17852
rect 13764 -17908 13768 -17852
rect 13704 -17912 13768 -17908
rect 13704 -18172 13768 -18168
rect 13704 -18228 13708 -18172
rect 13708 -18228 13764 -18172
rect 13764 -18228 13768 -18172
rect 13704 -18232 13768 -18228
rect 6238 -18492 6302 -18488
rect 6238 -18548 6242 -18492
rect 6242 -18548 6298 -18492
rect 6298 -18548 6302 -18492
rect 6238 -18552 6302 -18548
rect 13704 -18492 13768 -18488
rect 13704 -18548 13708 -18492
rect 13708 -18548 13764 -18492
rect 13764 -18548 13768 -18492
rect 13704 -18552 13768 -18548
rect 6608 -18702 6672 -18698
rect 6608 -18758 6612 -18702
rect 6612 -18758 6668 -18702
rect 6668 -18758 6672 -18702
rect 6608 -18762 6672 -18758
rect 6928 -18702 6992 -18698
rect 6928 -18758 6932 -18702
rect 6932 -18758 6988 -18702
rect 6988 -18758 6992 -18702
rect 6928 -18762 6992 -18758
rect 7248 -18702 7312 -18698
rect 7248 -18758 7252 -18702
rect 7252 -18758 7308 -18702
rect 7308 -18758 7312 -18702
rect 7248 -18762 7312 -18758
rect 7568 -18702 7632 -18698
rect 7568 -18758 7572 -18702
rect 7572 -18758 7628 -18702
rect 7628 -18758 7632 -18702
rect 7568 -18762 7632 -18758
rect 7888 -18702 7952 -18698
rect 7888 -18758 7892 -18702
rect 7892 -18758 7948 -18702
rect 7948 -18758 7952 -18702
rect 7888 -18762 7952 -18758
rect 8208 -18702 8272 -18698
rect 8208 -18758 8212 -18702
rect 8212 -18758 8268 -18702
rect 8268 -18758 8272 -18702
rect 8208 -18762 8272 -18758
rect 8528 -18702 8592 -18698
rect 8528 -18758 8532 -18702
rect 8532 -18758 8588 -18702
rect 8588 -18758 8592 -18702
rect 8528 -18762 8592 -18758
rect 8848 -18702 8912 -18698
rect 8848 -18758 8852 -18702
rect 8852 -18758 8908 -18702
rect 8908 -18758 8912 -18702
rect 8848 -18762 8912 -18758
rect 9168 -18702 9232 -18698
rect 9168 -18758 9172 -18702
rect 9172 -18758 9228 -18702
rect 9228 -18758 9232 -18702
rect 9168 -18762 9232 -18758
rect 9488 -18702 9552 -18698
rect 9488 -18758 9492 -18702
rect 9492 -18758 9548 -18702
rect 9548 -18758 9552 -18702
rect 9488 -18762 9552 -18758
rect 9808 -18702 9872 -18698
rect 9808 -18758 9812 -18702
rect 9812 -18758 9868 -18702
rect 9868 -18758 9872 -18702
rect 9808 -18762 9872 -18758
rect 10128 -18702 10192 -18698
rect 10128 -18758 10132 -18702
rect 10132 -18758 10188 -18702
rect 10188 -18758 10192 -18702
rect 10128 -18762 10192 -18758
rect 10448 -18702 10512 -18698
rect 10448 -18758 10452 -18702
rect 10452 -18758 10508 -18702
rect 10508 -18758 10512 -18702
rect 10448 -18762 10512 -18758
rect 10768 -18702 10832 -18698
rect 10768 -18758 10772 -18702
rect 10772 -18758 10828 -18702
rect 10828 -18758 10832 -18702
rect 10768 -18762 10832 -18758
rect 11088 -18702 11152 -18698
rect 11088 -18758 11092 -18702
rect 11092 -18758 11148 -18702
rect 11148 -18758 11152 -18702
rect 11088 -18762 11152 -18758
rect 11408 -18702 11472 -18698
rect 11408 -18758 11412 -18702
rect 11412 -18758 11468 -18702
rect 11468 -18758 11472 -18702
rect 11408 -18762 11472 -18758
rect 11728 -18702 11792 -18698
rect 11728 -18758 11732 -18702
rect 11732 -18758 11788 -18702
rect 11788 -18758 11792 -18702
rect 11728 -18762 11792 -18758
rect 12048 -18702 12112 -18698
rect 12048 -18758 12052 -18702
rect 12052 -18758 12108 -18702
rect 12108 -18758 12112 -18702
rect 12048 -18762 12112 -18758
rect 12368 -18702 12432 -18698
rect 12368 -18758 12372 -18702
rect 12372 -18758 12428 -18702
rect 12428 -18758 12432 -18702
rect 12368 -18762 12432 -18758
rect 12688 -18702 12752 -18698
rect 12688 -18758 12692 -18702
rect 12692 -18758 12748 -18702
rect 12748 -18758 12752 -18702
rect 12688 -18762 12752 -18758
rect 13008 -18702 13072 -18698
rect 13008 -18758 13012 -18702
rect 13012 -18758 13068 -18702
rect 13068 -18758 13072 -18702
rect 13008 -18762 13072 -18758
rect 13328 -18702 13392 -18698
rect 13328 -18758 13332 -18702
rect 13332 -18758 13388 -18702
rect 13388 -18758 13392 -18702
rect 13328 -18762 13392 -18758
rect 6608 -23246 6672 -23242
rect 6608 -23302 6612 -23246
rect 6612 -23302 6668 -23246
rect 6668 -23302 6672 -23246
rect 6608 -23306 6672 -23302
rect 6928 -23246 6992 -23242
rect 6928 -23302 6932 -23246
rect 6932 -23302 6988 -23246
rect 6988 -23302 6992 -23246
rect 6928 -23306 6992 -23302
rect 7248 -23246 7312 -23242
rect 7248 -23302 7252 -23246
rect 7252 -23302 7308 -23246
rect 7308 -23302 7312 -23246
rect 7248 -23306 7312 -23302
rect 7568 -23246 7632 -23242
rect 7568 -23302 7572 -23246
rect 7572 -23302 7628 -23246
rect 7628 -23302 7632 -23246
rect 7568 -23306 7632 -23302
rect 7888 -23246 7952 -23242
rect 7888 -23302 7892 -23246
rect 7892 -23302 7948 -23246
rect 7948 -23302 7952 -23246
rect 7888 -23306 7952 -23302
rect 8208 -23246 8272 -23242
rect 8208 -23302 8212 -23246
rect 8212 -23302 8268 -23246
rect 8268 -23302 8272 -23246
rect 8208 -23306 8272 -23302
rect 8528 -23246 8592 -23242
rect 8528 -23302 8532 -23246
rect 8532 -23302 8588 -23246
rect 8588 -23302 8592 -23246
rect 8528 -23306 8592 -23302
rect 8848 -23246 8912 -23242
rect 8848 -23302 8852 -23246
rect 8852 -23302 8908 -23246
rect 8908 -23302 8912 -23246
rect 8848 -23306 8912 -23302
rect 9168 -23246 9232 -23242
rect 9168 -23302 9172 -23246
rect 9172 -23302 9228 -23246
rect 9228 -23302 9232 -23246
rect 9168 -23306 9232 -23302
rect 9488 -23246 9552 -23242
rect 9488 -23302 9492 -23246
rect 9492 -23302 9548 -23246
rect 9548 -23302 9552 -23246
rect 9488 -23306 9552 -23302
rect 9808 -23246 9872 -23242
rect 9808 -23302 9812 -23246
rect 9812 -23302 9868 -23246
rect 9868 -23302 9872 -23246
rect 9808 -23306 9872 -23302
rect 10128 -23246 10192 -23242
rect 10128 -23302 10132 -23246
rect 10132 -23302 10188 -23246
rect 10188 -23302 10192 -23246
rect 10128 -23306 10192 -23302
rect 10448 -23246 10512 -23242
rect 10448 -23302 10452 -23246
rect 10452 -23302 10508 -23246
rect 10508 -23302 10512 -23246
rect 10448 -23306 10512 -23302
rect 10768 -23246 10832 -23242
rect 10768 -23302 10772 -23246
rect 10772 -23302 10828 -23246
rect 10828 -23302 10832 -23246
rect 10768 -23306 10832 -23302
rect 11088 -23246 11152 -23242
rect 11088 -23302 11092 -23246
rect 11092 -23302 11148 -23246
rect 11148 -23302 11152 -23246
rect 11088 -23306 11152 -23302
rect 11408 -23246 11472 -23242
rect 11408 -23302 11412 -23246
rect 11412 -23302 11468 -23246
rect 11468 -23302 11472 -23246
rect 11408 -23306 11472 -23302
rect 11728 -23246 11792 -23242
rect 11728 -23302 11732 -23246
rect 11732 -23302 11788 -23246
rect 11788 -23302 11792 -23246
rect 11728 -23306 11792 -23302
rect 12048 -23246 12112 -23242
rect 12048 -23302 12052 -23246
rect 12052 -23302 12108 -23246
rect 12108 -23302 12112 -23246
rect 12048 -23306 12112 -23302
rect 12368 -23246 12432 -23242
rect 12368 -23302 12372 -23246
rect 12372 -23302 12428 -23246
rect 12428 -23302 12432 -23246
rect 12368 -23306 12432 -23302
rect 12688 -23246 12752 -23242
rect 12688 -23302 12692 -23246
rect 12692 -23302 12748 -23246
rect 12748 -23302 12752 -23246
rect 12688 -23306 12752 -23302
rect 13008 -23246 13072 -23242
rect 13008 -23302 13012 -23246
rect 13012 -23302 13068 -23246
rect 13068 -23302 13072 -23246
rect 13008 -23306 13072 -23302
rect 13328 -23246 13392 -23242
rect 13328 -23302 13332 -23246
rect 13332 -23302 13388 -23246
rect 13388 -23302 13392 -23246
rect 13328 -23306 13392 -23302
rect 6238 -23452 6302 -23448
rect 6238 -23508 6242 -23452
rect 6242 -23508 6298 -23452
rect 6298 -23508 6302 -23452
rect 6238 -23512 6302 -23508
rect 13704 -23452 13768 -23448
rect 13704 -23508 13708 -23452
rect 13708 -23508 13764 -23452
rect 13764 -23508 13768 -23452
rect 13704 -23512 13768 -23508
rect 6238 -23772 6302 -23768
rect 6238 -23828 6242 -23772
rect 6242 -23828 6298 -23772
rect 6298 -23828 6302 -23772
rect 6238 -23832 6302 -23828
rect 6238 -24092 6302 -24088
rect 6238 -24148 6242 -24092
rect 6242 -24148 6298 -24092
rect 6298 -24148 6302 -24092
rect 6238 -24152 6302 -24148
rect 6238 -24412 6302 -24408
rect 6238 -24468 6242 -24412
rect 6242 -24468 6298 -24412
rect 6298 -24468 6302 -24412
rect 6238 -24472 6302 -24468
rect 6238 -24732 6302 -24728
rect 6238 -24788 6242 -24732
rect 6242 -24788 6298 -24732
rect 6298 -24788 6302 -24732
rect 6238 -24792 6302 -24788
rect 6238 -25052 6302 -25048
rect 6238 -25108 6242 -25052
rect 6242 -25108 6298 -25052
rect 6298 -25108 6302 -25052
rect 6238 -25112 6302 -25108
rect 6238 -25372 6302 -25368
rect 6238 -25428 6242 -25372
rect 6242 -25428 6298 -25372
rect 6298 -25428 6302 -25372
rect 6238 -25432 6302 -25428
rect 6238 -25692 6302 -25688
rect 6238 -25748 6242 -25692
rect 6242 -25748 6298 -25692
rect 6298 -25748 6302 -25692
rect 6238 -25752 6302 -25748
rect 6238 -26012 6302 -26008
rect 6238 -26068 6242 -26012
rect 6242 -26068 6298 -26012
rect 6298 -26068 6302 -26012
rect 6238 -26072 6302 -26068
rect 6238 -26332 6302 -26328
rect 6238 -26388 6242 -26332
rect 6242 -26388 6298 -26332
rect 6298 -26388 6302 -26332
rect 6238 -26392 6302 -26388
rect 6238 -26652 6302 -26648
rect 6238 -26708 6242 -26652
rect 6242 -26708 6298 -26652
rect 6298 -26708 6302 -26652
rect 6238 -26712 6302 -26708
rect 6238 -26972 6302 -26968
rect 6238 -27028 6242 -26972
rect 6242 -27028 6298 -26972
rect 6298 -27028 6302 -26972
rect 6238 -27032 6302 -27028
rect 6238 -27292 6302 -27288
rect 6238 -27348 6242 -27292
rect 6242 -27348 6298 -27292
rect 6298 -27348 6302 -27292
rect 6238 -27352 6302 -27348
rect 6238 -27612 6302 -27608
rect 6238 -27668 6242 -27612
rect 6242 -27668 6298 -27612
rect 6298 -27668 6302 -27612
rect 6238 -27672 6302 -27668
rect 6238 -27932 6302 -27928
rect 6238 -27988 6242 -27932
rect 6242 -27988 6298 -27932
rect 6298 -27988 6302 -27932
rect 6238 -27992 6302 -27988
rect 6238 -28252 6302 -28248
rect 6238 -28308 6242 -28252
rect 6242 -28308 6298 -28252
rect 6298 -28308 6302 -28252
rect 6238 -28312 6302 -28308
rect 6238 -28572 6302 -28568
rect 6238 -28628 6242 -28572
rect 6242 -28628 6298 -28572
rect 6298 -28628 6302 -28572
rect 6238 -28632 6302 -28628
rect 6238 -28892 6302 -28888
rect 6238 -28948 6242 -28892
rect 6242 -28948 6298 -28892
rect 6298 -28948 6302 -28892
rect 6238 -28952 6302 -28948
rect 6238 -29212 6302 -29208
rect 6238 -29268 6242 -29212
rect 6242 -29268 6298 -29212
rect 6298 -29268 6302 -29212
rect 6238 -29272 6302 -29268
rect 6238 -29532 6302 -29528
rect 6238 -29588 6242 -29532
rect 6242 -29588 6298 -29532
rect 6298 -29588 6302 -29532
rect 6238 -29592 6302 -29588
rect 6238 -29852 6302 -29848
rect 6238 -29908 6242 -29852
rect 6242 -29908 6298 -29852
rect 6298 -29908 6302 -29852
rect 6238 -29912 6302 -29908
rect 6238 -30172 6302 -30168
rect 6238 -30228 6242 -30172
rect 6242 -30228 6298 -30172
rect 6298 -30228 6302 -30172
rect 6238 -30232 6302 -30228
rect 13704 -23772 13768 -23768
rect 13704 -23828 13708 -23772
rect 13708 -23828 13764 -23772
rect 13764 -23828 13768 -23772
rect 13704 -23832 13768 -23828
rect 13704 -24092 13768 -24088
rect 13704 -24148 13708 -24092
rect 13708 -24148 13764 -24092
rect 13764 -24148 13768 -24092
rect 13704 -24152 13768 -24148
rect 13704 -24412 13768 -24408
rect 13704 -24468 13708 -24412
rect 13708 -24468 13764 -24412
rect 13764 -24468 13768 -24412
rect 13704 -24472 13768 -24468
rect 13704 -24732 13768 -24728
rect 13704 -24788 13708 -24732
rect 13708 -24788 13764 -24732
rect 13764 -24788 13768 -24732
rect 13704 -24792 13768 -24788
rect 13704 -25052 13768 -25048
rect 13704 -25108 13708 -25052
rect 13708 -25108 13764 -25052
rect 13764 -25108 13768 -25052
rect 13704 -25112 13768 -25108
rect 13704 -25372 13768 -25368
rect 13704 -25428 13708 -25372
rect 13708 -25428 13764 -25372
rect 13764 -25428 13768 -25372
rect 13704 -25432 13768 -25428
rect 13704 -25692 13768 -25688
rect 13704 -25748 13708 -25692
rect 13708 -25748 13764 -25692
rect 13764 -25748 13768 -25692
rect 13704 -25752 13768 -25748
rect 17700 -10200 18900 -9600
rect 20900 -10200 22100 -9600
rect 18608 -11246 18672 -11242
rect 18608 -11302 18612 -11246
rect 18612 -11302 18668 -11246
rect 18668 -11302 18672 -11246
rect 18608 -11306 18672 -11302
rect 18928 -11246 18992 -11242
rect 18928 -11302 18932 -11246
rect 18932 -11302 18988 -11246
rect 18988 -11302 18992 -11246
rect 18928 -11306 18992 -11302
rect 19248 -11246 19312 -11242
rect 19248 -11302 19252 -11246
rect 19252 -11302 19308 -11246
rect 19308 -11302 19312 -11246
rect 19248 -11306 19312 -11302
rect 19568 -11246 19632 -11242
rect 19568 -11302 19572 -11246
rect 19572 -11302 19628 -11246
rect 19628 -11302 19632 -11246
rect 19568 -11306 19632 -11302
rect 19888 -11246 19952 -11242
rect 19888 -11302 19892 -11246
rect 19892 -11302 19948 -11246
rect 19948 -11302 19952 -11246
rect 19888 -11306 19952 -11302
rect 20208 -11246 20272 -11242
rect 20208 -11302 20212 -11246
rect 20212 -11302 20268 -11246
rect 20268 -11302 20272 -11246
rect 20208 -11306 20272 -11302
rect 20528 -11246 20592 -11242
rect 20528 -11302 20532 -11246
rect 20532 -11302 20588 -11246
rect 20588 -11302 20592 -11246
rect 20528 -11306 20592 -11302
rect 20848 -11246 20912 -11242
rect 20848 -11302 20852 -11246
rect 20852 -11302 20908 -11246
rect 20908 -11302 20912 -11246
rect 20848 -11306 20912 -11302
rect 21168 -11246 21232 -11242
rect 21168 -11302 21172 -11246
rect 21172 -11302 21228 -11246
rect 21228 -11302 21232 -11246
rect 21168 -11306 21232 -11302
rect 21488 -11246 21552 -11242
rect 21488 -11302 21492 -11246
rect 21492 -11302 21548 -11246
rect 21548 -11302 21552 -11246
rect 21488 -11306 21552 -11302
rect 21808 -11246 21872 -11242
rect 21808 -11302 21812 -11246
rect 21812 -11302 21868 -11246
rect 21868 -11302 21872 -11246
rect 21808 -11306 21872 -11302
rect 22128 -11246 22192 -11242
rect 22128 -11302 22132 -11246
rect 22132 -11302 22188 -11246
rect 22188 -11302 22192 -11246
rect 22128 -11306 22192 -11302
rect 22448 -11246 22512 -11242
rect 22448 -11302 22452 -11246
rect 22452 -11302 22508 -11246
rect 22508 -11302 22512 -11246
rect 22448 -11306 22512 -11302
rect 22768 -11246 22832 -11242
rect 22768 -11302 22772 -11246
rect 22772 -11302 22828 -11246
rect 22828 -11302 22832 -11246
rect 22768 -11306 22832 -11302
rect 23088 -11246 23152 -11242
rect 23088 -11302 23092 -11246
rect 23092 -11302 23148 -11246
rect 23148 -11302 23152 -11246
rect 23088 -11306 23152 -11302
rect 23408 -11246 23472 -11242
rect 23408 -11302 23412 -11246
rect 23412 -11302 23468 -11246
rect 23468 -11302 23472 -11246
rect 23408 -11306 23472 -11302
rect 23728 -11246 23792 -11242
rect 23728 -11302 23732 -11246
rect 23732 -11302 23788 -11246
rect 23788 -11302 23792 -11246
rect 23728 -11306 23792 -11302
rect 24048 -11246 24112 -11242
rect 24048 -11302 24052 -11246
rect 24052 -11302 24108 -11246
rect 24108 -11302 24112 -11246
rect 24048 -11306 24112 -11302
rect 24368 -11246 24432 -11242
rect 24368 -11302 24372 -11246
rect 24372 -11302 24428 -11246
rect 24428 -11302 24432 -11246
rect 24368 -11306 24432 -11302
rect 24688 -11246 24752 -11242
rect 24688 -11302 24692 -11246
rect 24692 -11302 24748 -11246
rect 24748 -11302 24752 -11246
rect 24688 -11306 24752 -11302
rect 25008 -11246 25072 -11242
rect 25008 -11302 25012 -11246
rect 25012 -11302 25068 -11246
rect 25068 -11302 25072 -11246
rect 25008 -11306 25072 -11302
rect 25328 -11246 25392 -11242
rect 25328 -11302 25332 -11246
rect 25332 -11302 25388 -11246
rect 25388 -11302 25392 -11246
rect 25328 -11306 25392 -11302
rect 18238 -11452 18302 -11448
rect 18238 -11508 18242 -11452
rect 18242 -11508 18298 -11452
rect 18298 -11508 18302 -11452
rect 18238 -11512 18302 -11508
rect 25704 -11452 25768 -11448
rect 25704 -11508 25708 -11452
rect 25708 -11508 25764 -11452
rect 25764 -11508 25768 -11452
rect 25704 -11512 25768 -11508
rect 18238 -11772 18302 -11768
rect 18238 -11828 18242 -11772
rect 18242 -11828 18298 -11772
rect 18298 -11828 18302 -11772
rect 18238 -11832 18302 -11828
rect 18238 -12092 18302 -12088
rect 18238 -12148 18242 -12092
rect 18242 -12148 18298 -12092
rect 18298 -12148 18302 -12092
rect 18238 -12152 18302 -12148
rect 18238 -12412 18302 -12408
rect 18238 -12468 18242 -12412
rect 18242 -12468 18298 -12412
rect 18298 -12468 18302 -12412
rect 18238 -12472 18302 -12468
rect 18238 -12732 18302 -12728
rect 18238 -12788 18242 -12732
rect 18242 -12788 18298 -12732
rect 18298 -12788 18302 -12732
rect 18238 -12792 18302 -12788
rect 18238 -13052 18302 -13048
rect 18238 -13108 18242 -13052
rect 18242 -13108 18298 -13052
rect 18298 -13108 18302 -13052
rect 18238 -13112 18302 -13108
rect 18238 -13372 18302 -13368
rect 18238 -13428 18242 -13372
rect 18242 -13428 18298 -13372
rect 18298 -13428 18302 -13372
rect 18238 -13432 18302 -13428
rect 18238 -13692 18302 -13688
rect 18238 -13748 18242 -13692
rect 18242 -13748 18298 -13692
rect 18298 -13748 18302 -13692
rect 18238 -13752 18302 -13748
rect 18238 -14012 18302 -14008
rect 18238 -14068 18242 -14012
rect 18242 -14068 18298 -14012
rect 18298 -14068 18302 -14012
rect 18238 -14072 18302 -14068
rect 18238 -14332 18302 -14328
rect 18238 -14388 18242 -14332
rect 18242 -14388 18298 -14332
rect 18298 -14388 18302 -14332
rect 18238 -14392 18302 -14388
rect 18238 -14652 18302 -14648
rect 18238 -14708 18242 -14652
rect 18242 -14708 18298 -14652
rect 18298 -14708 18302 -14652
rect 18238 -14712 18302 -14708
rect 18238 -14972 18302 -14968
rect 18238 -15028 18242 -14972
rect 18242 -15028 18298 -14972
rect 18298 -15028 18302 -14972
rect 18238 -15032 18302 -15028
rect 18238 -15292 18302 -15288
rect 18238 -15348 18242 -15292
rect 18242 -15348 18298 -15292
rect 18298 -15348 18302 -15292
rect 18238 -15352 18302 -15348
rect 18238 -15612 18302 -15608
rect 18238 -15668 18242 -15612
rect 18242 -15668 18298 -15612
rect 18298 -15668 18302 -15612
rect 18238 -15672 18302 -15668
rect 18238 -15932 18302 -15928
rect 18238 -15988 18242 -15932
rect 18242 -15988 18298 -15932
rect 18298 -15988 18302 -15932
rect 18238 -15992 18302 -15988
rect 18238 -16252 18302 -16248
rect 18238 -16308 18242 -16252
rect 18242 -16308 18298 -16252
rect 18298 -16308 18302 -16252
rect 18238 -16312 18302 -16308
rect 18238 -16572 18302 -16568
rect 18238 -16628 18242 -16572
rect 18242 -16628 18298 -16572
rect 18298 -16628 18302 -16572
rect 18238 -16632 18302 -16628
rect 18238 -16892 18302 -16888
rect 18238 -16948 18242 -16892
rect 18242 -16948 18298 -16892
rect 18298 -16948 18302 -16892
rect 18238 -16952 18302 -16948
rect 18238 -17212 18302 -17208
rect 18238 -17268 18242 -17212
rect 18242 -17268 18298 -17212
rect 18298 -17268 18302 -17212
rect 18238 -17272 18302 -17268
rect 18238 -17532 18302 -17528
rect 18238 -17588 18242 -17532
rect 18242 -17588 18298 -17532
rect 18298 -17588 18302 -17532
rect 18238 -17592 18302 -17588
rect 18238 -17852 18302 -17848
rect 18238 -17908 18242 -17852
rect 18242 -17908 18298 -17852
rect 18298 -17908 18302 -17852
rect 18238 -17912 18302 -17908
rect 18238 -18172 18302 -18168
rect 18238 -18228 18242 -18172
rect 18242 -18228 18298 -18172
rect 18298 -18228 18302 -18172
rect 18238 -18232 18302 -18228
rect 25704 -11772 25768 -11768
rect 25704 -11828 25708 -11772
rect 25708 -11828 25764 -11772
rect 25764 -11828 25768 -11772
rect 25704 -11832 25768 -11828
rect 25704 -12092 25768 -12088
rect 25704 -12148 25708 -12092
rect 25708 -12148 25764 -12092
rect 25764 -12148 25768 -12092
rect 25704 -12152 25768 -12148
rect 25704 -12412 25768 -12408
rect 25704 -12468 25708 -12412
rect 25708 -12468 25764 -12412
rect 25764 -12468 25768 -12412
rect 25704 -12472 25768 -12468
rect 25704 -12732 25768 -12728
rect 25704 -12788 25708 -12732
rect 25708 -12788 25764 -12732
rect 25764 -12788 25768 -12732
rect 25704 -12792 25768 -12788
rect 25704 -13052 25768 -13048
rect 25704 -13108 25708 -13052
rect 25708 -13108 25764 -13052
rect 25764 -13108 25768 -13052
rect 25704 -13112 25768 -13108
rect 25704 -13372 25768 -13368
rect 25704 -13428 25708 -13372
rect 25708 -13428 25764 -13372
rect 25764 -13428 25768 -13372
rect 25704 -13432 25768 -13428
rect 25704 -13692 25768 -13688
rect 25704 -13748 25708 -13692
rect 25708 -13748 25764 -13692
rect 25764 -13748 25768 -13692
rect 25704 -13752 25768 -13748
rect 25704 -14012 25768 -14008
rect 25704 -14068 25708 -14012
rect 25708 -14068 25764 -14012
rect 25764 -14068 25768 -14012
rect 25704 -14072 25768 -14068
rect 25704 -14332 25768 -14328
rect 25704 -14388 25708 -14332
rect 25708 -14388 25764 -14332
rect 25764 -14388 25768 -14332
rect 25704 -14392 25768 -14388
rect 25704 -14652 25768 -14648
rect 25704 -14708 25708 -14652
rect 25708 -14708 25764 -14652
rect 25764 -14708 25768 -14652
rect 25704 -14712 25768 -14708
rect 25704 -14972 25768 -14968
rect 25704 -15028 25708 -14972
rect 25708 -15028 25764 -14972
rect 25764 -15028 25768 -14972
rect 25704 -15032 25768 -15028
rect 25704 -15292 25768 -15288
rect 25704 -15348 25708 -15292
rect 25708 -15348 25764 -15292
rect 25764 -15348 25768 -15292
rect 25704 -15352 25768 -15348
rect 25704 -15612 25768 -15608
rect 25704 -15668 25708 -15612
rect 25708 -15668 25764 -15612
rect 25764 -15668 25768 -15612
rect 25704 -15672 25768 -15668
rect 30608 -11246 30672 -11242
rect 30608 -11302 30612 -11246
rect 30612 -11302 30668 -11246
rect 30668 -11302 30672 -11246
rect 30608 -11306 30672 -11302
rect 30928 -11246 30992 -11242
rect 30928 -11302 30932 -11246
rect 30932 -11302 30988 -11246
rect 30988 -11302 30992 -11246
rect 30928 -11306 30992 -11302
rect 31248 -11246 31312 -11242
rect 31248 -11302 31252 -11246
rect 31252 -11302 31308 -11246
rect 31308 -11302 31312 -11246
rect 31248 -11306 31312 -11302
rect 31568 -11246 31632 -11242
rect 31568 -11302 31572 -11246
rect 31572 -11302 31628 -11246
rect 31628 -11302 31632 -11246
rect 31568 -11306 31632 -11302
rect 31888 -11246 31952 -11242
rect 31888 -11302 31892 -11246
rect 31892 -11302 31948 -11246
rect 31948 -11302 31952 -11246
rect 31888 -11306 31952 -11302
rect 32208 -11246 32272 -11242
rect 32208 -11302 32212 -11246
rect 32212 -11302 32268 -11246
rect 32268 -11302 32272 -11246
rect 32208 -11306 32272 -11302
rect 32528 -11246 32592 -11242
rect 32528 -11302 32532 -11246
rect 32532 -11302 32588 -11246
rect 32588 -11302 32592 -11246
rect 32528 -11306 32592 -11302
rect 32848 -11246 32912 -11242
rect 32848 -11302 32852 -11246
rect 32852 -11302 32908 -11246
rect 32908 -11302 32912 -11246
rect 32848 -11306 32912 -11302
rect 33168 -11246 33232 -11242
rect 33168 -11302 33172 -11246
rect 33172 -11302 33228 -11246
rect 33228 -11302 33232 -11246
rect 33168 -11306 33232 -11302
rect 33488 -11246 33552 -11242
rect 33488 -11302 33492 -11246
rect 33492 -11302 33548 -11246
rect 33548 -11302 33552 -11246
rect 33488 -11306 33552 -11302
rect 33808 -11246 33872 -11242
rect 33808 -11302 33812 -11246
rect 33812 -11302 33868 -11246
rect 33868 -11302 33872 -11246
rect 33808 -11306 33872 -11302
rect 34128 -11246 34192 -11242
rect 34128 -11302 34132 -11246
rect 34132 -11302 34188 -11246
rect 34188 -11302 34192 -11246
rect 34128 -11306 34192 -11302
rect 34448 -11246 34512 -11242
rect 34448 -11302 34452 -11246
rect 34452 -11302 34508 -11246
rect 34508 -11302 34512 -11246
rect 34448 -11306 34512 -11302
rect 34768 -11246 34832 -11242
rect 34768 -11302 34772 -11246
rect 34772 -11302 34828 -11246
rect 34828 -11302 34832 -11246
rect 34768 -11306 34832 -11302
rect 35088 -11246 35152 -11242
rect 35088 -11302 35092 -11246
rect 35092 -11302 35148 -11246
rect 35148 -11302 35152 -11246
rect 35088 -11306 35152 -11302
rect 35408 -11246 35472 -11242
rect 35408 -11302 35412 -11246
rect 35412 -11302 35468 -11246
rect 35468 -11302 35472 -11246
rect 35408 -11306 35472 -11302
rect 35728 -11246 35792 -11242
rect 35728 -11302 35732 -11246
rect 35732 -11302 35788 -11246
rect 35788 -11302 35792 -11246
rect 35728 -11306 35792 -11302
rect 36048 -11246 36112 -11242
rect 36048 -11302 36052 -11246
rect 36052 -11302 36108 -11246
rect 36108 -11302 36112 -11246
rect 36048 -11306 36112 -11302
rect 36368 -11246 36432 -11242
rect 36368 -11302 36372 -11246
rect 36372 -11302 36428 -11246
rect 36428 -11302 36432 -11246
rect 36368 -11306 36432 -11302
rect 36688 -11246 36752 -11242
rect 36688 -11302 36692 -11246
rect 36692 -11302 36748 -11246
rect 36748 -11302 36752 -11246
rect 36688 -11306 36752 -11302
rect 37008 -11246 37072 -11242
rect 37008 -11302 37012 -11246
rect 37012 -11302 37068 -11246
rect 37068 -11302 37072 -11246
rect 37008 -11306 37072 -11302
rect 37328 -11246 37392 -11242
rect 37328 -11302 37332 -11246
rect 37332 -11302 37388 -11246
rect 37388 -11302 37392 -11246
rect 37328 -11306 37392 -11302
rect 30238 -11452 30302 -11448
rect 30238 -11508 30242 -11452
rect 30242 -11508 30298 -11452
rect 30298 -11508 30302 -11452
rect 30238 -11512 30302 -11508
rect 37704 -11452 37768 -11448
rect 37704 -11508 37708 -11452
rect 37708 -11508 37764 -11452
rect 37764 -11508 37768 -11452
rect 37704 -11512 37768 -11508
rect 30238 -11772 30302 -11768
rect 30238 -11828 30242 -11772
rect 30242 -11828 30298 -11772
rect 30298 -11828 30302 -11772
rect 30238 -11832 30302 -11828
rect 30238 -12092 30302 -12088
rect 30238 -12148 30242 -12092
rect 30242 -12148 30298 -12092
rect 30298 -12148 30302 -12092
rect 30238 -12152 30302 -12148
rect 30238 -12412 30302 -12408
rect 30238 -12468 30242 -12412
rect 30242 -12468 30298 -12412
rect 30298 -12468 30302 -12412
rect 30238 -12472 30302 -12468
rect 30238 -12732 30302 -12728
rect 30238 -12788 30242 -12732
rect 30242 -12788 30298 -12732
rect 30298 -12788 30302 -12732
rect 30238 -12792 30302 -12788
rect 30238 -13052 30302 -13048
rect 30238 -13108 30242 -13052
rect 30242 -13108 30298 -13052
rect 30298 -13108 30302 -13052
rect 30238 -13112 30302 -13108
rect 30238 -13372 30302 -13368
rect 30238 -13428 30242 -13372
rect 30242 -13428 30298 -13372
rect 30298 -13428 30302 -13372
rect 30238 -13432 30302 -13428
rect 30238 -13692 30302 -13688
rect 30238 -13748 30242 -13692
rect 30242 -13748 30298 -13692
rect 30298 -13748 30302 -13692
rect 30238 -13752 30302 -13748
rect 30238 -14012 30302 -14008
rect 30238 -14068 30242 -14012
rect 30242 -14068 30298 -14012
rect 30298 -14068 30302 -14012
rect 30238 -14072 30302 -14068
rect 30238 -14332 30302 -14328
rect 30238 -14388 30242 -14332
rect 30242 -14388 30298 -14332
rect 30298 -14388 30302 -14332
rect 30238 -14392 30302 -14388
rect 30238 -14652 30302 -14648
rect 30238 -14708 30242 -14652
rect 30242 -14708 30298 -14652
rect 30298 -14708 30302 -14652
rect 30238 -14712 30302 -14708
rect 30238 -14972 30302 -14968
rect 30238 -15028 30242 -14972
rect 30242 -15028 30298 -14972
rect 30298 -15028 30302 -14972
rect 30238 -15032 30302 -15028
rect 30238 -15292 30302 -15288
rect 30238 -15348 30242 -15292
rect 30242 -15348 30298 -15292
rect 30298 -15348 30302 -15292
rect 30238 -15352 30302 -15348
rect 25704 -15932 25768 -15928
rect 25704 -15988 25708 -15932
rect 25708 -15988 25764 -15932
rect 25764 -15988 25768 -15932
rect 25704 -15992 25768 -15988
rect 25704 -16252 25768 -16248
rect 25704 -16308 25708 -16252
rect 25708 -16308 25764 -16252
rect 25764 -16308 25768 -16252
rect 25704 -16312 25768 -16308
rect 25704 -16572 25768 -16568
rect 25704 -16628 25708 -16572
rect 25708 -16628 25764 -16572
rect 25764 -16628 25768 -16572
rect 25704 -16632 25768 -16628
rect 25704 -16892 25768 -16888
rect 25704 -16948 25708 -16892
rect 25708 -16948 25764 -16892
rect 25764 -16948 25768 -16892
rect 25704 -16952 25768 -16948
rect 25704 -17212 25768 -17208
rect 25704 -17268 25708 -17212
rect 25708 -17268 25764 -17212
rect 25764 -17268 25768 -17212
rect 25704 -17272 25768 -17268
rect 25704 -17532 25768 -17528
rect 25704 -17588 25708 -17532
rect 25708 -17588 25764 -17532
rect 25764 -17588 25768 -17532
rect 25704 -17592 25768 -17588
rect 25704 -17852 25768 -17848
rect 25704 -17908 25708 -17852
rect 25708 -17908 25764 -17852
rect 25764 -17908 25768 -17852
rect 25704 -17912 25768 -17908
rect 25704 -18172 25768 -18168
rect 25704 -18228 25708 -18172
rect 25708 -18228 25764 -18172
rect 25764 -18228 25768 -18172
rect 25704 -18232 25768 -18228
rect 18238 -18492 18302 -18488
rect 18238 -18548 18242 -18492
rect 18242 -18548 18298 -18492
rect 18298 -18548 18302 -18492
rect 18238 -18552 18302 -18548
rect 25704 -18492 25768 -18488
rect 25704 -18548 25708 -18492
rect 25708 -18548 25764 -18492
rect 25764 -18548 25768 -18492
rect 25704 -18552 25768 -18548
rect 18608 -18702 18672 -18698
rect 18608 -18758 18612 -18702
rect 18612 -18758 18668 -18702
rect 18668 -18758 18672 -18702
rect 18608 -18762 18672 -18758
rect 18928 -18702 18992 -18698
rect 18928 -18758 18932 -18702
rect 18932 -18758 18988 -18702
rect 18988 -18758 18992 -18702
rect 18928 -18762 18992 -18758
rect 19248 -18702 19312 -18698
rect 19248 -18758 19252 -18702
rect 19252 -18758 19308 -18702
rect 19308 -18758 19312 -18702
rect 19248 -18762 19312 -18758
rect 19568 -18702 19632 -18698
rect 19568 -18758 19572 -18702
rect 19572 -18758 19628 -18702
rect 19628 -18758 19632 -18702
rect 19568 -18762 19632 -18758
rect 19888 -18702 19952 -18698
rect 19888 -18758 19892 -18702
rect 19892 -18758 19948 -18702
rect 19948 -18758 19952 -18702
rect 19888 -18762 19952 -18758
rect 20208 -18702 20272 -18698
rect 20208 -18758 20212 -18702
rect 20212 -18758 20268 -18702
rect 20268 -18758 20272 -18702
rect 20208 -18762 20272 -18758
rect 20528 -18702 20592 -18698
rect 20528 -18758 20532 -18702
rect 20532 -18758 20588 -18702
rect 20588 -18758 20592 -18702
rect 20528 -18762 20592 -18758
rect 20848 -18702 20912 -18698
rect 20848 -18758 20852 -18702
rect 20852 -18758 20908 -18702
rect 20908 -18758 20912 -18702
rect 20848 -18762 20912 -18758
rect 21168 -18702 21232 -18698
rect 21168 -18758 21172 -18702
rect 21172 -18758 21228 -18702
rect 21228 -18758 21232 -18702
rect 21168 -18762 21232 -18758
rect 21488 -18702 21552 -18698
rect 21488 -18758 21492 -18702
rect 21492 -18758 21548 -18702
rect 21548 -18758 21552 -18702
rect 21488 -18762 21552 -18758
rect 21808 -18702 21872 -18698
rect 21808 -18758 21812 -18702
rect 21812 -18758 21868 -18702
rect 21868 -18758 21872 -18702
rect 21808 -18762 21872 -18758
rect 22128 -18702 22192 -18698
rect 22128 -18758 22132 -18702
rect 22132 -18758 22188 -18702
rect 22188 -18758 22192 -18702
rect 22128 -18762 22192 -18758
rect 22448 -18702 22512 -18698
rect 22448 -18758 22452 -18702
rect 22452 -18758 22508 -18702
rect 22508 -18758 22512 -18702
rect 22448 -18762 22512 -18758
rect 22768 -18702 22832 -18698
rect 22768 -18758 22772 -18702
rect 22772 -18758 22828 -18702
rect 22828 -18758 22832 -18702
rect 22768 -18762 22832 -18758
rect 23088 -18702 23152 -18698
rect 23088 -18758 23092 -18702
rect 23092 -18758 23148 -18702
rect 23148 -18758 23152 -18702
rect 23088 -18762 23152 -18758
rect 23408 -18702 23472 -18698
rect 23408 -18758 23412 -18702
rect 23412 -18758 23468 -18702
rect 23468 -18758 23472 -18702
rect 23408 -18762 23472 -18758
rect 23728 -18702 23792 -18698
rect 23728 -18758 23732 -18702
rect 23732 -18758 23788 -18702
rect 23788 -18758 23792 -18702
rect 23728 -18762 23792 -18758
rect 24048 -18702 24112 -18698
rect 24048 -18758 24052 -18702
rect 24052 -18758 24108 -18702
rect 24108 -18758 24112 -18702
rect 24048 -18762 24112 -18758
rect 24368 -18702 24432 -18698
rect 24368 -18758 24372 -18702
rect 24372 -18758 24428 -18702
rect 24428 -18758 24432 -18702
rect 24368 -18762 24432 -18758
rect 24688 -18702 24752 -18698
rect 24688 -18758 24692 -18702
rect 24692 -18758 24748 -18702
rect 24748 -18758 24752 -18702
rect 24688 -18762 24752 -18758
rect 25008 -18702 25072 -18698
rect 25008 -18758 25012 -18702
rect 25012 -18758 25068 -18702
rect 25068 -18758 25072 -18702
rect 25008 -18762 25072 -18758
rect 25328 -18702 25392 -18698
rect 25328 -18758 25332 -18702
rect 25332 -18758 25388 -18702
rect 25388 -18758 25392 -18702
rect 25328 -18762 25392 -18758
rect 30238 -15612 30302 -15608
rect 30238 -15668 30242 -15612
rect 30242 -15668 30298 -15612
rect 30298 -15668 30302 -15612
rect 30238 -15672 30302 -15668
rect 30238 -15932 30302 -15928
rect 30238 -15988 30242 -15932
rect 30242 -15988 30298 -15932
rect 30298 -15988 30302 -15932
rect 30238 -15992 30302 -15988
rect 30238 -16252 30302 -16248
rect 30238 -16308 30242 -16252
rect 30242 -16308 30298 -16252
rect 30298 -16308 30302 -16252
rect 30238 -16312 30302 -16308
rect 30238 -16572 30302 -16568
rect 30238 -16628 30242 -16572
rect 30242 -16628 30298 -16572
rect 30298 -16628 30302 -16572
rect 30238 -16632 30302 -16628
rect 30238 -16892 30302 -16888
rect 30238 -16948 30242 -16892
rect 30242 -16948 30298 -16892
rect 30298 -16948 30302 -16892
rect 30238 -16952 30302 -16948
rect 30238 -17212 30302 -17208
rect 30238 -17268 30242 -17212
rect 30242 -17268 30298 -17212
rect 30298 -17268 30302 -17212
rect 30238 -17272 30302 -17268
rect 30238 -17532 30302 -17528
rect 30238 -17588 30242 -17532
rect 30242 -17588 30298 -17532
rect 30298 -17588 30302 -17532
rect 30238 -17592 30302 -17588
rect 30238 -17852 30302 -17848
rect 30238 -17908 30242 -17852
rect 30242 -17908 30298 -17852
rect 30298 -17908 30302 -17852
rect 30238 -17912 30302 -17908
rect 30238 -18172 30302 -18168
rect 30238 -18228 30242 -18172
rect 30242 -18228 30298 -18172
rect 30298 -18228 30302 -18172
rect 30238 -18232 30302 -18228
rect 37704 -11772 37768 -11768
rect 37704 -11828 37708 -11772
rect 37708 -11828 37764 -11772
rect 37764 -11828 37768 -11772
rect 37704 -11832 37768 -11828
rect 37704 -12092 37768 -12088
rect 37704 -12148 37708 -12092
rect 37708 -12148 37764 -12092
rect 37764 -12148 37768 -12092
rect 37704 -12152 37768 -12148
rect 37704 -12412 37768 -12408
rect 37704 -12468 37708 -12412
rect 37708 -12468 37764 -12412
rect 37764 -12468 37768 -12412
rect 37704 -12472 37768 -12468
rect 37704 -12732 37768 -12728
rect 37704 -12788 37708 -12732
rect 37708 -12788 37764 -12732
rect 37764 -12788 37768 -12732
rect 37704 -12792 37768 -12788
rect 37704 -13052 37768 -13048
rect 37704 -13108 37708 -13052
rect 37708 -13108 37764 -13052
rect 37764 -13108 37768 -13052
rect 37704 -13112 37768 -13108
rect 37704 -13372 37768 -13368
rect 37704 -13428 37708 -13372
rect 37708 -13428 37764 -13372
rect 37764 -13428 37768 -13372
rect 37704 -13432 37768 -13428
rect 37704 -13692 37768 -13688
rect 37704 -13748 37708 -13692
rect 37708 -13748 37764 -13692
rect 37764 -13748 37768 -13692
rect 37704 -13752 37768 -13748
rect 37704 -14012 37768 -14008
rect 37704 -14068 37708 -14012
rect 37708 -14068 37764 -14012
rect 37764 -14068 37768 -14012
rect 37704 -14072 37768 -14068
rect 37704 -14332 37768 -14328
rect 37704 -14388 37708 -14332
rect 37708 -14388 37764 -14332
rect 37764 -14388 37768 -14332
rect 37704 -14392 37768 -14388
rect 37704 -14652 37768 -14648
rect 37704 -14708 37708 -14652
rect 37708 -14708 37764 -14652
rect 37764 -14708 37768 -14652
rect 37704 -14712 37768 -14708
rect 37704 -14972 37768 -14968
rect 37704 -15028 37708 -14972
rect 37708 -15028 37764 -14972
rect 37764 -15028 37768 -14972
rect 37704 -15032 37768 -15028
rect 37704 -15292 37768 -15288
rect 37704 -15348 37708 -15292
rect 37708 -15348 37764 -15292
rect 37764 -15348 37768 -15292
rect 37704 -15352 37768 -15348
rect 37704 -15612 37768 -15608
rect 37704 -15668 37708 -15612
rect 37708 -15668 37764 -15612
rect 37764 -15668 37768 -15612
rect 37704 -15672 37768 -15668
rect 37704 -15932 37768 -15928
rect 37704 -15988 37708 -15932
rect 37708 -15988 37764 -15932
rect 37764 -15988 37768 -15932
rect 37704 -15992 37768 -15988
rect 37704 -16252 37768 -16248
rect 37704 -16308 37708 -16252
rect 37708 -16308 37764 -16252
rect 37764 -16308 37768 -16252
rect 37704 -16312 37768 -16308
rect 37704 -16572 37768 -16568
rect 37704 -16628 37708 -16572
rect 37708 -16628 37764 -16572
rect 37764 -16628 37768 -16572
rect 37704 -16632 37768 -16628
rect 37704 -16892 37768 -16888
rect 37704 -16948 37708 -16892
rect 37708 -16948 37764 -16892
rect 37764 -16948 37768 -16892
rect 37704 -16952 37768 -16948
rect 37704 -17212 37768 -17208
rect 37704 -17268 37708 -17212
rect 37708 -17268 37764 -17212
rect 37764 -17268 37768 -17212
rect 37704 -17272 37768 -17268
rect 37704 -17532 37768 -17528
rect 37704 -17588 37708 -17532
rect 37708 -17588 37764 -17532
rect 37764 -17588 37768 -17532
rect 37704 -17592 37768 -17588
rect 37704 -17852 37768 -17848
rect 37704 -17908 37708 -17852
rect 37708 -17908 37764 -17852
rect 37764 -17908 37768 -17852
rect 37704 -17912 37768 -17908
rect 37704 -18172 37768 -18168
rect 37704 -18228 37708 -18172
rect 37708 -18228 37764 -18172
rect 37764 -18228 37768 -18172
rect 37704 -18232 37768 -18228
rect 30238 -18492 30302 -18488
rect 30238 -18548 30242 -18492
rect 30242 -18548 30298 -18492
rect 30298 -18548 30302 -18492
rect 30238 -18552 30302 -18548
rect 37704 -18492 37768 -18488
rect 37704 -18548 37708 -18492
rect 37708 -18548 37764 -18492
rect 37764 -18548 37768 -18492
rect 37704 -18552 37768 -18548
rect 30608 -18702 30672 -18698
rect 30608 -18758 30612 -18702
rect 30612 -18758 30668 -18702
rect 30668 -18758 30672 -18702
rect 30608 -18762 30672 -18758
rect 30928 -18702 30992 -18698
rect 30928 -18758 30932 -18702
rect 30932 -18758 30988 -18702
rect 30988 -18758 30992 -18702
rect 30928 -18762 30992 -18758
rect 31248 -18702 31312 -18698
rect 31248 -18758 31252 -18702
rect 31252 -18758 31308 -18702
rect 31308 -18758 31312 -18702
rect 31248 -18762 31312 -18758
rect 31568 -18702 31632 -18698
rect 31568 -18758 31572 -18702
rect 31572 -18758 31628 -18702
rect 31628 -18758 31632 -18702
rect 31568 -18762 31632 -18758
rect 31888 -18702 31952 -18698
rect 31888 -18758 31892 -18702
rect 31892 -18758 31948 -18702
rect 31948 -18758 31952 -18702
rect 31888 -18762 31952 -18758
rect 32208 -18702 32272 -18698
rect 32208 -18758 32212 -18702
rect 32212 -18758 32268 -18702
rect 32268 -18758 32272 -18702
rect 32208 -18762 32272 -18758
rect 32528 -18702 32592 -18698
rect 32528 -18758 32532 -18702
rect 32532 -18758 32588 -18702
rect 32588 -18758 32592 -18702
rect 32528 -18762 32592 -18758
rect 32848 -18702 32912 -18698
rect 32848 -18758 32852 -18702
rect 32852 -18758 32908 -18702
rect 32908 -18758 32912 -18702
rect 32848 -18762 32912 -18758
rect 33168 -18702 33232 -18698
rect 33168 -18758 33172 -18702
rect 33172 -18758 33228 -18702
rect 33228 -18758 33232 -18702
rect 33168 -18762 33232 -18758
rect 33488 -18702 33552 -18698
rect 33488 -18758 33492 -18702
rect 33492 -18758 33548 -18702
rect 33548 -18758 33552 -18702
rect 33488 -18762 33552 -18758
rect 33808 -18702 33872 -18698
rect 33808 -18758 33812 -18702
rect 33812 -18758 33868 -18702
rect 33868 -18758 33872 -18702
rect 33808 -18762 33872 -18758
rect 34128 -18702 34192 -18698
rect 34128 -18758 34132 -18702
rect 34132 -18758 34188 -18702
rect 34188 -18758 34192 -18702
rect 34128 -18762 34192 -18758
rect 34448 -18702 34512 -18698
rect 34448 -18758 34452 -18702
rect 34452 -18758 34508 -18702
rect 34508 -18758 34512 -18702
rect 34448 -18762 34512 -18758
rect 34768 -18702 34832 -18698
rect 34768 -18758 34772 -18702
rect 34772 -18758 34828 -18702
rect 34828 -18758 34832 -18702
rect 34768 -18762 34832 -18758
rect 35088 -18702 35152 -18698
rect 35088 -18758 35092 -18702
rect 35092 -18758 35148 -18702
rect 35148 -18758 35152 -18702
rect 35088 -18762 35152 -18758
rect 35408 -18702 35472 -18698
rect 35408 -18758 35412 -18702
rect 35412 -18758 35468 -18702
rect 35468 -18758 35472 -18702
rect 35408 -18762 35472 -18758
rect 35728 -18702 35792 -18698
rect 35728 -18758 35732 -18702
rect 35732 -18758 35788 -18702
rect 35788 -18758 35792 -18702
rect 35728 -18762 35792 -18758
rect 36048 -18702 36112 -18698
rect 36048 -18758 36052 -18702
rect 36052 -18758 36108 -18702
rect 36108 -18758 36112 -18702
rect 36048 -18762 36112 -18758
rect 36368 -18702 36432 -18698
rect 36368 -18758 36372 -18702
rect 36372 -18758 36428 -18702
rect 36428 -18758 36432 -18702
rect 36368 -18762 36432 -18758
rect 36688 -18702 36752 -18698
rect 36688 -18758 36692 -18702
rect 36692 -18758 36748 -18702
rect 36748 -18758 36752 -18702
rect 36688 -18762 36752 -18758
rect 37008 -18702 37072 -18698
rect 37008 -18758 37012 -18702
rect 37012 -18758 37068 -18702
rect 37068 -18758 37072 -18702
rect 37008 -18762 37072 -18758
rect 37328 -18702 37392 -18698
rect 37328 -18758 37332 -18702
rect 37332 -18758 37388 -18702
rect 37388 -18758 37392 -18702
rect 37328 -18762 37392 -18758
rect 42608 -11246 42672 -11242
rect 42608 -11302 42612 -11246
rect 42612 -11302 42668 -11246
rect 42668 -11302 42672 -11246
rect 42608 -11306 42672 -11302
rect 42928 -11246 42992 -11242
rect 42928 -11302 42932 -11246
rect 42932 -11302 42988 -11246
rect 42988 -11302 42992 -11246
rect 42928 -11306 42992 -11302
rect 43248 -11246 43312 -11242
rect 43248 -11302 43252 -11246
rect 43252 -11302 43308 -11246
rect 43308 -11302 43312 -11246
rect 43248 -11306 43312 -11302
rect 43568 -11246 43632 -11242
rect 43568 -11302 43572 -11246
rect 43572 -11302 43628 -11246
rect 43628 -11302 43632 -11246
rect 43568 -11306 43632 -11302
rect 43888 -11246 43952 -11242
rect 43888 -11302 43892 -11246
rect 43892 -11302 43948 -11246
rect 43948 -11302 43952 -11246
rect 43888 -11306 43952 -11302
rect 44208 -11246 44272 -11242
rect 44208 -11302 44212 -11246
rect 44212 -11302 44268 -11246
rect 44268 -11302 44272 -11246
rect 44208 -11306 44272 -11302
rect 44528 -11246 44592 -11242
rect 44528 -11302 44532 -11246
rect 44532 -11302 44588 -11246
rect 44588 -11302 44592 -11246
rect 44528 -11306 44592 -11302
rect 44848 -11246 44912 -11242
rect 44848 -11302 44852 -11246
rect 44852 -11302 44908 -11246
rect 44908 -11302 44912 -11246
rect 44848 -11306 44912 -11302
rect 45168 -11246 45232 -11242
rect 45168 -11302 45172 -11246
rect 45172 -11302 45228 -11246
rect 45228 -11302 45232 -11246
rect 45168 -11306 45232 -11302
rect 45488 -11246 45552 -11242
rect 45488 -11302 45492 -11246
rect 45492 -11302 45548 -11246
rect 45548 -11302 45552 -11246
rect 45488 -11306 45552 -11302
rect 45808 -11246 45872 -11242
rect 45808 -11302 45812 -11246
rect 45812 -11302 45868 -11246
rect 45868 -11302 45872 -11246
rect 45808 -11306 45872 -11302
rect 46128 -11246 46192 -11242
rect 46128 -11302 46132 -11246
rect 46132 -11302 46188 -11246
rect 46188 -11302 46192 -11246
rect 46128 -11306 46192 -11302
rect 46448 -11246 46512 -11242
rect 46448 -11302 46452 -11246
rect 46452 -11302 46508 -11246
rect 46508 -11302 46512 -11246
rect 46448 -11306 46512 -11302
rect 46768 -11246 46832 -11242
rect 46768 -11302 46772 -11246
rect 46772 -11302 46828 -11246
rect 46828 -11302 46832 -11246
rect 46768 -11306 46832 -11302
rect 47088 -11246 47152 -11242
rect 47088 -11302 47092 -11246
rect 47092 -11302 47148 -11246
rect 47148 -11302 47152 -11246
rect 47088 -11306 47152 -11302
rect 47408 -11246 47472 -11242
rect 47408 -11302 47412 -11246
rect 47412 -11302 47468 -11246
rect 47468 -11302 47472 -11246
rect 47408 -11306 47472 -11302
rect 47728 -11246 47792 -11242
rect 47728 -11302 47732 -11246
rect 47732 -11302 47788 -11246
rect 47788 -11302 47792 -11246
rect 47728 -11306 47792 -11302
rect 48048 -11246 48112 -11242
rect 48048 -11302 48052 -11246
rect 48052 -11302 48108 -11246
rect 48108 -11302 48112 -11246
rect 48048 -11306 48112 -11302
rect 48368 -11246 48432 -11242
rect 48368 -11302 48372 -11246
rect 48372 -11302 48428 -11246
rect 48428 -11302 48432 -11246
rect 48368 -11306 48432 -11302
rect 48688 -11246 48752 -11242
rect 48688 -11302 48692 -11246
rect 48692 -11302 48748 -11246
rect 48748 -11302 48752 -11246
rect 48688 -11306 48752 -11302
rect 49008 -11246 49072 -11242
rect 49008 -11302 49012 -11246
rect 49012 -11302 49068 -11246
rect 49068 -11302 49072 -11246
rect 49008 -11306 49072 -11302
rect 49328 -11246 49392 -11242
rect 49328 -11302 49332 -11246
rect 49332 -11302 49388 -11246
rect 49388 -11302 49392 -11246
rect 49328 -11306 49392 -11302
rect 42238 -11452 42302 -11448
rect 42238 -11508 42242 -11452
rect 42242 -11508 42298 -11452
rect 42298 -11508 42302 -11452
rect 42238 -11512 42302 -11508
rect 49704 -11452 49768 -11448
rect 49704 -11508 49708 -11452
rect 49708 -11508 49764 -11452
rect 49764 -11508 49768 -11452
rect 49704 -11512 49768 -11508
rect 42238 -11772 42302 -11768
rect 42238 -11828 42242 -11772
rect 42242 -11828 42298 -11772
rect 42298 -11828 42302 -11772
rect 42238 -11832 42302 -11828
rect 42238 -12092 42302 -12088
rect 42238 -12148 42242 -12092
rect 42242 -12148 42298 -12092
rect 42298 -12148 42302 -12092
rect 42238 -12152 42302 -12148
rect 42238 -12412 42302 -12408
rect 42238 -12468 42242 -12412
rect 42242 -12468 42298 -12412
rect 42298 -12468 42302 -12412
rect 42238 -12472 42302 -12468
rect 42238 -12732 42302 -12728
rect 42238 -12788 42242 -12732
rect 42242 -12788 42298 -12732
rect 42298 -12788 42302 -12732
rect 42238 -12792 42302 -12788
rect 42238 -13052 42302 -13048
rect 42238 -13108 42242 -13052
rect 42242 -13108 42298 -13052
rect 42298 -13108 42302 -13052
rect 42238 -13112 42302 -13108
rect 42238 -13372 42302 -13368
rect 42238 -13428 42242 -13372
rect 42242 -13428 42298 -13372
rect 42298 -13428 42302 -13372
rect 42238 -13432 42302 -13428
rect 42238 -13692 42302 -13688
rect 42238 -13748 42242 -13692
rect 42242 -13748 42298 -13692
rect 42298 -13748 42302 -13692
rect 42238 -13752 42302 -13748
rect 42238 -14012 42302 -14008
rect 42238 -14068 42242 -14012
rect 42242 -14068 42298 -14012
rect 42298 -14068 42302 -14012
rect 42238 -14072 42302 -14068
rect 42238 -14332 42302 -14328
rect 42238 -14388 42242 -14332
rect 42242 -14388 42298 -14332
rect 42298 -14388 42302 -14332
rect 42238 -14392 42302 -14388
rect 42238 -14652 42302 -14648
rect 42238 -14708 42242 -14652
rect 42242 -14708 42298 -14652
rect 42298 -14708 42302 -14652
rect 42238 -14712 42302 -14708
rect 42238 -14972 42302 -14968
rect 42238 -15028 42242 -14972
rect 42242 -15028 42298 -14972
rect 42298 -15028 42302 -14972
rect 42238 -15032 42302 -15028
rect 42238 -15292 42302 -15288
rect 42238 -15348 42242 -15292
rect 42242 -15348 42298 -15292
rect 42298 -15348 42302 -15292
rect 42238 -15352 42302 -15348
rect 42238 -15612 42302 -15608
rect 42238 -15668 42242 -15612
rect 42242 -15668 42298 -15612
rect 42298 -15668 42302 -15612
rect 42238 -15672 42302 -15668
rect 42238 -15932 42302 -15928
rect 42238 -15988 42242 -15932
rect 42242 -15988 42298 -15932
rect 42298 -15988 42302 -15932
rect 42238 -15992 42302 -15988
rect 42238 -16252 42302 -16248
rect 42238 -16308 42242 -16252
rect 42242 -16308 42298 -16252
rect 42298 -16308 42302 -16252
rect 42238 -16312 42302 -16308
rect 42238 -16572 42302 -16568
rect 42238 -16628 42242 -16572
rect 42242 -16628 42298 -16572
rect 42298 -16628 42302 -16572
rect 42238 -16632 42302 -16628
rect 42238 -16892 42302 -16888
rect 42238 -16948 42242 -16892
rect 42242 -16948 42298 -16892
rect 42298 -16948 42302 -16892
rect 42238 -16952 42302 -16948
rect 42238 -17212 42302 -17208
rect 42238 -17268 42242 -17212
rect 42242 -17268 42298 -17212
rect 42298 -17268 42302 -17212
rect 42238 -17272 42302 -17268
rect 42238 -17532 42302 -17528
rect 42238 -17588 42242 -17532
rect 42242 -17588 42298 -17532
rect 42298 -17588 42302 -17532
rect 42238 -17592 42302 -17588
rect 42238 -17852 42302 -17848
rect 42238 -17908 42242 -17852
rect 42242 -17908 42298 -17852
rect 42298 -17908 42302 -17852
rect 42238 -17912 42302 -17908
rect 42238 -18172 42302 -18168
rect 42238 -18228 42242 -18172
rect 42242 -18228 42298 -18172
rect 42298 -18228 42302 -18172
rect 42238 -18232 42302 -18228
rect 49704 -11772 49768 -11768
rect 49704 -11828 49708 -11772
rect 49708 -11828 49764 -11772
rect 49764 -11828 49768 -11772
rect 49704 -11832 49768 -11828
rect 49704 -12092 49768 -12088
rect 49704 -12148 49708 -12092
rect 49708 -12148 49764 -12092
rect 49764 -12148 49768 -12092
rect 49704 -12152 49768 -12148
rect 49704 -12412 49768 -12408
rect 49704 -12468 49708 -12412
rect 49708 -12468 49764 -12412
rect 49764 -12468 49768 -12412
rect 49704 -12472 49768 -12468
rect 49704 -12732 49768 -12728
rect 49704 -12788 49708 -12732
rect 49708 -12788 49764 -12732
rect 49764 -12788 49768 -12732
rect 49704 -12792 49768 -12788
rect 49704 -13052 49768 -13048
rect 49704 -13108 49708 -13052
rect 49708 -13108 49764 -13052
rect 49764 -13108 49768 -13052
rect 49704 -13112 49768 -13108
rect 49704 -13372 49768 -13368
rect 49704 -13428 49708 -13372
rect 49708 -13428 49764 -13372
rect 49764 -13428 49768 -13372
rect 49704 -13432 49768 -13428
rect 49704 -13692 49768 -13688
rect 49704 -13748 49708 -13692
rect 49708 -13748 49764 -13692
rect 49764 -13748 49768 -13692
rect 49704 -13752 49768 -13748
rect 49704 -14012 49768 -14008
rect 49704 -14068 49708 -14012
rect 49708 -14068 49764 -14012
rect 49764 -14068 49768 -14012
rect 49704 -14072 49768 -14068
rect 49704 -14332 49768 -14328
rect 49704 -14388 49708 -14332
rect 49708 -14388 49764 -14332
rect 49764 -14388 49768 -14332
rect 49704 -14392 49768 -14388
rect 49704 -14652 49768 -14648
rect 49704 -14708 49708 -14652
rect 49708 -14708 49764 -14652
rect 49764 -14708 49768 -14652
rect 49704 -14712 49768 -14708
rect 49704 -14972 49768 -14968
rect 49704 -15028 49708 -14972
rect 49708 -15028 49764 -14972
rect 49764 -15028 49768 -14972
rect 49704 -15032 49768 -15028
rect 49704 -15292 49768 -15288
rect 49704 -15348 49708 -15292
rect 49708 -15348 49764 -15292
rect 49764 -15348 49768 -15292
rect 49704 -15352 49768 -15348
rect 49704 -15612 49768 -15608
rect 49704 -15668 49708 -15612
rect 49708 -15668 49764 -15612
rect 49764 -15668 49768 -15612
rect 49704 -15672 49768 -15668
rect 49704 -15932 49768 -15928
rect 49704 -15988 49708 -15932
rect 49708 -15988 49764 -15932
rect 49764 -15988 49768 -15932
rect 49704 -15992 49768 -15988
rect 49704 -16252 49768 -16248
rect 49704 -16308 49708 -16252
rect 49708 -16308 49764 -16252
rect 49764 -16308 49768 -16252
rect 49704 -16312 49768 -16308
rect 49704 -16572 49768 -16568
rect 49704 -16628 49708 -16572
rect 49708 -16628 49764 -16572
rect 49764 -16628 49768 -16572
rect 49704 -16632 49768 -16628
rect 49704 -16892 49768 -16888
rect 49704 -16948 49708 -16892
rect 49708 -16948 49764 -16892
rect 49764 -16948 49768 -16892
rect 49704 -16952 49768 -16948
rect 49704 -17212 49768 -17208
rect 49704 -17268 49708 -17212
rect 49708 -17268 49764 -17212
rect 49764 -17268 49768 -17212
rect 49704 -17272 49768 -17268
rect 49704 -17532 49768 -17528
rect 49704 -17588 49708 -17532
rect 49708 -17588 49764 -17532
rect 49764 -17588 49768 -17532
rect 49704 -17592 49768 -17588
rect 49704 -17852 49768 -17848
rect 49704 -17908 49708 -17852
rect 49708 -17908 49764 -17852
rect 49764 -17908 49768 -17852
rect 49704 -17912 49768 -17908
rect 49704 -18172 49768 -18168
rect 49704 -18228 49708 -18172
rect 49708 -18228 49764 -18172
rect 49764 -18228 49768 -18172
rect 49704 -18232 49768 -18228
rect 42238 -18492 42302 -18488
rect 42238 -18548 42242 -18492
rect 42242 -18548 42298 -18492
rect 42298 -18548 42302 -18492
rect 42238 -18552 42302 -18548
rect 49704 -18492 49768 -18488
rect 49704 -18548 49708 -18492
rect 49708 -18548 49764 -18492
rect 49764 -18548 49768 -18492
rect 49704 -18552 49768 -18548
rect 42608 -18702 42672 -18698
rect 42608 -18758 42612 -18702
rect 42612 -18758 42668 -18702
rect 42668 -18758 42672 -18702
rect 42608 -18762 42672 -18758
rect 42928 -18702 42992 -18698
rect 42928 -18758 42932 -18702
rect 42932 -18758 42988 -18702
rect 42988 -18758 42992 -18702
rect 42928 -18762 42992 -18758
rect 43248 -18702 43312 -18698
rect 43248 -18758 43252 -18702
rect 43252 -18758 43308 -18702
rect 43308 -18758 43312 -18702
rect 43248 -18762 43312 -18758
rect 43568 -18702 43632 -18698
rect 43568 -18758 43572 -18702
rect 43572 -18758 43628 -18702
rect 43628 -18758 43632 -18702
rect 43568 -18762 43632 -18758
rect 43888 -18702 43952 -18698
rect 43888 -18758 43892 -18702
rect 43892 -18758 43948 -18702
rect 43948 -18758 43952 -18702
rect 43888 -18762 43952 -18758
rect 44208 -18702 44272 -18698
rect 44208 -18758 44212 -18702
rect 44212 -18758 44268 -18702
rect 44268 -18758 44272 -18702
rect 44208 -18762 44272 -18758
rect 44528 -18702 44592 -18698
rect 44528 -18758 44532 -18702
rect 44532 -18758 44588 -18702
rect 44588 -18758 44592 -18702
rect 44528 -18762 44592 -18758
rect 44848 -18702 44912 -18698
rect 44848 -18758 44852 -18702
rect 44852 -18758 44908 -18702
rect 44908 -18758 44912 -18702
rect 44848 -18762 44912 -18758
rect 45168 -18702 45232 -18698
rect 45168 -18758 45172 -18702
rect 45172 -18758 45228 -18702
rect 45228 -18758 45232 -18702
rect 45168 -18762 45232 -18758
rect 45488 -18702 45552 -18698
rect 45488 -18758 45492 -18702
rect 45492 -18758 45548 -18702
rect 45548 -18758 45552 -18702
rect 45488 -18762 45552 -18758
rect 45808 -18702 45872 -18698
rect 45808 -18758 45812 -18702
rect 45812 -18758 45868 -18702
rect 45868 -18758 45872 -18702
rect 45808 -18762 45872 -18758
rect 46128 -18702 46192 -18698
rect 46128 -18758 46132 -18702
rect 46132 -18758 46188 -18702
rect 46188 -18758 46192 -18702
rect 46128 -18762 46192 -18758
rect 46448 -18702 46512 -18698
rect 46448 -18758 46452 -18702
rect 46452 -18758 46508 -18702
rect 46508 -18758 46512 -18702
rect 46448 -18762 46512 -18758
rect 46768 -18702 46832 -18698
rect 46768 -18758 46772 -18702
rect 46772 -18758 46828 -18702
rect 46828 -18758 46832 -18702
rect 46768 -18762 46832 -18758
rect 47088 -18702 47152 -18698
rect 47088 -18758 47092 -18702
rect 47092 -18758 47148 -18702
rect 47148 -18758 47152 -18702
rect 47088 -18762 47152 -18758
rect 47408 -18702 47472 -18698
rect 47408 -18758 47412 -18702
rect 47412 -18758 47468 -18702
rect 47468 -18758 47472 -18702
rect 47408 -18762 47472 -18758
rect 47728 -18702 47792 -18698
rect 47728 -18758 47732 -18702
rect 47732 -18758 47788 -18702
rect 47788 -18758 47792 -18702
rect 47728 -18762 47792 -18758
rect 48048 -18702 48112 -18698
rect 48048 -18758 48052 -18702
rect 48052 -18758 48108 -18702
rect 48108 -18758 48112 -18702
rect 48048 -18762 48112 -18758
rect 48368 -18702 48432 -18698
rect 48368 -18758 48372 -18702
rect 48372 -18758 48428 -18702
rect 48428 -18758 48432 -18702
rect 48368 -18762 48432 -18758
rect 48688 -18702 48752 -18698
rect 48688 -18758 48692 -18702
rect 48692 -18758 48748 -18702
rect 48748 -18758 48752 -18702
rect 48688 -18762 48752 -18758
rect 49008 -18702 49072 -18698
rect 49008 -18758 49012 -18702
rect 49012 -18758 49068 -18702
rect 49068 -18758 49072 -18702
rect 49008 -18762 49072 -18758
rect 49328 -18702 49392 -18698
rect 49328 -18758 49332 -18702
rect 49332 -18758 49388 -18702
rect 49388 -18758 49392 -18702
rect 49328 -18762 49392 -18758
rect 18608 -23246 18672 -23242
rect 18608 -23302 18612 -23246
rect 18612 -23302 18668 -23246
rect 18668 -23302 18672 -23246
rect 18608 -23306 18672 -23302
rect 18928 -23246 18992 -23242
rect 18928 -23302 18932 -23246
rect 18932 -23302 18988 -23246
rect 18988 -23302 18992 -23246
rect 18928 -23306 18992 -23302
rect 19248 -23246 19312 -23242
rect 19248 -23302 19252 -23246
rect 19252 -23302 19308 -23246
rect 19308 -23302 19312 -23246
rect 19248 -23306 19312 -23302
rect 19568 -23246 19632 -23242
rect 19568 -23302 19572 -23246
rect 19572 -23302 19628 -23246
rect 19628 -23302 19632 -23246
rect 19568 -23306 19632 -23302
rect 19888 -23246 19952 -23242
rect 19888 -23302 19892 -23246
rect 19892 -23302 19948 -23246
rect 19948 -23302 19952 -23246
rect 19888 -23306 19952 -23302
rect 20208 -23246 20272 -23242
rect 20208 -23302 20212 -23246
rect 20212 -23302 20268 -23246
rect 20268 -23302 20272 -23246
rect 20208 -23306 20272 -23302
rect 20528 -23246 20592 -23242
rect 20528 -23302 20532 -23246
rect 20532 -23302 20588 -23246
rect 20588 -23302 20592 -23246
rect 20528 -23306 20592 -23302
rect 20848 -23246 20912 -23242
rect 20848 -23302 20852 -23246
rect 20852 -23302 20908 -23246
rect 20908 -23302 20912 -23246
rect 20848 -23306 20912 -23302
rect 21168 -23246 21232 -23242
rect 21168 -23302 21172 -23246
rect 21172 -23302 21228 -23246
rect 21228 -23302 21232 -23246
rect 21168 -23306 21232 -23302
rect 21488 -23246 21552 -23242
rect 21488 -23302 21492 -23246
rect 21492 -23302 21548 -23246
rect 21548 -23302 21552 -23246
rect 21488 -23306 21552 -23302
rect 21808 -23246 21872 -23242
rect 21808 -23302 21812 -23246
rect 21812 -23302 21868 -23246
rect 21868 -23302 21872 -23246
rect 21808 -23306 21872 -23302
rect 22128 -23246 22192 -23242
rect 22128 -23302 22132 -23246
rect 22132 -23302 22188 -23246
rect 22188 -23302 22192 -23246
rect 22128 -23306 22192 -23302
rect 22448 -23246 22512 -23242
rect 22448 -23302 22452 -23246
rect 22452 -23302 22508 -23246
rect 22508 -23302 22512 -23246
rect 22448 -23306 22512 -23302
rect 22768 -23246 22832 -23242
rect 22768 -23302 22772 -23246
rect 22772 -23302 22828 -23246
rect 22828 -23302 22832 -23246
rect 22768 -23306 22832 -23302
rect 23088 -23246 23152 -23242
rect 23088 -23302 23092 -23246
rect 23092 -23302 23148 -23246
rect 23148 -23302 23152 -23246
rect 23088 -23306 23152 -23302
rect 23408 -23246 23472 -23242
rect 23408 -23302 23412 -23246
rect 23412 -23302 23468 -23246
rect 23468 -23302 23472 -23246
rect 23408 -23306 23472 -23302
rect 23728 -23246 23792 -23242
rect 23728 -23302 23732 -23246
rect 23732 -23302 23788 -23246
rect 23788 -23302 23792 -23246
rect 23728 -23306 23792 -23302
rect 24048 -23246 24112 -23242
rect 24048 -23302 24052 -23246
rect 24052 -23302 24108 -23246
rect 24108 -23302 24112 -23246
rect 24048 -23306 24112 -23302
rect 24368 -23246 24432 -23242
rect 24368 -23302 24372 -23246
rect 24372 -23302 24428 -23246
rect 24428 -23302 24432 -23246
rect 24368 -23306 24432 -23302
rect 24688 -23246 24752 -23242
rect 24688 -23302 24692 -23246
rect 24692 -23302 24748 -23246
rect 24748 -23302 24752 -23246
rect 24688 -23306 24752 -23302
rect 25008 -23246 25072 -23242
rect 25008 -23302 25012 -23246
rect 25012 -23302 25068 -23246
rect 25068 -23302 25072 -23246
rect 25008 -23306 25072 -23302
rect 25328 -23246 25392 -23242
rect 25328 -23302 25332 -23246
rect 25332 -23302 25388 -23246
rect 25388 -23302 25392 -23246
rect 25328 -23306 25392 -23302
rect 18238 -23452 18302 -23448
rect 18238 -23508 18242 -23452
rect 18242 -23508 18298 -23452
rect 18298 -23508 18302 -23452
rect 18238 -23512 18302 -23508
rect 25704 -23452 25768 -23448
rect 25704 -23508 25708 -23452
rect 25708 -23508 25764 -23452
rect 25764 -23508 25768 -23452
rect 25704 -23512 25768 -23508
rect 18238 -23772 18302 -23768
rect 18238 -23828 18242 -23772
rect 18242 -23828 18298 -23772
rect 18298 -23828 18302 -23772
rect 18238 -23832 18302 -23828
rect 18238 -24092 18302 -24088
rect 18238 -24148 18242 -24092
rect 18242 -24148 18298 -24092
rect 18298 -24148 18302 -24092
rect 18238 -24152 18302 -24148
rect 18238 -24412 18302 -24408
rect 18238 -24468 18242 -24412
rect 18242 -24468 18298 -24412
rect 18298 -24468 18302 -24412
rect 18238 -24472 18302 -24468
rect 18238 -24732 18302 -24728
rect 18238 -24788 18242 -24732
rect 18242 -24788 18298 -24732
rect 18298 -24788 18302 -24732
rect 18238 -24792 18302 -24788
rect 18238 -25052 18302 -25048
rect 18238 -25108 18242 -25052
rect 18242 -25108 18298 -25052
rect 18298 -25108 18302 -25052
rect 18238 -25112 18302 -25108
rect 18238 -25372 18302 -25368
rect 18238 -25428 18242 -25372
rect 18242 -25428 18298 -25372
rect 18298 -25428 18302 -25372
rect 18238 -25432 18302 -25428
rect 18238 -25692 18302 -25688
rect 18238 -25748 18242 -25692
rect 18242 -25748 18298 -25692
rect 18298 -25748 18302 -25692
rect 18238 -25752 18302 -25748
rect 13704 -26012 13768 -26008
rect 13704 -26068 13708 -26012
rect 13708 -26068 13764 -26012
rect 13764 -26068 13768 -26012
rect 13704 -26072 13768 -26068
rect 13704 -26332 13768 -26328
rect 13704 -26388 13708 -26332
rect 13708 -26388 13764 -26332
rect 13764 -26388 13768 -26332
rect 13704 -26392 13768 -26388
rect 13704 -26652 13768 -26648
rect 13704 -26708 13708 -26652
rect 13708 -26708 13764 -26652
rect 13764 -26708 13768 -26652
rect 13704 -26712 13768 -26708
rect 13704 -26972 13768 -26968
rect 13704 -27028 13708 -26972
rect 13708 -27028 13764 -26972
rect 13764 -27028 13768 -26972
rect 13704 -27032 13768 -27028
rect 13704 -27292 13768 -27288
rect 13704 -27348 13708 -27292
rect 13708 -27348 13764 -27292
rect 13764 -27348 13768 -27292
rect 13704 -27352 13768 -27348
rect 13704 -27612 13768 -27608
rect 13704 -27668 13708 -27612
rect 13708 -27668 13764 -27612
rect 13764 -27668 13768 -27612
rect 13704 -27672 13768 -27668
rect 13704 -27932 13768 -27928
rect 13704 -27988 13708 -27932
rect 13708 -27988 13764 -27932
rect 13764 -27988 13768 -27932
rect 13704 -27992 13768 -27988
rect 13704 -28252 13768 -28248
rect 13704 -28308 13708 -28252
rect 13708 -28308 13764 -28252
rect 13764 -28308 13768 -28252
rect 13704 -28312 13768 -28308
rect 13704 -28572 13768 -28568
rect 13704 -28628 13708 -28572
rect 13708 -28628 13764 -28572
rect 13764 -28628 13768 -28572
rect 13704 -28632 13768 -28628
rect 13704 -28892 13768 -28888
rect 13704 -28948 13708 -28892
rect 13708 -28948 13764 -28892
rect 13764 -28948 13768 -28892
rect 13704 -28952 13768 -28948
rect 13704 -29212 13768 -29208
rect 13704 -29268 13708 -29212
rect 13708 -29268 13764 -29212
rect 13764 -29268 13768 -29212
rect 13704 -29272 13768 -29268
rect 13704 -29532 13768 -29528
rect 13704 -29588 13708 -29532
rect 13708 -29588 13764 -29532
rect 13764 -29588 13768 -29532
rect 13704 -29592 13768 -29588
rect 13704 -29852 13768 -29848
rect 13704 -29908 13708 -29852
rect 13708 -29908 13764 -29852
rect 13764 -29908 13768 -29852
rect 13704 -29912 13768 -29908
rect 13704 -30172 13768 -30168
rect 13704 -30228 13708 -30172
rect 13708 -30228 13764 -30172
rect 13764 -30228 13768 -30172
rect 13704 -30232 13768 -30228
rect 6238 -30492 6302 -30488
rect 6238 -30548 6242 -30492
rect 6242 -30548 6298 -30492
rect 6298 -30548 6302 -30492
rect 6238 -30552 6302 -30548
rect 13704 -30492 13768 -30488
rect 13704 -30548 13708 -30492
rect 13708 -30548 13764 -30492
rect 13764 -30548 13768 -30492
rect 13704 -30552 13768 -30548
rect 6608 -30702 6672 -30698
rect 6608 -30758 6612 -30702
rect 6612 -30758 6668 -30702
rect 6668 -30758 6672 -30702
rect 6608 -30762 6672 -30758
rect 6928 -30702 6992 -30698
rect 6928 -30758 6932 -30702
rect 6932 -30758 6988 -30702
rect 6988 -30758 6992 -30702
rect 6928 -30762 6992 -30758
rect 7248 -30702 7312 -30698
rect 7248 -30758 7252 -30702
rect 7252 -30758 7308 -30702
rect 7308 -30758 7312 -30702
rect 7248 -30762 7312 -30758
rect 7568 -30702 7632 -30698
rect 7568 -30758 7572 -30702
rect 7572 -30758 7628 -30702
rect 7628 -30758 7632 -30702
rect 7568 -30762 7632 -30758
rect 7888 -30702 7952 -30698
rect 7888 -30758 7892 -30702
rect 7892 -30758 7948 -30702
rect 7948 -30758 7952 -30702
rect 7888 -30762 7952 -30758
rect 8208 -30702 8272 -30698
rect 8208 -30758 8212 -30702
rect 8212 -30758 8268 -30702
rect 8268 -30758 8272 -30702
rect 8208 -30762 8272 -30758
rect 8528 -30702 8592 -30698
rect 8528 -30758 8532 -30702
rect 8532 -30758 8588 -30702
rect 8588 -30758 8592 -30702
rect 8528 -30762 8592 -30758
rect 8848 -30702 8912 -30698
rect 8848 -30758 8852 -30702
rect 8852 -30758 8908 -30702
rect 8908 -30758 8912 -30702
rect 8848 -30762 8912 -30758
rect 9168 -30702 9232 -30698
rect 9168 -30758 9172 -30702
rect 9172 -30758 9228 -30702
rect 9228 -30758 9232 -30702
rect 9168 -30762 9232 -30758
rect 9488 -30702 9552 -30698
rect 9488 -30758 9492 -30702
rect 9492 -30758 9548 -30702
rect 9548 -30758 9552 -30702
rect 9488 -30762 9552 -30758
rect 9808 -30702 9872 -30698
rect 9808 -30758 9812 -30702
rect 9812 -30758 9868 -30702
rect 9868 -30758 9872 -30702
rect 9808 -30762 9872 -30758
rect 10128 -30702 10192 -30698
rect 10128 -30758 10132 -30702
rect 10132 -30758 10188 -30702
rect 10188 -30758 10192 -30702
rect 10128 -30762 10192 -30758
rect 10448 -30702 10512 -30698
rect 10448 -30758 10452 -30702
rect 10452 -30758 10508 -30702
rect 10508 -30758 10512 -30702
rect 10448 -30762 10512 -30758
rect 10768 -30702 10832 -30698
rect 10768 -30758 10772 -30702
rect 10772 -30758 10828 -30702
rect 10828 -30758 10832 -30702
rect 10768 -30762 10832 -30758
rect 11088 -30702 11152 -30698
rect 11088 -30758 11092 -30702
rect 11092 -30758 11148 -30702
rect 11148 -30758 11152 -30702
rect 11088 -30762 11152 -30758
rect 11408 -30702 11472 -30698
rect 11408 -30758 11412 -30702
rect 11412 -30758 11468 -30702
rect 11468 -30758 11472 -30702
rect 11408 -30762 11472 -30758
rect 11728 -30702 11792 -30698
rect 11728 -30758 11732 -30702
rect 11732 -30758 11788 -30702
rect 11788 -30758 11792 -30702
rect 11728 -30762 11792 -30758
rect 12048 -30702 12112 -30698
rect 12048 -30758 12052 -30702
rect 12052 -30758 12108 -30702
rect 12108 -30758 12112 -30702
rect 12048 -30762 12112 -30758
rect 12368 -30702 12432 -30698
rect 12368 -30758 12372 -30702
rect 12372 -30758 12428 -30702
rect 12428 -30758 12432 -30702
rect 12368 -30762 12432 -30758
rect 12688 -30702 12752 -30698
rect 12688 -30758 12692 -30702
rect 12692 -30758 12748 -30702
rect 12748 -30758 12752 -30702
rect 12688 -30762 12752 -30758
rect 13008 -30702 13072 -30698
rect 13008 -30758 13012 -30702
rect 13012 -30758 13068 -30702
rect 13068 -30758 13072 -30702
rect 13008 -30762 13072 -30758
rect 13328 -30702 13392 -30698
rect 13328 -30758 13332 -30702
rect 13332 -30758 13388 -30702
rect 13388 -30758 13392 -30702
rect 13328 -30762 13392 -30758
rect 18238 -26012 18302 -26008
rect 18238 -26068 18242 -26012
rect 18242 -26068 18298 -26012
rect 18298 -26068 18302 -26012
rect 18238 -26072 18302 -26068
rect 18238 -26332 18302 -26328
rect 18238 -26388 18242 -26332
rect 18242 -26388 18298 -26332
rect 18298 -26388 18302 -26332
rect 18238 -26392 18302 -26388
rect 18238 -26652 18302 -26648
rect 18238 -26708 18242 -26652
rect 18242 -26708 18298 -26652
rect 18298 -26708 18302 -26652
rect 18238 -26712 18302 -26708
rect 18238 -26972 18302 -26968
rect 18238 -27028 18242 -26972
rect 18242 -27028 18298 -26972
rect 18298 -27028 18302 -26972
rect 18238 -27032 18302 -27028
rect 18238 -27292 18302 -27288
rect 18238 -27348 18242 -27292
rect 18242 -27348 18298 -27292
rect 18298 -27348 18302 -27292
rect 18238 -27352 18302 -27348
rect 18238 -27612 18302 -27608
rect 18238 -27668 18242 -27612
rect 18242 -27668 18298 -27612
rect 18298 -27668 18302 -27612
rect 18238 -27672 18302 -27668
rect 18238 -27932 18302 -27928
rect 18238 -27988 18242 -27932
rect 18242 -27988 18298 -27932
rect 18298 -27988 18302 -27932
rect 18238 -27992 18302 -27988
rect 18238 -28252 18302 -28248
rect 18238 -28308 18242 -28252
rect 18242 -28308 18298 -28252
rect 18298 -28308 18302 -28252
rect 18238 -28312 18302 -28308
rect 18238 -28572 18302 -28568
rect 18238 -28628 18242 -28572
rect 18242 -28628 18298 -28572
rect 18298 -28628 18302 -28572
rect 18238 -28632 18302 -28628
rect 18238 -28892 18302 -28888
rect 18238 -28948 18242 -28892
rect 18242 -28948 18298 -28892
rect 18298 -28948 18302 -28892
rect 18238 -28952 18302 -28948
rect 18238 -29212 18302 -29208
rect 18238 -29268 18242 -29212
rect 18242 -29268 18298 -29212
rect 18298 -29268 18302 -29212
rect 18238 -29272 18302 -29268
rect 18238 -29532 18302 -29528
rect 18238 -29588 18242 -29532
rect 18242 -29588 18298 -29532
rect 18298 -29588 18302 -29532
rect 18238 -29592 18302 -29588
rect 18238 -29852 18302 -29848
rect 18238 -29908 18242 -29852
rect 18242 -29908 18298 -29852
rect 18298 -29908 18302 -29852
rect 18238 -29912 18302 -29908
rect 18238 -30172 18302 -30168
rect 18238 -30228 18242 -30172
rect 18242 -30228 18298 -30172
rect 18298 -30228 18302 -30172
rect 18238 -30232 18302 -30228
rect 25704 -23772 25768 -23768
rect 25704 -23828 25708 -23772
rect 25708 -23828 25764 -23772
rect 25764 -23828 25768 -23772
rect 25704 -23832 25768 -23828
rect 25704 -24092 25768 -24088
rect 25704 -24148 25708 -24092
rect 25708 -24148 25764 -24092
rect 25764 -24148 25768 -24092
rect 25704 -24152 25768 -24148
rect 25704 -24412 25768 -24408
rect 25704 -24468 25708 -24412
rect 25708 -24468 25764 -24412
rect 25764 -24468 25768 -24412
rect 25704 -24472 25768 -24468
rect 25704 -24732 25768 -24728
rect 25704 -24788 25708 -24732
rect 25708 -24788 25764 -24732
rect 25764 -24788 25768 -24732
rect 25704 -24792 25768 -24788
rect 25704 -25052 25768 -25048
rect 25704 -25108 25708 -25052
rect 25708 -25108 25764 -25052
rect 25764 -25108 25768 -25052
rect 25704 -25112 25768 -25108
rect 25704 -25372 25768 -25368
rect 25704 -25428 25708 -25372
rect 25708 -25428 25764 -25372
rect 25764 -25428 25768 -25372
rect 25704 -25432 25768 -25428
rect 25704 -25692 25768 -25688
rect 25704 -25748 25708 -25692
rect 25708 -25748 25764 -25692
rect 25764 -25748 25768 -25692
rect 25704 -25752 25768 -25748
rect 30608 -23246 30672 -23242
rect 30608 -23302 30612 -23246
rect 30612 -23302 30668 -23246
rect 30668 -23302 30672 -23246
rect 30608 -23306 30672 -23302
rect 30928 -23246 30992 -23242
rect 30928 -23302 30932 -23246
rect 30932 -23302 30988 -23246
rect 30988 -23302 30992 -23246
rect 30928 -23306 30992 -23302
rect 31248 -23246 31312 -23242
rect 31248 -23302 31252 -23246
rect 31252 -23302 31308 -23246
rect 31308 -23302 31312 -23246
rect 31248 -23306 31312 -23302
rect 31568 -23246 31632 -23242
rect 31568 -23302 31572 -23246
rect 31572 -23302 31628 -23246
rect 31628 -23302 31632 -23246
rect 31568 -23306 31632 -23302
rect 31888 -23246 31952 -23242
rect 31888 -23302 31892 -23246
rect 31892 -23302 31948 -23246
rect 31948 -23302 31952 -23246
rect 31888 -23306 31952 -23302
rect 32208 -23246 32272 -23242
rect 32208 -23302 32212 -23246
rect 32212 -23302 32268 -23246
rect 32268 -23302 32272 -23246
rect 32208 -23306 32272 -23302
rect 32528 -23246 32592 -23242
rect 32528 -23302 32532 -23246
rect 32532 -23302 32588 -23246
rect 32588 -23302 32592 -23246
rect 32528 -23306 32592 -23302
rect 32848 -23246 32912 -23242
rect 32848 -23302 32852 -23246
rect 32852 -23302 32908 -23246
rect 32908 -23302 32912 -23246
rect 32848 -23306 32912 -23302
rect 33168 -23246 33232 -23242
rect 33168 -23302 33172 -23246
rect 33172 -23302 33228 -23246
rect 33228 -23302 33232 -23246
rect 33168 -23306 33232 -23302
rect 33488 -23246 33552 -23242
rect 33488 -23302 33492 -23246
rect 33492 -23302 33548 -23246
rect 33548 -23302 33552 -23246
rect 33488 -23306 33552 -23302
rect 33808 -23246 33872 -23242
rect 33808 -23302 33812 -23246
rect 33812 -23302 33868 -23246
rect 33868 -23302 33872 -23246
rect 33808 -23306 33872 -23302
rect 34128 -23246 34192 -23242
rect 34128 -23302 34132 -23246
rect 34132 -23302 34188 -23246
rect 34188 -23302 34192 -23246
rect 34128 -23306 34192 -23302
rect 34448 -23246 34512 -23242
rect 34448 -23302 34452 -23246
rect 34452 -23302 34508 -23246
rect 34508 -23302 34512 -23246
rect 34448 -23306 34512 -23302
rect 34768 -23246 34832 -23242
rect 34768 -23302 34772 -23246
rect 34772 -23302 34828 -23246
rect 34828 -23302 34832 -23246
rect 34768 -23306 34832 -23302
rect 35088 -23246 35152 -23242
rect 35088 -23302 35092 -23246
rect 35092 -23302 35148 -23246
rect 35148 -23302 35152 -23246
rect 35088 -23306 35152 -23302
rect 35408 -23246 35472 -23242
rect 35408 -23302 35412 -23246
rect 35412 -23302 35468 -23246
rect 35468 -23302 35472 -23246
rect 35408 -23306 35472 -23302
rect 35728 -23246 35792 -23242
rect 35728 -23302 35732 -23246
rect 35732 -23302 35788 -23246
rect 35788 -23302 35792 -23246
rect 35728 -23306 35792 -23302
rect 36048 -23246 36112 -23242
rect 36048 -23302 36052 -23246
rect 36052 -23302 36108 -23246
rect 36108 -23302 36112 -23246
rect 36048 -23306 36112 -23302
rect 36368 -23246 36432 -23242
rect 36368 -23302 36372 -23246
rect 36372 -23302 36428 -23246
rect 36428 -23302 36432 -23246
rect 36368 -23306 36432 -23302
rect 36688 -23246 36752 -23242
rect 36688 -23302 36692 -23246
rect 36692 -23302 36748 -23246
rect 36748 -23302 36752 -23246
rect 36688 -23306 36752 -23302
rect 37008 -23246 37072 -23242
rect 37008 -23302 37012 -23246
rect 37012 -23302 37068 -23246
rect 37068 -23302 37072 -23246
rect 37008 -23306 37072 -23302
rect 37328 -23246 37392 -23242
rect 37328 -23302 37332 -23246
rect 37332 -23302 37388 -23246
rect 37388 -23302 37392 -23246
rect 37328 -23306 37392 -23302
rect 30238 -23452 30302 -23448
rect 30238 -23508 30242 -23452
rect 30242 -23508 30298 -23452
rect 30298 -23508 30302 -23452
rect 30238 -23512 30302 -23508
rect 37704 -23452 37768 -23448
rect 37704 -23508 37708 -23452
rect 37708 -23508 37764 -23452
rect 37764 -23508 37768 -23452
rect 37704 -23512 37768 -23508
rect 30238 -23772 30302 -23768
rect 30238 -23828 30242 -23772
rect 30242 -23828 30298 -23772
rect 30298 -23828 30302 -23772
rect 30238 -23832 30302 -23828
rect 30238 -24092 30302 -24088
rect 30238 -24148 30242 -24092
rect 30242 -24148 30298 -24092
rect 30298 -24148 30302 -24092
rect 30238 -24152 30302 -24148
rect 30238 -24412 30302 -24408
rect 30238 -24468 30242 -24412
rect 30242 -24468 30298 -24412
rect 30298 -24468 30302 -24412
rect 30238 -24472 30302 -24468
rect 30238 -24732 30302 -24728
rect 30238 -24788 30242 -24732
rect 30242 -24788 30298 -24732
rect 30298 -24788 30302 -24732
rect 30238 -24792 30302 -24788
rect 30238 -25052 30302 -25048
rect 30238 -25108 30242 -25052
rect 30242 -25108 30298 -25052
rect 30298 -25108 30302 -25052
rect 30238 -25112 30302 -25108
rect 30238 -25372 30302 -25368
rect 30238 -25428 30242 -25372
rect 30242 -25428 30298 -25372
rect 30298 -25428 30302 -25372
rect 30238 -25432 30302 -25428
rect 30238 -25692 30302 -25688
rect 30238 -25748 30242 -25692
rect 30242 -25748 30298 -25692
rect 30298 -25748 30302 -25692
rect 30238 -25752 30302 -25748
rect 25704 -26012 25768 -26008
rect 25704 -26068 25708 -26012
rect 25708 -26068 25764 -26012
rect 25764 -26068 25768 -26012
rect 25704 -26072 25768 -26068
rect 25704 -26332 25768 -26328
rect 25704 -26388 25708 -26332
rect 25708 -26388 25764 -26332
rect 25764 -26388 25768 -26332
rect 25704 -26392 25768 -26388
rect 25704 -26652 25768 -26648
rect 25704 -26708 25708 -26652
rect 25708 -26708 25764 -26652
rect 25764 -26708 25768 -26652
rect 25704 -26712 25768 -26708
rect 25704 -26972 25768 -26968
rect 25704 -27028 25708 -26972
rect 25708 -27028 25764 -26972
rect 25764 -27028 25768 -26972
rect 25704 -27032 25768 -27028
rect 25704 -27292 25768 -27288
rect 25704 -27348 25708 -27292
rect 25708 -27348 25764 -27292
rect 25764 -27348 25768 -27292
rect 25704 -27352 25768 -27348
rect 25704 -27612 25768 -27608
rect 25704 -27668 25708 -27612
rect 25708 -27668 25764 -27612
rect 25764 -27668 25768 -27612
rect 25704 -27672 25768 -27668
rect 25704 -27932 25768 -27928
rect 25704 -27988 25708 -27932
rect 25708 -27988 25764 -27932
rect 25764 -27988 25768 -27932
rect 25704 -27992 25768 -27988
rect 25704 -28252 25768 -28248
rect 25704 -28308 25708 -28252
rect 25708 -28308 25764 -28252
rect 25764 -28308 25768 -28252
rect 25704 -28312 25768 -28308
rect 25704 -28572 25768 -28568
rect 25704 -28628 25708 -28572
rect 25708 -28628 25764 -28572
rect 25764 -28628 25768 -28572
rect 25704 -28632 25768 -28628
rect 25704 -28892 25768 -28888
rect 25704 -28948 25708 -28892
rect 25708 -28948 25764 -28892
rect 25764 -28948 25768 -28892
rect 25704 -28952 25768 -28948
rect 25704 -29212 25768 -29208
rect 25704 -29268 25708 -29212
rect 25708 -29268 25764 -29212
rect 25764 -29268 25768 -29212
rect 25704 -29272 25768 -29268
rect 25704 -29532 25768 -29528
rect 25704 -29588 25708 -29532
rect 25708 -29588 25764 -29532
rect 25764 -29588 25768 -29532
rect 25704 -29592 25768 -29588
rect 25704 -29852 25768 -29848
rect 25704 -29908 25708 -29852
rect 25708 -29908 25764 -29852
rect 25764 -29908 25768 -29852
rect 25704 -29912 25768 -29908
rect 25704 -30172 25768 -30168
rect 25704 -30228 25708 -30172
rect 25708 -30228 25764 -30172
rect 25764 -30228 25768 -30172
rect 25704 -30232 25768 -30228
rect 18238 -30492 18302 -30488
rect 18238 -30548 18242 -30492
rect 18242 -30548 18298 -30492
rect 18298 -30548 18302 -30492
rect 18238 -30552 18302 -30548
rect 25704 -30492 25768 -30488
rect 25704 -30548 25708 -30492
rect 25708 -30548 25764 -30492
rect 25764 -30548 25768 -30492
rect 25704 -30552 25768 -30548
rect 18608 -30702 18672 -30698
rect 18608 -30758 18612 -30702
rect 18612 -30758 18668 -30702
rect 18668 -30758 18672 -30702
rect 18608 -30762 18672 -30758
rect 18928 -30702 18992 -30698
rect 18928 -30758 18932 -30702
rect 18932 -30758 18988 -30702
rect 18988 -30758 18992 -30702
rect 18928 -30762 18992 -30758
rect 19248 -30702 19312 -30698
rect 19248 -30758 19252 -30702
rect 19252 -30758 19308 -30702
rect 19308 -30758 19312 -30702
rect 19248 -30762 19312 -30758
rect 19568 -30702 19632 -30698
rect 19568 -30758 19572 -30702
rect 19572 -30758 19628 -30702
rect 19628 -30758 19632 -30702
rect 19568 -30762 19632 -30758
rect 19888 -30702 19952 -30698
rect 19888 -30758 19892 -30702
rect 19892 -30758 19948 -30702
rect 19948 -30758 19952 -30702
rect 19888 -30762 19952 -30758
rect 20208 -30702 20272 -30698
rect 20208 -30758 20212 -30702
rect 20212 -30758 20268 -30702
rect 20268 -30758 20272 -30702
rect 20208 -30762 20272 -30758
rect 20528 -30702 20592 -30698
rect 20528 -30758 20532 -30702
rect 20532 -30758 20588 -30702
rect 20588 -30758 20592 -30702
rect 20528 -30762 20592 -30758
rect 20848 -30702 20912 -30698
rect 20848 -30758 20852 -30702
rect 20852 -30758 20908 -30702
rect 20908 -30758 20912 -30702
rect 20848 -30762 20912 -30758
rect 21168 -30702 21232 -30698
rect 21168 -30758 21172 -30702
rect 21172 -30758 21228 -30702
rect 21228 -30758 21232 -30702
rect 21168 -30762 21232 -30758
rect 21488 -30702 21552 -30698
rect 21488 -30758 21492 -30702
rect 21492 -30758 21548 -30702
rect 21548 -30758 21552 -30702
rect 21488 -30762 21552 -30758
rect 21808 -30702 21872 -30698
rect 21808 -30758 21812 -30702
rect 21812 -30758 21868 -30702
rect 21868 -30758 21872 -30702
rect 21808 -30762 21872 -30758
rect 22128 -30702 22192 -30698
rect 22128 -30758 22132 -30702
rect 22132 -30758 22188 -30702
rect 22188 -30758 22192 -30702
rect 22128 -30762 22192 -30758
rect 22448 -30702 22512 -30698
rect 22448 -30758 22452 -30702
rect 22452 -30758 22508 -30702
rect 22508 -30758 22512 -30702
rect 22448 -30762 22512 -30758
rect 22768 -30702 22832 -30698
rect 22768 -30758 22772 -30702
rect 22772 -30758 22828 -30702
rect 22828 -30758 22832 -30702
rect 22768 -30762 22832 -30758
rect 23088 -30702 23152 -30698
rect 23088 -30758 23092 -30702
rect 23092 -30758 23148 -30702
rect 23148 -30758 23152 -30702
rect 23088 -30762 23152 -30758
rect 23408 -30702 23472 -30698
rect 23408 -30758 23412 -30702
rect 23412 -30758 23468 -30702
rect 23468 -30758 23472 -30702
rect 23408 -30762 23472 -30758
rect 23728 -30702 23792 -30698
rect 23728 -30758 23732 -30702
rect 23732 -30758 23788 -30702
rect 23788 -30758 23792 -30702
rect 23728 -30762 23792 -30758
rect 24048 -30702 24112 -30698
rect 24048 -30758 24052 -30702
rect 24052 -30758 24108 -30702
rect 24108 -30758 24112 -30702
rect 24048 -30762 24112 -30758
rect 24368 -30702 24432 -30698
rect 24368 -30758 24372 -30702
rect 24372 -30758 24428 -30702
rect 24428 -30758 24432 -30702
rect 24368 -30762 24432 -30758
rect 24688 -30702 24752 -30698
rect 24688 -30758 24692 -30702
rect 24692 -30758 24748 -30702
rect 24748 -30758 24752 -30702
rect 24688 -30762 24752 -30758
rect 25008 -30702 25072 -30698
rect 25008 -30758 25012 -30702
rect 25012 -30758 25068 -30702
rect 25068 -30758 25072 -30702
rect 25008 -30762 25072 -30758
rect 25328 -30702 25392 -30698
rect 25328 -30758 25332 -30702
rect 25332 -30758 25388 -30702
rect 25388 -30758 25392 -30702
rect 25328 -30762 25392 -30758
rect 30238 -26012 30302 -26008
rect 30238 -26068 30242 -26012
rect 30242 -26068 30298 -26012
rect 30298 -26068 30302 -26012
rect 30238 -26072 30302 -26068
rect 30238 -26332 30302 -26328
rect 30238 -26388 30242 -26332
rect 30242 -26388 30298 -26332
rect 30298 -26388 30302 -26332
rect 30238 -26392 30302 -26388
rect 30238 -26652 30302 -26648
rect 30238 -26708 30242 -26652
rect 30242 -26708 30298 -26652
rect 30298 -26708 30302 -26652
rect 30238 -26712 30302 -26708
rect 30238 -26972 30302 -26968
rect 30238 -27028 30242 -26972
rect 30242 -27028 30298 -26972
rect 30298 -27028 30302 -26972
rect 30238 -27032 30302 -27028
rect 30238 -27292 30302 -27288
rect 30238 -27348 30242 -27292
rect 30242 -27348 30298 -27292
rect 30298 -27348 30302 -27292
rect 30238 -27352 30302 -27348
rect 30238 -27612 30302 -27608
rect 30238 -27668 30242 -27612
rect 30242 -27668 30298 -27612
rect 30298 -27668 30302 -27612
rect 30238 -27672 30302 -27668
rect 30238 -27932 30302 -27928
rect 30238 -27988 30242 -27932
rect 30242 -27988 30298 -27932
rect 30298 -27988 30302 -27932
rect 30238 -27992 30302 -27988
rect 30238 -28252 30302 -28248
rect 30238 -28308 30242 -28252
rect 30242 -28308 30298 -28252
rect 30298 -28308 30302 -28252
rect 30238 -28312 30302 -28308
rect 30238 -28572 30302 -28568
rect 30238 -28628 30242 -28572
rect 30242 -28628 30298 -28572
rect 30298 -28628 30302 -28572
rect 30238 -28632 30302 -28628
rect 30238 -28892 30302 -28888
rect 30238 -28948 30242 -28892
rect 30242 -28948 30298 -28892
rect 30298 -28948 30302 -28892
rect 30238 -28952 30302 -28948
rect 30238 -29212 30302 -29208
rect 30238 -29268 30242 -29212
rect 30242 -29268 30298 -29212
rect 30298 -29268 30302 -29212
rect 30238 -29272 30302 -29268
rect 30238 -29532 30302 -29528
rect 30238 -29588 30242 -29532
rect 30242 -29588 30298 -29532
rect 30298 -29588 30302 -29532
rect 30238 -29592 30302 -29588
rect 30238 -29852 30302 -29848
rect 30238 -29908 30242 -29852
rect 30242 -29908 30298 -29852
rect 30298 -29908 30302 -29852
rect 30238 -29912 30302 -29908
rect 30238 -30172 30302 -30168
rect 30238 -30228 30242 -30172
rect 30242 -30228 30298 -30172
rect 30298 -30228 30302 -30172
rect 30238 -30232 30302 -30228
rect 37704 -23772 37768 -23768
rect 37704 -23828 37708 -23772
rect 37708 -23828 37764 -23772
rect 37764 -23828 37768 -23772
rect 37704 -23832 37768 -23828
rect 37704 -24092 37768 -24088
rect 37704 -24148 37708 -24092
rect 37708 -24148 37764 -24092
rect 37764 -24148 37768 -24092
rect 37704 -24152 37768 -24148
rect 37704 -24412 37768 -24408
rect 37704 -24468 37708 -24412
rect 37708 -24468 37764 -24412
rect 37764 -24468 37768 -24412
rect 37704 -24472 37768 -24468
rect 37704 -24732 37768 -24728
rect 37704 -24788 37708 -24732
rect 37708 -24788 37764 -24732
rect 37764 -24788 37768 -24732
rect 37704 -24792 37768 -24788
rect 37704 -25052 37768 -25048
rect 37704 -25108 37708 -25052
rect 37708 -25108 37764 -25052
rect 37764 -25108 37768 -25052
rect 37704 -25112 37768 -25108
rect 37704 -25372 37768 -25368
rect 37704 -25428 37708 -25372
rect 37708 -25428 37764 -25372
rect 37764 -25428 37768 -25372
rect 37704 -25432 37768 -25428
rect 37704 -25692 37768 -25688
rect 37704 -25748 37708 -25692
rect 37708 -25748 37764 -25692
rect 37764 -25748 37768 -25692
rect 37704 -25752 37768 -25748
rect 37704 -26012 37768 -26008
rect 37704 -26068 37708 -26012
rect 37708 -26068 37764 -26012
rect 37764 -26068 37768 -26012
rect 37704 -26072 37768 -26068
rect 37704 -26332 37768 -26328
rect 37704 -26388 37708 -26332
rect 37708 -26388 37764 -26332
rect 37764 -26388 37768 -26332
rect 37704 -26392 37768 -26388
rect 37704 -26652 37768 -26648
rect 37704 -26708 37708 -26652
rect 37708 -26708 37764 -26652
rect 37764 -26708 37768 -26652
rect 37704 -26712 37768 -26708
rect 37704 -26972 37768 -26968
rect 37704 -27028 37708 -26972
rect 37708 -27028 37764 -26972
rect 37764 -27028 37768 -26972
rect 37704 -27032 37768 -27028
rect 37704 -27292 37768 -27288
rect 37704 -27348 37708 -27292
rect 37708 -27348 37764 -27292
rect 37764 -27348 37768 -27292
rect 37704 -27352 37768 -27348
rect 37704 -27612 37768 -27608
rect 37704 -27668 37708 -27612
rect 37708 -27668 37764 -27612
rect 37764 -27668 37768 -27612
rect 37704 -27672 37768 -27668
rect 37704 -27932 37768 -27928
rect 37704 -27988 37708 -27932
rect 37708 -27988 37764 -27932
rect 37764 -27988 37768 -27932
rect 37704 -27992 37768 -27988
rect 37704 -28252 37768 -28248
rect 37704 -28308 37708 -28252
rect 37708 -28308 37764 -28252
rect 37764 -28308 37768 -28252
rect 37704 -28312 37768 -28308
rect 37704 -28572 37768 -28568
rect 37704 -28628 37708 -28572
rect 37708 -28628 37764 -28572
rect 37764 -28628 37768 -28572
rect 37704 -28632 37768 -28628
rect 37704 -28892 37768 -28888
rect 37704 -28948 37708 -28892
rect 37708 -28948 37764 -28892
rect 37764 -28948 37768 -28892
rect 37704 -28952 37768 -28948
rect 37704 -29212 37768 -29208
rect 37704 -29268 37708 -29212
rect 37708 -29268 37764 -29212
rect 37764 -29268 37768 -29212
rect 37704 -29272 37768 -29268
rect 37704 -29532 37768 -29528
rect 37704 -29588 37708 -29532
rect 37708 -29588 37764 -29532
rect 37764 -29588 37768 -29532
rect 37704 -29592 37768 -29588
rect 37704 -29852 37768 -29848
rect 37704 -29908 37708 -29852
rect 37708 -29908 37764 -29852
rect 37764 -29908 37768 -29852
rect 37704 -29912 37768 -29908
rect 37704 -30172 37768 -30168
rect 37704 -30228 37708 -30172
rect 37708 -30228 37764 -30172
rect 37764 -30228 37768 -30172
rect 37704 -30232 37768 -30228
rect 30238 -30492 30302 -30488
rect 30238 -30548 30242 -30492
rect 30242 -30548 30298 -30492
rect 30298 -30548 30302 -30492
rect 30238 -30552 30302 -30548
rect 37704 -30492 37768 -30488
rect 37704 -30548 37708 -30492
rect 37708 -30548 37764 -30492
rect 37764 -30548 37768 -30492
rect 37704 -30552 37768 -30548
rect 30608 -30702 30672 -30698
rect 30608 -30758 30612 -30702
rect 30612 -30758 30668 -30702
rect 30668 -30758 30672 -30702
rect 30608 -30762 30672 -30758
rect 30928 -30702 30992 -30698
rect 30928 -30758 30932 -30702
rect 30932 -30758 30988 -30702
rect 30988 -30758 30992 -30702
rect 30928 -30762 30992 -30758
rect 31248 -30702 31312 -30698
rect 31248 -30758 31252 -30702
rect 31252 -30758 31308 -30702
rect 31308 -30758 31312 -30702
rect 31248 -30762 31312 -30758
rect 31568 -30702 31632 -30698
rect 31568 -30758 31572 -30702
rect 31572 -30758 31628 -30702
rect 31628 -30758 31632 -30702
rect 31568 -30762 31632 -30758
rect 31888 -30702 31952 -30698
rect 31888 -30758 31892 -30702
rect 31892 -30758 31948 -30702
rect 31948 -30758 31952 -30702
rect 31888 -30762 31952 -30758
rect 32208 -30702 32272 -30698
rect 32208 -30758 32212 -30702
rect 32212 -30758 32268 -30702
rect 32268 -30758 32272 -30702
rect 32208 -30762 32272 -30758
rect 32528 -30702 32592 -30698
rect 32528 -30758 32532 -30702
rect 32532 -30758 32588 -30702
rect 32588 -30758 32592 -30702
rect 32528 -30762 32592 -30758
rect 32848 -30702 32912 -30698
rect 32848 -30758 32852 -30702
rect 32852 -30758 32908 -30702
rect 32908 -30758 32912 -30702
rect 32848 -30762 32912 -30758
rect 33168 -30702 33232 -30698
rect 33168 -30758 33172 -30702
rect 33172 -30758 33228 -30702
rect 33228 -30758 33232 -30702
rect 33168 -30762 33232 -30758
rect 33488 -30702 33552 -30698
rect 33488 -30758 33492 -30702
rect 33492 -30758 33548 -30702
rect 33548 -30758 33552 -30702
rect 33488 -30762 33552 -30758
rect 33808 -30702 33872 -30698
rect 33808 -30758 33812 -30702
rect 33812 -30758 33868 -30702
rect 33868 -30758 33872 -30702
rect 33808 -30762 33872 -30758
rect 34128 -30702 34192 -30698
rect 34128 -30758 34132 -30702
rect 34132 -30758 34188 -30702
rect 34188 -30758 34192 -30702
rect 34128 -30762 34192 -30758
rect 34448 -30702 34512 -30698
rect 34448 -30758 34452 -30702
rect 34452 -30758 34508 -30702
rect 34508 -30758 34512 -30702
rect 34448 -30762 34512 -30758
rect 34768 -30702 34832 -30698
rect 34768 -30758 34772 -30702
rect 34772 -30758 34828 -30702
rect 34828 -30758 34832 -30702
rect 34768 -30762 34832 -30758
rect 35088 -30702 35152 -30698
rect 35088 -30758 35092 -30702
rect 35092 -30758 35148 -30702
rect 35148 -30758 35152 -30702
rect 35088 -30762 35152 -30758
rect 35408 -30702 35472 -30698
rect 35408 -30758 35412 -30702
rect 35412 -30758 35468 -30702
rect 35468 -30758 35472 -30702
rect 35408 -30762 35472 -30758
rect 35728 -30702 35792 -30698
rect 35728 -30758 35732 -30702
rect 35732 -30758 35788 -30702
rect 35788 -30758 35792 -30702
rect 35728 -30762 35792 -30758
rect 36048 -30702 36112 -30698
rect 36048 -30758 36052 -30702
rect 36052 -30758 36108 -30702
rect 36108 -30758 36112 -30702
rect 36048 -30762 36112 -30758
rect 36368 -30702 36432 -30698
rect 36368 -30758 36372 -30702
rect 36372 -30758 36428 -30702
rect 36428 -30758 36432 -30702
rect 36368 -30762 36432 -30758
rect 36688 -30702 36752 -30698
rect 36688 -30758 36692 -30702
rect 36692 -30758 36748 -30702
rect 36748 -30758 36752 -30702
rect 36688 -30762 36752 -30758
rect 37008 -30702 37072 -30698
rect 37008 -30758 37012 -30702
rect 37012 -30758 37068 -30702
rect 37068 -30758 37072 -30702
rect 37008 -30762 37072 -30758
rect 37328 -30702 37392 -30698
rect 37328 -30758 37332 -30702
rect 37332 -30758 37388 -30702
rect 37388 -30758 37392 -30702
rect 37328 -30762 37392 -30758
rect 42608 -23246 42672 -23242
rect 42608 -23302 42612 -23246
rect 42612 -23302 42668 -23246
rect 42668 -23302 42672 -23246
rect 42608 -23306 42672 -23302
rect 42928 -23246 42992 -23242
rect 42928 -23302 42932 -23246
rect 42932 -23302 42988 -23246
rect 42988 -23302 42992 -23246
rect 42928 -23306 42992 -23302
rect 43248 -23246 43312 -23242
rect 43248 -23302 43252 -23246
rect 43252 -23302 43308 -23246
rect 43308 -23302 43312 -23246
rect 43248 -23306 43312 -23302
rect 43568 -23246 43632 -23242
rect 43568 -23302 43572 -23246
rect 43572 -23302 43628 -23246
rect 43628 -23302 43632 -23246
rect 43568 -23306 43632 -23302
rect 43888 -23246 43952 -23242
rect 43888 -23302 43892 -23246
rect 43892 -23302 43948 -23246
rect 43948 -23302 43952 -23246
rect 43888 -23306 43952 -23302
rect 44208 -23246 44272 -23242
rect 44208 -23302 44212 -23246
rect 44212 -23302 44268 -23246
rect 44268 -23302 44272 -23246
rect 44208 -23306 44272 -23302
rect 44528 -23246 44592 -23242
rect 44528 -23302 44532 -23246
rect 44532 -23302 44588 -23246
rect 44588 -23302 44592 -23246
rect 44528 -23306 44592 -23302
rect 44848 -23246 44912 -23242
rect 44848 -23302 44852 -23246
rect 44852 -23302 44908 -23246
rect 44908 -23302 44912 -23246
rect 44848 -23306 44912 -23302
rect 45168 -23246 45232 -23242
rect 45168 -23302 45172 -23246
rect 45172 -23302 45228 -23246
rect 45228 -23302 45232 -23246
rect 45168 -23306 45232 -23302
rect 45488 -23246 45552 -23242
rect 45488 -23302 45492 -23246
rect 45492 -23302 45548 -23246
rect 45548 -23302 45552 -23246
rect 45488 -23306 45552 -23302
rect 45808 -23246 45872 -23242
rect 45808 -23302 45812 -23246
rect 45812 -23302 45868 -23246
rect 45868 -23302 45872 -23246
rect 45808 -23306 45872 -23302
rect 46128 -23246 46192 -23242
rect 46128 -23302 46132 -23246
rect 46132 -23302 46188 -23246
rect 46188 -23302 46192 -23246
rect 46128 -23306 46192 -23302
rect 46448 -23246 46512 -23242
rect 46448 -23302 46452 -23246
rect 46452 -23302 46508 -23246
rect 46508 -23302 46512 -23246
rect 46448 -23306 46512 -23302
rect 46768 -23246 46832 -23242
rect 46768 -23302 46772 -23246
rect 46772 -23302 46828 -23246
rect 46828 -23302 46832 -23246
rect 46768 -23306 46832 -23302
rect 47088 -23246 47152 -23242
rect 47088 -23302 47092 -23246
rect 47092 -23302 47148 -23246
rect 47148 -23302 47152 -23246
rect 47088 -23306 47152 -23302
rect 47408 -23246 47472 -23242
rect 47408 -23302 47412 -23246
rect 47412 -23302 47468 -23246
rect 47468 -23302 47472 -23246
rect 47408 -23306 47472 -23302
rect 47728 -23246 47792 -23242
rect 47728 -23302 47732 -23246
rect 47732 -23302 47788 -23246
rect 47788 -23302 47792 -23246
rect 47728 -23306 47792 -23302
rect 48048 -23246 48112 -23242
rect 48048 -23302 48052 -23246
rect 48052 -23302 48108 -23246
rect 48108 -23302 48112 -23246
rect 48048 -23306 48112 -23302
rect 48368 -23246 48432 -23242
rect 48368 -23302 48372 -23246
rect 48372 -23302 48428 -23246
rect 48428 -23302 48432 -23246
rect 48368 -23306 48432 -23302
rect 48688 -23246 48752 -23242
rect 48688 -23302 48692 -23246
rect 48692 -23302 48748 -23246
rect 48748 -23302 48752 -23246
rect 48688 -23306 48752 -23302
rect 49008 -23246 49072 -23242
rect 49008 -23302 49012 -23246
rect 49012 -23302 49068 -23246
rect 49068 -23302 49072 -23246
rect 49008 -23306 49072 -23302
rect 49328 -23246 49392 -23242
rect 49328 -23302 49332 -23246
rect 49332 -23302 49388 -23246
rect 49388 -23302 49392 -23246
rect 49328 -23306 49392 -23302
rect 42238 -23452 42302 -23448
rect 42238 -23508 42242 -23452
rect 42242 -23508 42298 -23452
rect 42298 -23508 42302 -23452
rect 42238 -23512 42302 -23508
rect 49704 -23452 49768 -23448
rect 49704 -23508 49708 -23452
rect 49708 -23508 49764 -23452
rect 49764 -23508 49768 -23452
rect 49704 -23512 49768 -23508
rect 42238 -23772 42302 -23768
rect 42238 -23828 42242 -23772
rect 42242 -23828 42298 -23772
rect 42298 -23828 42302 -23772
rect 42238 -23832 42302 -23828
rect 42238 -24092 42302 -24088
rect 42238 -24148 42242 -24092
rect 42242 -24148 42298 -24092
rect 42298 -24148 42302 -24092
rect 42238 -24152 42302 -24148
rect 42238 -24412 42302 -24408
rect 42238 -24468 42242 -24412
rect 42242 -24468 42298 -24412
rect 42298 -24468 42302 -24412
rect 42238 -24472 42302 -24468
rect 42238 -24732 42302 -24728
rect 42238 -24788 42242 -24732
rect 42242 -24788 42298 -24732
rect 42298 -24788 42302 -24732
rect 42238 -24792 42302 -24788
rect 42238 -25052 42302 -25048
rect 42238 -25108 42242 -25052
rect 42242 -25108 42298 -25052
rect 42298 -25108 42302 -25052
rect 42238 -25112 42302 -25108
rect 42238 -25372 42302 -25368
rect 42238 -25428 42242 -25372
rect 42242 -25428 42298 -25372
rect 42298 -25428 42302 -25372
rect 42238 -25432 42302 -25428
rect 42238 -25692 42302 -25688
rect 42238 -25748 42242 -25692
rect 42242 -25748 42298 -25692
rect 42298 -25748 42302 -25692
rect 42238 -25752 42302 -25748
rect 42238 -26012 42302 -26008
rect 42238 -26068 42242 -26012
rect 42242 -26068 42298 -26012
rect 42298 -26068 42302 -26012
rect 42238 -26072 42302 -26068
rect 42238 -26332 42302 -26328
rect 42238 -26388 42242 -26332
rect 42242 -26388 42298 -26332
rect 42298 -26388 42302 -26332
rect 42238 -26392 42302 -26388
rect 42238 -26652 42302 -26648
rect 42238 -26708 42242 -26652
rect 42242 -26708 42298 -26652
rect 42298 -26708 42302 -26652
rect 42238 -26712 42302 -26708
rect 42238 -26972 42302 -26968
rect 42238 -27028 42242 -26972
rect 42242 -27028 42298 -26972
rect 42298 -27028 42302 -26972
rect 42238 -27032 42302 -27028
rect 42238 -27292 42302 -27288
rect 42238 -27348 42242 -27292
rect 42242 -27348 42298 -27292
rect 42298 -27348 42302 -27292
rect 42238 -27352 42302 -27348
rect 42238 -27612 42302 -27608
rect 42238 -27668 42242 -27612
rect 42242 -27668 42298 -27612
rect 42298 -27668 42302 -27612
rect 42238 -27672 42302 -27668
rect 42238 -27932 42302 -27928
rect 42238 -27988 42242 -27932
rect 42242 -27988 42298 -27932
rect 42298 -27988 42302 -27932
rect 42238 -27992 42302 -27988
rect 42238 -28252 42302 -28248
rect 42238 -28308 42242 -28252
rect 42242 -28308 42298 -28252
rect 42298 -28308 42302 -28252
rect 42238 -28312 42302 -28308
rect 42238 -28572 42302 -28568
rect 42238 -28628 42242 -28572
rect 42242 -28628 42298 -28572
rect 42298 -28628 42302 -28572
rect 42238 -28632 42302 -28628
rect 42238 -28892 42302 -28888
rect 42238 -28948 42242 -28892
rect 42242 -28948 42298 -28892
rect 42298 -28948 42302 -28892
rect 42238 -28952 42302 -28948
rect 42238 -29212 42302 -29208
rect 42238 -29268 42242 -29212
rect 42242 -29268 42298 -29212
rect 42298 -29268 42302 -29212
rect 42238 -29272 42302 -29268
rect 42238 -29532 42302 -29528
rect 42238 -29588 42242 -29532
rect 42242 -29588 42298 -29532
rect 42298 -29588 42302 -29532
rect 42238 -29592 42302 -29588
rect 42238 -29852 42302 -29848
rect 42238 -29908 42242 -29852
rect 42242 -29908 42298 -29852
rect 42298 -29908 42302 -29852
rect 42238 -29912 42302 -29908
rect 42238 -30172 42302 -30168
rect 42238 -30228 42242 -30172
rect 42242 -30228 42298 -30172
rect 42298 -30228 42302 -30172
rect 42238 -30232 42302 -30228
rect 49704 -23772 49768 -23768
rect 49704 -23828 49708 -23772
rect 49708 -23828 49764 -23772
rect 49764 -23828 49768 -23772
rect 49704 -23832 49768 -23828
rect 49704 -24092 49768 -24088
rect 49704 -24148 49708 -24092
rect 49708 -24148 49764 -24092
rect 49764 -24148 49768 -24092
rect 49704 -24152 49768 -24148
rect 49704 -24412 49768 -24408
rect 49704 -24468 49708 -24412
rect 49708 -24468 49764 -24412
rect 49764 -24468 49768 -24412
rect 49704 -24472 49768 -24468
rect 49704 -24732 49768 -24728
rect 49704 -24788 49708 -24732
rect 49708 -24788 49764 -24732
rect 49764 -24788 49768 -24732
rect 49704 -24792 49768 -24788
rect 49704 -25052 49768 -25048
rect 49704 -25108 49708 -25052
rect 49708 -25108 49764 -25052
rect 49764 -25108 49768 -25052
rect 49704 -25112 49768 -25108
rect 49704 -25372 49768 -25368
rect 49704 -25428 49708 -25372
rect 49708 -25428 49764 -25372
rect 49764 -25428 49768 -25372
rect 49704 -25432 49768 -25428
rect 49704 -25692 49768 -25688
rect 49704 -25748 49708 -25692
rect 49708 -25748 49764 -25692
rect 49764 -25748 49768 -25692
rect 49704 -25752 49768 -25748
rect 49704 -26012 49768 -26008
rect 49704 -26068 49708 -26012
rect 49708 -26068 49764 -26012
rect 49764 -26068 49768 -26012
rect 49704 -26072 49768 -26068
rect 49704 -26332 49768 -26328
rect 49704 -26388 49708 -26332
rect 49708 -26388 49764 -26332
rect 49764 -26388 49768 -26332
rect 49704 -26392 49768 -26388
rect 49704 -26652 49768 -26648
rect 49704 -26708 49708 -26652
rect 49708 -26708 49764 -26652
rect 49764 -26708 49768 -26652
rect 49704 -26712 49768 -26708
rect 49704 -26972 49768 -26968
rect 49704 -27028 49708 -26972
rect 49708 -27028 49764 -26972
rect 49764 -27028 49768 -26972
rect 49704 -27032 49768 -27028
rect 49704 -27292 49768 -27288
rect 49704 -27348 49708 -27292
rect 49708 -27348 49764 -27292
rect 49764 -27348 49768 -27292
rect 49704 -27352 49768 -27348
rect 49704 -27612 49768 -27608
rect 49704 -27668 49708 -27612
rect 49708 -27668 49764 -27612
rect 49764 -27668 49768 -27612
rect 49704 -27672 49768 -27668
rect 49704 -27932 49768 -27928
rect 49704 -27988 49708 -27932
rect 49708 -27988 49764 -27932
rect 49764 -27988 49768 -27932
rect 49704 -27992 49768 -27988
rect 49704 -28252 49768 -28248
rect 49704 -28308 49708 -28252
rect 49708 -28308 49764 -28252
rect 49764 -28308 49768 -28252
rect 49704 -28312 49768 -28308
rect 49704 -28572 49768 -28568
rect 49704 -28628 49708 -28572
rect 49708 -28628 49764 -28572
rect 49764 -28628 49768 -28572
rect 49704 -28632 49768 -28628
rect 49704 -28892 49768 -28888
rect 49704 -28948 49708 -28892
rect 49708 -28948 49764 -28892
rect 49764 -28948 49768 -28892
rect 49704 -28952 49768 -28948
rect 49704 -29212 49768 -29208
rect 49704 -29268 49708 -29212
rect 49708 -29268 49764 -29212
rect 49764 -29268 49768 -29212
rect 49704 -29272 49768 -29268
rect 49704 -29532 49768 -29528
rect 49704 -29588 49708 -29532
rect 49708 -29588 49764 -29532
rect 49764 -29588 49768 -29532
rect 49704 -29592 49768 -29588
rect 49704 -29852 49768 -29848
rect 49704 -29908 49708 -29852
rect 49708 -29908 49764 -29852
rect 49764 -29908 49768 -29852
rect 49704 -29912 49768 -29908
rect 49704 -30172 49768 -30168
rect 49704 -30228 49708 -30172
rect 49708 -30228 49764 -30172
rect 49764 -30228 49768 -30172
rect 49704 -30232 49768 -30228
rect 42238 -30492 42302 -30488
rect 42238 -30548 42242 -30492
rect 42242 -30548 42298 -30492
rect 42298 -30548 42302 -30492
rect 42238 -30552 42302 -30548
rect 49704 -30492 49768 -30488
rect 49704 -30548 49708 -30492
rect 49708 -30548 49764 -30492
rect 49764 -30548 49768 -30492
rect 49704 -30552 49768 -30548
rect 42608 -30702 42672 -30698
rect 42608 -30758 42612 -30702
rect 42612 -30758 42668 -30702
rect 42668 -30758 42672 -30702
rect 42608 -30762 42672 -30758
rect 42928 -30702 42992 -30698
rect 42928 -30758 42932 -30702
rect 42932 -30758 42988 -30702
rect 42988 -30758 42992 -30702
rect 42928 -30762 42992 -30758
rect 43248 -30702 43312 -30698
rect 43248 -30758 43252 -30702
rect 43252 -30758 43308 -30702
rect 43308 -30758 43312 -30702
rect 43248 -30762 43312 -30758
rect 43568 -30702 43632 -30698
rect 43568 -30758 43572 -30702
rect 43572 -30758 43628 -30702
rect 43628 -30758 43632 -30702
rect 43568 -30762 43632 -30758
rect 43888 -30702 43952 -30698
rect 43888 -30758 43892 -30702
rect 43892 -30758 43948 -30702
rect 43948 -30758 43952 -30702
rect 43888 -30762 43952 -30758
rect 44208 -30702 44272 -30698
rect 44208 -30758 44212 -30702
rect 44212 -30758 44268 -30702
rect 44268 -30758 44272 -30702
rect 44208 -30762 44272 -30758
rect 44528 -30702 44592 -30698
rect 44528 -30758 44532 -30702
rect 44532 -30758 44588 -30702
rect 44588 -30758 44592 -30702
rect 44528 -30762 44592 -30758
rect 44848 -30702 44912 -30698
rect 44848 -30758 44852 -30702
rect 44852 -30758 44908 -30702
rect 44908 -30758 44912 -30702
rect 44848 -30762 44912 -30758
rect 45168 -30702 45232 -30698
rect 45168 -30758 45172 -30702
rect 45172 -30758 45228 -30702
rect 45228 -30758 45232 -30702
rect 45168 -30762 45232 -30758
rect 45488 -30702 45552 -30698
rect 45488 -30758 45492 -30702
rect 45492 -30758 45548 -30702
rect 45548 -30758 45552 -30702
rect 45488 -30762 45552 -30758
rect 45808 -30702 45872 -30698
rect 45808 -30758 45812 -30702
rect 45812 -30758 45868 -30702
rect 45868 -30758 45872 -30702
rect 45808 -30762 45872 -30758
rect 46128 -30702 46192 -30698
rect 46128 -30758 46132 -30702
rect 46132 -30758 46188 -30702
rect 46188 -30758 46192 -30702
rect 46128 -30762 46192 -30758
rect 46448 -30702 46512 -30698
rect 46448 -30758 46452 -30702
rect 46452 -30758 46508 -30702
rect 46508 -30758 46512 -30702
rect 46448 -30762 46512 -30758
rect 46768 -30702 46832 -30698
rect 46768 -30758 46772 -30702
rect 46772 -30758 46828 -30702
rect 46828 -30758 46832 -30702
rect 46768 -30762 46832 -30758
rect 47088 -30702 47152 -30698
rect 47088 -30758 47092 -30702
rect 47092 -30758 47148 -30702
rect 47148 -30758 47152 -30702
rect 47088 -30762 47152 -30758
rect 47408 -30702 47472 -30698
rect 47408 -30758 47412 -30702
rect 47412 -30758 47468 -30702
rect 47468 -30758 47472 -30702
rect 47408 -30762 47472 -30758
rect 47728 -30702 47792 -30698
rect 47728 -30758 47732 -30702
rect 47732 -30758 47788 -30702
rect 47788 -30758 47792 -30702
rect 47728 -30762 47792 -30758
rect 48048 -30702 48112 -30698
rect 48048 -30758 48052 -30702
rect 48052 -30758 48108 -30702
rect 48108 -30758 48112 -30702
rect 48048 -30762 48112 -30758
rect 48368 -30702 48432 -30698
rect 48368 -30758 48372 -30702
rect 48372 -30758 48428 -30702
rect 48428 -30758 48432 -30702
rect 48368 -30762 48432 -30758
rect 48688 -30702 48752 -30698
rect 48688 -30758 48692 -30702
rect 48692 -30758 48748 -30702
rect 48748 -30758 48752 -30702
rect 48688 -30762 48752 -30758
rect 49008 -30702 49072 -30698
rect 49008 -30758 49012 -30702
rect 49012 -30758 49068 -30702
rect 49068 -30758 49072 -30702
rect 49008 -30762 49072 -30758
rect 49328 -30702 49392 -30698
rect 49328 -30758 49332 -30702
rect 49332 -30758 49388 -30702
rect 49388 -30758 49392 -30702
rect 49328 -30762 49392 -30758
<< mimcap >>
rect 16500 -2788 17600 -2748
rect 13300 -2840 15900 -2800
rect 13300 -8960 13340 -2840
rect 15860 -8960 15900 -2840
rect 16500 -8108 16540 -2788
rect 17560 -8108 17600 -2788
rect 22232 -2950 22972 -2930
rect 22232 -5550 22252 -2950
rect 22952 -5550 22972 -2950
rect 22232 -5570 22972 -5550
rect 16500 -8148 17600 -8108
rect 13300 -9000 15900 -8960
<< mimcapcontact >>
rect 13340 -8960 15860 -2840
rect 16540 -8108 17560 -2788
rect 22252 -5550 22952 -2950
<< metal4 >>
rect 13400 -2400 21600 -1900
rect 13400 -2700 15800 -2400
rect 18200 -2500 21600 -2400
rect 13200 -2840 16000 -2700
rect 13200 -7900 13340 -2840
rect 11000 -8960 13340 -7900
rect 15860 -8960 16000 -2840
rect 16400 -2788 17700 -2648
rect 16400 -8108 16540 -2788
rect 17560 -8108 17700 -2788
rect 18200 -3000 18300 -2500
rect 21500 -3000 21600 -2500
rect 18200 -3100 21600 -3000
rect 22202 -2950 23002 -2900
rect 22202 -5540 22252 -2950
rect 21872 -5550 22252 -5540
rect 22952 -5540 23002 -2950
rect 23500 -5540 24900 -5500
rect 22952 -5550 24900 -5540
rect 21872 -5560 24900 -5550
rect 21872 -5650 21882 -5560
rect 21992 -5600 24900 -5560
rect 21992 -5650 22002 -5600
rect 21872 -5660 22002 -5650
rect 23500 -5700 24900 -5600
rect 22402 -5720 23002 -5700
rect 22402 -5880 22422 -5720
rect 22402 -5960 22432 -5880
rect 22982 -5880 23002 -5720
rect 22972 -5960 23002 -5880
rect 22402 -5990 23002 -5960
rect 16400 -8248 17700 -8108
rect 17460 -8440 17700 -8248
rect 11000 -9100 16000 -8960
rect 16400 -8748 17300 -8648
rect 11000 -11000 12300 -9100
rect 16400 -9148 16500 -8748
rect 17200 -9148 17300 -8748
rect 16400 -9248 17300 -9148
rect 17460 -9360 17480 -8440
rect 17680 -9360 17700 -8440
rect 17460 -9380 17700 -9360
rect 17460 -9500 17699 -9380
rect 13200 -9600 16000 -9500
rect 13200 -10200 13300 -9600
rect 15900 -9800 16000 -9600
rect 17460 -9600 22200 -9500
rect 17460 -9800 17700 -9600
rect 15900 -10200 17700 -9800
rect 18900 -10200 20900 -9600
rect 22100 -10200 22200 -9600
rect 13200 -10300 22200 -10200
rect 18000 -11000 22200 -10300
rect 24700 -10300 24900 -5700
rect 24700 -10500 27100 -10300
rect 26900 -10700 27100 -10500
rect 26900 -10900 38700 -10700
rect 6000 -11156 14000 -11000
rect 6000 -11362 6522 -11156
rect 6000 -11598 6152 -11362
rect 6388 -11392 6522 -11362
rect 6758 -11392 6842 -11156
rect 7078 -11392 7162 -11156
rect 7398 -11392 7482 -11156
rect 7718 -11392 7802 -11156
rect 8038 -11392 8122 -11156
rect 8358 -11392 8442 -11156
rect 8678 -11392 8762 -11156
rect 8998 -11392 9082 -11156
rect 9318 -11392 9402 -11156
rect 9638 -11392 9722 -11156
rect 9958 -11392 10042 -11156
rect 10278 -11392 10362 -11156
rect 10598 -11392 10682 -11156
rect 10918 -11392 11002 -11156
rect 11238 -11392 11322 -11156
rect 11558 -11392 11642 -11156
rect 11878 -11392 11962 -11156
rect 12198 -11392 12282 -11156
rect 12518 -11392 12602 -11156
rect 12838 -11392 12922 -11156
rect 13158 -11392 13242 -11156
rect 13478 -11362 14000 -11156
rect 13478 -11392 13618 -11362
rect 6388 -11540 13618 -11392
rect 6388 -11598 6540 -11540
rect 6000 -11682 6540 -11598
rect 6000 -11918 6152 -11682
rect 6388 -11918 6540 -11682
rect 6000 -12002 6540 -11918
rect 6000 -12238 6152 -12002
rect 6388 -12238 6540 -12002
rect 6000 -12322 6540 -12238
rect 6000 -12558 6152 -12322
rect 6388 -12558 6540 -12322
rect 6000 -12642 6540 -12558
rect 6000 -12878 6152 -12642
rect 6388 -12878 6540 -12642
rect 6000 -12962 6540 -12878
rect 6000 -13198 6152 -12962
rect 6388 -13198 6540 -12962
rect 6000 -13282 6540 -13198
rect 6000 -13518 6152 -13282
rect 6388 -13518 6540 -13282
rect 6000 -13602 6540 -13518
rect 6000 -13838 6152 -13602
rect 6388 -13838 6540 -13602
rect 6000 -13922 6540 -13838
rect 6000 -14158 6152 -13922
rect 6388 -14158 6540 -13922
rect 6000 -14242 6540 -14158
rect 6000 -14478 6152 -14242
rect 6388 -14478 6540 -14242
rect 6000 -14562 6540 -14478
rect 6000 -14798 6152 -14562
rect 6388 -14798 6540 -14562
rect 6000 -14882 6540 -14798
rect 6000 -15118 6152 -14882
rect 6388 -15118 6540 -14882
rect 6000 -15202 6540 -15118
rect 6000 -15438 6152 -15202
rect 6388 -15438 6540 -15202
rect 6000 -15522 6540 -15438
rect 6000 -15758 6152 -15522
rect 6388 -15758 6540 -15522
rect 6000 -15842 6540 -15758
rect 6000 -16078 6152 -15842
rect 6388 -16078 6540 -15842
rect 6000 -16162 6540 -16078
rect 6000 -16398 6152 -16162
rect 6388 -16398 6540 -16162
rect 6000 -16482 6540 -16398
rect 6000 -16718 6152 -16482
rect 6388 -16718 6540 -16482
rect 6000 -16802 6540 -16718
rect 6000 -17038 6152 -16802
rect 6388 -17038 6540 -16802
rect 6000 -17122 6540 -17038
rect 6000 -17358 6152 -17122
rect 6388 -17358 6540 -17122
rect 6000 -17442 6540 -17358
rect 6000 -17678 6152 -17442
rect 6388 -17678 6540 -17442
rect 6000 -17762 6540 -17678
rect 6000 -17998 6152 -17762
rect 6388 -17998 6540 -17762
rect 6000 -18082 6540 -17998
rect 6000 -18318 6152 -18082
rect 6388 -18318 6540 -18082
rect 6000 -18402 6540 -18318
rect 6000 -18638 6152 -18402
rect 6388 -18460 6540 -18402
rect 13460 -11598 13618 -11540
rect 13854 -11598 14000 -11362
rect 13460 -11682 14000 -11598
rect 13460 -11918 13618 -11682
rect 13854 -11918 14000 -11682
rect 13460 -12002 14000 -11918
rect 13460 -12238 13618 -12002
rect 13854 -12238 14000 -12002
rect 13460 -12322 14000 -12238
rect 13460 -12558 13618 -12322
rect 13854 -12558 14000 -12322
rect 13460 -12642 14000 -12558
rect 13460 -12878 13618 -12642
rect 13854 -12878 14000 -12642
rect 13460 -12962 14000 -12878
rect 13460 -13198 13618 -12962
rect 13854 -13198 14000 -12962
rect 13460 -13282 14000 -13198
rect 13460 -13518 13618 -13282
rect 13854 -13518 14000 -13282
rect 13460 -13602 14000 -13518
rect 13460 -13838 13618 -13602
rect 13854 -13838 14000 -13602
rect 13460 -13922 14000 -13838
rect 13460 -14158 13618 -13922
rect 13854 -14158 14000 -13922
rect 13460 -14242 14000 -14158
rect 13460 -14478 13618 -14242
rect 13854 -14478 14000 -14242
rect 13460 -14562 14000 -14478
rect 13460 -14798 13618 -14562
rect 13854 -14798 14000 -14562
rect 13460 -14882 14000 -14798
rect 13460 -15118 13618 -14882
rect 13854 -15118 14000 -14882
rect 13460 -15202 14000 -15118
rect 13460 -15438 13618 -15202
rect 13854 -15438 14000 -15202
rect 13460 -15522 14000 -15438
rect 13460 -15758 13618 -15522
rect 13854 -15758 14000 -15522
rect 13460 -15842 14000 -15758
rect 13460 -16078 13618 -15842
rect 13854 -16078 14000 -15842
rect 13460 -16162 14000 -16078
rect 13460 -16398 13618 -16162
rect 13854 -16398 14000 -16162
rect 13460 -16482 14000 -16398
rect 13460 -16718 13618 -16482
rect 13854 -16718 14000 -16482
rect 13460 -16802 14000 -16718
rect 13460 -17038 13618 -16802
rect 13854 -17038 14000 -16802
rect 13460 -17122 14000 -17038
rect 13460 -17358 13618 -17122
rect 13854 -17358 14000 -17122
rect 13460 -17442 14000 -17358
rect 13460 -17678 13618 -17442
rect 13854 -17678 14000 -17442
rect 13460 -17762 14000 -17678
rect 13460 -17998 13618 -17762
rect 13854 -17998 14000 -17762
rect 13460 -18082 14000 -17998
rect 13460 -18318 13618 -18082
rect 13854 -18318 14000 -18082
rect 13460 -18402 14000 -18318
rect 13460 -18460 13618 -18402
rect 6388 -18612 13618 -18460
rect 6388 -18638 6522 -18612
rect 6000 -18848 6522 -18638
rect 6758 -18848 6842 -18612
rect 7078 -18848 7162 -18612
rect 7398 -18848 7482 -18612
rect 7718 -18848 7802 -18612
rect 8038 -18848 8122 -18612
rect 8358 -18848 8442 -18612
rect 8678 -18848 8762 -18612
rect 8998 -18848 9082 -18612
rect 9318 -18848 9402 -18612
rect 9638 -18848 9722 -18612
rect 9958 -18848 10042 -18612
rect 10278 -18848 10362 -18612
rect 10598 -18848 10682 -18612
rect 10918 -18848 11002 -18612
rect 11238 -18848 11322 -18612
rect 11558 -18848 11642 -18612
rect 11878 -18848 11962 -18612
rect 12198 -18848 12282 -18612
rect 12518 -18848 12602 -18612
rect 12838 -18848 12922 -18612
rect 13158 -18848 13242 -18612
rect 13478 -18638 13618 -18612
rect 13854 -18638 14000 -18402
rect 13478 -18848 14000 -18638
rect 6000 -19000 14000 -18848
rect 18000 -11156 26000 -11000
rect 18000 -11362 18522 -11156
rect 18000 -11598 18152 -11362
rect 18388 -11392 18522 -11362
rect 18758 -11392 18842 -11156
rect 19078 -11392 19162 -11156
rect 19398 -11392 19482 -11156
rect 19718 -11392 19802 -11156
rect 20038 -11392 20122 -11156
rect 20358 -11392 20442 -11156
rect 20678 -11392 20762 -11156
rect 20998 -11392 21082 -11156
rect 21318 -11392 21402 -11156
rect 21638 -11392 21722 -11156
rect 21958 -11392 22042 -11156
rect 22278 -11392 22362 -11156
rect 22598 -11392 22682 -11156
rect 22918 -11392 23002 -11156
rect 23238 -11392 23322 -11156
rect 23558 -11392 23642 -11156
rect 23878 -11392 23962 -11156
rect 24198 -11392 24282 -11156
rect 24518 -11392 24602 -11156
rect 24838 -11392 24922 -11156
rect 25158 -11392 25242 -11156
rect 25478 -11362 26000 -11156
rect 25478 -11392 25618 -11362
rect 18388 -11540 25618 -11392
rect 18388 -11598 18540 -11540
rect 18000 -11682 18540 -11598
rect 18000 -11918 18152 -11682
rect 18388 -11918 18540 -11682
rect 18000 -12002 18540 -11918
rect 18000 -12238 18152 -12002
rect 18388 -12238 18540 -12002
rect 18000 -12322 18540 -12238
rect 18000 -12558 18152 -12322
rect 18388 -12558 18540 -12322
rect 18000 -12642 18540 -12558
rect 18000 -12878 18152 -12642
rect 18388 -12878 18540 -12642
rect 18000 -12962 18540 -12878
rect 18000 -13198 18152 -12962
rect 18388 -13198 18540 -12962
rect 18000 -13282 18540 -13198
rect 18000 -13518 18152 -13282
rect 18388 -13518 18540 -13282
rect 18000 -13602 18540 -13518
rect 18000 -13838 18152 -13602
rect 18388 -13838 18540 -13602
rect 18000 -13922 18540 -13838
rect 18000 -14158 18152 -13922
rect 18388 -14158 18540 -13922
rect 18000 -14242 18540 -14158
rect 18000 -14478 18152 -14242
rect 18388 -14478 18540 -14242
rect 18000 -14562 18540 -14478
rect 18000 -14798 18152 -14562
rect 18388 -14798 18540 -14562
rect 18000 -14882 18540 -14798
rect 18000 -15118 18152 -14882
rect 18388 -15118 18540 -14882
rect 18000 -15202 18540 -15118
rect 18000 -15438 18152 -15202
rect 18388 -15438 18540 -15202
rect 18000 -15522 18540 -15438
rect 18000 -15758 18152 -15522
rect 18388 -15758 18540 -15522
rect 18000 -15842 18540 -15758
rect 18000 -16078 18152 -15842
rect 18388 -16078 18540 -15842
rect 18000 -16162 18540 -16078
rect 18000 -16398 18152 -16162
rect 18388 -16398 18540 -16162
rect 18000 -16482 18540 -16398
rect 18000 -16718 18152 -16482
rect 18388 -16718 18540 -16482
rect 18000 -16802 18540 -16718
rect 18000 -17038 18152 -16802
rect 18388 -17038 18540 -16802
rect 18000 -17122 18540 -17038
rect 18000 -17358 18152 -17122
rect 18388 -17358 18540 -17122
rect 18000 -17442 18540 -17358
rect 18000 -17678 18152 -17442
rect 18388 -17678 18540 -17442
rect 18000 -17762 18540 -17678
rect 18000 -17998 18152 -17762
rect 18388 -17998 18540 -17762
rect 18000 -18082 18540 -17998
rect 18000 -18318 18152 -18082
rect 18388 -18318 18540 -18082
rect 18000 -18402 18540 -18318
rect 18000 -18638 18152 -18402
rect 18388 -18460 18540 -18402
rect 25460 -11598 25618 -11540
rect 25854 -11598 26000 -11362
rect 25460 -11682 26000 -11598
rect 25460 -11918 25618 -11682
rect 25854 -11918 26000 -11682
rect 25460 -12002 26000 -11918
rect 25460 -12238 25618 -12002
rect 25854 -12238 26000 -12002
rect 25460 -12322 26000 -12238
rect 25460 -12558 25618 -12322
rect 25854 -12558 26000 -12322
rect 25460 -12642 26000 -12558
rect 25460 -12878 25618 -12642
rect 25854 -12878 26000 -12642
rect 25460 -12962 26000 -12878
rect 25460 -13198 25618 -12962
rect 25854 -13198 26000 -12962
rect 25460 -13282 26000 -13198
rect 25460 -13518 25618 -13282
rect 25854 -13518 26000 -13282
rect 25460 -13602 26000 -13518
rect 25460 -13838 25618 -13602
rect 25854 -13838 26000 -13602
rect 25460 -13922 26000 -13838
rect 25460 -14158 25618 -13922
rect 25854 -14158 26000 -13922
rect 25460 -14242 26000 -14158
rect 25460 -14478 25618 -14242
rect 25854 -14478 26000 -14242
rect 25460 -14562 26000 -14478
rect 25460 -14798 25618 -14562
rect 25854 -14798 26000 -14562
rect 25460 -14882 26000 -14798
rect 25460 -15118 25618 -14882
rect 25854 -15118 26000 -14882
rect 25460 -15202 26000 -15118
rect 25460 -15438 25618 -15202
rect 25854 -15438 26000 -15202
rect 25460 -15522 26000 -15438
rect 25460 -15758 25618 -15522
rect 25854 -15758 26000 -15522
rect 25460 -15842 26000 -15758
rect 25460 -16078 25618 -15842
rect 25854 -16078 26000 -15842
rect 25460 -16162 26000 -16078
rect 25460 -16398 25618 -16162
rect 25854 -16398 26000 -16162
rect 25460 -16482 26000 -16398
rect 25460 -16718 25618 -16482
rect 25854 -16718 26000 -16482
rect 25460 -16802 26000 -16718
rect 25460 -17038 25618 -16802
rect 25854 -17038 26000 -16802
rect 25460 -17122 26000 -17038
rect 25460 -17358 25618 -17122
rect 25854 -17358 26000 -17122
rect 25460 -17442 26000 -17358
rect 25460 -17678 25618 -17442
rect 25854 -17678 26000 -17442
rect 25460 -17762 26000 -17678
rect 25460 -17998 25618 -17762
rect 25854 -17998 26000 -17762
rect 25460 -18082 26000 -17998
rect 25460 -18318 25618 -18082
rect 25854 -18318 26000 -18082
rect 25460 -18402 26000 -18318
rect 25460 -18460 25618 -18402
rect 18388 -18612 25618 -18460
rect 18388 -18638 18522 -18612
rect 18000 -18848 18522 -18638
rect 18758 -18848 18842 -18612
rect 19078 -18848 19162 -18612
rect 19398 -18848 19482 -18612
rect 19718 -18848 19802 -18612
rect 20038 -18848 20122 -18612
rect 20358 -18848 20442 -18612
rect 20678 -18848 20762 -18612
rect 20998 -18848 21082 -18612
rect 21318 -18848 21402 -18612
rect 21638 -18848 21722 -18612
rect 21958 -18848 22042 -18612
rect 22278 -18848 22362 -18612
rect 22598 -18848 22682 -18612
rect 22918 -18848 23002 -18612
rect 23238 -18848 23322 -18612
rect 23558 -18848 23642 -18612
rect 23878 -18848 23962 -18612
rect 24198 -18848 24282 -18612
rect 24518 -18848 24602 -18612
rect 24838 -18848 24922 -18612
rect 25158 -18848 25242 -18612
rect 25478 -18638 25618 -18612
rect 25854 -18638 26000 -18402
rect 25478 -18848 26000 -18638
rect 18000 -19000 26000 -18848
rect 30000 -11156 38000 -11000
rect 30000 -11362 30522 -11156
rect 30000 -11598 30152 -11362
rect 30388 -11392 30522 -11362
rect 30758 -11392 30842 -11156
rect 31078 -11392 31162 -11156
rect 31398 -11392 31482 -11156
rect 31718 -11392 31802 -11156
rect 32038 -11392 32122 -11156
rect 32358 -11392 32442 -11156
rect 32678 -11392 32762 -11156
rect 32998 -11392 33082 -11156
rect 33318 -11392 33402 -11156
rect 33638 -11392 33722 -11156
rect 33958 -11392 34042 -11156
rect 34278 -11392 34362 -11156
rect 34598 -11392 34682 -11156
rect 34918 -11392 35002 -11156
rect 35238 -11392 35322 -11156
rect 35558 -11392 35642 -11156
rect 35878 -11392 35962 -11156
rect 36198 -11392 36282 -11156
rect 36518 -11392 36602 -11156
rect 36838 -11392 36922 -11156
rect 37158 -11392 37242 -11156
rect 37478 -11362 38000 -11156
rect 37478 -11392 37618 -11362
rect 30388 -11540 37618 -11392
rect 30388 -11598 30540 -11540
rect 30000 -11682 30540 -11598
rect 30000 -11918 30152 -11682
rect 30388 -11918 30540 -11682
rect 30000 -12002 30540 -11918
rect 30000 -12238 30152 -12002
rect 30388 -12238 30540 -12002
rect 30000 -12322 30540 -12238
rect 30000 -12558 30152 -12322
rect 30388 -12558 30540 -12322
rect 30000 -12642 30540 -12558
rect 30000 -12878 30152 -12642
rect 30388 -12878 30540 -12642
rect 30000 -12962 30540 -12878
rect 30000 -13198 30152 -12962
rect 30388 -13198 30540 -12962
rect 30000 -13282 30540 -13198
rect 30000 -13518 30152 -13282
rect 30388 -13518 30540 -13282
rect 30000 -13602 30540 -13518
rect 30000 -13838 30152 -13602
rect 30388 -13838 30540 -13602
rect 30000 -13922 30540 -13838
rect 30000 -14158 30152 -13922
rect 30388 -14158 30540 -13922
rect 30000 -14242 30540 -14158
rect 30000 -14478 30152 -14242
rect 30388 -14478 30540 -14242
rect 30000 -14562 30540 -14478
rect 30000 -14798 30152 -14562
rect 30388 -14798 30540 -14562
rect 30000 -14882 30540 -14798
rect 30000 -15118 30152 -14882
rect 30388 -15118 30540 -14882
rect 30000 -15202 30540 -15118
rect 30000 -15438 30152 -15202
rect 30388 -15438 30540 -15202
rect 30000 -15522 30540 -15438
rect 30000 -15758 30152 -15522
rect 30388 -15758 30540 -15522
rect 30000 -15842 30540 -15758
rect 30000 -16078 30152 -15842
rect 30388 -16078 30540 -15842
rect 30000 -16162 30540 -16078
rect 30000 -16398 30152 -16162
rect 30388 -16398 30540 -16162
rect 30000 -16482 30540 -16398
rect 30000 -16718 30152 -16482
rect 30388 -16718 30540 -16482
rect 30000 -16802 30540 -16718
rect 30000 -17038 30152 -16802
rect 30388 -17038 30540 -16802
rect 30000 -17122 30540 -17038
rect 30000 -17358 30152 -17122
rect 30388 -17358 30540 -17122
rect 30000 -17442 30540 -17358
rect 30000 -17678 30152 -17442
rect 30388 -17678 30540 -17442
rect 30000 -17762 30540 -17678
rect 30000 -17998 30152 -17762
rect 30388 -17998 30540 -17762
rect 30000 -18082 30540 -17998
rect 30000 -18318 30152 -18082
rect 30388 -18318 30540 -18082
rect 30000 -18402 30540 -18318
rect 30000 -18638 30152 -18402
rect 30388 -18460 30540 -18402
rect 37460 -11598 37618 -11540
rect 37854 -11598 38000 -11362
rect 38500 -11300 38700 -10900
rect 42000 -11156 50000 -11000
rect 42000 -11300 42522 -11156
rect 38500 -11362 42522 -11300
rect 38500 -11500 42152 -11362
rect 42388 -11392 42522 -11362
rect 42758 -11392 42842 -11156
rect 43078 -11392 43162 -11156
rect 43398 -11392 43482 -11156
rect 43718 -11392 43802 -11156
rect 44038 -11392 44122 -11156
rect 44358 -11392 44442 -11156
rect 44678 -11392 44762 -11156
rect 44998 -11392 45082 -11156
rect 45318 -11392 45402 -11156
rect 45638 -11392 45722 -11156
rect 45958 -11392 46042 -11156
rect 46278 -11392 46362 -11156
rect 46598 -11392 46682 -11156
rect 46918 -11392 47002 -11156
rect 47238 -11392 47322 -11156
rect 47558 -11392 47642 -11156
rect 47878 -11392 47962 -11156
rect 48198 -11392 48282 -11156
rect 48518 -11392 48602 -11156
rect 48838 -11392 48922 -11156
rect 49158 -11392 49242 -11156
rect 49478 -11362 50000 -11156
rect 49478 -11392 49618 -11362
rect 37460 -11682 38000 -11598
rect 37460 -11918 37618 -11682
rect 37854 -11918 38000 -11682
rect 37460 -12002 38000 -11918
rect 37460 -12238 37618 -12002
rect 37854 -12238 38000 -12002
rect 37460 -12322 38000 -12238
rect 37460 -12558 37618 -12322
rect 37854 -12558 38000 -12322
rect 37460 -12642 38000 -12558
rect 37460 -12878 37618 -12642
rect 37854 -12878 38000 -12642
rect 37460 -12962 38000 -12878
rect 37460 -13198 37618 -12962
rect 37854 -13198 38000 -12962
rect 37460 -13282 38000 -13198
rect 37460 -13518 37618 -13282
rect 37854 -13518 38000 -13282
rect 37460 -13602 38000 -13518
rect 37460 -13838 37618 -13602
rect 37854 -13838 38000 -13602
rect 37460 -13922 38000 -13838
rect 37460 -14158 37618 -13922
rect 37854 -14158 38000 -13922
rect 37460 -14242 38000 -14158
rect 37460 -14478 37618 -14242
rect 37854 -14478 38000 -14242
rect 37460 -14562 38000 -14478
rect 37460 -14798 37618 -14562
rect 37854 -14798 38000 -14562
rect 37460 -14882 38000 -14798
rect 37460 -15118 37618 -14882
rect 37854 -15118 38000 -14882
rect 37460 -15202 38000 -15118
rect 37460 -15438 37618 -15202
rect 37854 -15438 38000 -15202
rect 37460 -15522 38000 -15438
rect 37460 -15758 37618 -15522
rect 37854 -15758 38000 -15522
rect 37460 -15842 38000 -15758
rect 37460 -16078 37618 -15842
rect 37854 -16078 38000 -15842
rect 37460 -16162 38000 -16078
rect 37460 -16398 37618 -16162
rect 37854 -16398 38000 -16162
rect 37460 -16482 38000 -16398
rect 37460 -16718 37618 -16482
rect 37854 -16718 38000 -16482
rect 37460 -16802 38000 -16718
rect 37460 -17038 37618 -16802
rect 37854 -17038 38000 -16802
rect 37460 -17122 38000 -17038
rect 37460 -17358 37618 -17122
rect 37854 -17358 38000 -17122
rect 37460 -17442 38000 -17358
rect 37460 -17678 37618 -17442
rect 37854 -17678 38000 -17442
rect 37460 -17762 38000 -17678
rect 37460 -17998 37618 -17762
rect 37854 -17998 38000 -17762
rect 37460 -18082 38000 -17998
rect 37460 -18318 37618 -18082
rect 37854 -18318 38000 -18082
rect 37460 -18402 38000 -18318
rect 37460 -18460 37618 -18402
rect 30388 -18612 37618 -18460
rect 30388 -18638 30522 -18612
rect 30000 -18848 30522 -18638
rect 30758 -18848 30842 -18612
rect 31078 -18848 31162 -18612
rect 31398 -18848 31482 -18612
rect 31718 -18848 31802 -18612
rect 32038 -18848 32122 -18612
rect 32358 -18848 32442 -18612
rect 32678 -18848 32762 -18612
rect 32998 -18848 33082 -18612
rect 33318 -18848 33402 -18612
rect 33638 -18848 33722 -18612
rect 33958 -18848 34042 -18612
rect 34278 -18848 34362 -18612
rect 34598 -18848 34682 -18612
rect 34918 -18848 35002 -18612
rect 35238 -18848 35322 -18612
rect 35558 -18848 35642 -18612
rect 35878 -18848 35962 -18612
rect 36198 -18848 36282 -18612
rect 36518 -18848 36602 -18612
rect 36838 -18848 36922 -18612
rect 37158 -18848 37242 -18612
rect 37478 -18638 37618 -18612
rect 37854 -18638 38000 -18402
rect 37478 -18848 38000 -18638
rect 30000 -19000 38000 -18848
rect 42000 -11598 42152 -11500
rect 42388 -11540 49618 -11392
rect 42388 -11598 42540 -11540
rect 42000 -11682 42540 -11598
rect 42000 -11918 42152 -11682
rect 42388 -11918 42540 -11682
rect 42000 -12002 42540 -11918
rect 42000 -12238 42152 -12002
rect 42388 -12238 42540 -12002
rect 42000 -12322 42540 -12238
rect 42000 -12558 42152 -12322
rect 42388 -12558 42540 -12322
rect 42000 -12642 42540 -12558
rect 42000 -12878 42152 -12642
rect 42388 -12878 42540 -12642
rect 42000 -12962 42540 -12878
rect 42000 -13198 42152 -12962
rect 42388 -13198 42540 -12962
rect 42000 -13282 42540 -13198
rect 42000 -13518 42152 -13282
rect 42388 -13518 42540 -13282
rect 42000 -13602 42540 -13518
rect 42000 -13838 42152 -13602
rect 42388 -13838 42540 -13602
rect 42000 -13922 42540 -13838
rect 42000 -14158 42152 -13922
rect 42388 -14158 42540 -13922
rect 42000 -14242 42540 -14158
rect 42000 -14478 42152 -14242
rect 42388 -14478 42540 -14242
rect 42000 -14562 42540 -14478
rect 42000 -14798 42152 -14562
rect 42388 -14798 42540 -14562
rect 42000 -14882 42540 -14798
rect 42000 -15118 42152 -14882
rect 42388 -15118 42540 -14882
rect 42000 -15202 42540 -15118
rect 42000 -15438 42152 -15202
rect 42388 -15438 42540 -15202
rect 42000 -15522 42540 -15438
rect 42000 -15758 42152 -15522
rect 42388 -15758 42540 -15522
rect 42000 -15842 42540 -15758
rect 42000 -16078 42152 -15842
rect 42388 -16078 42540 -15842
rect 42000 -16162 42540 -16078
rect 42000 -16398 42152 -16162
rect 42388 -16398 42540 -16162
rect 42000 -16482 42540 -16398
rect 42000 -16718 42152 -16482
rect 42388 -16718 42540 -16482
rect 42000 -16802 42540 -16718
rect 42000 -17038 42152 -16802
rect 42388 -17038 42540 -16802
rect 42000 -17122 42540 -17038
rect 42000 -17358 42152 -17122
rect 42388 -17358 42540 -17122
rect 42000 -17442 42540 -17358
rect 42000 -17678 42152 -17442
rect 42388 -17678 42540 -17442
rect 42000 -17762 42540 -17678
rect 42000 -17998 42152 -17762
rect 42388 -17998 42540 -17762
rect 42000 -18082 42540 -17998
rect 42000 -18318 42152 -18082
rect 42388 -18318 42540 -18082
rect 42000 -18402 42540 -18318
rect 42000 -18638 42152 -18402
rect 42388 -18460 42540 -18402
rect 49460 -11598 49618 -11540
rect 49854 -11598 50000 -11362
rect 49460 -11682 50000 -11598
rect 49460 -11918 49618 -11682
rect 49854 -11918 50000 -11682
rect 49460 -12002 50000 -11918
rect 49460 -12238 49618 -12002
rect 49854 -12238 50000 -12002
rect 49460 -12322 50000 -12238
rect 49460 -12558 49618 -12322
rect 49854 -12558 50000 -12322
rect 49460 -12642 50000 -12558
rect 49460 -12878 49618 -12642
rect 49854 -12878 50000 -12642
rect 49460 -12962 50000 -12878
rect 49460 -13198 49618 -12962
rect 49854 -13198 50000 -12962
rect 49460 -13282 50000 -13198
rect 49460 -13518 49618 -13282
rect 49854 -13518 50000 -13282
rect 49460 -13602 50000 -13518
rect 49460 -13838 49618 -13602
rect 49854 -13838 50000 -13602
rect 49460 -13922 50000 -13838
rect 49460 -14158 49618 -13922
rect 49854 -14158 50000 -13922
rect 49460 -14242 50000 -14158
rect 49460 -14478 49618 -14242
rect 49854 -14478 50000 -14242
rect 49460 -14562 50000 -14478
rect 49460 -14798 49618 -14562
rect 49854 -14798 50000 -14562
rect 49460 -14882 50000 -14798
rect 49460 -15118 49618 -14882
rect 49854 -15118 50000 -14882
rect 49460 -15202 50000 -15118
rect 49460 -15438 49618 -15202
rect 49854 -15438 50000 -15202
rect 49460 -15522 50000 -15438
rect 49460 -15758 49618 -15522
rect 49854 -15758 50000 -15522
rect 49460 -15842 50000 -15758
rect 49460 -16078 49618 -15842
rect 49854 -16078 50000 -15842
rect 49460 -16162 50000 -16078
rect 49460 -16398 49618 -16162
rect 49854 -16398 50000 -16162
rect 49460 -16482 50000 -16398
rect 49460 -16718 49618 -16482
rect 49854 -16718 50000 -16482
rect 49460 -16802 50000 -16718
rect 49460 -17038 49618 -16802
rect 49854 -17038 50000 -16802
rect 49460 -17122 50000 -17038
rect 49460 -17358 49618 -17122
rect 49854 -17358 50000 -17122
rect 49460 -17442 50000 -17358
rect 49460 -17678 49618 -17442
rect 49854 -17678 50000 -17442
rect 49460 -17762 50000 -17678
rect 49460 -17998 49618 -17762
rect 49854 -17998 50000 -17762
rect 49460 -18082 50000 -17998
rect 49460 -18318 49618 -18082
rect 49854 -18318 50000 -18082
rect 49460 -18402 50000 -18318
rect 49460 -18460 49618 -18402
rect 42388 -18612 49618 -18460
rect 42388 -18638 42522 -18612
rect 42000 -18848 42522 -18638
rect 42758 -18848 42842 -18612
rect 43078 -18848 43162 -18612
rect 43398 -18848 43482 -18612
rect 43718 -18848 43802 -18612
rect 44038 -18848 44122 -18612
rect 44358 -18848 44442 -18612
rect 44678 -18848 44762 -18612
rect 44998 -18848 45082 -18612
rect 45318 -18848 45402 -18612
rect 45638 -18848 45722 -18612
rect 45958 -18848 46042 -18612
rect 46278 -18848 46362 -18612
rect 46598 -18848 46682 -18612
rect 46918 -18848 47002 -18612
rect 47238 -18848 47322 -18612
rect 47558 -18848 47642 -18612
rect 47878 -18848 47962 -18612
rect 48198 -18848 48282 -18612
rect 48518 -18848 48602 -18612
rect 48838 -18848 48922 -18612
rect 49158 -18848 49242 -18612
rect 49478 -18638 49618 -18612
rect 49854 -18638 50000 -18402
rect 49478 -18848 50000 -18638
rect 42000 -19000 50000 -18848
rect 6100 -19600 6300 -19100
rect 6500 -19600 6700 -19100
rect 6100 -19700 6700 -19600
rect 6900 -19200 7400 -19100
rect 7700 -19200 8200 -19100
rect 6900 -19300 7500 -19200
rect 6900 -19700 7100 -19300
rect 7300 -19700 7500 -19300
rect 6200 -19800 6600 -19700
rect 6900 -19800 7500 -19700
rect 7700 -19300 8300 -19200
rect 7700 -19700 7900 -19300
rect 8100 -19700 8300 -19300
rect 18100 -19600 18300 -19100
rect 18500 -19600 18700 -19100
rect 18900 -19300 19500 -19100
rect 19700 -19300 20300 -19100
rect 18900 -19400 19100 -19300
rect 19700 -19400 19900 -19300
rect 18900 -19500 19400 -19400
rect 19700 -19500 20200 -19400
rect 19000 -19600 19500 -19500
rect 19800 -19600 20300 -19500
rect 18100 -19700 18700 -19600
rect 19300 -19700 19500 -19600
rect 20100 -19700 20300 -19600
rect 30100 -19600 30300 -19100
rect 30500 -19600 30700 -19100
rect 30900 -19300 31500 -19100
rect 30100 -19700 30700 -19600
rect 31100 -19700 31300 -19300
rect 31900 -19400 32100 -19200
rect 31700 -19600 32300 -19400
rect 42100 -19600 42300 -19100
rect 42500 -19600 42700 -19100
rect 43000 -19200 43400 -19100
rect 7700 -19800 8300 -19700
rect 18200 -19800 18600 -19700
rect 6300 -19900 6500 -19800
rect 6900 -19900 7400 -19800
rect 7700 -19900 8200 -19800
rect 18300 -19900 18500 -19800
rect 18900 -19900 19500 -19700
rect 19700 -19900 20300 -19700
rect 30200 -19800 30600 -19700
rect 30300 -19900 30500 -19800
rect 30900 -19900 31500 -19700
rect 31900 -19800 32100 -19600
rect 42100 -19700 42700 -19600
rect 42900 -19300 43500 -19200
rect 42900 -19700 43100 -19300
rect 43300 -19700 43500 -19300
rect 43900 -19400 44100 -19200
rect 43700 -19600 44300 -19400
rect 42200 -19800 42600 -19700
rect 42900 -19800 43500 -19700
rect 43900 -19800 44100 -19600
rect 42300 -19900 42500 -19800
rect 43000 -19900 43400 -19800
rect 18100 -22000 18700 -21900
rect 6100 -22300 6700 -22100
rect 18100 -22300 18700 -22100
rect 6100 -22400 6300 -22300
rect 18100 -22400 18300 -22300
rect 6100 -22500 6600 -22400
rect 18100 -22500 18600 -22400
rect 6200 -22600 6700 -22500
rect 18200 -22600 18700 -22500
rect 6500 -22700 6700 -22600
rect 18500 -22700 18700 -22600
rect 30100 -22600 30300 -22100
rect 30500 -22600 30700 -22100
rect 30100 -22700 30700 -22600
rect 30900 -22200 31400 -22100
rect 30900 -22300 31500 -22200
rect 30900 -22500 31100 -22300
rect 31300 -22500 31500 -22300
rect 31700 -22300 32300 -22100
rect 32500 -22300 33100 -22100
rect 31700 -22400 31900 -22300
rect 32500 -22400 32700 -22300
rect 30900 -22700 31400 -22500
rect 31700 -22600 32200 -22400
rect 32500 -22600 33000 -22400
rect 42100 -22600 42300 -22100
rect 42500 -22600 42700 -22100
rect 42900 -22300 43500 -22100
rect 31700 -22700 31900 -22600
rect 6100 -22900 6700 -22700
rect 18100 -22900 18700 -22700
rect 30200 -22800 30600 -22700
rect 30300 -22900 30500 -22800
rect 30900 -22900 31100 -22700
rect 31300 -22900 31500 -22700
rect 31700 -22900 32300 -22700
rect 32500 -22900 32700 -22600
rect 42100 -22700 42700 -22600
rect 43100 -22700 43300 -22300
rect 43700 -22600 44300 -22400
rect 42200 -22800 42600 -22700
rect 42300 -22900 42500 -22800
rect 42900 -22900 43500 -22700
rect 6000 -23156 14000 -23000
rect 6000 -23362 6522 -23156
rect 6000 -23598 6152 -23362
rect 6388 -23392 6522 -23362
rect 6758 -23392 6842 -23156
rect 7078 -23392 7162 -23156
rect 7398 -23392 7482 -23156
rect 7718 -23392 7802 -23156
rect 8038 -23392 8122 -23156
rect 8358 -23392 8442 -23156
rect 8678 -23392 8762 -23156
rect 8998 -23392 9082 -23156
rect 9318 -23392 9402 -23156
rect 9638 -23392 9722 -23156
rect 9958 -23392 10042 -23156
rect 10278 -23392 10362 -23156
rect 10598 -23392 10682 -23156
rect 10918 -23392 11002 -23156
rect 11238 -23392 11322 -23156
rect 11558 -23392 11642 -23156
rect 11878 -23392 11962 -23156
rect 12198 -23392 12282 -23156
rect 12518 -23392 12602 -23156
rect 12838 -23392 12922 -23156
rect 13158 -23392 13242 -23156
rect 13478 -23362 14000 -23156
rect 13478 -23392 13618 -23362
rect 6388 -23540 13618 -23392
rect 6388 -23598 6540 -23540
rect 6000 -23682 6540 -23598
rect 6000 -23918 6152 -23682
rect 6388 -23918 6540 -23682
rect 6000 -24002 6540 -23918
rect 6000 -24238 6152 -24002
rect 6388 -24238 6540 -24002
rect 6000 -24322 6540 -24238
rect 6000 -24558 6152 -24322
rect 6388 -24558 6540 -24322
rect 6000 -24642 6540 -24558
rect 6000 -24878 6152 -24642
rect 6388 -24878 6540 -24642
rect 6000 -24962 6540 -24878
rect 6000 -25198 6152 -24962
rect 6388 -25198 6540 -24962
rect 6000 -25282 6540 -25198
rect 6000 -25518 6152 -25282
rect 6388 -25518 6540 -25282
rect 6000 -25602 6540 -25518
rect 6000 -25838 6152 -25602
rect 6388 -25838 6540 -25602
rect 6000 -25922 6540 -25838
rect 6000 -26158 6152 -25922
rect 6388 -26158 6540 -25922
rect 6000 -26242 6540 -26158
rect 6000 -26478 6152 -26242
rect 6388 -26478 6540 -26242
rect 6000 -26562 6540 -26478
rect 6000 -26798 6152 -26562
rect 6388 -26798 6540 -26562
rect 6000 -26882 6540 -26798
rect 6000 -27118 6152 -26882
rect 6388 -27118 6540 -26882
rect 6000 -27202 6540 -27118
rect 6000 -27438 6152 -27202
rect 6388 -27438 6540 -27202
rect 6000 -27522 6540 -27438
rect 6000 -27758 6152 -27522
rect 6388 -27758 6540 -27522
rect 6000 -27842 6540 -27758
rect 6000 -28078 6152 -27842
rect 6388 -28078 6540 -27842
rect 6000 -28162 6540 -28078
rect 6000 -28398 6152 -28162
rect 6388 -28398 6540 -28162
rect 6000 -28482 6540 -28398
rect 6000 -28718 6152 -28482
rect 6388 -28718 6540 -28482
rect 6000 -28802 6540 -28718
rect 6000 -29038 6152 -28802
rect 6388 -29038 6540 -28802
rect 6000 -29122 6540 -29038
rect 6000 -29358 6152 -29122
rect 6388 -29358 6540 -29122
rect 6000 -29442 6540 -29358
rect 6000 -29678 6152 -29442
rect 6388 -29678 6540 -29442
rect 6000 -29762 6540 -29678
rect 6000 -29998 6152 -29762
rect 6388 -29998 6540 -29762
rect 6000 -30082 6540 -29998
rect 6000 -30318 6152 -30082
rect 6388 -30318 6540 -30082
rect 6000 -30402 6540 -30318
rect 6000 -30638 6152 -30402
rect 6388 -30460 6540 -30402
rect 13460 -23598 13618 -23540
rect 13854 -23598 14000 -23362
rect 13460 -23682 14000 -23598
rect 13460 -23918 13618 -23682
rect 13854 -23918 14000 -23682
rect 13460 -24002 14000 -23918
rect 13460 -24238 13618 -24002
rect 13854 -24238 14000 -24002
rect 13460 -24322 14000 -24238
rect 13460 -24558 13618 -24322
rect 13854 -24558 14000 -24322
rect 13460 -24642 14000 -24558
rect 13460 -24878 13618 -24642
rect 13854 -24878 14000 -24642
rect 13460 -24962 14000 -24878
rect 13460 -25198 13618 -24962
rect 13854 -25198 14000 -24962
rect 13460 -25282 14000 -25198
rect 13460 -25518 13618 -25282
rect 13854 -25518 14000 -25282
rect 13460 -25602 14000 -25518
rect 13460 -25838 13618 -25602
rect 13854 -25838 14000 -25602
rect 13460 -25922 14000 -25838
rect 13460 -26158 13618 -25922
rect 13854 -26158 14000 -25922
rect 13460 -26242 14000 -26158
rect 13460 -26478 13618 -26242
rect 13854 -26478 14000 -26242
rect 13460 -26562 14000 -26478
rect 13460 -26798 13618 -26562
rect 13854 -26798 14000 -26562
rect 13460 -26882 14000 -26798
rect 13460 -27118 13618 -26882
rect 13854 -27118 14000 -26882
rect 13460 -27202 14000 -27118
rect 13460 -27438 13618 -27202
rect 13854 -27438 14000 -27202
rect 13460 -27522 14000 -27438
rect 13460 -27758 13618 -27522
rect 13854 -27758 14000 -27522
rect 13460 -27842 14000 -27758
rect 13460 -28078 13618 -27842
rect 13854 -28078 14000 -27842
rect 13460 -28162 14000 -28078
rect 13460 -28398 13618 -28162
rect 13854 -28398 14000 -28162
rect 13460 -28482 14000 -28398
rect 13460 -28718 13618 -28482
rect 13854 -28718 14000 -28482
rect 13460 -28802 14000 -28718
rect 13460 -29038 13618 -28802
rect 13854 -29038 14000 -28802
rect 13460 -29122 14000 -29038
rect 13460 -29358 13618 -29122
rect 13854 -29358 14000 -29122
rect 13460 -29442 14000 -29358
rect 13460 -29678 13618 -29442
rect 13854 -29678 14000 -29442
rect 13460 -29762 14000 -29678
rect 13460 -29998 13618 -29762
rect 13854 -29998 14000 -29762
rect 13460 -30082 14000 -29998
rect 13460 -30318 13618 -30082
rect 13854 -30318 14000 -30082
rect 13460 -30402 14000 -30318
rect 13460 -30460 13618 -30402
rect 6388 -30612 13618 -30460
rect 6388 -30638 6522 -30612
rect 6000 -30848 6522 -30638
rect 6758 -30848 6842 -30612
rect 7078 -30848 7162 -30612
rect 7398 -30848 7482 -30612
rect 7718 -30848 7802 -30612
rect 8038 -30848 8122 -30612
rect 8358 -30848 8442 -30612
rect 8678 -30848 8762 -30612
rect 8998 -30848 9082 -30612
rect 9318 -30848 9402 -30612
rect 9638 -30848 9722 -30612
rect 9958 -30848 10042 -30612
rect 10278 -30848 10362 -30612
rect 10598 -30848 10682 -30612
rect 10918 -30848 11002 -30612
rect 11238 -30848 11322 -30612
rect 11558 -30848 11642 -30612
rect 11878 -30848 11962 -30612
rect 12198 -30848 12282 -30612
rect 12518 -30848 12602 -30612
rect 12838 -30848 12922 -30612
rect 13158 -30848 13242 -30612
rect 13478 -30638 13618 -30612
rect 13854 -30638 14000 -30402
rect 13478 -30848 14000 -30638
rect 6000 -31000 14000 -30848
rect 18000 -23156 26000 -23000
rect 18000 -23362 18522 -23156
rect 18000 -23598 18152 -23362
rect 18388 -23392 18522 -23362
rect 18758 -23392 18842 -23156
rect 19078 -23392 19162 -23156
rect 19398 -23392 19482 -23156
rect 19718 -23392 19802 -23156
rect 20038 -23392 20122 -23156
rect 20358 -23392 20442 -23156
rect 20678 -23392 20762 -23156
rect 20998 -23392 21082 -23156
rect 21318 -23392 21402 -23156
rect 21638 -23392 21722 -23156
rect 21958 -23392 22042 -23156
rect 22278 -23392 22362 -23156
rect 22598 -23392 22682 -23156
rect 22918 -23392 23002 -23156
rect 23238 -23392 23322 -23156
rect 23558 -23392 23642 -23156
rect 23878 -23392 23962 -23156
rect 24198 -23392 24282 -23156
rect 24518 -23392 24602 -23156
rect 24838 -23392 24922 -23156
rect 25158 -23392 25242 -23156
rect 25478 -23362 26000 -23156
rect 25478 -23392 25618 -23362
rect 18388 -23540 25618 -23392
rect 18388 -23598 18540 -23540
rect 18000 -23682 18540 -23598
rect 18000 -23918 18152 -23682
rect 18388 -23918 18540 -23682
rect 18000 -24002 18540 -23918
rect 18000 -24238 18152 -24002
rect 18388 -24238 18540 -24002
rect 18000 -24322 18540 -24238
rect 18000 -24558 18152 -24322
rect 18388 -24558 18540 -24322
rect 18000 -24642 18540 -24558
rect 18000 -24878 18152 -24642
rect 18388 -24878 18540 -24642
rect 18000 -24962 18540 -24878
rect 18000 -25198 18152 -24962
rect 18388 -25198 18540 -24962
rect 18000 -25282 18540 -25198
rect 18000 -25518 18152 -25282
rect 18388 -25518 18540 -25282
rect 18000 -25602 18540 -25518
rect 18000 -25838 18152 -25602
rect 18388 -25838 18540 -25602
rect 18000 -25922 18540 -25838
rect 18000 -26158 18152 -25922
rect 18388 -26158 18540 -25922
rect 18000 -26242 18540 -26158
rect 18000 -26478 18152 -26242
rect 18388 -26478 18540 -26242
rect 18000 -26562 18540 -26478
rect 18000 -26798 18152 -26562
rect 18388 -26798 18540 -26562
rect 18000 -26882 18540 -26798
rect 18000 -27118 18152 -26882
rect 18388 -27118 18540 -26882
rect 18000 -27202 18540 -27118
rect 18000 -27438 18152 -27202
rect 18388 -27438 18540 -27202
rect 18000 -27522 18540 -27438
rect 18000 -27758 18152 -27522
rect 18388 -27758 18540 -27522
rect 18000 -27842 18540 -27758
rect 18000 -28078 18152 -27842
rect 18388 -28078 18540 -27842
rect 18000 -28162 18540 -28078
rect 18000 -28398 18152 -28162
rect 18388 -28398 18540 -28162
rect 18000 -28482 18540 -28398
rect 18000 -28718 18152 -28482
rect 18388 -28718 18540 -28482
rect 18000 -28802 18540 -28718
rect 18000 -29038 18152 -28802
rect 18388 -29038 18540 -28802
rect 18000 -29122 18540 -29038
rect 18000 -29358 18152 -29122
rect 18388 -29358 18540 -29122
rect 18000 -29442 18540 -29358
rect 18000 -29678 18152 -29442
rect 18388 -29678 18540 -29442
rect 18000 -29762 18540 -29678
rect 18000 -29998 18152 -29762
rect 18388 -29998 18540 -29762
rect 18000 -30082 18540 -29998
rect 18000 -30318 18152 -30082
rect 18388 -30318 18540 -30082
rect 18000 -30402 18540 -30318
rect 18000 -30638 18152 -30402
rect 18388 -30460 18540 -30402
rect 25460 -23598 25618 -23540
rect 25854 -23598 26000 -23362
rect 25460 -23682 26000 -23598
rect 25460 -23918 25618 -23682
rect 25854 -23918 26000 -23682
rect 25460 -24002 26000 -23918
rect 25460 -24238 25618 -24002
rect 25854 -24238 26000 -24002
rect 25460 -24322 26000 -24238
rect 25460 -24558 25618 -24322
rect 25854 -24558 26000 -24322
rect 25460 -24642 26000 -24558
rect 25460 -24878 25618 -24642
rect 25854 -24878 26000 -24642
rect 25460 -24962 26000 -24878
rect 25460 -25198 25618 -24962
rect 25854 -25198 26000 -24962
rect 25460 -25282 26000 -25198
rect 25460 -25518 25618 -25282
rect 25854 -25518 26000 -25282
rect 25460 -25602 26000 -25518
rect 25460 -25838 25618 -25602
rect 25854 -25838 26000 -25602
rect 25460 -25922 26000 -25838
rect 25460 -26158 25618 -25922
rect 25854 -26158 26000 -25922
rect 25460 -26242 26000 -26158
rect 25460 -26478 25618 -26242
rect 25854 -26478 26000 -26242
rect 25460 -26562 26000 -26478
rect 25460 -26798 25618 -26562
rect 25854 -26798 26000 -26562
rect 25460 -26882 26000 -26798
rect 25460 -27118 25618 -26882
rect 25854 -27118 26000 -26882
rect 25460 -27202 26000 -27118
rect 25460 -27438 25618 -27202
rect 25854 -27438 26000 -27202
rect 25460 -27522 26000 -27438
rect 25460 -27758 25618 -27522
rect 25854 -27758 26000 -27522
rect 25460 -27842 26000 -27758
rect 25460 -28078 25618 -27842
rect 25854 -28078 26000 -27842
rect 25460 -28162 26000 -28078
rect 25460 -28398 25618 -28162
rect 25854 -28398 26000 -28162
rect 25460 -28482 26000 -28398
rect 25460 -28718 25618 -28482
rect 25854 -28718 26000 -28482
rect 25460 -28802 26000 -28718
rect 25460 -29038 25618 -28802
rect 25854 -29038 26000 -28802
rect 25460 -29122 26000 -29038
rect 25460 -29358 25618 -29122
rect 25854 -29358 26000 -29122
rect 25460 -29442 26000 -29358
rect 25460 -29678 25618 -29442
rect 25854 -29678 26000 -29442
rect 25460 -29762 26000 -29678
rect 25460 -29998 25618 -29762
rect 25854 -29998 26000 -29762
rect 25460 -30082 26000 -29998
rect 25460 -30318 25618 -30082
rect 25854 -30318 26000 -30082
rect 25460 -30402 26000 -30318
rect 25460 -30460 25618 -30402
rect 18388 -30612 25618 -30460
rect 18388 -30638 18522 -30612
rect 18000 -30848 18522 -30638
rect 18758 -30848 18842 -30612
rect 19078 -30848 19162 -30612
rect 19398 -30848 19482 -30612
rect 19718 -30848 19802 -30612
rect 20038 -30848 20122 -30612
rect 20358 -30848 20442 -30612
rect 20678 -30848 20762 -30612
rect 20998 -30848 21082 -30612
rect 21318 -30848 21402 -30612
rect 21638 -30848 21722 -30612
rect 21958 -30848 22042 -30612
rect 22278 -30848 22362 -30612
rect 22598 -30848 22682 -30612
rect 22918 -30848 23002 -30612
rect 23238 -30848 23322 -30612
rect 23558 -30848 23642 -30612
rect 23878 -30848 23962 -30612
rect 24198 -30848 24282 -30612
rect 24518 -30848 24602 -30612
rect 24838 -30848 24922 -30612
rect 25158 -30848 25242 -30612
rect 25478 -30638 25618 -30612
rect 25854 -30638 26000 -30402
rect 25478 -30848 26000 -30638
rect 18000 -31000 26000 -30848
rect 30000 -23156 38000 -23000
rect 30000 -23362 30522 -23156
rect 30000 -23598 30152 -23362
rect 30388 -23392 30522 -23362
rect 30758 -23392 30842 -23156
rect 31078 -23392 31162 -23156
rect 31398 -23392 31482 -23156
rect 31718 -23392 31802 -23156
rect 32038 -23392 32122 -23156
rect 32358 -23392 32442 -23156
rect 32678 -23392 32762 -23156
rect 32998 -23392 33082 -23156
rect 33318 -23392 33402 -23156
rect 33638 -23392 33722 -23156
rect 33958 -23392 34042 -23156
rect 34278 -23392 34362 -23156
rect 34598 -23392 34682 -23156
rect 34918 -23392 35002 -23156
rect 35238 -23392 35322 -23156
rect 35558 -23392 35642 -23156
rect 35878 -23392 35962 -23156
rect 36198 -23392 36282 -23156
rect 36518 -23392 36602 -23156
rect 36838 -23392 36922 -23156
rect 37158 -23392 37242 -23156
rect 37478 -23362 38000 -23156
rect 37478 -23392 37618 -23362
rect 30388 -23540 37618 -23392
rect 30388 -23598 30540 -23540
rect 30000 -23682 30540 -23598
rect 30000 -23918 30152 -23682
rect 30388 -23918 30540 -23682
rect 30000 -24002 30540 -23918
rect 30000 -24238 30152 -24002
rect 30388 -24238 30540 -24002
rect 30000 -24322 30540 -24238
rect 30000 -24558 30152 -24322
rect 30388 -24558 30540 -24322
rect 30000 -24642 30540 -24558
rect 30000 -24878 30152 -24642
rect 30388 -24878 30540 -24642
rect 30000 -24962 30540 -24878
rect 30000 -25198 30152 -24962
rect 30388 -25198 30540 -24962
rect 30000 -25282 30540 -25198
rect 30000 -25518 30152 -25282
rect 30388 -25518 30540 -25282
rect 30000 -25602 30540 -25518
rect 30000 -25838 30152 -25602
rect 30388 -25838 30540 -25602
rect 30000 -25922 30540 -25838
rect 30000 -26158 30152 -25922
rect 30388 -26158 30540 -25922
rect 30000 -26242 30540 -26158
rect 30000 -26478 30152 -26242
rect 30388 -26478 30540 -26242
rect 30000 -26562 30540 -26478
rect 30000 -26798 30152 -26562
rect 30388 -26798 30540 -26562
rect 30000 -26882 30540 -26798
rect 30000 -27118 30152 -26882
rect 30388 -27118 30540 -26882
rect 30000 -27202 30540 -27118
rect 30000 -27438 30152 -27202
rect 30388 -27438 30540 -27202
rect 30000 -27522 30540 -27438
rect 30000 -27758 30152 -27522
rect 30388 -27758 30540 -27522
rect 30000 -27842 30540 -27758
rect 30000 -28078 30152 -27842
rect 30388 -28078 30540 -27842
rect 30000 -28162 30540 -28078
rect 30000 -28398 30152 -28162
rect 30388 -28398 30540 -28162
rect 30000 -28482 30540 -28398
rect 30000 -28718 30152 -28482
rect 30388 -28718 30540 -28482
rect 30000 -28802 30540 -28718
rect 30000 -29038 30152 -28802
rect 30388 -29038 30540 -28802
rect 30000 -29122 30540 -29038
rect 30000 -29358 30152 -29122
rect 30388 -29358 30540 -29122
rect 30000 -29442 30540 -29358
rect 30000 -29678 30152 -29442
rect 30388 -29678 30540 -29442
rect 30000 -29762 30540 -29678
rect 30000 -29998 30152 -29762
rect 30388 -29998 30540 -29762
rect 30000 -30082 30540 -29998
rect 30000 -30318 30152 -30082
rect 30388 -30318 30540 -30082
rect 30000 -30402 30540 -30318
rect 30000 -30638 30152 -30402
rect 30388 -30460 30540 -30402
rect 37460 -23598 37618 -23540
rect 37854 -23598 38000 -23362
rect 37460 -23682 38000 -23598
rect 37460 -23918 37618 -23682
rect 37854 -23918 38000 -23682
rect 37460 -24002 38000 -23918
rect 37460 -24238 37618 -24002
rect 37854 -24238 38000 -24002
rect 37460 -24322 38000 -24238
rect 37460 -24558 37618 -24322
rect 37854 -24558 38000 -24322
rect 37460 -24642 38000 -24558
rect 37460 -24878 37618 -24642
rect 37854 -24878 38000 -24642
rect 37460 -24962 38000 -24878
rect 37460 -25198 37618 -24962
rect 37854 -25198 38000 -24962
rect 37460 -25282 38000 -25198
rect 37460 -25518 37618 -25282
rect 37854 -25518 38000 -25282
rect 37460 -25602 38000 -25518
rect 37460 -25838 37618 -25602
rect 37854 -25838 38000 -25602
rect 37460 -25922 38000 -25838
rect 37460 -26158 37618 -25922
rect 37854 -26158 38000 -25922
rect 37460 -26242 38000 -26158
rect 37460 -26478 37618 -26242
rect 37854 -26478 38000 -26242
rect 37460 -26562 38000 -26478
rect 37460 -26798 37618 -26562
rect 37854 -26798 38000 -26562
rect 37460 -26882 38000 -26798
rect 37460 -27118 37618 -26882
rect 37854 -27118 38000 -26882
rect 37460 -27202 38000 -27118
rect 37460 -27438 37618 -27202
rect 37854 -27438 38000 -27202
rect 37460 -27522 38000 -27438
rect 37460 -27758 37618 -27522
rect 37854 -27758 38000 -27522
rect 37460 -27842 38000 -27758
rect 37460 -28078 37618 -27842
rect 37854 -28078 38000 -27842
rect 37460 -28162 38000 -28078
rect 37460 -28398 37618 -28162
rect 37854 -28398 38000 -28162
rect 37460 -28482 38000 -28398
rect 37460 -28718 37618 -28482
rect 37854 -28718 38000 -28482
rect 37460 -28802 38000 -28718
rect 37460 -29038 37618 -28802
rect 37854 -29038 38000 -28802
rect 37460 -29122 38000 -29038
rect 37460 -29358 37618 -29122
rect 37854 -29358 38000 -29122
rect 37460 -29442 38000 -29358
rect 37460 -29678 37618 -29442
rect 37854 -29678 38000 -29442
rect 37460 -29762 38000 -29678
rect 37460 -29998 37618 -29762
rect 37854 -29998 38000 -29762
rect 37460 -30082 38000 -29998
rect 37460 -30318 37618 -30082
rect 37854 -30318 38000 -30082
rect 37460 -30402 38000 -30318
rect 37460 -30460 37618 -30402
rect 30388 -30612 37618 -30460
rect 30388 -30638 30522 -30612
rect 30000 -30848 30522 -30638
rect 30758 -30848 30842 -30612
rect 31078 -30848 31162 -30612
rect 31398 -30848 31482 -30612
rect 31718 -30848 31802 -30612
rect 32038 -30848 32122 -30612
rect 32358 -30848 32442 -30612
rect 32678 -30848 32762 -30612
rect 32998 -30848 33082 -30612
rect 33318 -30848 33402 -30612
rect 33638 -30848 33722 -30612
rect 33958 -30848 34042 -30612
rect 34278 -30848 34362 -30612
rect 34598 -30848 34682 -30612
rect 34918 -30848 35002 -30612
rect 35238 -30848 35322 -30612
rect 35558 -30848 35642 -30612
rect 35878 -30848 35962 -30612
rect 36198 -30848 36282 -30612
rect 36518 -30848 36602 -30612
rect 36838 -30848 36922 -30612
rect 37158 -30848 37242 -30612
rect 37478 -30638 37618 -30612
rect 37854 -30638 38000 -30402
rect 37478 -30848 38000 -30638
rect 30000 -31000 38000 -30848
rect 42000 -23156 50000 -23000
rect 42000 -23362 42522 -23156
rect 42000 -23598 42152 -23362
rect 42388 -23392 42522 -23362
rect 42758 -23392 42842 -23156
rect 43078 -23392 43162 -23156
rect 43398 -23392 43482 -23156
rect 43718 -23392 43802 -23156
rect 44038 -23392 44122 -23156
rect 44358 -23392 44442 -23156
rect 44678 -23392 44762 -23156
rect 44998 -23392 45082 -23156
rect 45318 -23392 45402 -23156
rect 45638 -23392 45722 -23156
rect 45958 -23392 46042 -23156
rect 46278 -23392 46362 -23156
rect 46598 -23392 46682 -23156
rect 46918 -23392 47002 -23156
rect 47238 -23392 47322 -23156
rect 47558 -23392 47642 -23156
rect 47878 -23392 47962 -23156
rect 48198 -23392 48282 -23156
rect 48518 -23392 48602 -23156
rect 48838 -23392 48922 -23156
rect 49158 -23392 49242 -23156
rect 49478 -23362 50000 -23156
rect 49478 -23392 49618 -23362
rect 42388 -23540 49618 -23392
rect 42388 -23598 42540 -23540
rect 42000 -23682 42540 -23598
rect 42000 -23918 42152 -23682
rect 42388 -23918 42540 -23682
rect 42000 -24002 42540 -23918
rect 42000 -24238 42152 -24002
rect 42388 -24238 42540 -24002
rect 42000 -24322 42540 -24238
rect 42000 -24558 42152 -24322
rect 42388 -24558 42540 -24322
rect 42000 -24642 42540 -24558
rect 42000 -24878 42152 -24642
rect 42388 -24878 42540 -24642
rect 42000 -24962 42540 -24878
rect 42000 -25198 42152 -24962
rect 42388 -25198 42540 -24962
rect 42000 -25282 42540 -25198
rect 42000 -25518 42152 -25282
rect 42388 -25518 42540 -25282
rect 42000 -25602 42540 -25518
rect 42000 -25838 42152 -25602
rect 42388 -25838 42540 -25602
rect 42000 -25922 42540 -25838
rect 42000 -26158 42152 -25922
rect 42388 -26158 42540 -25922
rect 42000 -26242 42540 -26158
rect 42000 -26478 42152 -26242
rect 42388 -26478 42540 -26242
rect 42000 -26562 42540 -26478
rect 42000 -26798 42152 -26562
rect 42388 -26798 42540 -26562
rect 42000 -26882 42540 -26798
rect 42000 -27118 42152 -26882
rect 42388 -27118 42540 -26882
rect 42000 -27202 42540 -27118
rect 42000 -27438 42152 -27202
rect 42388 -27438 42540 -27202
rect 42000 -27522 42540 -27438
rect 42000 -27758 42152 -27522
rect 42388 -27758 42540 -27522
rect 42000 -27842 42540 -27758
rect 42000 -28078 42152 -27842
rect 42388 -28078 42540 -27842
rect 42000 -28162 42540 -28078
rect 42000 -28398 42152 -28162
rect 42388 -28398 42540 -28162
rect 42000 -28482 42540 -28398
rect 42000 -28718 42152 -28482
rect 42388 -28718 42540 -28482
rect 42000 -28802 42540 -28718
rect 42000 -29038 42152 -28802
rect 42388 -29038 42540 -28802
rect 42000 -29122 42540 -29038
rect 42000 -29358 42152 -29122
rect 42388 -29358 42540 -29122
rect 42000 -29442 42540 -29358
rect 42000 -29678 42152 -29442
rect 42388 -29678 42540 -29442
rect 42000 -29762 42540 -29678
rect 42000 -29998 42152 -29762
rect 42388 -29998 42540 -29762
rect 42000 -30082 42540 -29998
rect 42000 -30318 42152 -30082
rect 42388 -30318 42540 -30082
rect 42000 -30402 42540 -30318
rect 42000 -30638 42152 -30402
rect 42388 -30460 42540 -30402
rect 49460 -23598 49618 -23540
rect 49854 -23598 50000 -23362
rect 49460 -23682 50000 -23598
rect 49460 -23918 49618 -23682
rect 49854 -23918 50000 -23682
rect 49460 -24002 50000 -23918
rect 49460 -24238 49618 -24002
rect 49854 -24238 50000 -24002
rect 49460 -24322 50000 -24238
rect 49460 -24558 49618 -24322
rect 49854 -24558 50000 -24322
rect 49460 -24642 50000 -24558
rect 49460 -24878 49618 -24642
rect 49854 -24878 50000 -24642
rect 49460 -24962 50000 -24878
rect 49460 -25198 49618 -24962
rect 49854 -25198 50000 -24962
rect 49460 -25282 50000 -25198
rect 49460 -25518 49618 -25282
rect 49854 -25518 50000 -25282
rect 49460 -25602 50000 -25518
rect 49460 -25838 49618 -25602
rect 49854 -25838 50000 -25602
rect 49460 -25922 50000 -25838
rect 49460 -26158 49618 -25922
rect 49854 -26158 50000 -25922
rect 49460 -26242 50000 -26158
rect 49460 -26478 49618 -26242
rect 49854 -26478 50000 -26242
rect 49460 -26562 50000 -26478
rect 49460 -26798 49618 -26562
rect 49854 -26798 50000 -26562
rect 49460 -26882 50000 -26798
rect 49460 -27118 49618 -26882
rect 49854 -27118 50000 -26882
rect 49460 -27202 50000 -27118
rect 49460 -27438 49618 -27202
rect 49854 -27438 50000 -27202
rect 49460 -27522 50000 -27438
rect 49460 -27758 49618 -27522
rect 49854 -27758 50000 -27522
rect 49460 -27842 50000 -27758
rect 49460 -28078 49618 -27842
rect 49854 -28078 50000 -27842
rect 49460 -28162 50000 -28078
rect 49460 -28398 49618 -28162
rect 49854 -28398 50000 -28162
rect 49460 -28482 50000 -28398
rect 49460 -28718 49618 -28482
rect 49854 -28718 50000 -28482
rect 49460 -28802 50000 -28718
rect 49460 -29038 49618 -28802
rect 49854 -29038 50000 -28802
rect 49460 -29122 50000 -29038
rect 49460 -29358 49618 -29122
rect 49854 -29358 50000 -29122
rect 49460 -29442 50000 -29358
rect 49460 -29678 49618 -29442
rect 49854 -29678 50000 -29442
rect 49460 -29762 50000 -29678
rect 49460 -29998 49618 -29762
rect 49854 -29998 50000 -29762
rect 49460 -30082 50000 -29998
rect 49460 -30318 49618 -30082
rect 49854 -30318 50000 -30082
rect 49460 -30402 50000 -30318
rect 49460 -30460 49618 -30402
rect 42388 -30612 49618 -30460
rect 42388 -30638 42522 -30612
rect 42000 -30848 42522 -30638
rect 42758 -30848 42842 -30612
rect 43078 -30848 43162 -30612
rect 43398 -30848 43482 -30612
rect 43718 -30848 43802 -30612
rect 44038 -30848 44122 -30612
rect 44358 -30848 44442 -30612
rect 44678 -30848 44762 -30612
rect 44998 -30848 45082 -30612
rect 45318 -30848 45402 -30612
rect 45638 -30848 45722 -30612
rect 45958 -30848 46042 -30612
rect 46278 -30848 46362 -30612
rect 46598 -30848 46682 -30612
rect 46918 -30848 47002 -30612
rect 47238 -30848 47322 -30612
rect 47558 -30848 47642 -30612
rect 47878 -30848 47962 -30612
rect 48198 -30848 48282 -30612
rect 48518 -30848 48602 -30612
rect 48838 -30848 48922 -30612
rect 49158 -30848 49242 -30612
rect 49478 -30638 49618 -30612
rect 49854 -30638 50000 -30402
rect 49478 -30848 50000 -30638
rect 42000 -31000 50000 -30848
<< via4 >>
rect 22432 -5960 22972 -5720
rect 16500 -9148 17200 -8748
rect 13300 -10200 15900 -9600
rect 6522 -11242 6758 -11156
rect 6522 -11306 6608 -11242
rect 6608 -11306 6672 -11242
rect 6672 -11306 6758 -11242
rect 6152 -11448 6388 -11362
rect 6522 -11392 6758 -11306
rect 6842 -11242 7078 -11156
rect 6842 -11306 6928 -11242
rect 6928 -11306 6992 -11242
rect 6992 -11306 7078 -11242
rect 6842 -11392 7078 -11306
rect 7162 -11242 7398 -11156
rect 7162 -11306 7248 -11242
rect 7248 -11306 7312 -11242
rect 7312 -11306 7398 -11242
rect 7162 -11392 7398 -11306
rect 7482 -11242 7718 -11156
rect 7482 -11306 7568 -11242
rect 7568 -11306 7632 -11242
rect 7632 -11306 7718 -11242
rect 7482 -11392 7718 -11306
rect 7802 -11242 8038 -11156
rect 7802 -11306 7888 -11242
rect 7888 -11306 7952 -11242
rect 7952 -11306 8038 -11242
rect 7802 -11392 8038 -11306
rect 8122 -11242 8358 -11156
rect 8122 -11306 8208 -11242
rect 8208 -11306 8272 -11242
rect 8272 -11306 8358 -11242
rect 8122 -11392 8358 -11306
rect 8442 -11242 8678 -11156
rect 8442 -11306 8528 -11242
rect 8528 -11306 8592 -11242
rect 8592 -11306 8678 -11242
rect 8442 -11392 8678 -11306
rect 8762 -11242 8998 -11156
rect 8762 -11306 8848 -11242
rect 8848 -11306 8912 -11242
rect 8912 -11306 8998 -11242
rect 8762 -11392 8998 -11306
rect 9082 -11242 9318 -11156
rect 9082 -11306 9168 -11242
rect 9168 -11306 9232 -11242
rect 9232 -11306 9318 -11242
rect 9082 -11392 9318 -11306
rect 9402 -11242 9638 -11156
rect 9402 -11306 9488 -11242
rect 9488 -11306 9552 -11242
rect 9552 -11306 9638 -11242
rect 9402 -11392 9638 -11306
rect 9722 -11242 9958 -11156
rect 9722 -11306 9808 -11242
rect 9808 -11306 9872 -11242
rect 9872 -11306 9958 -11242
rect 9722 -11392 9958 -11306
rect 10042 -11242 10278 -11156
rect 10042 -11306 10128 -11242
rect 10128 -11306 10192 -11242
rect 10192 -11306 10278 -11242
rect 10042 -11392 10278 -11306
rect 10362 -11242 10598 -11156
rect 10362 -11306 10448 -11242
rect 10448 -11306 10512 -11242
rect 10512 -11306 10598 -11242
rect 10362 -11392 10598 -11306
rect 10682 -11242 10918 -11156
rect 10682 -11306 10768 -11242
rect 10768 -11306 10832 -11242
rect 10832 -11306 10918 -11242
rect 10682 -11392 10918 -11306
rect 11002 -11242 11238 -11156
rect 11002 -11306 11088 -11242
rect 11088 -11306 11152 -11242
rect 11152 -11306 11238 -11242
rect 11002 -11392 11238 -11306
rect 11322 -11242 11558 -11156
rect 11322 -11306 11408 -11242
rect 11408 -11306 11472 -11242
rect 11472 -11306 11558 -11242
rect 11322 -11392 11558 -11306
rect 11642 -11242 11878 -11156
rect 11642 -11306 11728 -11242
rect 11728 -11306 11792 -11242
rect 11792 -11306 11878 -11242
rect 11642 -11392 11878 -11306
rect 11962 -11242 12198 -11156
rect 11962 -11306 12048 -11242
rect 12048 -11306 12112 -11242
rect 12112 -11306 12198 -11242
rect 11962 -11392 12198 -11306
rect 12282 -11242 12518 -11156
rect 12282 -11306 12368 -11242
rect 12368 -11306 12432 -11242
rect 12432 -11306 12518 -11242
rect 12282 -11392 12518 -11306
rect 12602 -11242 12838 -11156
rect 12602 -11306 12688 -11242
rect 12688 -11306 12752 -11242
rect 12752 -11306 12838 -11242
rect 12602 -11392 12838 -11306
rect 12922 -11242 13158 -11156
rect 12922 -11306 13008 -11242
rect 13008 -11306 13072 -11242
rect 13072 -11306 13158 -11242
rect 12922 -11392 13158 -11306
rect 13242 -11242 13478 -11156
rect 13242 -11306 13328 -11242
rect 13328 -11306 13392 -11242
rect 13392 -11306 13478 -11242
rect 13242 -11392 13478 -11306
rect 6152 -11512 6238 -11448
rect 6238 -11512 6302 -11448
rect 6302 -11512 6388 -11448
rect 6152 -11598 6388 -11512
rect 13618 -11448 13854 -11362
rect 13618 -11512 13704 -11448
rect 13704 -11512 13768 -11448
rect 13768 -11512 13854 -11448
rect 6152 -11768 6388 -11682
rect 6152 -11832 6238 -11768
rect 6238 -11832 6302 -11768
rect 6302 -11832 6388 -11768
rect 6152 -11918 6388 -11832
rect 6152 -12088 6388 -12002
rect 6152 -12152 6238 -12088
rect 6238 -12152 6302 -12088
rect 6302 -12152 6388 -12088
rect 6152 -12238 6388 -12152
rect 6152 -12408 6388 -12322
rect 6152 -12472 6238 -12408
rect 6238 -12472 6302 -12408
rect 6302 -12472 6388 -12408
rect 6152 -12558 6388 -12472
rect 6152 -12728 6388 -12642
rect 6152 -12792 6238 -12728
rect 6238 -12792 6302 -12728
rect 6302 -12792 6388 -12728
rect 6152 -12878 6388 -12792
rect 6152 -13048 6388 -12962
rect 6152 -13112 6238 -13048
rect 6238 -13112 6302 -13048
rect 6302 -13112 6388 -13048
rect 6152 -13198 6388 -13112
rect 6152 -13368 6388 -13282
rect 6152 -13432 6238 -13368
rect 6238 -13432 6302 -13368
rect 6302 -13432 6388 -13368
rect 6152 -13518 6388 -13432
rect 6152 -13688 6388 -13602
rect 6152 -13752 6238 -13688
rect 6238 -13752 6302 -13688
rect 6302 -13752 6388 -13688
rect 6152 -13838 6388 -13752
rect 6152 -14008 6388 -13922
rect 6152 -14072 6238 -14008
rect 6238 -14072 6302 -14008
rect 6302 -14072 6388 -14008
rect 6152 -14158 6388 -14072
rect 6152 -14328 6388 -14242
rect 6152 -14392 6238 -14328
rect 6238 -14392 6302 -14328
rect 6302 -14392 6388 -14328
rect 6152 -14478 6388 -14392
rect 6152 -14648 6388 -14562
rect 6152 -14712 6238 -14648
rect 6238 -14712 6302 -14648
rect 6302 -14712 6388 -14648
rect 6152 -14798 6388 -14712
rect 6152 -14968 6388 -14882
rect 6152 -15032 6238 -14968
rect 6238 -15032 6302 -14968
rect 6302 -15032 6388 -14968
rect 6152 -15118 6388 -15032
rect 6152 -15288 6388 -15202
rect 6152 -15352 6238 -15288
rect 6238 -15352 6302 -15288
rect 6302 -15352 6388 -15288
rect 6152 -15438 6388 -15352
rect 6152 -15608 6388 -15522
rect 6152 -15672 6238 -15608
rect 6238 -15672 6302 -15608
rect 6302 -15672 6388 -15608
rect 6152 -15758 6388 -15672
rect 6152 -15928 6388 -15842
rect 6152 -15992 6238 -15928
rect 6238 -15992 6302 -15928
rect 6302 -15992 6388 -15928
rect 6152 -16078 6388 -15992
rect 6152 -16248 6388 -16162
rect 6152 -16312 6238 -16248
rect 6238 -16312 6302 -16248
rect 6302 -16312 6388 -16248
rect 6152 -16398 6388 -16312
rect 6152 -16568 6388 -16482
rect 6152 -16632 6238 -16568
rect 6238 -16632 6302 -16568
rect 6302 -16632 6388 -16568
rect 6152 -16718 6388 -16632
rect 6152 -16888 6388 -16802
rect 6152 -16952 6238 -16888
rect 6238 -16952 6302 -16888
rect 6302 -16952 6388 -16888
rect 6152 -17038 6388 -16952
rect 6152 -17208 6388 -17122
rect 6152 -17272 6238 -17208
rect 6238 -17272 6302 -17208
rect 6302 -17272 6388 -17208
rect 6152 -17358 6388 -17272
rect 6152 -17528 6388 -17442
rect 6152 -17592 6238 -17528
rect 6238 -17592 6302 -17528
rect 6302 -17592 6388 -17528
rect 6152 -17678 6388 -17592
rect 6152 -17848 6388 -17762
rect 6152 -17912 6238 -17848
rect 6238 -17912 6302 -17848
rect 6302 -17912 6388 -17848
rect 6152 -17998 6388 -17912
rect 6152 -18168 6388 -18082
rect 6152 -18232 6238 -18168
rect 6238 -18232 6302 -18168
rect 6302 -18232 6388 -18168
rect 6152 -18318 6388 -18232
rect 6152 -18488 6388 -18402
rect 13618 -11598 13854 -11512
rect 13618 -11768 13854 -11682
rect 13618 -11832 13704 -11768
rect 13704 -11832 13768 -11768
rect 13768 -11832 13854 -11768
rect 13618 -11918 13854 -11832
rect 13618 -12088 13854 -12002
rect 13618 -12152 13704 -12088
rect 13704 -12152 13768 -12088
rect 13768 -12152 13854 -12088
rect 13618 -12238 13854 -12152
rect 13618 -12408 13854 -12322
rect 13618 -12472 13704 -12408
rect 13704 -12472 13768 -12408
rect 13768 -12472 13854 -12408
rect 13618 -12558 13854 -12472
rect 13618 -12728 13854 -12642
rect 13618 -12792 13704 -12728
rect 13704 -12792 13768 -12728
rect 13768 -12792 13854 -12728
rect 13618 -12878 13854 -12792
rect 13618 -13048 13854 -12962
rect 13618 -13112 13704 -13048
rect 13704 -13112 13768 -13048
rect 13768 -13112 13854 -13048
rect 13618 -13198 13854 -13112
rect 13618 -13368 13854 -13282
rect 13618 -13432 13704 -13368
rect 13704 -13432 13768 -13368
rect 13768 -13432 13854 -13368
rect 13618 -13518 13854 -13432
rect 13618 -13688 13854 -13602
rect 13618 -13752 13704 -13688
rect 13704 -13752 13768 -13688
rect 13768 -13752 13854 -13688
rect 13618 -13838 13854 -13752
rect 13618 -14008 13854 -13922
rect 13618 -14072 13704 -14008
rect 13704 -14072 13768 -14008
rect 13768 -14072 13854 -14008
rect 13618 -14158 13854 -14072
rect 13618 -14328 13854 -14242
rect 13618 -14392 13704 -14328
rect 13704 -14392 13768 -14328
rect 13768 -14392 13854 -14328
rect 13618 -14478 13854 -14392
rect 13618 -14648 13854 -14562
rect 13618 -14712 13704 -14648
rect 13704 -14712 13768 -14648
rect 13768 -14712 13854 -14648
rect 13618 -14798 13854 -14712
rect 13618 -14968 13854 -14882
rect 13618 -15032 13704 -14968
rect 13704 -15032 13768 -14968
rect 13768 -15032 13854 -14968
rect 13618 -15118 13854 -15032
rect 13618 -15288 13854 -15202
rect 13618 -15352 13704 -15288
rect 13704 -15352 13768 -15288
rect 13768 -15352 13854 -15288
rect 13618 -15438 13854 -15352
rect 13618 -15608 13854 -15522
rect 13618 -15672 13704 -15608
rect 13704 -15672 13768 -15608
rect 13768 -15672 13854 -15608
rect 13618 -15758 13854 -15672
rect 13618 -15928 13854 -15842
rect 13618 -15992 13704 -15928
rect 13704 -15992 13768 -15928
rect 13768 -15992 13854 -15928
rect 13618 -16078 13854 -15992
rect 13618 -16248 13854 -16162
rect 13618 -16312 13704 -16248
rect 13704 -16312 13768 -16248
rect 13768 -16312 13854 -16248
rect 13618 -16398 13854 -16312
rect 13618 -16568 13854 -16482
rect 13618 -16632 13704 -16568
rect 13704 -16632 13768 -16568
rect 13768 -16632 13854 -16568
rect 13618 -16718 13854 -16632
rect 13618 -16888 13854 -16802
rect 13618 -16952 13704 -16888
rect 13704 -16952 13768 -16888
rect 13768 -16952 13854 -16888
rect 13618 -17038 13854 -16952
rect 13618 -17208 13854 -17122
rect 13618 -17272 13704 -17208
rect 13704 -17272 13768 -17208
rect 13768 -17272 13854 -17208
rect 13618 -17358 13854 -17272
rect 13618 -17528 13854 -17442
rect 13618 -17592 13704 -17528
rect 13704 -17592 13768 -17528
rect 13768 -17592 13854 -17528
rect 13618 -17678 13854 -17592
rect 13618 -17848 13854 -17762
rect 13618 -17912 13704 -17848
rect 13704 -17912 13768 -17848
rect 13768 -17912 13854 -17848
rect 13618 -17998 13854 -17912
rect 13618 -18168 13854 -18082
rect 13618 -18232 13704 -18168
rect 13704 -18232 13768 -18168
rect 13768 -18232 13854 -18168
rect 13618 -18318 13854 -18232
rect 6152 -18552 6238 -18488
rect 6238 -18552 6302 -18488
rect 6302 -18552 6388 -18488
rect 6152 -18638 6388 -18552
rect 13618 -18488 13854 -18402
rect 13618 -18552 13704 -18488
rect 13704 -18552 13768 -18488
rect 13768 -18552 13854 -18488
rect 6522 -18698 6758 -18612
rect 6522 -18762 6608 -18698
rect 6608 -18762 6672 -18698
rect 6672 -18762 6758 -18698
rect 6522 -18848 6758 -18762
rect 6842 -18698 7078 -18612
rect 6842 -18762 6928 -18698
rect 6928 -18762 6992 -18698
rect 6992 -18762 7078 -18698
rect 6842 -18848 7078 -18762
rect 7162 -18698 7398 -18612
rect 7162 -18762 7248 -18698
rect 7248 -18762 7312 -18698
rect 7312 -18762 7398 -18698
rect 7162 -18848 7398 -18762
rect 7482 -18698 7718 -18612
rect 7482 -18762 7568 -18698
rect 7568 -18762 7632 -18698
rect 7632 -18762 7718 -18698
rect 7482 -18848 7718 -18762
rect 7802 -18698 8038 -18612
rect 7802 -18762 7888 -18698
rect 7888 -18762 7952 -18698
rect 7952 -18762 8038 -18698
rect 7802 -18848 8038 -18762
rect 8122 -18698 8358 -18612
rect 8122 -18762 8208 -18698
rect 8208 -18762 8272 -18698
rect 8272 -18762 8358 -18698
rect 8122 -18848 8358 -18762
rect 8442 -18698 8678 -18612
rect 8442 -18762 8528 -18698
rect 8528 -18762 8592 -18698
rect 8592 -18762 8678 -18698
rect 8442 -18848 8678 -18762
rect 8762 -18698 8998 -18612
rect 8762 -18762 8848 -18698
rect 8848 -18762 8912 -18698
rect 8912 -18762 8998 -18698
rect 8762 -18848 8998 -18762
rect 9082 -18698 9318 -18612
rect 9082 -18762 9168 -18698
rect 9168 -18762 9232 -18698
rect 9232 -18762 9318 -18698
rect 9082 -18848 9318 -18762
rect 9402 -18698 9638 -18612
rect 9402 -18762 9488 -18698
rect 9488 -18762 9552 -18698
rect 9552 -18762 9638 -18698
rect 9402 -18848 9638 -18762
rect 9722 -18698 9958 -18612
rect 9722 -18762 9808 -18698
rect 9808 -18762 9872 -18698
rect 9872 -18762 9958 -18698
rect 9722 -18848 9958 -18762
rect 10042 -18698 10278 -18612
rect 10042 -18762 10128 -18698
rect 10128 -18762 10192 -18698
rect 10192 -18762 10278 -18698
rect 10042 -18848 10278 -18762
rect 10362 -18698 10598 -18612
rect 10362 -18762 10448 -18698
rect 10448 -18762 10512 -18698
rect 10512 -18762 10598 -18698
rect 10362 -18848 10598 -18762
rect 10682 -18698 10918 -18612
rect 10682 -18762 10768 -18698
rect 10768 -18762 10832 -18698
rect 10832 -18762 10918 -18698
rect 10682 -18848 10918 -18762
rect 11002 -18698 11238 -18612
rect 11002 -18762 11088 -18698
rect 11088 -18762 11152 -18698
rect 11152 -18762 11238 -18698
rect 11002 -18848 11238 -18762
rect 11322 -18698 11558 -18612
rect 11322 -18762 11408 -18698
rect 11408 -18762 11472 -18698
rect 11472 -18762 11558 -18698
rect 11322 -18848 11558 -18762
rect 11642 -18698 11878 -18612
rect 11642 -18762 11728 -18698
rect 11728 -18762 11792 -18698
rect 11792 -18762 11878 -18698
rect 11642 -18848 11878 -18762
rect 11962 -18698 12198 -18612
rect 11962 -18762 12048 -18698
rect 12048 -18762 12112 -18698
rect 12112 -18762 12198 -18698
rect 11962 -18848 12198 -18762
rect 12282 -18698 12518 -18612
rect 12282 -18762 12368 -18698
rect 12368 -18762 12432 -18698
rect 12432 -18762 12518 -18698
rect 12282 -18848 12518 -18762
rect 12602 -18698 12838 -18612
rect 12602 -18762 12688 -18698
rect 12688 -18762 12752 -18698
rect 12752 -18762 12838 -18698
rect 12602 -18848 12838 -18762
rect 12922 -18698 13158 -18612
rect 12922 -18762 13008 -18698
rect 13008 -18762 13072 -18698
rect 13072 -18762 13158 -18698
rect 12922 -18848 13158 -18762
rect 13242 -18698 13478 -18612
rect 13618 -18638 13854 -18552
rect 13242 -18762 13328 -18698
rect 13328 -18762 13392 -18698
rect 13392 -18762 13478 -18698
rect 13242 -18848 13478 -18762
rect 18522 -11242 18758 -11156
rect 18522 -11306 18608 -11242
rect 18608 -11306 18672 -11242
rect 18672 -11306 18758 -11242
rect 18152 -11448 18388 -11362
rect 18522 -11392 18758 -11306
rect 18842 -11242 19078 -11156
rect 18842 -11306 18928 -11242
rect 18928 -11306 18992 -11242
rect 18992 -11306 19078 -11242
rect 18842 -11392 19078 -11306
rect 19162 -11242 19398 -11156
rect 19162 -11306 19248 -11242
rect 19248 -11306 19312 -11242
rect 19312 -11306 19398 -11242
rect 19162 -11392 19398 -11306
rect 19482 -11242 19718 -11156
rect 19482 -11306 19568 -11242
rect 19568 -11306 19632 -11242
rect 19632 -11306 19718 -11242
rect 19482 -11392 19718 -11306
rect 19802 -11242 20038 -11156
rect 19802 -11306 19888 -11242
rect 19888 -11306 19952 -11242
rect 19952 -11306 20038 -11242
rect 19802 -11392 20038 -11306
rect 20122 -11242 20358 -11156
rect 20122 -11306 20208 -11242
rect 20208 -11306 20272 -11242
rect 20272 -11306 20358 -11242
rect 20122 -11392 20358 -11306
rect 20442 -11242 20678 -11156
rect 20442 -11306 20528 -11242
rect 20528 -11306 20592 -11242
rect 20592 -11306 20678 -11242
rect 20442 -11392 20678 -11306
rect 20762 -11242 20998 -11156
rect 20762 -11306 20848 -11242
rect 20848 -11306 20912 -11242
rect 20912 -11306 20998 -11242
rect 20762 -11392 20998 -11306
rect 21082 -11242 21318 -11156
rect 21082 -11306 21168 -11242
rect 21168 -11306 21232 -11242
rect 21232 -11306 21318 -11242
rect 21082 -11392 21318 -11306
rect 21402 -11242 21638 -11156
rect 21402 -11306 21488 -11242
rect 21488 -11306 21552 -11242
rect 21552 -11306 21638 -11242
rect 21402 -11392 21638 -11306
rect 21722 -11242 21958 -11156
rect 21722 -11306 21808 -11242
rect 21808 -11306 21872 -11242
rect 21872 -11306 21958 -11242
rect 21722 -11392 21958 -11306
rect 22042 -11242 22278 -11156
rect 22042 -11306 22128 -11242
rect 22128 -11306 22192 -11242
rect 22192 -11306 22278 -11242
rect 22042 -11392 22278 -11306
rect 22362 -11242 22598 -11156
rect 22362 -11306 22448 -11242
rect 22448 -11306 22512 -11242
rect 22512 -11306 22598 -11242
rect 22362 -11392 22598 -11306
rect 22682 -11242 22918 -11156
rect 22682 -11306 22768 -11242
rect 22768 -11306 22832 -11242
rect 22832 -11306 22918 -11242
rect 22682 -11392 22918 -11306
rect 23002 -11242 23238 -11156
rect 23002 -11306 23088 -11242
rect 23088 -11306 23152 -11242
rect 23152 -11306 23238 -11242
rect 23002 -11392 23238 -11306
rect 23322 -11242 23558 -11156
rect 23322 -11306 23408 -11242
rect 23408 -11306 23472 -11242
rect 23472 -11306 23558 -11242
rect 23322 -11392 23558 -11306
rect 23642 -11242 23878 -11156
rect 23642 -11306 23728 -11242
rect 23728 -11306 23792 -11242
rect 23792 -11306 23878 -11242
rect 23642 -11392 23878 -11306
rect 23962 -11242 24198 -11156
rect 23962 -11306 24048 -11242
rect 24048 -11306 24112 -11242
rect 24112 -11306 24198 -11242
rect 23962 -11392 24198 -11306
rect 24282 -11242 24518 -11156
rect 24282 -11306 24368 -11242
rect 24368 -11306 24432 -11242
rect 24432 -11306 24518 -11242
rect 24282 -11392 24518 -11306
rect 24602 -11242 24838 -11156
rect 24602 -11306 24688 -11242
rect 24688 -11306 24752 -11242
rect 24752 -11306 24838 -11242
rect 24602 -11392 24838 -11306
rect 24922 -11242 25158 -11156
rect 24922 -11306 25008 -11242
rect 25008 -11306 25072 -11242
rect 25072 -11306 25158 -11242
rect 24922 -11392 25158 -11306
rect 25242 -11242 25478 -11156
rect 25242 -11306 25328 -11242
rect 25328 -11306 25392 -11242
rect 25392 -11306 25478 -11242
rect 25242 -11392 25478 -11306
rect 18152 -11512 18238 -11448
rect 18238 -11512 18302 -11448
rect 18302 -11512 18388 -11448
rect 18152 -11598 18388 -11512
rect 25618 -11448 25854 -11362
rect 25618 -11512 25704 -11448
rect 25704 -11512 25768 -11448
rect 25768 -11512 25854 -11448
rect 18152 -11768 18388 -11682
rect 18152 -11832 18238 -11768
rect 18238 -11832 18302 -11768
rect 18302 -11832 18388 -11768
rect 18152 -11918 18388 -11832
rect 18152 -12088 18388 -12002
rect 18152 -12152 18238 -12088
rect 18238 -12152 18302 -12088
rect 18302 -12152 18388 -12088
rect 18152 -12238 18388 -12152
rect 18152 -12408 18388 -12322
rect 18152 -12472 18238 -12408
rect 18238 -12472 18302 -12408
rect 18302 -12472 18388 -12408
rect 18152 -12558 18388 -12472
rect 18152 -12728 18388 -12642
rect 18152 -12792 18238 -12728
rect 18238 -12792 18302 -12728
rect 18302 -12792 18388 -12728
rect 18152 -12878 18388 -12792
rect 18152 -13048 18388 -12962
rect 18152 -13112 18238 -13048
rect 18238 -13112 18302 -13048
rect 18302 -13112 18388 -13048
rect 18152 -13198 18388 -13112
rect 18152 -13368 18388 -13282
rect 18152 -13432 18238 -13368
rect 18238 -13432 18302 -13368
rect 18302 -13432 18388 -13368
rect 18152 -13518 18388 -13432
rect 18152 -13688 18388 -13602
rect 18152 -13752 18238 -13688
rect 18238 -13752 18302 -13688
rect 18302 -13752 18388 -13688
rect 18152 -13838 18388 -13752
rect 18152 -14008 18388 -13922
rect 18152 -14072 18238 -14008
rect 18238 -14072 18302 -14008
rect 18302 -14072 18388 -14008
rect 18152 -14158 18388 -14072
rect 18152 -14328 18388 -14242
rect 18152 -14392 18238 -14328
rect 18238 -14392 18302 -14328
rect 18302 -14392 18388 -14328
rect 18152 -14478 18388 -14392
rect 18152 -14648 18388 -14562
rect 18152 -14712 18238 -14648
rect 18238 -14712 18302 -14648
rect 18302 -14712 18388 -14648
rect 18152 -14798 18388 -14712
rect 18152 -14968 18388 -14882
rect 18152 -15032 18238 -14968
rect 18238 -15032 18302 -14968
rect 18302 -15032 18388 -14968
rect 18152 -15118 18388 -15032
rect 18152 -15288 18388 -15202
rect 18152 -15352 18238 -15288
rect 18238 -15352 18302 -15288
rect 18302 -15352 18388 -15288
rect 18152 -15438 18388 -15352
rect 18152 -15608 18388 -15522
rect 18152 -15672 18238 -15608
rect 18238 -15672 18302 -15608
rect 18302 -15672 18388 -15608
rect 18152 -15758 18388 -15672
rect 18152 -15928 18388 -15842
rect 18152 -15992 18238 -15928
rect 18238 -15992 18302 -15928
rect 18302 -15992 18388 -15928
rect 18152 -16078 18388 -15992
rect 18152 -16248 18388 -16162
rect 18152 -16312 18238 -16248
rect 18238 -16312 18302 -16248
rect 18302 -16312 18388 -16248
rect 18152 -16398 18388 -16312
rect 18152 -16568 18388 -16482
rect 18152 -16632 18238 -16568
rect 18238 -16632 18302 -16568
rect 18302 -16632 18388 -16568
rect 18152 -16718 18388 -16632
rect 18152 -16888 18388 -16802
rect 18152 -16952 18238 -16888
rect 18238 -16952 18302 -16888
rect 18302 -16952 18388 -16888
rect 18152 -17038 18388 -16952
rect 18152 -17208 18388 -17122
rect 18152 -17272 18238 -17208
rect 18238 -17272 18302 -17208
rect 18302 -17272 18388 -17208
rect 18152 -17358 18388 -17272
rect 18152 -17528 18388 -17442
rect 18152 -17592 18238 -17528
rect 18238 -17592 18302 -17528
rect 18302 -17592 18388 -17528
rect 18152 -17678 18388 -17592
rect 18152 -17848 18388 -17762
rect 18152 -17912 18238 -17848
rect 18238 -17912 18302 -17848
rect 18302 -17912 18388 -17848
rect 18152 -17998 18388 -17912
rect 18152 -18168 18388 -18082
rect 18152 -18232 18238 -18168
rect 18238 -18232 18302 -18168
rect 18302 -18232 18388 -18168
rect 18152 -18318 18388 -18232
rect 18152 -18488 18388 -18402
rect 25618 -11598 25854 -11512
rect 25618 -11768 25854 -11682
rect 25618 -11832 25704 -11768
rect 25704 -11832 25768 -11768
rect 25768 -11832 25854 -11768
rect 25618 -11918 25854 -11832
rect 25618 -12088 25854 -12002
rect 25618 -12152 25704 -12088
rect 25704 -12152 25768 -12088
rect 25768 -12152 25854 -12088
rect 25618 -12238 25854 -12152
rect 25618 -12408 25854 -12322
rect 25618 -12472 25704 -12408
rect 25704 -12472 25768 -12408
rect 25768 -12472 25854 -12408
rect 25618 -12558 25854 -12472
rect 25618 -12728 25854 -12642
rect 25618 -12792 25704 -12728
rect 25704 -12792 25768 -12728
rect 25768 -12792 25854 -12728
rect 25618 -12878 25854 -12792
rect 25618 -13048 25854 -12962
rect 25618 -13112 25704 -13048
rect 25704 -13112 25768 -13048
rect 25768 -13112 25854 -13048
rect 25618 -13198 25854 -13112
rect 25618 -13368 25854 -13282
rect 25618 -13432 25704 -13368
rect 25704 -13432 25768 -13368
rect 25768 -13432 25854 -13368
rect 25618 -13518 25854 -13432
rect 25618 -13688 25854 -13602
rect 25618 -13752 25704 -13688
rect 25704 -13752 25768 -13688
rect 25768 -13752 25854 -13688
rect 25618 -13838 25854 -13752
rect 25618 -14008 25854 -13922
rect 25618 -14072 25704 -14008
rect 25704 -14072 25768 -14008
rect 25768 -14072 25854 -14008
rect 25618 -14158 25854 -14072
rect 25618 -14328 25854 -14242
rect 25618 -14392 25704 -14328
rect 25704 -14392 25768 -14328
rect 25768 -14392 25854 -14328
rect 25618 -14478 25854 -14392
rect 25618 -14648 25854 -14562
rect 25618 -14712 25704 -14648
rect 25704 -14712 25768 -14648
rect 25768 -14712 25854 -14648
rect 25618 -14798 25854 -14712
rect 25618 -14968 25854 -14882
rect 25618 -15032 25704 -14968
rect 25704 -15032 25768 -14968
rect 25768 -15032 25854 -14968
rect 25618 -15118 25854 -15032
rect 25618 -15288 25854 -15202
rect 25618 -15352 25704 -15288
rect 25704 -15352 25768 -15288
rect 25768 -15352 25854 -15288
rect 25618 -15438 25854 -15352
rect 25618 -15608 25854 -15522
rect 25618 -15672 25704 -15608
rect 25704 -15672 25768 -15608
rect 25768 -15672 25854 -15608
rect 25618 -15758 25854 -15672
rect 25618 -15928 25854 -15842
rect 25618 -15992 25704 -15928
rect 25704 -15992 25768 -15928
rect 25768 -15992 25854 -15928
rect 25618 -16078 25854 -15992
rect 25618 -16248 25854 -16162
rect 25618 -16312 25704 -16248
rect 25704 -16312 25768 -16248
rect 25768 -16312 25854 -16248
rect 25618 -16398 25854 -16312
rect 25618 -16568 25854 -16482
rect 25618 -16632 25704 -16568
rect 25704 -16632 25768 -16568
rect 25768 -16632 25854 -16568
rect 25618 -16718 25854 -16632
rect 25618 -16888 25854 -16802
rect 25618 -16952 25704 -16888
rect 25704 -16952 25768 -16888
rect 25768 -16952 25854 -16888
rect 25618 -17038 25854 -16952
rect 25618 -17208 25854 -17122
rect 25618 -17272 25704 -17208
rect 25704 -17272 25768 -17208
rect 25768 -17272 25854 -17208
rect 25618 -17358 25854 -17272
rect 25618 -17528 25854 -17442
rect 25618 -17592 25704 -17528
rect 25704 -17592 25768 -17528
rect 25768 -17592 25854 -17528
rect 25618 -17678 25854 -17592
rect 25618 -17848 25854 -17762
rect 25618 -17912 25704 -17848
rect 25704 -17912 25768 -17848
rect 25768 -17912 25854 -17848
rect 25618 -17998 25854 -17912
rect 25618 -18168 25854 -18082
rect 25618 -18232 25704 -18168
rect 25704 -18232 25768 -18168
rect 25768 -18232 25854 -18168
rect 25618 -18318 25854 -18232
rect 18152 -18552 18238 -18488
rect 18238 -18552 18302 -18488
rect 18302 -18552 18388 -18488
rect 18152 -18638 18388 -18552
rect 25618 -18488 25854 -18402
rect 25618 -18552 25704 -18488
rect 25704 -18552 25768 -18488
rect 25768 -18552 25854 -18488
rect 18522 -18698 18758 -18612
rect 18522 -18762 18608 -18698
rect 18608 -18762 18672 -18698
rect 18672 -18762 18758 -18698
rect 18522 -18848 18758 -18762
rect 18842 -18698 19078 -18612
rect 18842 -18762 18928 -18698
rect 18928 -18762 18992 -18698
rect 18992 -18762 19078 -18698
rect 18842 -18848 19078 -18762
rect 19162 -18698 19398 -18612
rect 19162 -18762 19248 -18698
rect 19248 -18762 19312 -18698
rect 19312 -18762 19398 -18698
rect 19162 -18848 19398 -18762
rect 19482 -18698 19718 -18612
rect 19482 -18762 19568 -18698
rect 19568 -18762 19632 -18698
rect 19632 -18762 19718 -18698
rect 19482 -18848 19718 -18762
rect 19802 -18698 20038 -18612
rect 19802 -18762 19888 -18698
rect 19888 -18762 19952 -18698
rect 19952 -18762 20038 -18698
rect 19802 -18848 20038 -18762
rect 20122 -18698 20358 -18612
rect 20122 -18762 20208 -18698
rect 20208 -18762 20272 -18698
rect 20272 -18762 20358 -18698
rect 20122 -18848 20358 -18762
rect 20442 -18698 20678 -18612
rect 20442 -18762 20528 -18698
rect 20528 -18762 20592 -18698
rect 20592 -18762 20678 -18698
rect 20442 -18848 20678 -18762
rect 20762 -18698 20998 -18612
rect 20762 -18762 20848 -18698
rect 20848 -18762 20912 -18698
rect 20912 -18762 20998 -18698
rect 20762 -18848 20998 -18762
rect 21082 -18698 21318 -18612
rect 21082 -18762 21168 -18698
rect 21168 -18762 21232 -18698
rect 21232 -18762 21318 -18698
rect 21082 -18848 21318 -18762
rect 21402 -18698 21638 -18612
rect 21402 -18762 21488 -18698
rect 21488 -18762 21552 -18698
rect 21552 -18762 21638 -18698
rect 21402 -18848 21638 -18762
rect 21722 -18698 21958 -18612
rect 21722 -18762 21808 -18698
rect 21808 -18762 21872 -18698
rect 21872 -18762 21958 -18698
rect 21722 -18848 21958 -18762
rect 22042 -18698 22278 -18612
rect 22042 -18762 22128 -18698
rect 22128 -18762 22192 -18698
rect 22192 -18762 22278 -18698
rect 22042 -18848 22278 -18762
rect 22362 -18698 22598 -18612
rect 22362 -18762 22448 -18698
rect 22448 -18762 22512 -18698
rect 22512 -18762 22598 -18698
rect 22362 -18848 22598 -18762
rect 22682 -18698 22918 -18612
rect 22682 -18762 22768 -18698
rect 22768 -18762 22832 -18698
rect 22832 -18762 22918 -18698
rect 22682 -18848 22918 -18762
rect 23002 -18698 23238 -18612
rect 23002 -18762 23088 -18698
rect 23088 -18762 23152 -18698
rect 23152 -18762 23238 -18698
rect 23002 -18848 23238 -18762
rect 23322 -18698 23558 -18612
rect 23322 -18762 23408 -18698
rect 23408 -18762 23472 -18698
rect 23472 -18762 23558 -18698
rect 23322 -18848 23558 -18762
rect 23642 -18698 23878 -18612
rect 23642 -18762 23728 -18698
rect 23728 -18762 23792 -18698
rect 23792 -18762 23878 -18698
rect 23642 -18848 23878 -18762
rect 23962 -18698 24198 -18612
rect 23962 -18762 24048 -18698
rect 24048 -18762 24112 -18698
rect 24112 -18762 24198 -18698
rect 23962 -18848 24198 -18762
rect 24282 -18698 24518 -18612
rect 24282 -18762 24368 -18698
rect 24368 -18762 24432 -18698
rect 24432 -18762 24518 -18698
rect 24282 -18848 24518 -18762
rect 24602 -18698 24838 -18612
rect 24602 -18762 24688 -18698
rect 24688 -18762 24752 -18698
rect 24752 -18762 24838 -18698
rect 24602 -18848 24838 -18762
rect 24922 -18698 25158 -18612
rect 24922 -18762 25008 -18698
rect 25008 -18762 25072 -18698
rect 25072 -18762 25158 -18698
rect 24922 -18848 25158 -18762
rect 25242 -18698 25478 -18612
rect 25618 -18638 25854 -18552
rect 25242 -18762 25328 -18698
rect 25328 -18762 25392 -18698
rect 25392 -18762 25478 -18698
rect 25242 -18848 25478 -18762
rect 30522 -11242 30758 -11156
rect 30522 -11306 30608 -11242
rect 30608 -11306 30672 -11242
rect 30672 -11306 30758 -11242
rect 30152 -11448 30388 -11362
rect 30522 -11392 30758 -11306
rect 30842 -11242 31078 -11156
rect 30842 -11306 30928 -11242
rect 30928 -11306 30992 -11242
rect 30992 -11306 31078 -11242
rect 30842 -11392 31078 -11306
rect 31162 -11242 31398 -11156
rect 31162 -11306 31248 -11242
rect 31248 -11306 31312 -11242
rect 31312 -11306 31398 -11242
rect 31162 -11392 31398 -11306
rect 31482 -11242 31718 -11156
rect 31482 -11306 31568 -11242
rect 31568 -11306 31632 -11242
rect 31632 -11306 31718 -11242
rect 31482 -11392 31718 -11306
rect 31802 -11242 32038 -11156
rect 31802 -11306 31888 -11242
rect 31888 -11306 31952 -11242
rect 31952 -11306 32038 -11242
rect 31802 -11392 32038 -11306
rect 32122 -11242 32358 -11156
rect 32122 -11306 32208 -11242
rect 32208 -11306 32272 -11242
rect 32272 -11306 32358 -11242
rect 32122 -11392 32358 -11306
rect 32442 -11242 32678 -11156
rect 32442 -11306 32528 -11242
rect 32528 -11306 32592 -11242
rect 32592 -11306 32678 -11242
rect 32442 -11392 32678 -11306
rect 32762 -11242 32998 -11156
rect 32762 -11306 32848 -11242
rect 32848 -11306 32912 -11242
rect 32912 -11306 32998 -11242
rect 32762 -11392 32998 -11306
rect 33082 -11242 33318 -11156
rect 33082 -11306 33168 -11242
rect 33168 -11306 33232 -11242
rect 33232 -11306 33318 -11242
rect 33082 -11392 33318 -11306
rect 33402 -11242 33638 -11156
rect 33402 -11306 33488 -11242
rect 33488 -11306 33552 -11242
rect 33552 -11306 33638 -11242
rect 33402 -11392 33638 -11306
rect 33722 -11242 33958 -11156
rect 33722 -11306 33808 -11242
rect 33808 -11306 33872 -11242
rect 33872 -11306 33958 -11242
rect 33722 -11392 33958 -11306
rect 34042 -11242 34278 -11156
rect 34042 -11306 34128 -11242
rect 34128 -11306 34192 -11242
rect 34192 -11306 34278 -11242
rect 34042 -11392 34278 -11306
rect 34362 -11242 34598 -11156
rect 34362 -11306 34448 -11242
rect 34448 -11306 34512 -11242
rect 34512 -11306 34598 -11242
rect 34362 -11392 34598 -11306
rect 34682 -11242 34918 -11156
rect 34682 -11306 34768 -11242
rect 34768 -11306 34832 -11242
rect 34832 -11306 34918 -11242
rect 34682 -11392 34918 -11306
rect 35002 -11242 35238 -11156
rect 35002 -11306 35088 -11242
rect 35088 -11306 35152 -11242
rect 35152 -11306 35238 -11242
rect 35002 -11392 35238 -11306
rect 35322 -11242 35558 -11156
rect 35322 -11306 35408 -11242
rect 35408 -11306 35472 -11242
rect 35472 -11306 35558 -11242
rect 35322 -11392 35558 -11306
rect 35642 -11242 35878 -11156
rect 35642 -11306 35728 -11242
rect 35728 -11306 35792 -11242
rect 35792 -11306 35878 -11242
rect 35642 -11392 35878 -11306
rect 35962 -11242 36198 -11156
rect 35962 -11306 36048 -11242
rect 36048 -11306 36112 -11242
rect 36112 -11306 36198 -11242
rect 35962 -11392 36198 -11306
rect 36282 -11242 36518 -11156
rect 36282 -11306 36368 -11242
rect 36368 -11306 36432 -11242
rect 36432 -11306 36518 -11242
rect 36282 -11392 36518 -11306
rect 36602 -11242 36838 -11156
rect 36602 -11306 36688 -11242
rect 36688 -11306 36752 -11242
rect 36752 -11306 36838 -11242
rect 36602 -11392 36838 -11306
rect 36922 -11242 37158 -11156
rect 36922 -11306 37008 -11242
rect 37008 -11306 37072 -11242
rect 37072 -11306 37158 -11242
rect 36922 -11392 37158 -11306
rect 37242 -11242 37478 -11156
rect 37242 -11306 37328 -11242
rect 37328 -11306 37392 -11242
rect 37392 -11306 37478 -11242
rect 37242 -11392 37478 -11306
rect 30152 -11512 30238 -11448
rect 30238 -11512 30302 -11448
rect 30302 -11512 30388 -11448
rect 30152 -11598 30388 -11512
rect 37618 -11448 37854 -11362
rect 37618 -11512 37704 -11448
rect 37704 -11512 37768 -11448
rect 37768 -11512 37854 -11448
rect 30152 -11768 30388 -11682
rect 30152 -11832 30238 -11768
rect 30238 -11832 30302 -11768
rect 30302 -11832 30388 -11768
rect 30152 -11918 30388 -11832
rect 30152 -12088 30388 -12002
rect 30152 -12152 30238 -12088
rect 30238 -12152 30302 -12088
rect 30302 -12152 30388 -12088
rect 30152 -12238 30388 -12152
rect 30152 -12408 30388 -12322
rect 30152 -12472 30238 -12408
rect 30238 -12472 30302 -12408
rect 30302 -12472 30388 -12408
rect 30152 -12558 30388 -12472
rect 30152 -12728 30388 -12642
rect 30152 -12792 30238 -12728
rect 30238 -12792 30302 -12728
rect 30302 -12792 30388 -12728
rect 30152 -12878 30388 -12792
rect 30152 -13048 30388 -12962
rect 30152 -13112 30238 -13048
rect 30238 -13112 30302 -13048
rect 30302 -13112 30388 -13048
rect 30152 -13198 30388 -13112
rect 30152 -13368 30388 -13282
rect 30152 -13432 30238 -13368
rect 30238 -13432 30302 -13368
rect 30302 -13432 30388 -13368
rect 30152 -13518 30388 -13432
rect 30152 -13688 30388 -13602
rect 30152 -13752 30238 -13688
rect 30238 -13752 30302 -13688
rect 30302 -13752 30388 -13688
rect 30152 -13838 30388 -13752
rect 30152 -14008 30388 -13922
rect 30152 -14072 30238 -14008
rect 30238 -14072 30302 -14008
rect 30302 -14072 30388 -14008
rect 30152 -14158 30388 -14072
rect 30152 -14328 30388 -14242
rect 30152 -14392 30238 -14328
rect 30238 -14392 30302 -14328
rect 30302 -14392 30388 -14328
rect 30152 -14478 30388 -14392
rect 30152 -14648 30388 -14562
rect 30152 -14712 30238 -14648
rect 30238 -14712 30302 -14648
rect 30302 -14712 30388 -14648
rect 30152 -14798 30388 -14712
rect 30152 -14968 30388 -14882
rect 30152 -15032 30238 -14968
rect 30238 -15032 30302 -14968
rect 30302 -15032 30388 -14968
rect 30152 -15118 30388 -15032
rect 30152 -15288 30388 -15202
rect 30152 -15352 30238 -15288
rect 30238 -15352 30302 -15288
rect 30302 -15352 30388 -15288
rect 30152 -15438 30388 -15352
rect 30152 -15608 30388 -15522
rect 30152 -15672 30238 -15608
rect 30238 -15672 30302 -15608
rect 30302 -15672 30388 -15608
rect 30152 -15758 30388 -15672
rect 30152 -15928 30388 -15842
rect 30152 -15992 30238 -15928
rect 30238 -15992 30302 -15928
rect 30302 -15992 30388 -15928
rect 30152 -16078 30388 -15992
rect 30152 -16248 30388 -16162
rect 30152 -16312 30238 -16248
rect 30238 -16312 30302 -16248
rect 30302 -16312 30388 -16248
rect 30152 -16398 30388 -16312
rect 30152 -16568 30388 -16482
rect 30152 -16632 30238 -16568
rect 30238 -16632 30302 -16568
rect 30302 -16632 30388 -16568
rect 30152 -16718 30388 -16632
rect 30152 -16888 30388 -16802
rect 30152 -16952 30238 -16888
rect 30238 -16952 30302 -16888
rect 30302 -16952 30388 -16888
rect 30152 -17038 30388 -16952
rect 30152 -17208 30388 -17122
rect 30152 -17272 30238 -17208
rect 30238 -17272 30302 -17208
rect 30302 -17272 30388 -17208
rect 30152 -17358 30388 -17272
rect 30152 -17528 30388 -17442
rect 30152 -17592 30238 -17528
rect 30238 -17592 30302 -17528
rect 30302 -17592 30388 -17528
rect 30152 -17678 30388 -17592
rect 30152 -17848 30388 -17762
rect 30152 -17912 30238 -17848
rect 30238 -17912 30302 -17848
rect 30302 -17912 30388 -17848
rect 30152 -17998 30388 -17912
rect 30152 -18168 30388 -18082
rect 30152 -18232 30238 -18168
rect 30238 -18232 30302 -18168
rect 30302 -18232 30388 -18168
rect 30152 -18318 30388 -18232
rect 30152 -18488 30388 -18402
rect 37618 -11598 37854 -11512
rect 42522 -11242 42758 -11156
rect 42522 -11306 42608 -11242
rect 42608 -11306 42672 -11242
rect 42672 -11306 42758 -11242
rect 42152 -11448 42388 -11362
rect 42522 -11392 42758 -11306
rect 42842 -11242 43078 -11156
rect 42842 -11306 42928 -11242
rect 42928 -11306 42992 -11242
rect 42992 -11306 43078 -11242
rect 42842 -11392 43078 -11306
rect 43162 -11242 43398 -11156
rect 43162 -11306 43248 -11242
rect 43248 -11306 43312 -11242
rect 43312 -11306 43398 -11242
rect 43162 -11392 43398 -11306
rect 43482 -11242 43718 -11156
rect 43482 -11306 43568 -11242
rect 43568 -11306 43632 -11242
rect 43632 -11306 43718 -11242
rect 43482 -11392 43718 -11306
rect 43802 -11242 44038 -11156
rect 43802 -11306 43888 -11242
rect 43888 -11306 43952 -11242
rect 43952 -11306 44038 -11242
rect 43802 -11392 44038 -11306
rect 44122 -11242 44358 -11156
rect 44122 -11306 44208 -11242
rect 44208 -11306 44272 -11242
rect 44272 -11306 44358 -11242
rect 44122 -11392 44358 -11306
rect 44442 -11242 44678 -11156
rect 44442 -11306 44528 -11242
rect 44528 -11306 44592 -11242
rect 44592 -11306 44678 -11242
rect 44442 -11392 44678 -11306
rect 44762 -11242 44998 -11156
rect 44762 -11306 44848 -11242
rect 44848 -11306 44912 -11242
rect 44912 -11306 44998 -11242
rect 44762 -11392 44998 -11306
rect 45082 -11242 45318 -11156
rect 45082 -11306 45168 -11242
rect 45168 -11306 45232 -11242
rect 45232 -11306 45318 -11242
rect 45082 -11392 45318 -11306
rect 45402 -11242 45638 -11156
rect 45402 -11306 45488 -11242
rect 45488 -11306 45552 -11242
rect 45552 -11306 45638 -11242
rect 45402 -11392 45638 -11306
rect 45722 -11242 45958 -11156
rect 45722 -11306 45808 -11242
rect 45808 -11306 45872 -11242
rect 45872 -11306 45958 -11242
rect 45722 -11392 45958 -11306
rect 46042 -11242 46278 -11156
rect 46042 -11306 46128 -11242
rect 46128 -11306 46192 -11242
rect 46192 -11306 46278 -11242
rect 46042 -11392 46278 -11306
rect 46362 -11242 46598 -11156
rect 46362 -11306 46448 -11242
rect 46448 -11306 46512 -11242
rect 46512 -11306 46598 -11242
rect 46362 -11392 46598 -11306
rect 46682 -11242 46918 -11156
rect 46682 -11306 46768 -11242
rect 46768 -11306 46832 -11242
rect 46832 -11306 46918 -11242
rect 46682 -11392 46918 -11306
rect 47002 -11242 47238 -11156
rect 47002 -11306 47088 -11242
rect 47088 -11306 47152 -11242
rect 47152 -11306 47238 -11242
rect 47002 -11392 47238 -11306
rect 47322 -11242 47558 -11156
rect 47322 -11306 47408 -11242
rect 47408 -11306 47472 -11242
rect 47472 -11306 47558 -11242
rect 47322 -11392 47558 -11306
rect 47642 -11242 47878 -11156
rect 47642 -11306 47728 -11242
rect 47728 -11306 47792 -11242
rect 47792 -11306 47878 -11242
rect 47642 -11392 47878 -11306
rect 47962 -11242 48198 -11156
rect 47962 -11306 48048 -11242
rect 48048 -11306 48112 -11242
rect 48112 -11306 48198 -11242
rect 47962 -11392 48198 -11306
rect 48282 -11242 48518 -11156
rect 48282 -11306 48368 -11242
rect 48368 -11306 48432 -11242
rect 48432 -11306 48518 -11242
rect 48282 -11392 48518 -11306
rect 48602 -11242 48838 -11156
rect 48602 -11306 48688 -11242
rect 48688 -11306 48752 -11242
rect 48752 -11306 48838 -11242
rect 48602 -11392 48838 -11306
rect 48922 -11242 49158 -11156
rect 48922 -11306 49008 -11242
rect 49008 -11306 49072 -11242
rect 49072 -11306 49158 -11242
rect 48922 -11392 49158 -11306
rect 49242 -11242 49478 -11156
rect 49242 -11306 49328 -11242
rect 49328 -11306 49392 -11242
rect 49392 -11306 49478 -11242
rect 49242 -11392 49478 -11306
rect 37618 -11768 37854 -11682
rect 37618 -11832 37704 -11768
rect 37704 -11832 37768 -11768
rect 37768 -11832 37854 -11768
rect 37618 -11918 37854 -11832
rect 37618 -12088 37854 -12002
rect 37618 -12152 37704 -12088
rect 37704 -12152 37768 -12088
rect 37768 -12152 37854 -12088
rect 37618 -12238 37854 -12152
rect 37618 -12408 37854 -12322
rect 37618 -12472 37704 -12408
rect 37704 -12472 37768 -12408
rect 37768 -12472 37854 -12408
rect 37618 -12558 37854 -12472
rect 37618 -12728 37854 -12642
rect 37618 -12792 37704 -12728
rect 37704 -12792 37768 -12728
rect 37768 -12792 37854 -12728
rect 37618 -12878 37854 -12792
rect 37618 -13048 37854 -12962
rect 37618 -13112 37704 -13048
rect 37704 -13112 37768 -13048
rect 37768 -13112 37854 -13048
rect 37618 -13198 37854 -13112
rect 37618 -13368 37854 -13282
rect 37618 -13432 37704 -13368
rect 37704 -13432 37768 -13368
rect 37768 -13432 37854 -13368
rect 37618 -13518 37854 -13432
rect 37618 -13688 37854 -13602
rect 37618 -13752 37704 -13688
rect 37704 -13752 37768 -13688
rect 37768 -13752 37854 -13688
rect 37618 -13838 37854 -13752
rect 37618 -14008 37854 -13922
rect 37618 -14072 37704 -14008
rect 37704 -14072 37768 -14008
rect 37768 -14072 37854 -14008
rect 37618 -14158 37854 -14072
rect 37618 -14328 37854 -14242
rect 37618 -14392 37704 -14328
rect 37704 -14392 37768 -14328
rect 37768 -14392 37854 -14328
rect 37618 -14478 37854 -14392
rect 37618 -14648 37854 -14562
rect 37618 -14712 37704 -14648
rect 37704 -14712 37768 -14648
rect 37768 -14712 37854 -14648
rect 37618 -14798 37854 -14712
rect 37618 -14968 37854 -14882
rect 37618 -15032 37704 -14968
rect 37704 -15032 37768 -14968
rect 37768 -15032 37854 -14968
rect 37618 -15118 37854 -15032
rect 37618 -15288 37854 -15202
rect 37618 -15352 37704 -15288
rect 37704 -15352 37768 -15288
rect 37768 -15352 37854 -15288
rect 37618 -15438 37854 -15352
rect 37618 -15608 37854 -15522
rect 37618 -15672 37704 -15608
rect 37704 -15672 37768 -15608
rect 37768 -15672 37854 -15608
rect 37618 -15758 37854 -15672
rect 37618 -15928 37854 -15842
rect 37618 -15992 37704 -15928
rect 37704 -15992 37768 -15928
rect 37768 -15992 37854 -15928
rect 37618 -16078 37854 -15992
rect 37618 -16248 37854 -16162
rect 37618 -16312 37704 -16248
rect 37704 -16312 37768 -16248
rect 37768 -16312 37854 -16248
rect 37618 -16398 37854 -16312
rect 37618 -16568 37854 -16482
rect 37618 -16632 37704 -16568
rect 37704 -16632 37768 -16568
rect 37768 -16632 37854 -16568
rect 37618 -16718 37854 -16632
rect 37618 -16888 37854 -16802
rect 37618 -16952 37704 -16888
rect 37704 -16952 37768 -16888
rect 37768 -16952 37854 -16888
rect 37618 -17038 37854 -16952
rect 37618 -17208 37854 -17122
rect 37618 -17272 37704 -17208
rect 37704 -17272 37768 -17208
rect 37768 -17272 37854 -17208
rect 37618 -17358 37854 -17272
rect 37618 -17528 37854 -17442
rect 37618 -17592 37704 -17528
rect 37704 -17592 37768 -17528
rect 37768 -17592 37854 -17528
rect 37618 -17678 37854 -17592
rect 37618 -17848 37854 -17762
rect 37618 -17912 37704 -17848
rect 37704 -17912 37768 -17848
rect 37768 -17912 37854 -17848
rect 37618 -17998 37854 -17912
rect 37618 -18168 37854 -18082
rect 37618 -18232 37704 -18168
rect 37704 -18232 37768 -18168
rect 37768 -18232 37854 -18168
rect 37618 -18318 37854 -18232
rect 30152 -18552 30238 -18488
rect 30238 -18552 30302 -18488
rect 30302 -18552 30388 -18488
rect 30152 -18638 30388 -18552
rect 37618 -18488 37854 -18402
rect 37618 -18552 37704 -18488
rect 37704 -18552 37768 -18488
rect 37768 -18552 37854 -18488
rect 30522 -18698 30758 -18612
rect 30522 -18762 30608 -18698
rect 30608 -18762 30672 -18698
rect 30672 -18762 30758 -18698
rect 30522 -18848 30758 -18762
rect 30842 -18698 31078 -18612
rect 30842 -18762 30928 -18698
rect 30928 -18762 30992 -18698
rect 30992 -18762 31078 -18698
rect 30842 -18848 31078 -18762
rect 31162 -18698 31398 -18612
rect 31162 -18762 31248 -18698
rect 31248 -18762 31312 -18698
rect 31312 -18762 31398 -18698
rect 31162 -18848 31398 -18762
rect 31482 -18698 31718 -18612
rect 31482 -18762 31568 -18698
rect 31568 -18762 31632 -18698
rect 31632 -18762 31718 -18698
rect 31482 -18848 31718 -18762
rect 31802 -18698 32038 -18612
rect 31802 -18762 31888 -18698
rect 31888 -18762 31952 -18698
rect 31952 -18762 32038 -18698
rect 31802 -18848 32038 -18762
rect 32122 -18698 32358 -18612
rect 32122 -18762 32208 -18698
rect 32208 -18762 32272 -18698
rect 32272 -18762 32358 -18698
rect 32122 -18848 32358 -18762
rect 32442 -18698 32678 -18612
rect 32442 -18762 32528 -18698
rect 32528 -18762 32592 -18698
rect 32592 -18762 32678 -18698
rect 32442 -18848 32678 -18762
rect 32762 -18698 32998 -18612
rect 32762 -18762 32848 -18698
rect 32848 -18762 32912 -18698
rect 32912 -18762 32998 -18698
rect 32762 -18848 32998 -18762
rect 33082 -18698 33318 -18612
rect 33082 -18762 33168 -18698
rect 33168 -18762 33232 -18698
rect 33232 -18762 33318 -18698
rect 33082 -18848 33318 -18762
rect 33402 -18698 33638 -18612
rect 33402 -18762 33488 -18698
rect 33488 -18762 33552 -18698
rect 33552 -18762 33638 -18698
rect 33402 -18848 33638 -18762
rect 33722 -18698 33958 -18612
rect 33722 -18762 33808 -18698
rect 33808 -18762 33872 -18698
rect 33872 -18762 33958 -18698
rect 33722 -18848 33958 -18762
rect 34042 -18698 34278 -18612
rect 34042 -18762 34128 -18698
rect 34128 -18762 34192 -18698
rect 34192 -18762 34278 -18698
rect 34042 -18848 34278 -18762
rect 34362 -18698 34598 -18612
rect 34362 -18762 34448 -18698
rect 34448 -18762 34512 -18698
rect 34512 -18762 34598 -18698
rect 34362 -18848 34598 -18762
rect 34682 -18698 34918 -18612
rect 34682 -18762 34768 -18698
rect 34768 -18762 34832 -18698
rect 34832 -18762 34918 -18698
rect 34682 -18848 34918 -18762
rect 35002 -18698 35238 -18612
rect 35002 -18762 35088 -18698
rect 35088 -18762 35152 -18698
rect 35152 -18762 35238 -18698
rect 35002 -18848 35238 -18762
rect 35322 -18698 35558 -18612
rect 35322 -18762 35408 -18698
rect 35408 -18762 35472 -18698
rect 35472 -18762 35558 -18698
rect 35322 -18848 35558 -18762
rect 35642 -18698 35878 -18612
rect 35642 -18762 35728 -18698
rect 35728 -18762 35792 -18698
rect 35792 -18762 35878 -18698
rect 35642 -18848 35878 -18762
rect 35962 -18698 36198 -18612
rect 35962 -18762 36048 -18698
rect 36048 -18762 36112 -18698
rect 36112 -18762 36198 -18698
rect 35962 -18848 36198 -18762
rect 36282 -18698 36518 -18612
rect 36282 -18762 36368 -18698
rect 36368 -18762 36432 -18698
rect 36432 -18762 36518 -18698
rect 36282 -18848 36518 -18762
rect 36602 -18698 36838 -18612
rect 36602 -18762 36688 -18698
rect 36688 -18762 36752 -18698
rect 36752 -18762 36838 -18698
rect 36602 -18848 36838 -18762
rect 36922 -18698 37158 -18612
rect 36922 -18762 37008 -18698
rect 37008 -18762 37072 -18698
rect 37072 -18762 37158 -18698
rect 36922 -18848 37158 -18762
rect 37242 -18698 37478 -18612
rect 37618 -18638 37854 -18552
rect 37242 -18762 37328 -18698
rect 37328 -18762 37392 -18698
rect 37392 -18762 37478 -18698
rect 37242 -18848 37478 -18762
rect 42152 -11512 42238 -11448
rect 42238 -11512 42302 -11448
rect 42302 -11512 42388 -11448
rect 42152 -11598 42388 -11512
rect 49618 -11448 49854 -11362
rect 49618 -11512 49704 -11448
rect 49704 -11512 49768 -11448
rect 49768 -11512 49854 -11448
rect 42152 -11768 42388 -11682
rect 42152 -11832 42238 -11768
rect 42238 -11832 42302 -11768
rect 42302 -11832 42388 -11768
rect 42152 -11918 42388 -11832
rect 42152 -12088 42388 -12002
rect 42152 -12152 42238 -12088
rect 42238 -12152 42302 -12088
rect 42302 -12152 42388 -12088
rect 42152 -12238 42388 -12152
rect 42152 -12408 42388 -12322
rect 42152 -12472 42238 -12408
rect 42238 -12472 42302 -12408
rect 42302 -12472 42388 -12408
rect 42152 -12558 42388 -12472
rect 42152 -12728 42388 -12642
rect 42152 -12792 42238 -12728
rect 42238 -12792 42302 -12728
rect 42302 -12792 42388 -12728
rect 42152 -12878 42388 -12792
rect 42152 -13048 42388 -12962
rect 42152 -13112 42238 -13048
rect 42238 -13112 42302 -13048
rect 42302 -13112 42388 -13048
rect 42152 -13198 42388 -13112
rect 42152 -13368 42388 -13282
rect 42152 -13432 42238 -13368
rect 42238 -13432 42302 -13368
rect 42302 -13432 42388 -13368
rect 42152 -13518 42388 -13432
rect 42152 -13688 42388 -13602
rect 42152 -13752 42238 -13688
rect 42238 -13752 42302 -13688
rect 42302 -13752 42388 -13688
rect 42152 -13838 42388 -13752
rect 42152 -14008 42388 -13922
rect 42152 -14072 42238 -14008
rect 42238 -14072 42302 -14008
rect 42302 -14072 42388 -14008
rect 42152 -14158 42388 -14072
rect 42152 -14328 42388 -14242
rect 42152 -14392 42238 -14328
rect 42238 -14392 42302 -14328
rect 42302 -14392 42388 -14328
rect 42152 -14478 42388 -14392
rect 42152 -14648 42388 -14562
rect 42152 -14712 42238 -14648
rect 42238 -14712 42302 -14648
rect 42302 -14712 42388 -14648
rect 42152 -14798 42388 -14712
rect 42152 -14968 42388 -14882
rect 42152 -15032 42238 -14968
rect 42238 -15032 42302 -14968
rect 42302 -15032 42388 -14968
rect 42152 -15118 42388 -15032
rect 42152 -15288 42388 -15202
rect 42152 -15352 42238 -15288
rect 42238 -15352 42302 -15288
rect 42302 -15352 42388 -15288
rect 42152 -15438 42388 -15352
rect 42152 -15608 42388 -15522
rect 42152 -15672 42238 -15608
rect 42238 -15672 42302 -15608
rect 42302 -15672 42388 -15608
rect 42152 -15758 42388 -15672
rect 42152 -15928 42388 -15842
rect 42152 -15992 42238 -15928
rect 42238 -15992 42302 -15928
rect 42302 -15992 42388 -15928
rect 42152 -16078 42388 -15992
rect 42152 -16248 42388 -16162
rect 42152 -16312 42238 -16248
rect 42238 -16312 42302 -16248
rect 42302 -16312 42388 -16248
rect 42152 -16398 42388 -16312
rect 42152 -16568 42388 -16482
rect 42152 -16632 42238 -16568
rect 42238 -16632 42302 -16568
rect 42302 -16632 42388 -16568
rect 42152 -16718 42388 -16632
rect 42152 -16888 42388 -16802
rect 42152 -16952 42238 -16888
rect 42238 -16952 42302 -16888
rect 42302 -16952 42388 -16888
rect 42152 -17038 42388 -16952
rect 42152 -17208 42388 -17122
rect 42152 -17272 42238 -17208
rect 42238 -17272 42302 -17208
rect 42302 -17272 42388 -17208
rect 42152 -17358 42388 -17272
rect 42152 -17528 42388 -17442
rect 42152 -17592 42238 -17528
rect 42238 -17592 42302 -17528
rect 42302 -17592 42388 -17528
rect 42152 -17678 42388 -17592
rect 42152 -17848 42388 -17762
rect 42152 -17912 42238 -17848
rect 42238 -17912 42302 -17848
rect 42302 -17912 42388 -17848
rect 42152 -17998 42388 -17912
rect 42152 -18168 42388 -18082
rect 42152 -18232 42238 -18168
rect 42238 -18232 42302 -18168
rect 42302 -18232 42388 -18168
rect 42152 -18318 42388 -18232
rect 42152 -18488 42388 -18402
rect 49618 -11598 49854 -11512
rect 49618 -11768 49854 -11682
rect 49618 -11832 49704 -11768
rect 49704 -11832 49768 -11768
rect 49768 -11832 49854 -11768
rect 49618 -11918 49854 -11832
rect 49618 -12088 49854 -12002
rect 49618 -12152 49704 -12088
rect 49704 -12152 49768 -12088
rect 49768 -12152 49854 -12088
rect 49618 -12238 49854 -12152
rect 49618 -12408 49854 -12322
rect 49618 -12472 49704 -12408
rect 49704 -12472 49768 -12408
rect 49768 -12472 49854 -12408
rect 49618 -12558 49854 -12472
rect 49618 -12728 49854 -12642
rect 49618 -12792 49704 -12728
rect 49704 -12792 49768 -12728
rect 49768 -12792 49854 -12728
rect 49618 -12878 49854 -12792
rect 49618 -13048 49854 -12962
rect 49618 -13112 49704 -13048
rect 49704 -13112 49768 -13048
rect 49768 -13112 49854 -13048
rect 49618 -13198 49854 -13112
rect 49618 -13368 49854 -13282
rect 49618 -13432 49704 -13368
rect 49704 -13432 49768 -13368
rect 49768 -13432 49854 -13368
rect 49618 -13518 49854 -13432
rect 49618 -13688 49854 -13602
rect 49618 -13752 49704 -13688
rect 49704 -13752 49768 -13688
rect 49768 -13752 49854 -13688
rect 49618 -13838 49854 -13752
rect 49618 -14008 49854 -13922
rect 49618 -14072 49704 -14008
rect 49704 -14072 49768 -14008
rect 49768 -14072 49854 -14008
rect 49618 -14158 49854 -14072
rect 49618 -14328 49854 -14242
rect 49618 -14392 49704 -14328
rect 49704 -14392 49768 -14328
rect 49768 -14392 49854 -14328
rect 49618 -14478 49854 -14392
rect 49618 -14648 49854 -14562
rect 49618 -14712 49704 -14648
rect 49704 -14712 49768 -14648
rect 49768 -14712 49854 -14648
rect 49618 -14798 49854 -14712
rect 49618 -14968 49854 -14882
rect 49618 -15032 49704 -14968
rect 49704 -15032 49768 -14968
rect 49768 -15032 49854 -14968
rect 49618 -15118 49854 -15032
rect 49618 -15288 49854 -15202
rect 49618 -15352 49704 -15288
rect 49704 -15352 49768 -15288
rect 49768 -15352 49854 -15288
rect 49618 -15438 49854 -15352
rect 49618 -15608 49854 -15522
rect 49618 -15672 49704 -15608
rect 49704 -15672 49768 -15608
rect 49768 -15672 49854 -15608
rect 49618 -15758 49854 -15672
rect 49618 -15928 49854 -15842
rect 49618 -15992 49704 -15928
rect 49704 -15992 49768 -15928
rect 49768 -15992 49854 -15928
rect 49618 -16078 49854 -15992
rect 49618 -16248 49854 -16162
rect 49618 -16312 49704 -16248
rect 49704 -16312 49768 -16248
rect 49768 -16312 49854 -16248
rect 49618 -16398 49854 -16312
rect 49618 -16568 49854 -16482
rect 49618 -16632 49704 -16568
rect 49704 -16632 49768 -16568
rect 49768 -16632 49854 -16568
rect 49618 -16718 49854 -16632
rect 49618 -16888 49854 -16802
rect 49618 -16952 49704 -16888
rect 49704 -16952 49768 -16888
rect 49768 -16952 49854 -16888
rect 49618 -17038 49854 -16952
rect 49618 -17208 49854 -17122
rect 49618 -17272 49704 -17208
rect 49704 -17272 49768 -17208
rect 49768 -17272 49854 -17208
rect 49618 -17358 49854 -17272
rect 49618 -17528 49854 -17442
rect 49618 -17592 49704 -17528
rect 49704 -17592 49768 -17528
rect 49768 -17592 49854 -17528
rect 49618 -17678 49854 -17592
rect 49618 -17848 49854 -17762
rect 49618 -17912 49704 -17848
rect 49704 -17912 49768 -17848
rect 49768 -17912 49854 -17848
rect 49618 -17998 49854 -17912
rect 49618 -18168 49854 -18082
rect 49618 -18232 49704 -18168
rect 49704 -18232 49768 -18168
rect 49768 -18232 49854 -18168
rect 49618 -18318 49854 -18232
rect 42152 -18552 42238 -18488
rect 42238 -18552 42302 -18488
rect 42302 -18552 42388 -18488
rect 42152 -18638 42388 -18552
rect 49618 -18488 49854 -18402
rect 49618 -18552 49704 -18488
rect 49704 -18552 49768 -18488
rect 49768 -18552 49854 -18488
rect 42522 -18698 42758 -18612
rect 42522 -18762 42608 -18698
rect 42608 -18762 42672 -18698
rect 42672 -18762 42758 -18698
rect 42522 -18848 42758 -18762
rect 42842 -18698 43078 -18612
rect 42842 -18762 42928 -18698
rect 42928 -18762 42992 -18698
rect 42992 -18762 43078 -18698
rect 42842 -18848 43078 -18762
rect 43162 -18698 43398 -18612
rect 43162 -18762 43248 -18698
rect 43248 -18762 43312 -18698
rect 43312 -18762 43398 -18698
rect 43162 -18848 43398 -18762
rect 43482 -18698 43718 -18612
rect 43482 -18762 43568 -18698
rect 43568 -18762 43632 -18698
rect 43632 -18762 43718 -18698
rect 43482 -18848 43718 -18762
rect 43802 -18698 44038 -18612
rect 43802 -18762 43888 -18698
rect 43888 -18762 43952 -18698
rect 43952 -18762 44038 -18698
rect 43802 -18848 44038 -18762
rect 44122 -18698 44358 -18612
rect 44122 -18762 44208 -18698
rect 44208 -18762 44272 -18698
rect 44272 -18762 44358 -18698
rect 44122 -18848 44358 -18762
rect 44442 -18698 44678 -18612
rect 44442 -18762 44528 -18698
rect 44528 -18762 44592 -18698
rect 44592 -18762 44678 -18698
rect 44442 -18848 44678 -18762
rect 44762 -18698 44998 -18612
rect 44762 -18762 44848 -18698
rect 44848 -18762 44912 -18698
rect 44912 -18762 44998 -18698
rect 44762 -18848 44998 -18762
rect 45082 -18698 45318 -18612
rect 45082 -18762 45168 -18698
rect 45168 -18762 45232 -18698
rect 45232 -18762 45318 -18698
rect 45082 -18848 45318 -18762
rect 45402 -18698 45638 -18612
rect 45402 -18762 45488 -18698
rect 45488 -18762 45552 -18698
rect 45552 -18762 45638 -18698
rect 45402 -18848 45638 -18762
rect 45722 -18698 45958 -18612
rect 45722 -18762 45808 -18698
rect 45808 -18762 45872 -18698
rect 45872 -18762 45958 -18698
rect 45722 -18848 45958 -18762
rect 46042 -18698 46278 -18612
rect 46042 -18762 46128 -18698
rect 46128 -18762 46192 -18698
rect 46192 -18762 46278 -18698
rect 46042 -18848 46278 -18762
rect 46362 -18698 46598 -18612
rect 46362 -18762 46448 -18698
rect 46448 -18762 46512 -18698
rect 46512 -18762 46598 -18698
rect 46362 -18848 46598 -18762
rect 46682 -18698 46918 -18612
rect 46682 -18762 46768 -18698
rect 46768 -18762 46832 -18698
rect 46832 -18762 46918 -18698
rect 46682 -18848 46918 -18762
rect 47002 -18698 47238 -18612
rect 47002 -18762 47088 -18698
rect 47088 -18762 47152 -18698
rect 47152 -18762 47238 -18698
rect 47002 -18848 47238 -18762
rect 47322 -18698 47558 -18612
rect 47322 -18762 47408 -18698
rect 47408 -18762 47472 -18698
rect 47472 -18762 47558 -18698
rect 47322 -18848 47558 -18762
rect 47642 -18698 47878 -18612
rect 47642 -18762 47728 -18698
rect 47728 -18762 47792 -18698
rect 47792 -18762 47878 -18698
rect 47642 -18848 47878 -18762
rect 47962 -18698 48198 -18612
rect 47962 -18762 48048 -18698
rect 48048 -18762 48112 -18698
rect 48112 -18762 48198 -18698
rect 47962 -18848 48198 -18762
rect 48282 -18698 48518 -18612
rect 48282 -18762 48368 -18698
rect 48368 -18762 48432 -18698
rect 48432 -18762 48518 -18698
rect 48282 -18848 48518 -18762
rect 48602 -18698 48838 -18612
rect 48602 -18762 48688 -18698
rect 48688 -18762 48752 -18698
rect 48752 -18762 48838 -18698
rect 48602 -18848 48838 -18762
rect 48922 -18698 49158 -18612
rect 48922 -18762 49008 -18698
rect 49008 -18762 49072 -18698
rect 49072 -18762 49158 -18698
rect 48922 -18848 49158 -18762
rect 49242 -18698 49478 -18612
rect 49618 -18638 49854 -18552
rect 49242 -18762 49328 -18698
rect 49328 -18762 49392 -18698
rect 49392 -18762 49478 -18698
rect 49242 -18848 49478 -18762
rect 6522 -23242 6758 -23156
rect 6522 -23306 6608 -23242
rect 6608 -23306 6672 -23242
rect 6672 -23306 6758 -23242
rect 6152 -23448 6388 -23362
rect 6522 -23392 6758 -23306
rect 6842 -23242 7078 -23156
rect 6842 -23306 6928 -23242
rect 6928 -23306 6992 -23242
rect 6992 -23306 7078 -23242
rect 6842 -23392 7078 -23306
rect 7162 -23242 7398 -23156
rect 7162 -23306 7248 -23242
rect 7248 -23306 7312 -23242
rect 7312 -23306 7398 -23242
rect 7162 -23392 7398 -23306
rect 7482 -23242 7718 -23156
rect 7482 -23306 7568 -23242
rect 7568 -23306 7632 -23242
rect 7632 -23306 7718 -23242
rect 7482 -23392 7718 -23306
rect 7802 -23242 8038 -23156
rect 7802 -23306 7888 -23242
rect 7888 -23306 7952 -23242
rect 7952 -23306 8038 -23242
rect 7802 -23392 8038 -23306
rect 8122 -23242 8358 -23156
rect 8122 -23306 8208 -23242
rect 8208 -23306 8272 -23242
rect 8272 -23306 8358 -23242
rect 8122 -23392 8358 -23306
rect 8442 -23242 8678 -23156
rect 8442 -23306 8528 -23242
rect 8528 -23306 8592 -23242
rect 8592 -23306 8678 -23242
rect 8442 -23392 8678 -23306
rect 8762 -23242 8998 -23156
rect 8762 -23306 8848 -23242
rect 8848 -23306 8912 -23242
rect 8912 -23306 8998 -23242
rect 8762 -23392 8998 -23306
rect 9082 -23242 9318 -23156
rect 9082 -23306 9168 -23242
rect 9168 -23306 9232 -23242
rect 9232 -23306 9318 -23242
rect 9082 -23392 9318 -23306
rect 9402 -23242 9638 -23156
rect 9402 -23306 9488 -23242
rect 9488 -23306 9552 -23242
rect 9552 -23306 9638 -23242
rect 9402 -23392 9638 -23306
rect 9722 -23242 9958 -23156
rect 9722 -23306 9808 -23242
rect 9808 -23306 9872 -23242
rect 9872 -23306 9958 -23242
rect 9722 -23392 9958 -23306
rect 10042 -23242 10278 -23156
rect 10042 -23306 10128 -23242
rect 10128 -23306 10192 -23242
rect 10192 -23306 10278 -23242
rect 10042 -23392 10278 -23306
rect 10362 -23242 10598 -23156
rect 10362 -23306 10448 -23242
rect 10448 -23306 10512 -23242
rect 10512 -23306 10598 -23242
rect 10362 -23392 10598 -23306
rect 10682 -23242 10918 -23156
rect 10682 -23306 10768 -23242
rect 10768 -23306 10832 -23242
rect 10832 -23306 10918 -23242
rect 10682 -23392 10918 -23306
rect 11002 -23242 11238 -23156
rect 11002 -23306 11088 -23242
rect 11088 -23306 11152 -23242
rect 11152 -23306 11238 -23242
rect 11002 -23392 11238 -23306
rect 11322 -23242 11558 -23156
rect 11322 -23306 11408 -23242
rect 11408 -23306 11472 -23242
rect 11472 -23306 11558 -23242
rect 11322 -23392 11558 -23306
rect 11642 -23242 11878 -23156
rect 11642 -23306 11728 -23242
rect 11728 -23306 11792 -23242
rect 11792 -23306 11878 -23242
rect 11642 -23392 11878 -23306
rect 11962 -23242 12198 -23156
rect 11962 -23306 12048 -23242
rect 12048 -23306 12112 -23242
rect 12112 -23306 12198 -23242
rect 11962 -23392 12198 -23306
rect 12282 -23242 12518 -23156
rect 12282 -23306 12368 -23242
rect 12368 -23306 12432 -23242
rect 12432 -23306 12518 -23242
rect 12282 -23392 12518 -23306
rect 12602 -23242 12838 -23156
rect 12602 -23306 12688 -23242
rect 12688 -23306 12752 -23242
rect 12752 -23306 12838 -23242
rect 12602 -23392 12838 -23306
rect 12922 -23242 13158 -23156
rect 12922 -23306 13008 -23242
rect 13008 -23306 13072 -23242
rect 13072 -23306 13158 -23242
rect 12922 -23392 13158 -23306
rect 13242 -23242 13478 -23156
rect 13242 -23306 13328 -23242
rect 13328 -23306 13392 -23242
rect 13392 -23306 13478 -23242
rect 13242 -23392 13478 -23306
rect 6152 -23512 6238 -23448
rect 6238 -23512 6302 -23448
rect 6302 -23512 6388 -23448
rect 6152 -23598 6388 -23512
rect 13618 -23448 13854 -23362
rect 13618 -23512 13704 -23448
rect 13704 -23512 13768 -23448
rect 13768 -23512 13854 -23448
rect 6152 -23768 6388 -23682
rect 6152 -23832 6238 -23768
rect 6238 -23832 6302 -23768
rect 6302 -23832 6388 -23768
rect 6152 -23918 6388 -23832
rect 6152 -24088 6388 -24002
rect 6152 -24152 6238 -24088
rect 6238 -24152 6302 -24088
rect 6302 -24152 6388 -24088
rect 6152 -24238 6388 -24152
rect 6152 -24408 6388 -24322
rect 6152 -24472 6238 -24408
rect 6238 -24472 6302 -24408
rect 6302 -24472 6388 -24408
rect 6152 -24558 6388 -24472
rect 6152 -24728 6388 -24642
rect 6152 -24792 6238 -24728
rect 6238 -24792 6302 -24728
rect 6302 -24792 6388 -24728
rect 6152 -24878 6388 -24792
rect 6152 -25048 6388 -24962
rect 6152 -25112 6238 -25048
rect 6238 -25112 6302 -25048
rect 6302 -25112 6388 -25048
rect 6152 -25198 6388 -25112
rect 6152 -25368 6388 -25282
rect 6152 -25432 6238 -25368
rect 6238 -25432 6302 -25368
rect 6302 -25432 6388 -25368
rect 6152 -25518 6388 -25432
rect 6152 -25688 6388 -25602
rect 6152 -25752 6238 -25688
rect 6238 -25752 6302 -25688
rect 6302 -25752 6388 -25688
rect 6152 -25838 6388 -25752
rect 6152 -26008 6388 -25922
rect 6152 -26072 6238 -26008
rect 6238 -26072 6302 -26008
rect 6302 -26072 6388 -26008
rect 6152 -26158 6388 -26072
rect 6152 -26328 6388 -26242
rect 6152 -26392 6238 -26328
rect 6238 -26392 6302 -26328
rect 6302 -26392 6388 -26328
rect 6152 -26478 6388 -26392
rect 6152 -26648 6388 -26562
rect 6152 -26712 6238 -26648
rect 6238 -26712 6302 -26648
rect 6302 -26712 6388 -26648
rect 6152 -26798 6388 -26712
rect 6152 -26968 6388 -26882
rect 6152 -27032 6238 -26968
rect 6238 -27032 6302 -26968
rect 6302 -27032 6388 -26968
rect 6152 -27118 6388 -27032
rect 6152 -27288 6388 -27202
rect 6152 -27352 6238 -27288
rect 6238 -27352 6302 -27288
rect 6302 -27352 6388 -27288
rect 6152 -27438 6388 -27352
rect 6152 -27608 6388 -27522
rect 6152 -27672 6238 -27608
rect 6238 -27672 6302 -27608
rect 6302 -27672 6388 -27608
rect 6152 -27758 6388 -27672
rect 6152 -27928 6388 -27842
rect 6152 -27992 6238 -27928
rect 6238 -27992 6302 -27928
rect 6302 -27992 6388 -27928
rect 6152 -28078 6388 -27992
rect 6152 -28248 6388 -28162
rect 6152 -28312 6238 -28248
rect 6238 -28312 6302 -28248
rect 6302 -28312 6388 -28248
rect 6152 -28398 6388 -28312
rect 6152 -28568 6388 -28482
rect 6152 -28632 6238 -28568
rect 6238 -28632 6302 -28568
rect 6302 -28632 6388 -28568
rect 6152 -28718 6388 -28632
rect 6152 -28888 6388 -28802
rect 6152 -28952 6238 -28888
rect 6238 -28952 6302 -28888
rect 6302 -28952 6388 -28888
rect 6152 -29038 6388 -28952
rect 6152 -29208 6388 -29122
rect 6152 -29272 6238 -29208
rect 6238 -29272 6302 -29208
rect 6302 -29272 6388 -29208
rect 6152 -29358 6388 -29272
rect 6152 -29528 6388 -29442
rect 6152 -29592 6238 -29528
rect 6238 -29592 6302 -29528
rect 6302 -29592 6388 -29528
rect 6152 -29678 6388 -29592
rect 6152 -29848 6388 -29762
rect 6152 -29912 6238 -29848
rect 6238 -29912 6302 -29848
rect 6302 -29912 6388 -29848
rect 6152 -29998 6388 -29912
rect 6152 -30168 6388 -30082
rect 6152 -30232 6238 -30168
rect 6238 -30232 6302 -30168
rect 6302 -30232 6388 -30168
rect 6152 -30318 6388 -30232
rect 6152 -30488 6388 -30402
rect 13618 -23598 13854 -23512
rect 13618 -23768 13854 -23682
rect 13618 -23832 13704 -23768
rect 13704 -23832 13768 -23768
rect 13768 -23832 13854 -23768
rect 13618 -23918 13854 -23832
rect 13618 -24088 13854 -24002
rect 13618 -24152 13704 -24088
rect 13704 -24152 13768 -24088
rect 13768 -24152 13854 -24088
rect 13618 -24238 13854 -24152
rect 13618 -24408 13854 -24322
rect 13618 -24472 13704 -24408
rect 13704 -24472 13768 -24408
rect 13768 -24472 13854 -24408
rect 13618 -24558 13854 -24472
rect 13618 -24728 13854 -24642
rect 13618 -24792 13704 -24728
rect 13704 -24792 13768 -24728
rect 13768 -24792 13854 -24728
rect 13618 -24878 13854 -24792
rect 13618 -25048 13854 -24962
rect 13618 -25112 13704 -25048
rect 13704 -25112 13768 -25048
rect 13768 -25112 13854 -25048
rect 13618 -25198 13854 -25112
rect 13618 -25368 13854 -25282
rect 13618 -25432 13704 -25368
rect 13704 -25432 13768 -25368
rect 13768 -25432 13854 -25368
rect 13618 -25518 13854 -25432
rect 13618 -25688 13854 -25602
rect 13618 -25752 13704 -25688
rect 13704 -25752 13768 -25688
rect 13768 -25752 13854 -25688
rect 13618 -25838 13854 -25752
rect 13618 -26008 13854 -25922
rect 13618 -26072 13704 -26008
rect 13704 -26072 13768 -26008
rect 13768 -26072 13854 -26008
rect 13618 -26158 13854 -26072
rect 13618 -26328 13854 -26242
rect 13618 -26392 13704 -26328
rect 13704 -26392 13768 -26328
rect 13768 -26392 13854 -26328
rect 13618 -26478 13854 -26392
rect 13618 -26648 13854 -26562
rect 13618 -26712 13704 -26648
rect 13704 -26712 13768 -26648
rect 13768 -26712 13854 -26648
rect 13618 -26798 13854 -26712
rect 13618 -26968 13854 -26882
rect 13618 -27032 13704 -26968
rect 13704 -27032 13768 -26968
rect 13768 -27032 13854 -26968
rect 13618 -27118 13854 -27032
rect 13618 -27288 13854 -27202
rect 13618 -27352 13704 -27288
rect 13704 -27352 13768 -27288
rect 13768 -27352 13854 -27288
rect 13618 -27438 13854 -27352
rect 13618 -27608 13854 -27522
rect 13618 -27672 13704 -27608
rect 13704 -27672 13768 -27608
rect 13768 -27672 13854 -27608
rect 13618 -27758 13854 -27672
rect 13618 -27928 13854 -27842
rect 13618 -27992 13704 -27928
rect 13704 -27992 13768 -27928
rect 13768 -27992 13854 -27928
rect 13618 -28078 13854 -27992
rect 13618 -28248 13854 -28162
rect 13618 -28312 13704 -28248
rect 13704 -28312 13768 -28248
rect 13768 -28312 13854 -28248
rect 13618 -28398 13854 -28312
rect 13618 -28568 13854 -28482
rect 13618 -28632 13704 -28568
rect 13704 -28632 13768 -28568
rect 13768 -28632 13854 -28568
rect 13618 -28718 13854 -28632
rect 13618 -28888 13854 -28802
rect 13618 -28952 13704 -28888
rect 13704 -28952 13768 -28888
rect 13768 -28952 13854 -28888
rect 13618 -29038 13854 -28952
rect 13618 -29208 13854 -29122
rect 13618 -29272 13704 -29208
rect 13704 -29272 13768 -29208
rect 13768 -29272 13854 -29208
rect 13618 -29358 13854 -29272
rect 13618 -29528 13854 -29442
rect 13618 -29592 13704 -29528
rect 13704 -29592 13768 -29528
rect 13768 -29592 13854 -29528
rect 13618 -29678 13854 -29592
rect 13618 -29848 13854 -29762
rect 13618 -29912 13704 -29848
rect 13704 -29912 13768 -29848
rect 13768 -29912 13854 -29848
rect 13618 -29998 13854 -29912
rect 13618 -30168 13854 -30082
rect 13618 -30232 13704 -30168
rect 13704 -30232 13768 -30168
rect 13768 -30232 13854 -30168
rect 13618 -30318 13854 -30232
rect 6152 -30552 6238 -30488
rect 6238 -30552 6302 -30488
rect 6302 -30552 6388 -30488
rect 6152 -30638 6388 -30552
rect 13618 -30488 13854 -30402
rect 13618 -30552 13704 -30488
rect 13704 -30552 13768 -30488
rect 13768 -30552 13854 -30488
rect 6522 -30698 6758 -30612
rect 6522 -30762 6608 -30698
rect 6608 -30762 6672 -30698
rect 6672 -30762 6758 -30698
rect 6522 -30848 6758 -30762
rect 6842 -30698 7078 -30612
rect 6842 -30762 6928 -30698
rect 6928 -30762 6992 -30698
rect 6992 -30762 7078 -30698
rect 6842 -30848 7078 -30762
rect 7162 -30698 7398 -30612
rect 7162 -30762 7248 -30698
rect 7248 -30762 7312 -30698
rect 7312 -30762 7398 -30698
rect 7162 -30848 7398 -30762
rect 7482 -30698 7718 -30612
rect 7482 -30762 7568 -30698
rect 7568 -30762 7632 -30698
rect 7632 -30762 7718 -30698
rect 7482 -30848 7718 -30762
rect 7802 -30698 8038 -30612
rect 7802 -30762 7888 -30698
rect 7888 -30762 7952 -30698
rect 7952 -30762 8038 -30698
rect 7802 -30848 8038 -30762
rect 8122 -30698 8358 -30612
rect 8122 -30762 8208 -30698
rect 8208 -30762 8272 -30698
rect 8272 -30762 8358 -30698
rect 8122 -30848 8358 -30762
rect 8442 -30698 8678 -30612
rect 8442 -30762 8528 -30698
rect 8528 -30762 8592 -30698
rect 8592 -30762 8678 -30698
rect 8442 -30848 8678 -30762
rect 8762 -30698 8998 -30612
rect 8762 -30762 8848 -30698
rect 8848 -30762 8912 -30698
rect 8912 -30762 8998 -30698
rect 8762 -30848 8998 -30762
rect 9082 -30698 9318 -30612
rect 9082 -30762 9168 -30698
rect 9168 -30762 9232 -30698
rect 9232 -30762 9318 -30698
rect 9082 -30848 9318 -30762
rect 9402 -30698 9638 -30612
rect 9402 -30762 9488 -30698
rect 9488 -30762 9552 -30698
rect 9552 -30762 9638 -30698
rect 9402 -30848 9638 -30762
rect 9722 -30698 9958 -30612
rect 9722 -30762 9808 -30698
rect 9808 -30762 9872 -30698
rect 9872 -30762 9958 -30698
rect 9722 -30848 9958 -30762
rect 10042 -30698 10278 -30612
rect 10042 -30762 10128 -30698
rect 10128 -30762 10192 -30698
rect 10192 -30762 10278 -30698
rect 10042 -30848 10278 -30762
rect 10362 -30698 10598 -30612
rect 10362 -30762 10448 -30698
rect 10448 -30762 10512 -30698
rect 10512 -30762 10598 -30698
rect 10362 -30848 10598 -30762
rect 10682 -30698 10918 -30612
rect 10682 -30762 10768 -30698
rect 10768 -30762 10832 -30698
rect 10832 -30762 10918 -30698
rect 10682 -30848 10918 -30762
rect 11002 -30698 11238 -30612
rect 11002 -30762 11088 -30698
rect 11088 -30762 11152 -30698
rect 11152 -30762 11238 -30698
rect 11002 -30848 11238 -30762
rect 11322 -30698 11558 -30612
rect 11322 -30762 11408 -30698
rect 11408 -30762 11472 -30698
rect 11472 -30762 11558 -30698
rect 11322 -30848 11558 -30762
rect 11642 -30698 11878 -30612
rect 11642 -30762 11728 -30698
rect 11728 -30762 11792 -30698
rect 11792 -30762 11878 -30698
rect 11642 -30848 11878 -30762
rect 11962 -30698 12198 -30612
rect 11962 -30762 12048 -30698
rect 12048 -30762 12112 -30698
rect 12112 -30762 12198 -30698
rect 11962 -30848 12198 -30762
rect 12282 -30698 12518 -30612
rect 12282 -30762 12368 -30698
rect 12368 -30762 12432 -30698
rect 12432 -30762 12518 -30698
rect 12282 -30848 12518 -30762
rect 12602 -30698 12838 -30612
rect 12602 -30762 12688 -30698
rect 12688 -30762 12752 -30698
rect 12752 -30762 12838 -30698
rect 12602 -30848 12838 -30762
rect 12922 -30698 13158 -30612
rect 12922 -30762 13008 -30698
rect 13008 -30762 13072 -30698
rect 13072 -30762 13158 -30698
rect 12922 -30848 13158 -30762
rect 13242 -30698 13478 -30612
rect 13618 -30638 13854 -30552
rect 13242 -30762 13328 -30698
rect 13328 -30762 13392 -30698
rect 13392 -30762 13478 -30698
rect 13242 -30848 13478 -30762
rect 18522 -23242 18758 -23156
rect 18522 -23306 18608 -23242
rect 18608 -23306 18672 -23242
rect 18672 -23306 18758 -23242
rect 18152 -23448 18388 -23362
rect 18522 -23392 18758 -23306
rect 18842 -23242 19078 -23156
rect 18842 -23306 18928 -23242
rect 18928 -23306 18992 -23242
rect 18992 -23306 19078 -23242
rect 18842 -23392 19078 -23306
rect 19162 -23242 19398 -23156
rect 19162 -23306 19248 -23242
rect 19248 -23306 19312 -23242
rect 19312 -23306 19398 -23242
rect 19162 -23392 19398 -23306
rect 19482 -23242 19718 -23156
rect 19482 -23306 19568 -23242
rect 19568 -23306 19632 -23242
rect 19632 -23306 19718 -23242
rect 19482 -23392 19718 -23306
rect 19802 -23242 20038 -23156
rect 19802 -23306 19888 -23242
rect 19888 -23306 19952 -23242
rect 19952 -23306 20038 -23242
rect 19802 -23392 20038 -23306
rect 20122 -23242 20358 -23156
rect 20122 -23306 20208 -23242
rect 20208 -23306 20272 -23242
rect 20272 -23306 20358 -23242
rect 20122 -23392 20358 -23306
rect 20442 -23242 20678 -23156
rect 20442 -23306 20528 -23242
rect 20528 -23306 20592 -23242
rect 20592 -23306 20678 -23242
rect 20442 -23392 20678 -23306
rect 20762 -23242 20998 -23156
rect 20762 -23306 20848 -23242
rect 20848 -23306 20912 -23242
rect 20912 -23306 20998 -23242
rect 20762 -23392 20998 -23306
rect 21082 -23242 21318 -23156
rect 21082 -23306 21168 -23242
rect 21168 -23306 21232 -23242
rect 21232 -23306 21318 -23242
rect 21082 -23392 21318 -23306
rect 21402 -23242 21638 -23156
rect 21402 -23306 21488 -23242
rect 21488 -23306 21552 -23242
rect 21552 -23306 21638 -23242
rect 21402 -23392 21638 -23306
rect 21722 -23242 21958 -23156
rect 21722 -23306 21808 -23242
rect 21808 -23306 21872 -23242
rect 21872 -23306 21958 -23242
rect 21722 -23392 21958 -23306
rect 22042 -23242 22278 -23156
rect 22042 -23306 22128 -23242
rect 22128 -23306 22192 -23242
rect 22192 -23306 22278 -23242
rect 22042 -23392 22278 -23306
rect 22362 -23242 22598 -23156
rect 22362 -23306 22448 -23242
rect 22448 -23306 22512 -23242
rect 22512 -23306 22598 -23242
rect 22362 -23392 22598 -23306
rect 22682 -23242 22918 -23156
rect 22682 -23306 22768 -23242
rect 22768 -23306 22832 -23242
rect 22832 -23306 22918 -23242
rect 22682 -23392 22918 -23306
rect 23002 -23242 23238 -23156
rect 23002 -23306 23088 -23242
rect 23088 -23306 23152 -23242
rect 23152 -23306 23238 -23242
rect 23002 -23392 23238 -23306
rect 23322 -23242 23558 -23156
rect 23322 -23306 23408 -23242
rect 23408 -23306 23472 -23242
rect 23472 -23306 23558 -23242
rect 23322 -23392 23558 -23306
rect 23642 -23242 23878 -23156
rect 23642 -23306 23728 -23242
rect 23728 -23306 23792 -23242
rect 23792 -23306 23878 -23242
rect 23642 -23392 23878 -23306
rect 23962 -23242 24198 -23156
rect 23962 -23306 24048 -23242
rect 24048 -23306 24112 -23242
rect 24112 -23306 24198 -23242
rect 23962 -23392 24198 -23306
rect 24282 -23242 24518 -23156
rect 24282 -23306 24368 -23242
rect 24368 -23306 24432 -23242
rect 24432 -23306 24518 -23242
rect 24282 -23392 24518 -23306
rect 24602 -23242 24838 -23156
rect 24602 -23306 24688 -23242
rect 24688 -23306 24752 -23242
rect 24752 -23306 24838 -23242
rect 24602 -23392 24838 -23306
rect 24922 -23242 25158 -23156
rect 24922 -23306 25008 -23242
rect 25008 -23306 25072 -23242
rect 25072 -23306 25158 -23242
rect 24922 -23392 25158 -23306
rect 25242 -23242 25478 -23156
rect 25242 -23306 25328 -23242
rect 25328 -23306 25392 -23242
rect 25392 -23306 25478 -23242
rect 25242 -23392 25478 -23306
rect 18152 -23512 18238 -23448
rect 18238 -23512 18302 -23448
rect 18302 -23512 18388 -23448
rect 18152 -23598 18388 -23512
rect 25618 -23448 25854 -23362
rect 25618 -23512 25704 -23448
rect 25704 -23512 25768 -23448
rect 25768 -23512 25854 -23448
rect 18152 -23768 18388 -23682
rect 18152 -23832 18238 -23768
rect 18238 -23832 18302 -23768
rect 18302 -23832 18388 -23768
rect 18152 -23918 18388 -23832
rect 18152 -24088 18388 -24002
rect 18152 -24152 18238 -24088
rect 18238 -24152 18302 -24088
rect 18302 -24152 18388 -24088
rect 18152 -24238 18388 -24152
rect 18152 -24408 18388 -24322
rect 18152 -24472 18238 -24408
rect 18238 -24472 18302 -24408
rect 18302 -24472 18388 -24408
rect 18152 -24558 18388 -24472
rect 18152 -24728 18388 -24642
rect 18152 -24792 18238 -24728
rect 18238 -24792 18302 -24728
rect 18302 -24792 18388 -24728
rect 18152 -24878 18388 -24792
rect 18152 -25048 18388 -24962
rect 18152 -25112 18238 -25048
rect 18238 -25112 18302 -25048
rect 18302 -25112 18388 -25048
rect 18152 -25198 18388 -25112
rect 18152 -25368 18388 -25282
rect 18152 -25432 18238 -25368
rect 18238 -25432 18302 -25368
rect 18302 -25432 18388 -25368
rect 18152 -25518 18388 -25432
rect 18152 -25688 18388 -25602
rect 18152 -25752 18238 -25688
rect 18238 -25752 18302 -25688
rect 18302 -25752 18388 -25688
rect 18152 -25838 18388 -25752
rect 18152 -26008 18388 -25922
rect 18152 -26072 18238 -26008
rect 18238 -26072 18302 -26008
rect 18302 -26072 18388 -26008
rect 18152 -26158 18388 -26072
rect 18152 -26328 18388 -26242
rect 18152 -26392 18238 -26328
rect 18238 -26392 18302 -26328
rect 18302 -26392 18388 -26328
rect 18152 -26478 18388 -26392
rect 18152 -26648 18388 -26562
rect 18152 -26712 18238 -26648
rect 18238 -26712 18302 -26648
rect 18302 -26712 18388 -26648
rect 18152 -26798 18388 -26712
rect 18152 -26968 18388 -26882
rect 18152 -27032 18238 -26968
rect 18238 -27032 18302 -26968
rect 18302 -27032 18388 -26968
rect 18152 -27118 18388 -27032
rect 18152 -27288 18388 -27202
rect 18152 -27352 18238 -27288
rect 18238 -27352 18302 -27288
rect 18302 -27352 18388 -27288
rect 18152 -27438 18388 -27352
rect 18152 -27608 18388 -27522
rect 18152 -27672 18238 -27608
rect 18238 -27672 18302 -27608
rect 18302 -27672 18388 -27608
rect 18152 -27758 18388 -27672
rect 18152 -27928 18388 -27842
rect 18152 -27992 18238 -27928
rect 18238 -27992 18302 -27928
rect 18302 -27992 18388 -27928
rect 18152 -28078 18388 -27992
rect 18152 -28248 18388 -28162
rect 18152 -28312 18238 -28248
rect 18238 -28312 18302 -28248
rect 18302 -28312 18388 -28248
rect 18152 -28398 18388 -28312
rect 18152 -28568 18388 -28482
rect 18152 -28632 18238 -28568
rect 18238 -28632 18302 -28568
rect 18302 -28632 18388 -28568
rect 18152 -28718 18388 -28632
rect 18152 -28888 18388 -28802
rect 18152 -28952 18238 -28888
rect 18238 -28952 18302 -28888
rect 18302 -28952 18388 -28888
rect 18152 -29038 18388 -28952
rect 18152 -29208 18388 -29122
rect 18152 -29272 18238 -29208
rect 18238 -29272 18302 -29208
rect 18302 -29272 18388 -29208
rect 18152 -29358 18388 -29272
rect 18152 -29528 18388 -29442
rect 18152 -29592 18238 -29528
rect 18238 -29592 18302 -29528
rect 18302 -29592 18388 -29528
rect 18152 -29678 18388 -29592
rect 18152 -29848 18388 -29762
rect 18152 -29912 18238 -29848
rect 18238 -29912 18302 -29848
rect 18302 -29912 18388 -29848
rect 18152 -29998 18388 -29912
rect 18152 -30168 18388 -30082
rect 18152 -30232 18238 -30168
rect 18238 -30232 18302 -30168
rect 18302 -30232 18388 -30168
rect 18152 -30318 18388 -30232
rect 18152 -30488 18388 -30402
rect 25618 -23598 25854 -23512
rect 25618 -23768 25854 -23682
rect 25618 -23832 25704 -23768
rect 25704 -23832 25768 -23768
rect 25768 -23832 25854 -23768
rect 25618 -23918 25854 -23832
rect 25618 -24088 25854 -24002
rect 25618 -24152 25704 -24088
rect 25704 -24152 25768 -24088
rect 25768 -24152 25854 -24088
rect 25618 -24238 25854 -24152
rect 25618 -24408 25854 -24322
rect 25618 -24472 25704 -24408
rect 25704 -24472 25768 -24408
rect 25768 -24472 25854 -24408
rect 25618 -24558 25854 -24472
rect 25618 -24728 25854 -24642
rect 25618 -24792 25704 -24728
rect 25704 -24792 25768 -24728
rect 25768 -24792 25854 -24728
rect 25618 -24878 25854 -24792
rect 25618 -25048 25854 -24962
rect 25618 -25112 25704 -25048
rect 25704 -25112 25768 -25048
rect 25768 -25112 25854 -25048
rect 25618 -25198 25854 -25112
rect 25618 -25368 25854 -25282
rect 25618 -25432 25704 -25368
rect 25704 -25432 25768 -25368
rect 25768 -25432 25854 -25368
rect 25618 -25518 25854 -25432
rect 25618 -25688 25854 -25602
rect 25618 -25752 25704 -25688
rect 25704 -25752 25768 -25688
rect 25768 -25752 25854 -25688
rect 25618 -25838 25854 -25752
rect 25618 -26008 25854 -25922
rect 25618 -26072 25704 -26008
rect 25704 -26072 25768 -26008
rect 25768 -26072 25854 -26008
rect 25618 -26158 25854 -26072
rect 25618 -26328 25854 -26242
rect 25618 -26392 25704 -26328
rect 25704 -26392 25768 -26328
rect 25768 -26392 25854 -26328
rect 25618 -26478 25854 -26392
rect 25618 -26648 25854 -26562
rect 25618 -26712 25704 -26648
rect 25704 -26712 25768 -26648
rect 25768 -26712 25854 -26648
rect 25618 -26798 25854 -26712
rect 25618 -26968 25854 -26882
rect 25618 -27032 25704 -26968
rect 25704 -27032 25768 -26968
rect 25768 -27032 25854 -26968
rect 25618 -27118 25854 -27032
rect 25618 -27288 25854 -27202
rect 25618 -27352 25704 -27288
rect 25704 -27352 25768 -27288
rect 25768 -27352 25854 -27288
rect 25618 -27438 25854 -27352
rect 25618 -27608 25854 -27522
rect 25618 -27672 25704 -27608
rect 25704 -27672 25768 -27608
rect 25768 -27672 25854 -27608
rect 25618 -27758 25854 -27672
rect 25618 -27928 25854 -27842
rect 25618 -27992 25704 -27928
rect 25704 -27992 25768 -27928
rect 25768 -27992 25854 -27928
rect 25618 -28078 25854 -27992
rect 25618 -28248 25854 -28162
rect 25618 -28312 25704 -28248
rect 25704 -28312 25768 -28248
rect 25768 -28312 25854 -28248
rect 25618 -28398 25854 -28312
rect 25618 -28568 25854 -28482
rect 25618 -28632 25704 -28568
rect 25704 -28632 25768 -28568
rect 25768 -28632 25854 -28568
rect 25618 -28718 25854 -28632
rect 25618 -28888 25854 -28802
rect 25618 -28952 25704 -28888
rect 25704 -28952 25768 -28888
rect 25768 -28952 25854 -28888
rect 25618 -29038 25854 -28952
rect 25618 -29208 25854 -29122
rect 25618 -29272 25704 -29208
rect 25704 -29272 25768 -29208
rect 25768 -29272 25854 -29208
rect 25618 -29358 25854 -29272
rect 25618 -29528 25854 -29442
rect 25618 -29592 25704 -29528
rect 25704 -29592 25768 -29528
rect 25768 -29592 25854 -29528
rect 25618 -29678 25854 -29592
rect 25618 -29848 25854 -29762
rect 25618 -29912 25704 -29848
rect 25704 -29912 25768 -29848
rect 25768 -29912 25854 -29848
rect 25618 -29998 25854 -29912
rect 25618 -30168 25854 -30082
rect 25618 -30232 25704 -30168
rect 25704 -30232 25768 -30168
rect 25768 -30232 25854 -30168
rect 25618 -30318 25854 -30232
rect 18152 -30552 18238 -30488
rect 18238 -30552 18302 -30488
rect 18302 -30552 18388 -30488
rect 18152 -30638 18388 -30552
rect 25618 -30488 25854 -30402
rect 25618 -30552 25704 -30488
rect 25704 -30552 25768 -30488
rect 25768 -30552 25854 -30488
rect 18522 -30698 18758 -30612
rect 18522 -30762 18608 -30698
rect 18608 -30762 18672 -30698
rect 18672 -30762 18758 -30698
rect 18522 -30848 18758 -30762
rect 18842 -30698 19078 -30612
rect 18842 -30762 18928 -30698
rect 18928 -30762 18992 -30698
rect 18992 -30762 19078 -30698
rect 18842 -30848 19078 -30762
rect 19162 -30698 19398 -30612
rect 19162 -30762 19248 -30698
rect 19248 -30762 19312 -30698
rect 19312 -30762 19398 -30698
rect 19162 -30848 19398 -30762
rect 19482 -30698 19718 -30612
rect 19482 -30762 19568 -30698
rect 19568 -30762 19632 -30698
rect 19632 -30762 19718 -30698
rect 19482 -30848 19718 -30762
rect 19802 -30698 20038 -30612
rect 19802 -30762 19888 -30698
rect 19888 -30762 19952 -30698
rect 19952 -30762 20038 -30698
rect 19802 -30848 20038 -30762
rect 20122 -30698 20358 -30612
rect 20122 -30762 20208 -30698
rect 20208 -30762 20272 -30698
rect 20272 -30762 20358 -30698
rect 20122 -30848 20358 -30762
rect 20442 -30698 20678 -30612
rect 20442 -30762 20528 -30698
rect 20528 -30762 20592 -30698
rect 20592 -30762 20678 -30698
rect 20442 -30848 20678 -30762
rect 20762 -30698 20998 -30612
rect 20762 -30762 20848 -30698
rect 20848 -30762 20912 -30698
rect 20912 -30762 20998 -30698
rect 20762 -30848 20998 -30762
rect 21082 -30698 21318 -30612
rect 21082 -30762 21168 -30698
rect 21168 -30762 21232 -30698
rect 21232 -30762 21318 -30698
rect 21082 -30848 21318 -30762
rect 21402 -30698 21638 -30612
rect 21402 -30762 21488 -30698
rect 21488 -30762 21552 -30698
rect 21552 -30762 21638 -30698
rect 21402 -30848 21638 -30762
rect 21722 -30698 21958 -30612
rect 21722 -30762 21808 -30698
rect 21808 -30762 21872 -30698
rect 21872 -30762 21958 -30698
rect 21722 -30848 21958 -30762
rect 22042 -30698 22278 -30612
rect 22042 -30762 22128 -30698
rect 22128 -30762 22192 -30698
rect 22192 -30762 22278 -30698
rect 22042 -30848 22278 -30762
rect 22362 -30698 22598 -30612
rect 22362 -30762 22448 -30698
rect 22448 -30762 22512 -30698
rect 22512 -30762 22598 -30698
rect 22362 -30848 22598 -30762
rect 22682 -30698 22918 -30612
rect 22682 -30762 22768 -30698
rect 22768 -30762 22832 -30698
rect 22832 -30762 22918 -30698
rect 22682 -30848 22918 -30762
rect 23002 -30698 23238 -30612
rect 23002 -30762 23088 -30698
rect 23088 -30762 23152 -30698
rect 23152 -30762 23238 -30698
rect 23002 -30848 23238 -30762
rect 23322 -30698 23558 -30612
rect 23322 -30762 23408 -30698
rect 23408 -30762 23472 -30698
rect 23472 -30762 23558 -30698
rect 23322 -30848 23558 -30762
rect 23642 -30698 23878 -30612
rect 23642 -30762 23728 -30698
rect 23728 -30762 23792 -30698
rect 23792 -30762 23878 -30698
rect 23642 -30848 23878 -30762
rect 23962 -30698 24198 -30612
rect 23962 -30762 24048 -30698
rect 24048 -30762 24112 -30698
rect 24112 -30762 24198 -30698
rect 23962 -30848 24198 -30762
rect 24282 -30698 24518 -30612
rect 24282 -30762 24368 -30698
rect 24368 -30762 24432 -30698
rect 24432 -30762 24518 -30698
rect 24282 -30848 24518 -30762
rect 24602 -30698 24838 -30612
rect 24602 -30762 24688 -30698
rect 24688 -30762 24752 -30698
rect 24752 -30762 24838 -30698
rect 24602 -30848 24838 -30762
rect 24922 -30698 25158 -30612
rect 24922 -30762 25008 -30698
rect 25008 -30762 25072 -30698
rect 25072 -30762 25158 -30698
rect 24922 -30848 25158 -30762
rect 25242 -30698 25478 -30612
rect 25618 -30638 25854 -30552
rect 25242 -30762 25328 -30698
rect 25328 -30762 25392 -30698
rect 25392 -30762 25478 -30698
rect 25242 -30848 25478 -30762
rect 30522 -23242 30758 -23156
rect 30522 -23306 30608 -23242
rect 30608 -23306 30672 -23242
rect 30672 -23306 30758 -23242
rect 30152 -23448 30388 -23362
rect 30522 -23392 30758 -23306
rect 30842 -23242 31078 -23156
rect 30842 -23306 30928 -23242
rect 30928 -23306 30992 -23242
rect 30992 -23306 31078 -23242
rect 30842 -23392 31078 -23306
rect 31162 -23242 31398 -23156
rect 31162 -23306 31248 -23242
rect 31248 -23306 31312 -23242
rect 31312 -23306 31398 -23242
rect 31162 -23392 31398 -23306
rect 31482 -23242 31718 -23156
rect 31482 -23306 31568 -23242
rect 31568 -23306 31632 -23242
rect 31632 -23306 31718 -23242
rect 31482 -23392 31718 -23306
rect 31802 -23242 32038 -23156
rect 31802 -23306 31888 -23242
rect 31888 -23306 31952 -23242
rect 31952 -23306 32038 -23242
rect 31802 -23392 32038 -23306
rect 32122 -23242 32358 -23156
rect 32122 -23306 32208 -23242
rect 32208 -23306 32272 -23242
rect 32272 -23306 32358 -23242
rect 32122 -23392 32358 -23306
rect 32442 -23242 32678 -23156
rect 32442 -23306 32528 -23242
rect 32528 -23306 32592 -23242
rect 32592 -23306 32678 -23242
rect 32442 -23392 32678 -23306
rect 32762 -23242 32998 -23156
rect 32762 -23306 32848 -23242
rect 32848 -23306 32912 -23242
rect 32912 -23306 32998 -23242
rect 32762 -23392 32998 -23306
rect 33082 -23242 33318 -23156
rect 33082 -23306 33168 -23242
rect 33168 -23306 33232 -23242
rect 33232 -23306 33318 -23242
rect 33082 -23392 33318 -23306
rect 33402 -23242 33638 -23156
rect 33402 -23306 33488 -23242
rect 33488 -23306 33552 -23242
rect 33552 -23306 33638 -23242
rect 33402 -23392 33638 -23306
rect 33722 -23242 33958 -23156
rect 33722 -23306 33808 -23242
rect 33808 -23306 33872 -23242
rect 33872 -23306 33958 -23242
rect 33722 -23392 33958 -23306
rect 34042 -23242 34278 -23156
rect 34042 -23306 34128 -23242
rect 34128 -23306 34192 -23242
rect 34192 -23306 34278 -23242
rect 34042 -23392 34278 -23306
rect 34362 -23242 34598 -23156
rect 34362 -23306 34448 -23242
rect 34448 -23306 34512 -23242
rect 34512 -23306 34598 -23242
rect 34362 -23392 34598 -23306
rect 34682 -23242 34918 -23156
rect 34682 -23306 34768 -23242
rect 34768 -23306 34832 -23242
rect 34832 -23306 34918 -23242
rect 34682 -23392 34918 -23306
rect 35002 -23242 35238 -23156
rect 35002 -23306 35088 -23242
rect 35088 -23306 35152 -23242
rect 35152 -23306 35238 -23242
rect 35002 -23392 35238 -23306
rect 35322 -23242 35558 -23156
rect 35322 -23306 35408 -23242
rect 35408 -23306 35472 -23242
rect 35472 -23306 35558 -23242
rect 35322 -23392 35558 -23306
rect 35642 -23242 35878 -23156
rect 35642 -23306 35728 -23242
rect 35728 -23306 35792 -23242
rect 35792 -23306 35878 -23242
rect 35642 -23392 35878 -23306
rect 35962 -23242 36198 -23156
rect 35962 -23306 36048 -23242
rect 36048 -23306 36112 -23242
rect 36112 -23306 36198 -23242
rect 35962 -23392 36198 -23306
rect 36282 -23242 36518 -23156
rect 36282 -23306 36368 -23242
rect 36368 -23306 36432 -23242
rect 36432 -23306 36518 -23242
rect 36282 -23392 36518 -23306
rect 36602 -23242 36838 -23156
rect 36602 -23306 36688 -23242
rect 36688 -23306 36752 -23242
rect 36752 -23306 36838 -23242
rect 36602 -23392 36838 -23306
rect 36922 -23242 37158 -23156
rect 36922 -23306 37008 -23242
rect 37008 -23306 37072 -23242
rect 37072 -23306 37158 -23242
rect 36922 -23392 37158 -23306
rect 37242 -23242 37478 -23156
rect 37242 -23306 37328 -23242
rect 37328 -23306 37392 -23242
rect 37392 -23306 37478 -23242
rect 37242 -23392 37478 -23306
rect 30152 -23512 30238 -23448
rect 30238 -23512 30302 -23448
rect 30302 -23512 30388 -23448
rect 30152 -23598 30388 -23512
rect 37618 -23448 37854 -23362
rect 37618 -23512 37704 -23448
rect 37704 -23512 37768 -23448
rect 37768 -23512 37854 -23448
rect 30152 -23768 30388 -23682
rect 30152 -23832 30238 -23768
rect 30238 -23832 30302 -23768
rect 30302 -23832 30388 -23768
rect 30152 -23918 30388 -23832
rect 30152 -24088 30388 -24002
rect 30152 -24152 30238 -24088
rect 30238 -24152 30302 -24088
rect 30302 -24152 30388 -24088
rect 30152 -24238 30388 -24152
rect 30152 -24408 30388 -24322
rect 30152 -24472 30238 -24408
rect 30238 -24472 30302 -24408
rect 30302 -24472 30388 -24408
rect 30152 -24558 30388 -24472
rect 30152 -24728 30388 -24642
rect 30152 -24792 30238 -24728
rect 30238 -24792 30302 -24728
rect 30302 -24792 30388 -24728
rect 30152 -24878 30388 -24792
rect 30152 -25048 30388 -24962
rect 30152 -25112 30238 -25048
rect 30238 -25112 30302 -25048
rect 30302 -25112 30388 -25048
rect 30152 -25198 30388 -25112
rect 30152 -25368 30388 -25282
rect 30152 -25432 30238 -25368
rect 30238 -25432 30302 -25368
rect 30302 -25432 30388 -25368
rect 30152 -25518 30388 -25432
rect 30152 -25688 30388 -25602
rect 30152 -25752 30238 -25688
rect 30238 -25752 30302 -25688
rect 30302 -25752 30388 -25688
rect 30152 -25838 30388 -25752
rect 30152 -26008 30388 -25922
rect 30152 -26072 30238 -26008
rect 30238 -26072 30302 -26008
rect 30302 -26072 30388 -26008
rect 30152 -26158 30388 -26072
rect 30152 -26328 30388 -26242
rect 30152 -26392 30238 -26328
rect 30238 -26392 30302 -26328
rect 30302 -26392 30388 -26328
rect 30152 -26478 30388 -26392
rect 30152 -26648 30388 -26562
rect 30152 -26712 30238 -26648
rect 30238 -26712 30302 -26648
rect 30302 -26712 30388 -26648
rect 30152 -26798 30388 -26712
rect 30152 -26968 30388 -26882
rect 30152 -27032 30238 -26968
rect 30238 -27032 30302 -26968
rect 30302 -27032 30388 -26968
rect 30152 -27118 30388 -27032
rect 30152 -27288 30388 -27202
rect 30152 -27352 30238 -27288
rect 30238 -27352 30302 -27288
rect 30302 -27352 30388 -27288
rect 30152 -27438 30388 -27352
rect 30152 -27608 30388 -27522
rect 30152 -27672 30238 -27608
rect 30238 -27672 30302 -27608
rect 30302 -27672 30388 -27608
rect 30152 -27758 30388 -27672
rect 30152 -27928 30388 -27842
rect 30152 -27992 30238 -27928
rect 30238 -27992 30302 -27928
rect 30302 -27992 30388 -27928
rect 30152 -28078 30388 -27992
rect 30152 -28248 30388 -28162
rect 30152 -28312 30238 -28248
rect 30238 -28312 30302 -28248
rect 30302 -28312 30388 -28248
rect 30152 -28398 30388 -28312
rect 30152 -28568 30388 -28482
rect 30152 -28632 30238 -28568
rect 30238 -28632 30302 -28568
rect 30302 -28632 30388 -28568
rect 30152 -28718 30388 -28632
rect 30152 -28888 30388 -28802
rect 30152 -28952 30238 -28888
rect 30238 -28952 30302 -28888
rect 30302 -28952 30388 -28888
rect 30152 -29038 30388 -28952
rect 30152 -29208 30388 -29122
rect 30152 -29272 30238 -29208
rect 30238 -29272 30302 -29208
rect 30302 -29272 30388 -29208
rect 30152 -29358 30388 -29272
rect 30152 -29528 30388 -29442
rect 30152 -29592 30238 -29528
rect 30238 -29592 30302 -29528
rect 30302 -29592 30388 -29528
rect 30152 -29678 30388 -29592
rect 30152 -29848 30388 -29762
rect 30152 -29912 30238 -29848
rect 30238 -29912 30302 -29848
rect 30302 -29912 30388 -29848
rect 30152 -29998 30388 -29912
rect 30152 -30168 30388 -30082
rect 30152 -30232 30238 -30168
rect 30238 -30232 30302 -30168
rect 30302 -30232 30388 -30168
rect 30152 -30318 30388 -30232
rect 30152 -30488 30388 -30402
rect 37618 -23598 37854 -23512
rect 37618 -23768 37854 -23682
rect 37618 -23832 37704 -23768
rect 37704 -23832 37768 -23768
rect 37768 -23832 37854 -23768
rect 37618 -23918 37854 -23832
rect 37618 -24088 37854 -24002
rect 37618 -24152 37704 -24088
rect 37704 -24152 37768 -24088
rect 37768 -24152 37854 -24088
rect 37618 -24238 37854 -24152
rect 37618 -24408 37854 -24322
rect 37618 -24472 37704 -24408
rect 37704 -24472 37768 -24408
rect 37768 -24472 37854 -24408
rect 37618 -24558 37854 -24472
rect 37618 -24728 37854 -24642
rect 37618 -24792 37704 -24728
rect 37704 -24792 37768 -24728
rect 37768 -24792 37854 -24728
rect 37618 -24878 37854 -24792
rect 37618 -25048 37854 -24962
rect 37618 -25112 37704 -25048
rect 37704 -25112 37768 -25048
rect 37768 -25112 37854 -25048
rect 37618 -25198 37854 -25112
rect 37618 -25368 37854 -25282
rect 37618 -25432 37704 -25368
rect 37704 -25432 37768 -25368
rect 37768 -25432 37854 -25368
rect 37618 -25518 37854 -25432
rect 37618 -25688 37854 -25602
rect 37618 -25752 37704 -25688
rect 37704 -25752 37768 -25688
rect 37768 -25752 37854 -25688
rect 37618 -25838 37854 -25752
rect 37618 -26008 37854 -25922
rect 37618 -26072 37704 -26008
rect 37704 -26072 37768 -26008
rect 37768 -26072 37854 -26008
rect 37618 -26158 37854 -26072
rect 37618 -26328 37854 -26242
rect 37618 -26392 37704 -26328
rect 37704 -26392 37768 -26328
rect 37768 -26392 37854 -26328
rect 37618 -26478 37854 -26392
rect 37618 -26648 37854 -26562
rect 37618 -26712 37704 -26648
rect 37704 -26712 37768 -26648
rect 37768 -26712 37854 -26648
rect 37618 -26798 37854 -26712
rect 37618 -26968 37854 -26882
rect 37618 -27032 37704 -26968
rect 37704 -27032 37768 -26968
rect 37768 -27032 37854 -26968
rect 37618 -27118 37854 -27032
rect 37618 -27288 37854 -27202
rect 37618 -27352 37704 -27288
rect 37704 -27352 37768 -27288
rect 37768 -27352 37854 -27288
rect 37618 -27438 37854 -27352
rect 37618 -27608 37854 -27522
rect 37618 -27672 37704 -27608
rect 37704 -27672 37768 -27608
rect 37768 -27672 37854 -27608
rect 37618 -27758 37854 -27672
rect 37618 -27928 37854 -27842
rect 37618 -27992 37704 -27928
rect 37704 -27992 37768 -27928
rect 37768 -27992 37854 -27928
rect 37618 -28078 37854 -27992
rect 37618 -28248 37854 -28162
rect 37618 -28312 37704 -28248
rect 37704 -28312 37768 -28248
rect 37768 -28312 37854 -28248
rect 37618 -28398 37854 -28312
rect 37618 -28568 37854 -28482
rect 37618 -28632 37704 -28568
rect 37704 -28632 37768 -28568
rect 37768 -28632 37854 -28568
rect 37618 -28718 37854 -28632
rect 37618 -28888 37854 -28802
rect 37618 -28952 37704 -28888
rect 37704 -28952 37768 -28888
rect 37768 -28952 37854 -28888
rect 37618 -29038 37854 -28952
rect 37618 -29208 37854 -29122
rect 37618 -29272 37704 -29208
rect 37704 -29272 37768 -29208
rect 37768 -29272 37854 -29208
rect 37618 -29358 37854 -29272
rect 37618 -29528 37854 -29442
rect 37618 -29592 37704 -29528
rect 37704 -29592 37768 -29528
rect 37768 -29592 37854 -29528
rect 37618 -29678 37854 -29592
rect 37618 -29848 37854 -29762
rect 37618 -29912 37704 -29848
rect 37704 -29912 37768 -29848
rect 37768 -29912 37854 -29848
rect 37618 -29998 37854 -29912
rect 37618 -30168 37854 -30082
rect 37618 -30232 37704 -30168
rect 37704 -30232 37768 -30168
rect 37768 -30232 37854 -30168
rect 37618 -30318 37854 -30232
rect 30152 -30552 30238 -30488
rect 30238 -30552 30302 -30488
rect 30302 -30552 30388 -30488
rect 30152 -30638 30388 -30552
rect 37618 -30488 37854 -30402
rect 37618 -30552 37704 -30488
rect 37704 -30552 37768 -30488
rect 37768 -30552 37854 -30488
rect 30522 -30698 30758 -30612
rect 30522 -30762 30608 -30698
rect 30608 -30762 30672 -30698
rect 30672 -30762 30758 -30698
rect 30522 -30848 30758 -30762
rect 30842 -30698 31078 -30612
rect 30842 -30762 30928 -30698
rect 30928 -30762 30992 -30698
rect 30992 -30762 31078 -30698
rect 30842 -30848 31078 -30762
rect 31162 -30698 31398 -30612
rect 31162 -30762 31248 -30698
rect 31248 -30762 31312 -30698
rect 31312 -30762 31398 -30698
rect 31162 -30848 31398 -30762
rect 31482 -30698 31718 -30612
rect 31482 -30762 31568 -30698
rect 31568 -30762 31632 -30698
rect 31632 -30762 31718 -30698
rect 31482 -30848 31718 -30762
rect 31802 -30698 32038 -30612
rect 31802 -30762 31888 -30698
rect 31888 -30762 31952 -30698
rect 31952 -30762 32038 -30698
rect 31802 -30848 32038 -30762
rect 32122 -30698 32358 -30612
rect 32122 -30762 32208 -30698
rect 32208 -30762 32272 -30698
rect 32272 -30762 32358 -30698
rect 32122 -30848 32358 -30762
rect 32442 -30698 32678 -30612
rect 32442 -30762 32528 -30698
rect 32528 -30762 32592 -30698
rect 32592 -30762 32678 -30698
rect 32442 -30848 32678 -30762
rect 32762 -30698 32998 -30612
rect 32762 -30762 32848 -30698
rect 32848 -30762 32912 -30698
rect 32912 -30762 32998 -30698
rect 32762 -30848 32998 -30762
rect 33082 -30698 33318 -30612
rect 33082 -30762 33168 -30698
rect 33168 -30762 33232 -30698
rect 33232 -30762 33318 -30698
rect 33082 -30848 33318 -30762
rect 33402 -30698 33638 -30612
rect 33402 -30762 33488 -30698
rect 33488 -30762 33552 -30698
rect 33552 -30762 33638 -30698
rect 33402 -30848 33638 -30762
rect 33722 -30698 33958 -30612
rect 33722 -30762 33808 -30698
rect 33808 -30762 33872 -30698
rect 33872 -30762 33958 -30698
rect 33722 -30848 33958 -30762
rect 34042 -30698 34278 -30612
rect 34042 -30762 34128 -30698
rect 34128 -30762 34192 -30698
rect 34192 -30762 34278 -30698
rect 34042 -30848 34278 -30762
rect 34362 -30698 34598 -30612
rect 34362 -30762 34448 -30698
rect 34448 -30762 34512 -30698
rect 34512 -30762 34598 -30698
rect 34362 -30848 34598 -30762
rect 34682 -30698 34918 -30612
rect 34682 -30762 34768 -30698
rect 34768 -30762 34832 -30698
rect 34832 -30762 34918 -30698
rect 34682 -30848 34918 -30762
rect 35002 -30698 35238 -30612
rect 35002 -30762 35088 -30698
rect 35088 -30762 35152 -30698
rect 35152 -30762 35238 -30698
rect 35002 -30848 35238 -30762
rect 35322 -30698 35558 -30612
rect 35322 -30762 35408 -30698
rect 35408 -30762 35472 -30698
rect 35472 -30762 35558 -30698
rect 35322 -30848 35558 -30762
rect 35642 -30698 35878 -30612
rect 35642 -30762 35728 -30698
rect 35728 -30762 35792 -30698
rect 35792 -30762 35878 -30698
rect 35642 -30848 35878 -30762
rect 35962 -30698 36198 -30612
rect 35962 -30762 36048 -30698
rect 36048 -30762 36112 -30698
rect 36112 -30762 36198 -30698
rect 35962 -30848 36198 -30762
rect 36282 -30698 36518 -30612
rect 36282 -30762 36368 -30698
rect 36368 -30762 36432 -30698
rect 36432 -30762 36518 -30698
rect 36282 -30848 36518 -30762
rect 36602 -30698 36838 -30612
rect 36602 -30762 36688 -30698
rect 36688 -30762 36752 -30698
rect 36752 -30762 36838 -30698
rect 36602 -30848 36838 -30762
rect 36922 -30698 37158 -30612
rect 36922 -30762 37008 -30698
rect 37008 -30762 37072 -30698
rect 37072 -30762 37158 -30698
rect 36922 -30848 37158 -30762
rect 37242 -30698 37478 -30612
rect 37618 -30638 37854 -30552
rect 37242 -30762 37328 -30698
rect 37328 -30762 37392 -30698
rect 37392 -30762 37478 -30698
rect 37242 -30848 37478 -30762
rect 42522 -23242 42758 -23156
rect 42522 -23306 42608 -23242
rect 42608 -23306 42672 -23242
rect 42672 -23306 42758 -23242
rect 42152 -23448 42388 -23362
rect 42522 -23392 42758 -23306
rect 42842 -23242 43078 -23156
rect 42842 -23306 42928 -23242
rect 42928 -23306 42992 -23242
rect 42992 -23306 43078 -23242
rect 42842 -23392 43078 -23306
rect 43162 -23242 43398 -23156
rect 43162 -23306 43248 -23242
rect 43248 -23306 43312 -23242
rect 43312 -23306 43398 -23242
rect 43162 -23392 43398 -23306
rect 43482 -23242 43718 -23156
rect 43482 -23306 43568 -23242
rect 43568 -23306 43632 -23242
rect 43632 -23306 43718 -23242
rect 43482 -23392 43718 -23306
rect 43802 -23242 44038 -23156
rect 43802 -23306 43888 -23242
rect 43888 -23306 43952 -23242
rect 43952 -23306 44038 -23242
rect 43802 -23392 44038 -23306
rect 44122 -23242 44358 -23156
rect 44122 -23306 44208 -23242
rect 44208 -23306 44272 -23242
rect 44272 -23306 44358 -23242
rect 44122 -23392 44358 -23306
rect 44442 -23242 44678 -23156
rect 44442 -23306 44528 -23242
rect 44528 -23306 44592 -23242
rect 44592 -23306 44678 -23242
rect 44442 -23392 44678 -23306
rect 44762 -23242 44998 -23156
rect 44762 -23306 44848 -23242
rect 44848 -23306 44912 -23242
rect 44912 -23306 44998 -23242
rect 44762 -23392 44998 -23306
rect 45082 -23242 45318 -23156
rect 45082 -23306 45168 -23242
rect 45168 -23306 45232 -23242
rect 45232 -23306 45318 -23242
rect 45082 -23392 45318 -23306
rect 45402 -23242 45638 -23156
rect 45402 -23306 45488 -23242
rect 45488 -23306 45552 -23242
rect 45552 -23306 45638 -23242
rect 45402 -23392 45638 -23306
rect 45722 -23242 45958 -23156
rect 45722 -23306 45808 -23242
rect 45808 -23306 45872 -23242
rect 45872 -23306 45958 -23242
rect 45722 -23392 45958 -23306
rect 46042 -23242 46278 -23156
rect 46042 -23306 46128 -23242
rect 46128 -23306 46192 -23242
rect 46192 -23306 46278 -23242
rect 46042 -23392 46278 -23306
rect 46362 -23242 46598 -23156
rect 46362 -23306 46448 -23242
rect 46448 -23306 46512 -23242
rect 46512 -23306 46598 -23242
rect 46362 -23392 46598 -23306
rect 46682 -23242 46918 -23156
rect 46682 -23306 46768 -23242
rect 46768 -23306 46832 -23242
rect 46832 -23306 46918 -23242
rect 46682 -23392 46918 -23306
rect 47002 -23242 47238 -23156
rect 47002 -23306 47088 -23242
rect 47088 -23306 47152 -23242
rect 47152 -23306 47238 -23242
rect 47002 -23392 47238 -23306
rect 47322 -23242 47558 -23156
rect 47322 -23306 47408 -23242
rect 47408 -23306 47472 -23242
rect 47472 -23306 47558 -23242
rect 47322 -23392 47558 -23306
rect 47642 -23242 47878 -23156
rect 47642 -23306 47728 -23242
rect 47728 -23306 47792 -23242
rect 47792 -23306 47878 -23242
rect 47642 -23392 47878 -23306
rect 47962 -23242 48198 -23156
rect 47962 -23306 48048 -23242
rect 48048 -23306 48112 -23242
rect 48112 -23306 48198 -23242
rect 47962 -23392 48198 -23306
rect 48282 -23242 48518 -23156
rect 48282 -23306 48368 -23242
rect 48368 -23306 48432 -23242
rect 48432 -23306 48518 -23242
rect 48282 -23392 48518 -23306
rect 48602 -23242 48838 -23156
rect 48602 -23306 48688 -23242
rect 48688 -23306 48752 -23242
rect 48752 -23306 48838 -23242
rect 48602 -23392 48838 -23306
rect 48922 -23242 49158 -23156
rect 48922 -23306 49008 -23242
rect 49008 -23306 49072 -23242
rect 49072 -23306 49158 -23242
rect 48922 -23392 49158 -23306
rect 49242 -23242 49478 -23156
rect 49242 -23306 49328 -23242
rect 49328 -23306 49392 -23242
rect 49392 -23306 49478 -23242
rect 49242 -23392 49478 -23306
rect 42152 -23512 42238 -23448
rect 42238 -23512 42302 -23448
rect 42302 -23512 42388 -23448
rect 42152 -23598 42388 -23512
rect 49618 -23448 49854 -23362
rect 49618 -23512 49704 -23448
rect 49704 -23512 49768 -23448
rect 49768 -23512 49854 -23448
rect 42152 -23768 42388 -23682
rect 42152 -23832 42238 -23768
rect 42238 -23832 42302 -23768
rect 42302 -23832 42388 -23768
rect 42152 -23918 42388 -23832
rect 42152 -24088 42388 -24002
rect 42152 -24152 42238 -24088
rect 42238 -24152 42302 -24088
rect 42302 -24152 42388 -24088
rect 42152 -24238 42388 -24152
rect 42152 -24408 42388 -24322
rect 42152 -24472 42238 -24408
rect 42238 -24472 42302 -24408
rect 42302 -24472 42388 -24408
rect 42152 -24558 42388 -24472
rect 42152 -24728 42388 -24642
rect 42152 -24792 42238 -24728
rect 42238 -24792 42302 -24728
rect 42302 -24792 42388 -24728
rect 42152 -24878 42388 -24792
rect 42152 -25048 42388 -24962
rect 42152 -25112 42238 -25048
rect 42238 -25112 42302 -25048
rect 42302 -25112 42388 -25048
rect 42152 -25198 42388 -25112
rect 42152 -25368 42388 -25282
rect 42152 -25432 42238 -25368
rect 42238 -25432 42302 -25368
rect 42302 -25432 42388 -25368
rect 42152 -25518 42388 -25432
rect 42152 -25688 42388 -25602
rect 42152 -25752 42238 -25688
rect 42238 -25752 42302 -25688
rect 42302 -25752 42388 -25688
rect 42152 -25838 42388 -25752
rect 42152 -26008 42388 -25922
rect 42152 -26072 42238 -26008
rect 42238 -26072 42302 -26008
rect 42302 -26072 42388 -26008
rect 42152 -26158 42388 -26072
rect 42152 -26328 42388 -26242
rect 42152 -26392 42238 -26328
rect 42238 -26392 42302 -26328
rect 42302 -26392 42388 -26328
rect 42152 -26478 42388 -26392
rect 42152 -26648 42388 -26562
rect 42152 -26712 42238 -26648
rect 42238 -26712 42302 -26648
rect 42302 -26712 42388 -26648
rect 42152 -26798 42388 -26712
rect 42152 -26968 42388 -26882
rect 42152 -27032 42238 -26968
rect 42238 -27032 42302 -26968
rect 42302 -27032 42388 -26968
rect 42152 -27118 42388 -27032
rect 42152 -27288 42388 -27202
rect 42152 -27352 42238 -27288
rect 42238 -27352 42302 -27288
rect 42302 -27352 42388 -27288
rect 42152 -27438 42388 -27352
rect 42152 -27608 42388 -27522
rect 42152 -27672 42238 -27608
rect 42238 -27672 42302 -27608
rect 42302 -27672 42388 -27608
rect 42152 -27758 42388 -27672
rect 42152 -27928 42388 -27842
rect 42152 -27992 42238 -27928
rect 42238 -27992 42302 -27928
rect 42302 -27992 42388 -27928
rect 42152 -28078 42388 -27992
rect 42152 -28248 42388 -28162
rect 42152 -28312 42238 -28248
rect 42238 -28312 42302 -28248
rect 42302 -28312 42388 -28248
rect 42152 -28398 42388 -28312
rect 42152 -28568 42388 -28482
rect 42152 -28632 42238 -28568
rect 42238 -28632 42302 -28568
rect 42302 -28632 42388 -28568
rect 42152 -28718 42388 -28632
rect 42152 -28888 42388 -28802
rect 42152 -28952 42238 -28888
rect 42238 -28952 42302 -28888
rect 42302 -28952 42388 -28888
rect 42152 -29038 42388 -28952
rect 42152 -29208 42388 -29122
rect 42152 -29272 42238 -29208
rect 42238 -29272 42302 -29208
rect 42302 -29272 42388 -29208
rect 42152 -29358 42388 -29272
rect 42152 -29528 42388 -29442
rect 42152 -29592 42238 -29528
rect 42238 -29592 42302 -29528
rect 42302 -29592 42388 -29528
rect 42152 -29678 42388 -29592
rect 42152 -29848 42388 -29762
rect 42152 -29912 42238 -29848
rect 42238 -29912 42302 -29848
rect 42302 -29912 42388 -29848
rect 42152 -29998 42388 -29912
rect 42152 -30168 42388 -30082
rect 42152 -30232 42238 -30168
rect 42238 -30232 42302 -30168
rect 42302 -30232 42388 -30168
rect 42152 -30318 42388 -30232
rect 42152 -30488 42388 -30402
rect 49618 -23598 49854 -23512
rect 49618 -23768 49854 -23682
rect 49618 -23832 49704 -23768
rect 49704 -23832 49768 -23768
rect 49768 -23832 49854 -23768
rect 49618 -23918 49854 -23832
rect 49618 -24088 49854 -24002
rect 49618 -24152 49704 -24088
rect 49704 -24152 49768 -24088
rect 49768 -24152 49854 -24088
rect 49618 -24238 49854 -24152
rect 49618 -24408 49854 -24322
rect 49618 -24472 49704 -24408
rect 49704 -24472 49768 -24408
rect 49768 -24472 49854 -24408
rect 49618 -24558 49854 -24472
rect 49618 -24728 49854 -24642
rect 49618 -24792 49704 -24728
rect 49704 -24792 49768 -24728
rect 49768 -24792 49854 -24728
rect 49618 -24878 49854 -24792
rect 49618 -25048 49854 -24962
rect 49618 -25112 49704 -25048
rect 49704 -25112 49768 -25048
rect 49768 -25112 49854 -25048
rect 49618 -25198 49854 -25112
rect 49618 -25368 49854 -25282
rect 49618 -25432 49704 -25368
rect 49704 -25432 49768 -25368
rect 49768 -25432 49854 -25368
rect 49618 -25518 49854 -25432
rect 49618 -25688 49854 -25602
rect 49618 -25752 49704 -25688
rect 49704 -25752 49768 -25688
rect 49768 -25752 49854 -25688
rect 49618 -25838 49854 -25752
rect 49618 -26008 49854 -25922
rect 49618 -26072 49704 -26008
rect 49704 -26072 49768 -26008
rect 49768 -26072 49854 -26008
rect 49618 -26158 49854 -26072
rect 49618 -26328 49854 -26242
rect 49618 -26392 49704 -26328
rect 49704 -26392 49768 -26328
rect 49768 -26392 49854 -26328
rect 49618 -26478 49854 -26392
rect 49618 -26648 49854 -26562
rect 49618 -26712 49704 -26648
rect 49704 -26712 49768 -26648
rect 49768 -26712 49854 -26648
rect 49618 -26798 49854 -26712
rect 49618 -26968 49854 -26882
rect 49618 -27032 49704 -26968
rect 49704 -27032 49768 -26968
rect 49768 -27032 49854 -26968
rect 49618 -27118 49854 -27032
rect 49618 -27288 49854 -27202
rect 49618 -27352 49704 -27288
rect 49704 -27352 49768 -27288
rect 49768 -27352 49854 -27288
rect 49618 -27438 49854 -27352
rect 49618 -27608 49854 -27522
rect 49618 -27672 49704 -27608
rect 49704 -27672 49768 -27608
rect 49768 -27672 49854 -27608
rect 49618 -27758 49854 -27672
rect 49618 -27928 49854 -27842
rect 49618 -27992 49704 -27928
rect 49704 -27992 49768 -27928
rect 49768 -27992 49854 -27928
rect 49618 -28078 49854 -27992
rect 49618 -28248 49854 -28162
rect 49618 -28312 49704 -28248
rect 49704 -28312 49768 -28248
rect 49768 -28312 49854 -28248
rect 49618 -28398 49854 -28312
rect 49618 -28568 49854 -28482
rect 49618 -28632 49704 -28568
rect 49704 -28632 49768 -28568
rect 49768 -28632 49854 -28568
rect 49618 -28718 49854 -28632
rect 49618 -28888 49854 -28802
rect 49618 -28952 49704 -28888
rect 49704 -28952 49768 -28888
rect 49768 -28952 49854 -28888
rect 49618 -29038 49854 -28952
rect 49618 -29208 49854 -29122
rect 49618 -29272 49704 -29208
rect 49704 -29272 49768 -29208
rect 49768 -29272 49854 -29208
rect 49618 -29358 49854 -29272
rect 49618 -29528 49854 -29442
rect 49618 -29592 49704 -29528
rect 49704 -29592 49768 -29528
rect 49768 -29592 49854 -29528
rect 49618 -29678 49854 -29592
rect 49618 -29848 49854 -29762
rect 49618 -29912 49704 -29848
rect 49704 -29912 49768 -29848
rect 49768 -29912 49854 -29848
rect 49618 -29998 49854 -29912
rect 49618 -30168 49854 -30082
rect 49618 -30232 49704 -30168
rect 49704 -30232 49768 -30168
rect 49768 -30232 49854 -30168
rect 49618 -30318 49854 -30232
rect 42152 -30552 42238 -30488
rect 42238 -30552 42302 -30488
rect 42302 -30552 42388 -30488
rect 42152 -30638 42388 -30552
rect 49618 -30488 49854 -30402
rect 49618 -30552 49704 -30488
rect 49704 -30552 49768 -30488
rect 49768 -30552 49854 -30488
rect 42522 -30698 42758 -30612
rect 42522 -30762 42608 -30698
rect 42608 -30762 42672 -30698
rect 42672 -30762 42758 -30698
rect 42522 -30848 42758 -30762
rect 42842 -30698 43078 -30612
rect 42842 -30762 42928 -30698
rect 42928 -30762 42992 -30698
rect 42992 -30762 43078 -30698
rect 42842 -30848 43078 -30762
rect 43162 -30698 43398 -30612
rect 43162 -30762 43248 -30698
rect 43248 -30762 43312 -30698
rect 43312 -30762 43398 -30698
rect 43162 -30848 43398 -30762
rect 43482 -30698 43718 -30612
rect 43482 -30762 43568 -30698
rect 43568 -30762 43632 -30698
rect 43632 -30762 43718 -30698
rect 43482 -30848 43718 -30762
rect 43802 -30698 44038 -30612
rect 43802 -30762 43888 -30698
rect 43888 -30762 43952 -30698
rect 43952 -30762 44038 -30698
rect 43802 -30848 44038 -30762
rect 44122 -30698 44358 -30612
rect 44122 -30762 44208 -30698
rect 44208 -30762 44272 -30698
rect 44272 -30762 44358 -30698
rect 44122 -30848 44358 -30762
rect 44442 -30698 44678 -30612
rect 44442 -30762 44528 -30698
rect 44528 -30762 44592 -30698
rect 44592 -30762 44678 -30698
rect 44442 -30848 44678 -30762
rect 44762 -30698 44998 -30612
rect 44762 -30762 44848 -30698
rect 44848 -30762 44912 -30698
rect 44912 -30762 44998 -30698
rect 44762 -30848 44998 -30762
rect 45082 -30698 45318 -30612
rect 45082 -30762 45168 -30698
rect 45168 -30762 45232 -30698
rect 45232 -30762 45318 -30698
rect 45082 -30848 45318 -30762
rect 45402 -30698 45638 -30612
rect 45402 -30762 45488 -30698
rect 45488 -30762 45552 -30698
rect 45552 -30762 45638 -30698
rect 45402 -30848 45638 -30762
rect 45722 -30698 45958 -30612
rect 45722 -30762 45808 -30698
rect 45808 -30762 45872 -30698
rect 45872 -30762 45958 -30698
rect 45722 -30848 45958 -30762
rect 46042 -30698 46278 -30612
rect 46042 -30762 46128 -30698
rect 46128 -30762 46192 -30698
rect 46192 -30762 46278 -30698
rect 46042 -30848 46278 -30762
rect 46362 -30698 46598 -30612
rect 46362 -30762 46448 -30698
rect 46448 -30762 46512 -30698
rect 46512 -30762 46598 -30698
rect 46362 -30848 46598 -30762
rect 46682 -30698 46918 -30612
rect 46682 -30762 46768 -30698
rect 46768 -30762 46832 -30698
rect 46832 -30762 46918 -30698
rect 46682 -30848 46918 -30762
rect 47002 -30698 47238 -30612
rect 47002 -30762 47088 -30698
rect 47088 -30762 47152 -30698
rect 47152 -30762 47238 -30698
rect 47002 -30848 47238 -30762
rect 47322 -30698 47558 -30612
rect 47322 -30762 47408 -30698
rect 47408 -30762 47472 -30698
rect 47472 -30762 47558 -30698
rect 47322 -30848 47558 -30762
rect 47642 -30698 47878 -30612
rect 47642 -30762 47728 -30698
rect 47728 -30762 47792 -30698
rect 47792 -30762 47878 -30698
rect 47642 -30848 47878 -30762
rect 47962 -30698 48198 -30612
rect 47962 -30762 48048 -30698
rect 48048 -30762 48112 -30698
rect 48112 -30762 48198 -30698
rect 47962 -30848 48198 -30762
rect 48282 -30698 48518 -30612
rect 48282 -30762 48368 -30698
rect 48368 -30762 48432 -30698
rect 48432 -30762 48518 -30698
rect 48282 -30848 48518 -30762
rect 48602 -30698 48838 -30612
rect 48602 -30762 48688 -30698
rect 48688 -30762 48752 -30698
rect 48752 -30762 48838 -30698
rect 48602 -30848 48838 -30762
rect 48922 -30698 49158 -30612
rect 48922 -30762 49008 -30698
rect 49008 -30762 49072 -30698
rect 49072 -30762 49158 -30698
rect 48922 -30848 49158 -30762
rect 49242 -30698 49478 -30612
rect 49618 -30638 49854 -30552
rect 49242 -30762 49328 -30698
rect 49328 -30762 49392 -30698
rect 49392 -30762 49478 -30698
rect 49242 -30848 49478 -30762
<< mimcap2 >>
rect 16500 -2788 17600 -2748
rect 13300 -2840 15900 -2800
rect 13300 -8960 13340 -2840
rect 15860 -8960 15900 -2840
rect 16500 -8108 16540 -2788
rect 17560 -8108 17600 -2788
rect 22232 -2950 22972 -2930
rect 22232 -5550 22252 -2950
rect 22952 -5550 22972 -2950
rect 22232 -5570 22972 -5550
rect 16500 -8148 17600 -8108
rect 13300 -9000 15900 -8960
<< mimcap2contact >>
rect 13340 -8960 15860 -2840
rect 16540 -8108 17560 -2788
rect 22252 -5550 22952 -2950
<< metal5 >>
rect 13200 -2840 16000 -2700
rect 13200 -8960 13340 -2840
rect 15860 -8960 16000 -2840
rect 13200 -9600 16000 -8960
rect 16400 -2788 17700 -2648
rect 16400 -8108 16540 -2788
rect 17560 -8108 17700 -2788
rect 22202 -2950 23002 -2900
rect 22202 -5550 22252 -2950
rect 22952 -5550 23002 -2950
rect 22202 -5600 23002 -5550
rect 22402 -5720 23002 -5600
rect 22402 -5960 22432 -5720
rect 22972 -5960 23002 -5720
rect 22402 -5990 23002 -5960
rect 16400 -8248 17700 -8108
rect 16400 -8748 17300 -8248
rect 16400 -9148 16500 -8748
rect 17200 -9148 17300 -8748
rect 16400 -9248 17300 -9148
rect 13200 -10200 13300 -9600
rect 15900 -10200 16000 -9600
rect 13200 -10300 16000 -10200
rect 6000 -11156 14000 -11000
rect 6000 -11362 6522 -11156
rect 6000 -11598 6152 -11362
rect 6388 -11392 6522 -11362
rect 6758 -11392 6842 -11156
rect 7078 -11392 7162 -11156
rect 7398 -11392 7482 -11156
rect 7718 -11392 7802 -11156
rect 8038 -11392 8122 -11156
rect 8358 -11392 8442 -11156
rect 8678 -11392 8762 -11156
rect 8998 -11392 9082 -11156
rect 9318 -11392 9402 -11156
rect 9638 -11392 9722 -11156
rect 9958 -11392 10042 -11156
rect 10278 -11392 10362 -11156
rect 10598 -11392 10682 -11156
rect 10918 -11392 11002 -11156
rect 11238 -11392 11322 -11156
rect 11558 -11392 11642 -11156
rect 11878 -11392 11962 -11156
rect 12198 -11392 12282 -11156
rect 12518 -11392 12602 -11156
rect 12838 -11392 12922 -11156
rect 13158 -11392 13242 -11156
rect 13478 -11362 14000 -11156
rect 13478 -11392 13618 -11362
rect 6388 -11598 13618 -11392
rect 13854 -11598 14000 -11362
rect 6000 -11682 14000 -11598
rect 6000 -11918 6152 -11682
rect 6388 -11918 13618 -11682
rect 13854 -11918 14000 -11682
rect 6000 -12002 14000 -11918
rect 6000 -12238 6152 -12002
rect 6388 -12238 13618 -12002
rect 13854 -12238 14000 -12002
rect 6000 -12322 14000 -12238
rect 6000 -12558 6152 -12322
rect 6388 -12558 13618 -12322
rect 13854 -12558 14000 -12322
rect 6000 -12642 14000 -12558
rect 6000 -12878 6152 -12642
rect 6388 -12878 13618 -12642
rect 13854 -12878 14000 -12642
rect 6000 -12962 14000 -12878
rect 6000 -13198 6152 -12962
rect 6388 -13198 13618 -12962
rect 13854 -13198 14000 -12962
rect 6000 -13282 14000 -13198
rect 6000 -13518 6152 -13282
rect 6388 -13518 13618 -13282
rect 13854 -13518 14000 -13282
rect 6000 -13602 14000 -13518
rect 6000 -13838 6152 -13602
rect 6388 -13838 13618 -13602
rect 13854 -13838 14000 -13602
rect 6000 -13922 14000 -13838
rect 6000 -14158 6152 -13922
rect 6388 -14158 13618 -13922
rect 13854 -14158 14000 -13922
rect 6000 -14242 14000 -14158
rect 6000 -14478 6152 -14242
rect 6388 -14478 13618 -14242
rect 13854 -14478 14000 -14242
rect 6000 -14562 14000 -14478
rect 6000 -14798 6152 -14562
rect 6388 -14798 13618 -14562
rect 13854 -14798 14000 -14562
rect 6000 -14882 14000 -14798
rect 6000 -15118 6152 -14882
rect 6388 -15118 13618 -14882
rect 13854 -15118 14000 -14882
rect 6000 -15202 14000 -15118
rect 6000 -15438 6152 -15202
rect 6388 -15438 13618 -15202
rect 13854 -15438 14000 -15202
rect 6000 -15522 14000 -15438
rect 6000 -15758 6152 -15522
rect 6388 -15758 13618 -15522
rect 13854 -15758 14000 -15522
rect 6000 -15842 14000 -15758
rect 6000 -16078 6152 -15842
rect 6388 -16078 13618 -15842
rect 13854 -16078 14000 -15842
rect 6000 -16162 14000 -16078
rect 6000 -16398 6152 -16162
rect 6388 -16398 13618 -16162
rect 13854 -16398 14000 -16162
rect 6000 -16482 14000 -16398
rect 6000 -16718 6152 -16482
rect 6388 -16718 13618 -16482
rect 13854 -16718 14000 -16482
rect 6000 -16802 14000 -16718
rect 6000 -17038 6152 -16802
rect 6388 -17038 13618 -16802
rect 13854 -17038 14000 -16802
rect 6000 -17122 14000 -17038
rect 6000 -17358 6152 -17122
rect 6388 -17358 13618 -17122
rect 13854 -17358 14000 -17122
rect 6000 -17442 14000 -17358
rect 6000 -17678 6152 -17442
rect 6388 -17678 13618 -17442
rect 13854 -17678 14000 -17442
rect 6000 -17762 14000 -17678
rect 6000 -17998 6152 -17762
rect 6388 -17998 13618 -17762
rect 13854 -17998 14000 -17762
rect 6000 -18082 14000 -17998
rect 6000 -18318 6152 -18082
rect 6388 -18318 13618 -18082
rect 13854 -18318 14000 -18082
rect 6000 -18402 14000 -18318
rect 6000 -18638 6152 -18402
rect 6388 -18612 13618 -18402
rect 6388 -18638 6522 -18612
rect 6000 -18848 6522 -18638
rect 6758 -18848 6842 -18612
rect 7078 -18848 7162 -18612
rect 7398 -18848 7482 -18612
rect 7718 -18848 7802 -18612
rect 8038 -18848 8122 -18612
rect 8358 -18848 8442 -18612
rect 8678 -18848 8762 -18612
rect 8998 -18848 9082 -18612
rect 9318 -18848 9402 -18612
rect 9638 -18848 9722 -18612
rect 9958 -18848 10042 -18612
rect 10278 -18848 10362 -18612
rect 10598 -18848 10682 -18612
rect 10918 -18848 11002 -18612
rect 11238 -18848 11322 -18612
rect 11558 -18848 11642 -18612
rect 11878 -18848 11962 -18612
rect 12198 -18848 12282 -18612
rect 12518 -18848 12602 -18612
rect 12838 -18848 12922 -18612
rect 13158 -18848 13242 -18612
rect 13478 -18638 13618 -18612
rect 13854 -18638 14000 -18402
rect 13478 -18848 14000 -18638
rect 6000 -19000 14000 -18848
rect 18000 -11156 26000 -11000
rect 18000 -11362 18522 -11156
rect 18000 -11598 18152 -11362
rect 18388 -11392 18522 -11362
rect 18758 -11392 18842 -11156
rect 19078 -11392 19162 -11156
rect 19398 -11392 19482 -11156
rect 19718 -11392 19802 -11156
rect 20038 -11392 20122 -11156
rect 20358 -11392 20442 -11156
rect 20678 -11392 20762 -11156
rect 20998 -11392 21082 -11156
rect 21318 -11392 21402 -11156
rect 21638 -11392 21722 -11156
rect 21958 -11392 22042 -11156
rect 22278 -11392 22362 -11156
rect 22598 -11392 22682 -11156
rect 22918 -11392 23002 -11156
rect 23238 -11392 23322 -11156
rect 23558 -11392 23642 -11156
rect 23878 -11392 23962 -11156
rect 24198 -11392 24282 -11156
rect 24518 -11392 24602 -11156
rect 24838 -11392 24922 -11156
rect 25158 -11392 25242 -11156
rect 25478 -11362 26000 -11156
rect 25478 -11392 25618 -11362
rect 18388 -11598 25618 -11392
rect 25854 -11598 26000 -11362
rect 18000 -11682 26000 -11598
rect 18000 -11918 18152 -11682
rect 18388 -11918 25618 -11682
rect 25854 -11918 26000 -11682
rect 18000 -12002 26000 -11918
rect 18000 -12238 18152 -12002
rect 18388 -12238 25618 -12002
rect 25854 -12238 26000 -12002
rect 18000 -12322 26000 -12238
rect 18000 -12558 18152 -12322
rect 18388 -12558 25618 -12322
rect 25854 -12558 26000 -12322
rect 18000 -12642 26000 -12558
rect 18000 -12878 18152 -12642
rect 18388 -12878 25618 -12642
rect 25854 -12878 26000 -12642
rect 18000 -12962 26000 -12878
rect 18000 -13198 18152 -12962
rect 18388 -13198 25618 -12962
rect 25854 -13198 26000 -12962
rect 18000 -13282 26000 -13198
rect 18000 -13518 18152 -13282
rect 18388 -13518 25618 -13282
rect 25854 -13518 26000 -13282
rect 18000 -13602 26000 -13518
rect 18000 -13838 18152 -13602
rect 18388 -13838 25618 -13602
rect 25854 -13838 26000 -13602
rect 18000 -13922 26000 -13838
rect 18000 -14158 18152 -13922
rect 18388 -14158 25618 -13922
rect 25854 -14158 26000 -13922
rect 18000 -14242 26000 -14158
rect 18000 -14478 18152 -14242
rect 18388 -14478 25618 -14242
rect 25854 -14478 26000 -14242
rect 18000 -14562 26000 -14478
rect 18000 -14798 18152 -14562
rect 18388 -14798 25618 -14562
rect 25854 -14798 26000 -14562
rect 18000 -14882 26000 -14798
rect 18000 -15118 18152 -14882
rect 18388 -15118 25618 -14882
rect 25854 -15118 26000 -14882
rect 18000 -15202 26000 -15118
rect 18000 -15438 18152 -15202
rect 18388 -15438 25618 -15202
rect 25854 -15438 26000 -15202
rect 18000 -15522 26000 -15438
rect 18000 -15758 18152 -15522
rect 18388 -15758 25618 -15522
rect 25854 -15758 26000 -15522
rect 18000 -15842 26000 -15758
rect 18000 -16078 18152 -15842
rect 18388 -16078 25618 -15842
rect 25854 -16078 26000 -15842
rect 18000 -16162 26000 -16078
rect 18000 -16398 18152 -16162
rect 18388 -16398 25618 -16162
rect 25854 -16398 26000 -16162
rect 18000 -16482 26000 -16398
rect 18000 -16718 18152 -16482
rect 18388 -16718 25618 -16482
rect 25854 -16718 26000 -16482
rect 18000 -16802 26000 -16718
rect 18000 -17038 18152 -16802
rect 18388 -17038 25618 -16802
rect 25854 -17038 26000 -16802
rect 18000 -17122 26000 -17038
rect 18000 -17358 18152 -17122
rect 18388 -17358 25618 -17122
rect 25854 -17358 26000 -17122
rect 18000 -17442 26000 -17358
rect 18000 -17678 18152 -17442
rect 18388 -17678 25618 -17442
rect 25854 -17678 26000 -17442
rect 18000 -17762 26000 -17678
rect 18000 -17998 18152 -17762
rect 18388 -17998 25618 -17762
rect 25854 -17998 26000 -17762
rect 18000 -18082 26000 -17998
rect 18000 -18318 18152 -18082
rect 18388 -18318 25618 -18082
rect 25854 -18318 26000 -18082
rect 18000 -18402 26000 -18318
rect 18000 -18638 18152 -18402
rect 18388 -18612 25618 -18402
rect 18388 -18638 18522 -18612
rect 18000 -18848 18522 -18638
rect 18758 -18848 18842 -18612
rect 19078 -18848 19162 -18612
rect 19398 -18848 19482 -18612
rect 19718 -18848 19802 -18612
rect 20038 -18848 20122 -18612
rect 20358 -18848 20442 -18612
rect 20678 -18848 20762 -18612
rect 20998 -18848 21082 -18612
rect 21318 -18848 21402 -18612
rect 21638 -18848 21722 -18612
rect 21958 -18848 22042 -18612
rect 22278 -18848 22362 -18612
rect 22598 -18848 22682 -18612
rect 22918 -18848 23002 -18612
rect 23238 -18848 23322 -18612
rect 23558 -18848 23642 -18612
rect 23878 -18848 23962 -18612
rect 24198 -18848 24282 -18612
rect 24518 -18848 24602 -18612
rect 24838 -18848 24922 -18612
rect 25158 -18848 25242 -18612
rect 25478 -18638 25618 -18612
rect 25854 -18638 26000 -18402
rect 25478 -18848 26000 -18638
rect 18000 -19000 26000 -18848
rect 30000 -11156 38000 -11000
rect 30000 -11362 30522 -11156
rect 30000 -11598 30152 -11362
rect 30388 -11392 30522 -11362
rect 30758 -11392 30842 -11156
rect 31078 -11392 31162 -11156
rect 31398 -11392 31482 -11156
rect 31718 -11392 31802 -11156
rect 32038 -11392 32122 -11156
rect 32358 -11392 32442 -11156
rect 32678 -11392 32762 -11156
rect 32998 -11392 33082 -11156
rect 33318 -11392 33402 -11156
rect 33638 -11392 33722 -11156
rect 33958 -11392 34042 -11156
rect 34278 -11392 34362 -11156
rect 34598 -11392 34682 -11156
rect 34918 -11392 35002 -11156
rect 35238 -11392 35322 -11156
rect 35558 -11392 35642 -11156
rect 35878 -11392 35962 -11156
rect 36198 -11392 36282 -11156
rect 36518 -11392 36602 -11156
rect 36838 -11392 36922 -11156
rect 37158 -11392 37242 -11156
rect 37478 -11362 38000 -11156
rect 37478 -11392 37618 -11362
rect 30388 -11598 37618 -11392
rect 37854 -11598 38000 -11362
rect 30000 -11682 38000 -11598
rect 30000 -11918 30152 -11682
rect 30388 -11918 37618 -11682
rect 37854 -11918 38000 -11682
rect 30000 -12002 38000 -11918
rect 30000 -12238 30152 -12002
rect 30388 -12238 37618 -12002
rect 37854 -12238 38000 -12002
rect 30000 -12322 38000 -12238
rect 30000 -12558 30152 -12322
rect 30388 -12558 37618 -12322
rect 37854 -12558 38000 -12322
rect 30000 -12642 38000 -12558
rect 30000 -12878 30152 -12642
rect 30388 -12878 37618 -12642
rect 37854 -12878 38000 -12642
rect 30000 -12962 38000 -12878
rect 30000 -13198 30152 -12962
rect 30388 -13198 37618 -12962
rect 37854 -13198 38000 -12962
rect 30000 -13282 38000 -13198
rect 30000 -13518 30152 -13282
rect 30388 -13518 37618 -13282
rect 37854 -13518 38000 -13282
rect 30000 -13602 38000 -13518
rect 30000 -13838 30152 -13602
rect 30388 -13838 37618 -13602
rect 37854 -13838 38000 -13602
rect 30000 -13922 38000 -13838
rect 30000 -14158 30152 -13922
rect 30388 -14158 37618 -13922
rect 37854 -14158 38000 -13922
rect 30000 -14242 38000 -14158
rect 30000 -14478 30152 -14242
rect 30388 -14478 37618 -14242
rect 37854 -14478 38000 -14242
rect 30000 -14562 38000 -14478
rect 30000 -14798 30152 -14562
rect 30388 -14798 37618 -14562
rect 37854 -14798 38000 -14562
rect 30000 -14882 38000 -14798
rect 30000 -15118 30152 -14882
rect 30388 -15118 37618 -14882
rect 37854 -15118 38000 -14882
rect 30000 -15202 38000 -15118
rect 30000 -15438 30152 -15202
rect 30388 -15438 37618 -15202
rect 37854 -15438 38000 -15202
rect 30000 -15522 38000 -15438
rect 30000 -15758 30152 -15522
rect 30388 -15758 37618 -15522
rect 37854 -15758 38000 -15522
rect 30000 -15842 38000 -15758
rect 30000 -16078 30152 -15842
rect 30388 -16078 37618 -15842
rect 37854 -16078 38000 -15842
rect 30000 -16162 38000 -16078
rect 30000 -16398 30152 -16162
rect 30388 -16398 37618 -16162
rect 37854 -16398 38000 -16162
rect 30000 -16482 38000 -16398
rect 30000 -16718 30152 -16482
rect 30388 -16718 37618 -16482
rect 37854 -16718 38000 -16482
rect 30000 -16802 38000 -16718
rect 30000 -17038 30152 -16802
rect 30388 -17038 37618 -16802
rect 37854 -17038 38000 -16802
rect 30000 -17122 38000 -17038
rect 30000 -17358 30152 -17122
rect 30388 -17358 37618 -17122
rect 37854 -17358 38000 -17122
rect 30000 -17442 38000 -17358
rect 30000 -17678 30152 -17442
rect 30388 -17678 37618 -17442
rect 37854 -17678 38000 -17442
rect 30000 -17762 38000 -17678
rect 30000 -17998 30152 -17762
rect 30388 -17998 37618 -17762
rect 37854 -17998 38000 -17762
rect 30000 -18082 38000 -17998
rect 30000 -18318 30152 -18082
rect 30388 -18318 37618 -18082
rect 37854 -18318 38000 -18082
rect 30000 -18402 38000 -18318
rect 30000 -18638 30152 -18402
rect 30388 -18612 37618 -18402
rect 30388 -18638 30522 -18612
rect 30000 -18848 30522 -18638
rect 30758 -18848 30842 -18612
rect 31078 -18848 31162 -18612
rect 31398 -18848 31482 -18612
rect 31718 -18848 31802 -18612
rect 32038 -18848 32122 -18612
rect 32358 -18848 32442 -18612
rect 32678 -18848 32762 -18612
rect 32998 -18848 33082 -18612
rect 33318 -18848 33402 -18612
rect 33638 -18848 33722 -18612
rect 33958 -18848 34042 -18612
rect 34278 -18848 34362 -18612
rect 34598 -18848 34682 -18612
rect 34918 -18848 35002 -18612
rect 35238 -18848 35322 -18612
rect 35558 -18848 35642 -18612
rect 35878 -18848 35962 -18612
rect 36198 -18848 36282 -18612
rect 36518 -18848 36602 -18612
rect 36838 -18848 36922 -18612
rect 37158 -18848 37242 -18612
rect 37478 -18638 37618 -18612
rect 37854 -18638 38000 -18402
rect 37478 -18848 38000 -18638
rect 30000 -19000 38000 -18848
rect 42000 -11156 50000 -11000
rect 42000 -11362 42522 -11156
rect 42000 -11598 42152 -11362
rect 42388 -11392 42522 -11362
rect 42758 -11392 42842 -11156
rect 43078 -11392 43162 -11156
rect 43398 -11392 43482 -11156
rect 43718 -11392 43802 -11156
rect 44038 -11392 44122 -11156
rect 44358 -11392 44442 -11156
rect 44678 -11392 44762 -11156
rect 44998 -11392 45082 -11156
rect 45318 -11392 45402 -11156
rect 45638 -11392 45722 -11156
rect 45958 -11392 46042 -11156
rect 46278 -11392 46362 -11156
rect 46598 -11392 46682 -11156
rect 46918 -11392 47002 -11156
rect 47238 -11392 47322 -11156
rect 47558 -11392 47642 -11156
rect 47878 -11392 47962 -11156
rect 48198 -11392 48282 -11156
rect 48518 -11392 48602 -11156
rect 48838 -11392 48922 -11156
rect 49158 -11392 49242 -11156
rect 49478 -11362 50000 -11156
rect 49478 -11392 49618 -11362
rect 42388 -11598 49618 -11392
rect 49854 -11598 50000 -11362
rect 42000 -11682 50000 -11598
rect 42000 -11918 42152 -11682
rect 42388 -11918 49618 -11682
rect 49854 -11918 50000 -11682
rect 42000 -12002 50000 -11918
rect 42000 -12238 42152 -12002
rect 42388 -12238 49618 -12002
rect 49854 -12238 50000 -12002
rect 42000 -12322 50000 -12238
rect 42000 -12558 42152 -12322
rect 42388 -12558 49618 -12322
rect 49854 -12558 50000 -12322
rect 42000 -12642 50000 -12558
rect 42000 -12878 42152 -12642
rect 42388 -12878 49618 -12642
rect 49854 -12878 50000 -12642
rect 42000 -12962 50000 -12878
rect 42000 -13198 42152 -12962
rect 42388 -13198 49618 -12962
rect 49854 -13198 50000 -12962
rect 42000 -13282 50000 -13198
rect 42000 -13518 42152 -13282
rect 42388 -13518 49618 -13282
rect 49854 -13518 50000 -13282
rect 42000 -13602 50000 -13518
rect 42000 -13838 42152 -13602
rect 42388 -13838 49618 -13602
rect 49854 -13838 50000 -13602
rect 42000 -13922 50000 -13838
rect 42000 -14158 42152 -13922
rect 42388 -14158 49618 -13922
rect 49854 -14158 50000 -13922
rect 42000 -14242 50000 -14158
rect 42000 -14478 42152 -14242
rect 42388 -14478 49618 -14242
rect 49854 -14478 50000 -14242
rect 42000 -14562 50000 -14478
rect 42000 -14798 42152 -14562
rect 42388 -14798 49618 -14562
rect 49854 -14798 50000 -14562
rect 42000 -14882 50000 -14798
rect 42000 -15118 42152 -14882
rect 42388 -15118 49618 -14882
rect 49854 -15118 50000 -14882
rect 42000 -15202 50000 -15118
rect 42000 -15438 42152 -15202
rect 42388 -15438 49618 -15202
rect 49854 -15438 50000 -15202
rect 42000 -15522 50000 -15438
rect 42000 -15758 42152 -15522
rect 42388 -15758 49618 -15522
rect 49854 -15758 50000 -15522
rect 42000 -15842 50000 -15758
rect 42000 -16078 42152 -15842
rect 42388 -16078 49618 -15842
rect 49854 -16078 50000 -15842
rect 42000 -16162 50000 -16078
rect 42000 -16398 42152 -16162
rect 42388 -16398 49618 -16162
rect 49854 -16398 50000 -16162
rect 42000 -16482 50000 -16398
rect 42000 -16718 42152 -16482
rect 42388 -16718 49618 -16482
rect 49854 -16718 50000 -16482
rect 42000 -16802 50000 -16718
rect 42000 -17038 42152 -16802
rect 42388 -17038 49618 -16802
rect 49854 -17038 50000 -16802
rect 42000 -17122 50000 -17038
rect 42000 -17358 42152 -17122
rect 42388 -17358 49618 -17122
rect 49854 -17358 50000 -17122
rect 42000 -17442 50000 -17358
rect 42000 -17678 42152 -17442
rect 42388 -17678 49618 -17442
rect 49854 -17678 50000 -17442
rect 42000 -17762 50000 -17678
rect 42000 -17998 42152 -17762
rect 42388 -17998 49618 -17762
rect 49854 -17998 50000 -17762
rect 42000 -18082 50000 -17998
rect 42000 -18318 42152 -18082
rect 42388 -18318 49618 -18082
rect 49854 -18318 50000 -18082
rect 42000 -18402 50000 -18318
rect 42000 -18638 42152 -18402
rect 42388 -18612 49618 -18402
rect 42388 -18638 42522 -18612
rect 42000 -18848 42522 -18638
rect 42758 -18848 42842 -18612
rect 43078 -18848 43162 -18612
rect 43398 -18848 43482 -18612
rect 43718 -18848 43802 -18612
rect 44038 -18848 44122 -18612
rect 44358 -18848 44442 -18612
rect 44678 -18848 44762 -18612
rect 44998 -18848 45082 -18612
rect 45318 -18848 45402 -18612
rect 45638 -18848 45722 -18612
rect 45958 -18848 46042 -18612
rect 46278 -18848 46362 -18612
rect 46598 -18848 46682 -18612
rect 46918 -18848 47002 -18612
rect 47238 -18848 47322 -18612
rect 47558 -18848 47642 -18612
rect 47878 -18848 47962 -18612
rect 48198 -18848 48282 -18612
rect 48518 -18848 48602 -18612
rect 48838 -18848 48922 -18612
rect 49158 -18848 49242 -18612
rect 49478 -18638 49618 -18612
rect 49854 -18638 50000 -18402
rect 49478 -18848 50000 -18638
rect 42000 -19000 50000 -18848
rect 6000 -23156 14000 -23000
rect 6000 -23362 6522 -23156
rect 6000 -23598 6152 -23362
rect 6388 -23392 6522 -23362
rect 6758 -23392 6842 -23156
rect 7078 -23392 7162 -23156
rect 7398 -23392 7482 -23156
rect 7718 -23392 7802 -23156
rect 8038 -23392 8122 -23156
rect 8358 -23392 8442 -23156
rect 8678 -23392 8762 -23156
rect 8998 -23392 9082 -23156
rect 9318 -23392 9402 -23156
rect 9638 -23392 9722 -23156
rect 9958 -23392 10042 -23156
rect 10278 -23392 10362 -23156
rect 10598 -23392 10682 -23156
rect 10918 -23392 11002 -23156
rect 11238 -23392 11322 -23156
rect 11558 -23392 11642 -23156
rect 11878 -23392 11962 -23156
rect 12198 -23392 12282 -23156
rect 12518 -23392 12602 -23156
rect 12838 -23392 12922 -23156
rect 13158 -23392 13242 -23156
rect 13478 -23362 14000 -23156
rect 13478 -23392 13618 -23362
rect 6388 -23598 13618 -23392
rect 13854 -23598 14000 -23362
rect 6000 -23682 14000 -23598
rect 6000 -23918 6152 -23682
rect 6388 -23918 13618 -23682
rect 13854 -23918 14000 -23682
rect 6000 -24002 14000 -23918
rect 6000 -24238 6152 -24002
rect 6388 -24238 13618 -24002
rect 13854 -24238 14000 -24002
rect 6000 -24322 14000 -24238
rect 6000 -24558 6152 -24322
rect 6388 -24558 13618 -24322
rect 13854 -24558 14000 -24322
rect 6000 -24642 14000 -24558
rect 6000 -24878 6152 -24642
rect 6388 -24878 13618 -24642
rect 13854 -24878 14000 -24642
rect 6000 -24962 14000 -24878
rect 6000 -25198 6152 -24962
rect 6388 -25198 13618 -24962
rect 13854 -25198 14000 -24962
rect 6000 -25282 14000 -25198
rect 6000 -25518 6152 -25282
rect 6388 -25518 13618 -25282
rect 13854 -25518 14000 -25282
rect 6000 -25602 14000 -25518
rect 6000 -25838 6152 -25602
rect 6388 -25838 13618 -25602
rect 13854 -25838 14000 -25602
rect 6000 -25922 14000 -25838
rect 6000 -26158 6152 -25922
rect 6388 -26158 13618 -25922
rect 13854 -26158 14000 -25922
rect 6000 -26242 14000 -26158
rect 6000 -26478 6152 -26242
rect 6388 -26478 13618 -26242
rect 13854 -26478 14000 -26242
rect 6000 -26562 14000 -26478
rect 6000 -26798 6152 -26562
rect 6388 -26798 13618 -26562
rect 13854 -26798 14000 -26562
rect 6000 -26882 14000 -26798
rect 6000 -27118 6152 -26882
rect 6388 -27118 13618 -26882
rect 13854 -27118 14000 -26882
rect 6000 -27202 14000 -27118
rect 6000 -27438 6152 -27202
rect 6388 -27438 13618 -27202
rect 13854 -27438 14000 -27202
rect 6000 -27522 14000 -27438
rect 6000 -27758 6152 -27522
rect 6388 -27758 13618 -27522
rect 13854 -27758 14000 -27522
rect 6000 -27842 14000 -27758
rect 6000 -28078 6152 -27842
rect 6388 -28078 13618 -27842
rect 13854 -28078 14000 -27842
rect 6000 -28162 14000 -28078
rect 6000 -28398 6152 -28162
rect 6388 -28398 13618 -28162
rect 13854 -28398 14000 -28162
rect 6000 -28482 14000 -28398
rect 6000 -28718 6152 -28482
rect 6388 -28718 13618 -28482
rect 13854 -28718 14000 -28482
rect 6000 -28802 14000 -28718
rect 6000 -29038 6152 -28802
rect 6388 -29038 13618 -28802
rect 13854 -29038 14000 -28802
rect 6000 -29122 14000 -29038
rect 6000 -29358 6152 -29122
rect 6388 -29358 13618 -29122
rect 13854 -29358 14000 -29122
rect 6000 -29442 14000 -29358
rect 6000 -29678 6152 -29442
rect 6388 -29678 13618 -29442
rect 13854 -29678 14000 -29442
rect 6000 -29762 14000 -29678
rect 6000 -29998 6152 -29762
rect 6388 -29998 13618 -29762
rect 13854 -29998 14000 -29762
rect 6000 -30082 14000 -29998
rect 6000 -30318 6152 -30082
rect 6388 -30318 13618 -30082
rect 13854 -30318 14000 -30082
rect 6000 -30402 14000 -30318
rect 6000 -30638 6152 -30402
rect 6388 -30612 13618 -30402
rect 6388 -30638 6522 -30612
rect 6000 -30848 6522 -30638
rect 6758 -30848 6842 -30612
rect 7078 -30848 7162 -30612
rect 7398 -30848 7482 -30612
rect 7718 -30848 7802 -30612
rect 8038 -30848 8122 -30612
rect 8358 -30848 8442 -30612
rect 8678 -30848 8762 -30612
rect 8998 -30848 9082 -30612
rect 9318 -30848 9402 -30612
rect 9638 -30848 9722 -30612
rect 9958 -30848 10042 -30612
rect 10278 -30848 10362 -30612
rect 10598 -30848 10682 -30612
rect 10918 -30848 11002 -30612
rect 11238 -30848 11322 -30612
rect 11558 -30848 11642 -30612
rect 11878 -30848 11962 -30612
rect 12198 -30848 12282 -30612
rect 12518 -30848 12602 -30612
rect 12838 -30848 12922 -30612
rect 13158 -30848 13242 -30612
rect 13478 -30638 13618 -30612
rect 13854 -30638 14000 -30402
rect 13478 -30848 14000 -30638
rect 6000 -31000 14000 -30848
rect 18000 -23156 26000 -23000
rect 18000 -23362 18522 -23156
rect 18000 -23598 18152 -23362
rect 18388 -23392 18522 -23362
rect 18758 -23392 18842 -23156
rect 19078 -23392 19162 -23156
rect 19398 -23392 19482 -23156
rect 19718 -23392 19802 -23156
rect 20038 -23392 20122 -23156
rect 20358 -23392 20442 -23156
rect 20678 -23392 20762 -23156
rect 20998 -23392 21082 -23156
rect 21318 -23392 21402 -23156
rect 21638 -23392 21722 -23156
rect 21958 -23392 22042 -23156
rect 22278 -23392 22362 -23156
rect 22598 -23392 22682 -23156
rect 22918 -23392 23002 -23156
rect 23238 -23392 23322 -23156
rect 23558 -23392 23642 -23156
rect 23878 -23392 23962 -23156
rect 24198 -23392 24282 -23156
rect 24518 -23392 24602 -23156
rect 24838 -23392 24922 -23156
rect 25158 -23392 25242 -23156
rect 25478 -23362 26000 -23156
rect 25478 -23392 25618 -23362
rect 18388 -23598 25618 -23392
rect 25854 -23598 26000 -23362
rect 18000 -23682 26000 -23598
rect 18000 -23918 18152 -23682
rect 18388 -23918 25618 -23682
rect 25854 -23918 26000 -23682
rect 18000 -24002 26000 -23918
rect 18000 -24238 18152 -24002
rect 18388 -24238 25618 -24002
rect 25854 -24238 26000 -24002
rect 18000 -24322 26000 -24238
rect 18000 -24558 18152 -24322
rect 18388 -24558 25618 -24322
rect 25854 -24558 26000 -24322
rect 18000 -24642 26000 -24558
rect 18000 -24878 18152 -24642
rect 18388 -24878 25618 -24642
rect 25854 -24878 26000 -24642
rect 18000 -24962 26000 -24878
rect 18000 -25198 18152 -24962
rect 18388 -25198 25618 -24962
rect 25854 -25198 26000 -24962
rect 18000 -25282 26000 -25198
rect 18000 -25518 18152 -25282
rect 18388 -25518 25618 -25282
rect 25854 -25518 26000 -25282
rect 18000 -25602 26000 -25518
rect 18000 -25838 18152 -25602
rect 18388 -25838 25618 -25602
rect 25854 -25838 26000 -25602
rect 18000 -25922 26000 -25838
rect 18000 -26158 18152 -25922
rect 18388 -26158 25618 -25922
rect 25854 -26158 26000 -25922
rect 18000 -26242 26000 -26158
rect 18000 -26478 18152 -26242
rect 18388 -26478 25618 -26242
rect 25854 -26478 26000 -26242
rect 18000 -26562 26000 -26478
rect 18000 -26798 18152 -26562
rect 18388 -26798 25618 -26562
rect 25854 -26798 26000 -26562
rect 18000 -26882 26000 -26798
rect 18000 -27118 18152 -26882
rect 18388 -27118 25618 -26882
rect 25854 -27118 26000 -26882
rect 18000 -27202 26000 -27118
rect 18000 -27438 18152 -27202
rect 18388 -27438 25618 -27202
rect 25854 -27438 26000 -27202
rect 18000 -27522 26000 -27438
rect 18000 -27758 18152 -27522
rect 18388 -27758 25618 -27522
rect 25854 -27758 26000 -27522
rect 18000 -27842 26000 -27758
rect 18000 -28078 18152 -27842
rect 18388 -28078 25618 -27842
rect 25854 -28078 26000 -27842
rect 18000 -28162 26000 -28078
rect 18000 -28398 18152 -28162
rect 18388 -28398 25618 -28162
rect 25854 -28398 26000 -28162
rect 18000 -28482 26000 -28398
rect 18000 -28718 18152 -28482
rect 18388 -28718 25618 -28482
rect 25854 -28718 26000 -28482
rect 18000 -28802 26000 -28718
rect 18000 -29038 18152 -28802
rect 18388 -29038 25618 -28802
rect 25854 -29038 26000 -28802
rect 18000 -29122 26000 -29038
rect 18000 -29358 18152 -29122
rect 18388 -29358 25618 -29122
rect 25854 -29358 26000 -29122
rect 18000 -29442 26000 -29358
rect 18000 -29678 18152 -29442
rect 18388 -29678 25618 -29442
rect 25854 -29678 26000 -29442
rect 18000 -29762 26000 -29678
rect 18000 -29998 18152 -29762
rect 18388 -29998 25618 -29762
rect 25854 -29998 26000 -29762
rect 18000 -30082 26000 -29998
rect 18000 -30318 18152 -30082
rect 18388 -30318 25618 -30082
rect 25854 -30318 26000 -30082
rect 18000 -30402 26000 -30318
rect 18000 -30638 18152 -30402
rect 18388 -30612 25618 -30402
rect 18388 -30638 18522 -30612
rect 18000 -30848 18522 -30638
rect 18758 -30848 18842 -30612
rect 19078 -30848 19162 -30612
rect 19398 -30848 19482 -30612
rect 19718 -30848 19802 -30612
rect 20038 -30848 20122 -30612
rect 20358 -30848 20442 -30612
rect 20678 -30848 20762 -30612
rect 20998 -30848 21082 -30612
rect 21318 -30848 21402 -30612
rect 21638 -30848 21722 -30612
rect 21958 -30848 22042 -30612
rect 22278 -30848 22362 -30612
rect 22598 -30848 22682 -30612
rect 22918 -30848 23002 -30612
rect 23238 -30848 23322 -30612
rect 23558 -30848 23642 -30612
rect 23878 -30848 23962 -30612
rect 24198 -30848 24282 -30612
rect 24518 -30848 24602 -30612
rect 24838 -30848 24922 -30612
rect 25158 -30848 25242 -30612
rect 25478 -30638 25618 -30612
rect 25854 -30638 26000 -30402
rect 25478 -30848 26000 -30638
rect 18000 -31000 26000 -30848
rect 30000 -23156 38000 -23000
rect 30000 -23362 30522 -23156
rect 30000 -23598 30152 -23362
rect 30388 -23392 30522 -23362
rect 30758 -23392 30842 -23156
rect 31078 -23392 31162 -23156
rect 31398 -23392 31482 -23156
rect 31718 -23392 31802 -23156
rect 32038 -23392 32122 -23156
rect 32358 -23392 32442 -23156
rect 32678 -23392 32762 -23156
rect 32998 -23392 33082 -23156
rect 33318 -23392 33402 -23156
rect 33638 -23392 33722 -23156
rect 33958 -23392 34042 -23156
rect 34278 -23392 34362 -23156
rect 34598 -23392 34682 -23156
rect 34918 -23392 35002 -23156
rect 35238 -23392 35322 -23156
rect 35558 -23392 35642 -23156
rect 35878 -23392 35962 -23156
rect 36198 -23392 36282 -23156
rect 36518 -23392 36602 -23156
rect 36838 -23392 36922 -23156
rect 37158 -23392 37242 -23156
rect 37478 -23362 38000 -23156
rect 37478 -23392 37618 -23362
rect 30388 -23598 37618 -23392
rect 37854 -23598 38000 -23362
rect 30000 -23682 38000 -23598
rect 30000 -23918 30152 -23682
rect 30388 -23918 37618 -23682
rect 37854 -23918 38000 -23682
rect 30000 -24002 38000 -23918
rect 30000 -24238 30152 -24002
rect 30388 -24238 37618 -24002
rect 37854 -24238 38000 -24002
rect 30000 -24322 38000 -24238
rect 30000 -24558 30152 -24322
rect 30388 -24558 37618 -24322
rect 37854 -24558 38000 -24322
rect 30000 -24642 38000 -24558
rect 30000 -24878 30152 -24642
rect 30388 -24878 37618 -24642
rect 37854 -24878 38000 -24642
rect 30000 -24962 38000 -24878
rect 30000 -25198 30152 -24962
rect 30388 -25198 37618 -24962
rect 37854 -25198 38000 -24962
rect 30000 -25282 38000 -25198
rect 30000 -25518 30152 -25282
rect 30388 -25518 37618 -25282
rect 37854 -25518 38000 -25282
rect 30000 -25602 38000 -25518
rect 30000 -25838 30152 -25602
rect 30388 -25838 37618 -25602
rect 37854 -25838 38000 -25602
rect 30000 -25922 38000 -25838
rect 30000 -26158 30152 -25922
rect 30388 -26158 37618 -25922
rect 37854 -26158 38000 -25922
rect 30000 -26242 38000 -26158
rect 30000 -26478 30152 -26242
rect 30388 -26478 37618 -26242
rect 37854 -26478 38000 -26242
rect 30000 -26562 38000 -26478
rect 30000 -26798 30152 -26562
rect 30388 -26798 37618 -26562
rect 37854 -26798 38000 -26562
rect 30000 -26882 38000 -26798
rect 30000 -27118 30152 -26882
rect 30388 -27118 37618 -26882
rect 37854 -27118 38000 -26882
rect 30000 -27202 38000 -27118
rect 30000 -27438 30152 -27202
rect 30388 -27438 37618 -27202
rect 37854 -27438 38000 -27202
rect 30000 -27522 38000 -27438
rect 30000 -27758 30152 -27522
rect 30388 -27758 37618 -27522
rect 37854 -27758 38000 -27522
rect 30000 -27842 38000 -27758
rect 30000 -28078 30152 -27842
rect 30388 -28078 37618 -27842
rect 37854 -28078 38000 -27842
rect 30000 -28162 38000 -28078
rect 30000 -28398 30152 -28162
rect 30388 -28398 37618 -28162
rect 37854 -28398 38000 -28162
rect 30000 -28482 38000 -28398
rect 30000 -28718 30152 -28482
rect 30388 -28718 37618 -28482
rect 37854 -28718 38000 -28482
rect 30000 -28802 38000 -28718
rect 30000 -29038 30152 -28802
rect 30388 -29038 37618 -28802
rect 37854 -29038 38000 -28802
rect 30000 -29122 38000 -29038
rect 30000 -29358 30152 -29122
rect 30388 -29358 37618 -29122
rect 37854 -29358 38000 -29122
rect 30000 -29442 38000 -29358
rect 30000 -29678 30152 -29442
rect 30388 -29678 37618 -29442
rect 37854 -29678 38000 -29442
rect 30000 -29762 38000 -29678
rect 30000 -29998 30152 -29762
rect 30388 -29998 37618 -29762
rect 37854 -29998 38000 -29762
rect 30000 -30082 38000 -29998
rect 30000 -30318 30152 -30082
rect 30388 -30318 37618 -30082
rect 37854 -30318 38000 -30082
rect 30000 -30402 38000 -30318
rect 30000 -30638 30152 -30402
rect 30388 -30612 37618 -30402
rect 30388 -30638 30522 -30612
rect 30000 -30848 30522 -30638
rect 30758 -30848 30842 -30612
rect 31078 -30848 31162 -30612
rect 31398 -30848 31482 -30612
rect 31718 -30848 31802 -30612
rect 32038 -30848 32122 -30612
rect 32358 -30848 32442 -30612
rect 32678 -30848 32762 -30612
rect 32998 -30848 33082 -30612
rect 33318 -30848 33402 -30612
rect 33638 -30848 33722 -30612
rect 33958 -30848 34042 -30612
rect 34278 -30848 34362 -30612
rect 34598 -30848 34682 -30612
rect 34918 -30848 35002 -30612
rect 35238 -30848 35322 -30612
rect 35558 -30848 35642 -30612
rect 35878 -30848 35962 -30612
rect 36198 -30848 36282 -30612
rect 36518 -30848 36602 -30612
rect 36838 -30848 36922 -30612
rect 37158 -30848 37242 -30612
rect 37478 -30638 37618 -30612
rect 37854 -30638 38000 -30402
rect 37478 -30848 38000 -30638
rect 30000 -31000 38000 -30848
rect 42000 -23156 50000 -23000
rect 42000 -23362 42522 -23156
rect 42000 -23598 42152 -23362
rect 42388 -23392 42522 -23362
rect 42758 -23392 42842 -23156
rect 43078 -23392 43162 -23156
rect 43398 -23392 43482 -23156
rect 43718 -23392 43802 -23156
rect 44038 -23392 44122 -23156
rect 44358 -23392 44442 -23156
rect 44678 -23392 44762 -23156
rect 44998 -23392 45082 -23156
rect 45318 -23392 45402 -23156
rect 45638 -23392 45722 -23156
rect 45958 -23392 46042 -23156
rect 46278 -23392 46362 -23156
rect 46598 -23392 46682 -23156
rect 46918 -23392 47002 -23156
rect 47238 -23392 47322 -23156
rect 47558 -23392 47642 -23156
rect 47878 -23392 47962 -23156
rect 48198 -23392 48282 -23156
rect 48518 -23392 48602 -23156
rect 48838 -23392 48922 -23156
rect 49158 -23392 49242 -23156
rect 49478 -23362 50000 -23156
rect 49478 -23392 49618 -23362
rect 42388 -23598 49618 -23392
rect 49854 -23598 50000 -23362
rect 42000 -23682 50000 -23598
rect 42000 -23918 42152 -23682
rect 42388 -23918 49618 -23682
rect 49854 -23918 50000 -23682
rect 42000 -24002 50000 -23918
rect 42000 -24238 42152 -24002
rect 42388 -24238 49618 -24002
rect 49854 -24238 50000 -24002
rect 42000 -24322 50000 -24238
rect 42000 -24558 42152 -24322
rect 42388 -24558 49618 -24322
rect 49854 -24558 50000 -24322
rect 42000 -24642 50000 -24558
rect 42000 -24878 42152 -24642
rect 42388 -24878 49618 -24642
rect 49854 -24878 50000 -24642
rect 42000 -24962 50000 -24878
rect 42000 -25198 42152 -24962
rect 42388 -25198 49618 -24962
rect 49854 -25198 50000 -24962
rect 42000 -25282 50000 -25198
rect 42000 -25518 42152 -25282
rect 42388 -25518 49618 -25282
rect 49854 -25518 50000 -25282
rect 42000 -25602 50000 -25518
rect 42000 -25838 42152 -25602
rect 42388 -25838 49618 -25602
rect 49854 -25838 50000 -25602
rect 42000 -25922 50000 -25838
rect 42000 -26158 42152 -25922
rect 42388 -26158 49618 -25922
rect 49854 -26158 50000 -25922
rect 42000 -26242 50000 -26158
rect 42000 -26478 42152 -26242
rect 42388 -26478 49618 -26242
rect 49854 -26478 50000 -26242
rect 42000 -26562 50000 -26478
rect 42000 -26798 42152 -26562
rect 42388 -26798 49618 -26562
rect 49854 -26798 50000 -26562
rect 42000 -26882 50000 -26798
rect 42000 -27118 42152 -26882
rect 42388 -27118 49618 -26882
rect 49854 -27118 50000 -26882
rect 42000 -27202 50000 -27118
rect 42000 -27438 42152 -27202
rect 42388 -27438 49618 -27202
rect 49854 -27438 50000 -27202
rect 42000 -27522 50000 -27438
rect 42000 -27758 42152 -27522
rect 42388 -27758 49618 -27522
rect 49854 -27758 50000 -27522
rect 42000 -27842 50000 -27758
rect 42000 -28078 42152 -27842
rect 42388 -28078 49618 -27842
rect 49854 -28078 50000 -27842
rect 42000 -28162 50000 -28078
rect 42000 -28398 42152 -28162
rect 42388 -28398 49618 -28162
rect 49854 -28398 50000 -28162
rect 42000 -28482 50000 -28398
rect 42000 -28718 42152 -28482
rect 42388 -28718 49618 -28482
rect 49854 -28718 50000 -28482
rect 42000 -28802 50000 -28718
rect 42000 -29038 42152 -28802
rect 42388 -29038 49618 -28802
rect 49854 -29038 50000 -28802
rect 42000 -29122 50000 -29038
rect 42000 -29358 42152 -29122
rect 42388 -29358 49618 -29122
rect 49854 -29358 50000 -29122
rect 42000 -29442 50000 -29358
rect 42000 -29678 42152 -29442
rect 42388 -29678 49618 -29442
rect 49854 -29678 50000 -29442
rect 42000 -29762 50000 -29678
rect 42000 -29998 42152 -29762
rect 42388 -29998 49618 -29762
rect 49854 -29998 50000 -29762
rect 42000 -30082 50000 -29998
rect 42000 -30318 42152 -30082
rect 42388 -30318 49618 -30082
rect 49854 -30318 50000 -30082
rect 42000 -30402 50000 -30318
rect 42000 -30638 42152 -30402
rect 42388 -30612 49618 -30402
rect 42388 -30638 42522 -30612
rect 42000 -30848 42522 -30638
rect 42758 -30848 42842 -30612
rect 43078 -30848 43162 -30612
rect 43398 -30848 43482 -30612
rect 43718 -30848 43802 -30612
rect 44038 -30848 44122 -30612
rect 44358 -30848 44442 -30612
rect 44678 -30848 44762 -30612
rect 44998 -30848 45082 -30612
rect 45318 -30848 45402 -30612
rect 45638 -30848 45722 -30612
rect 45958 -30848 46042 -30612
rect 46278 -30848 46362 -30612
rect 46598 -30848 46682 -30612
rect 46918 -30848 47002 -30612
rect 47238 -30848 47322 -30612
rect 47558 -30848 47642 -30612
rect 47878 -30848 47962 -30612
rect 48198 -30848 48282 -30612
rect 48518 -30848 48602 -30612
rect 48838 -30848 48922 -30612
rect 49158 -30848 49242 -30612
rect 49478 -30638 49618 -30612
rect 49854 -30638 50000 -30402
rect 49478 -30848 50000 -30638
rect 42000 -31000 50000 -30848
<< fillblock >>
rect 6000 -20000 8400 -19000
rect 18000 -20000 20400 -19000
rect 30000 -20000 32400 -19000
rect 42000 -20000 44400 -19000
rect 6000 -23000 6800 -21800
rect 18000 -23000 18800 -21820
rect 30000 -23000 33200 -22000
rect 42000 -23000 44400 -22000
<< comment >>
rect 20002 -7600 20005 -3060
rect 1800 -19000 2000 -10600
<< labels >>
rlabel metal5 7200 -17600 12500 -13000 1 VHI
rlabel metal5 19500 -17400 24800 -12800 1 VLO
rlabel metal5 31300 -17400 36600 -12800 1 VIP
rlabel metal5 43300 -17400 48600 -12800 1 VOP
rlabel metal5 43300 -29200 48600 -24600 1 VIN
rlabel metal5 31300 -29300 36600 -24700 1 VREF
rlabel metal5 19400 -29300 24700 -24700 1 SBAR
rlabel metal5 7500 -29400 12800 -24800 1 S
<< end >>
