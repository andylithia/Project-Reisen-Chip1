magic
tech sky130A
timestamp 1672075913
<< metal4 >>
rect -10 285 130 295
rect -10 165 0 285
rect 120 165 130 285
rect -10 155 130 165
rect -10 115 130 125
rect -10 -5 0 115
rect 120 -5 130 115
rect -10 -15 130 -5
<< via4 >>
rect 0 165 120 285
rect 0 -5 120 115
<< metal5 >>
rect -20 285 140 305
rect -20 165 0 285
rect 120 165 140 285
rect -20 115 140 165
rect -20 -5 0 115
rect 120 -5 140 115
rect -20 -25 140 -5
<< end >>
