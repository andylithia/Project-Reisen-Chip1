** sch_path: /home/andylithia/openmpw/Project-Reisen-Chip1/xschem/untitled-2.sch
**.subckt untitled-2
x1 net5 net3 GND net2 net1 net6 net4 net7 net8 GND GND net9 GND net10 net11 GND GND net12 net13 GND
+ net14 GND net15 GND GND net16 GND net17 net18 net19 net20 net21 net22 net23 net24 net25 net26 net27 net28
+ daccon
V1 net1 GND PULSE(0 1.8 10n 1n 1n 100n 200n)
.save i(v1)
V2 net2 GND 1.8
.save i(v2)
V3 net3 GND 0
.save i(v3)
V4 net4 GND PULSE(1.8 0 10n 1n 1n 400n 1)
.save i(v4)
V5 net5 GND 1.8
.save i(v5)
**** begin user architecture code
.lib /home/andylithia/openmpw/pdk_1/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.include /home/andylithia/openmpw/pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice


*.ac dec 100 1e3 1e12
.tran 0.1ns 2500ns
.save all
.control
run
display
plot vout gn gp
.endc


**** end user architecture code
**.ends

* expanding   symbol:  daccon.sym # of pins=39
** sym_path: /home/andylithia/openmpw/Project-Reisen-Chip1/xschem/daccon.sym
** sch_path: /home/andylithia/openmpw/Project-Reisen-Chip1/xschem/daccon.sch
.subckt daccon vccd1 dummy vssd1 test_mode clk msb[15] rst_n msb[14] msb[13] dac_in[9] dac_in[8]
+ msb[12] dac_in[7] msb[11] msb[10] dac_in[6] dac_in[5] msb[9] msb[8] dac_in[4] msb[7] dac_in[3] msb[6]
+ dac_in[2] dac_in[1] msb[5] dac_in[0] msb[4] msb[3] msb[2] msb[1] msb[0] lsb[6] lsb[5] lsb[4] lsb[3] lsb[2]
+ lsb[1] lsb[0]
*.ipin test_mode
*.ipin clk
*.ipin rst_n
*.ipin dac_in[9]
*.ipin dac_in[8]
*.ipin dac_in[7]
*.ipin dac_in[6]
*.ipin dac_in[5]
*.ipin dac_in[4]
*.ipin dac_in[3]
*.ipin dac_in[2]
*.ipin dac_in[1]
*.ipin dac_in[0]
*.iopin vccd1
*.iopin vssd1
*.ipin dummy
*.opin msb[15]
*.opin msb[14]
*.opin msb[13]
*.opin msb[12]
*.opin msb[11]
*.opin msb[10]
*.opin msb[9]
*.opin msb[8]
*.opin msb[7]
*.opin msb[6]
*.opin msb[5]
*.opin msb[4]
*.opin msb[3]
*.opin msb[2]
*.opin msb[1]
*.opin msb[0]
*.opin lsb[6]
*.opin lsb[5]
*.opin lsb[4]
*.opin lsb[3]
*.opin lsb[2]
*.opin lsb[1]
*.opin lsb[0]
**** begin user architecture code

* NGSPICE file created from dac_con.ext - technology: sky130A

.subckt dac_con clk dac_in[0] dac_in[1] dac_in[2] dac_in[3] dac_in[4] dac_in[5] dac_in[6]  dac_in[7]
+ dac_in[8] dac_in[9] dummy llsb llsb_n lsb[0] lsb[1] lsb[2] lsb[3] lsb[4]  lsb[5] lsb_n[0] lsb_n[1] lsb_n[2]
+ lsb_n[3] lsb_n[4] lsb_n[5] msb[0] msb[10] msb[11]  msb[12] msb[13] msb[14] msb[15] msb[1] msb[2] msb[3]
+ msb[4] msb[5] msb[6] msb[7]  msb[8] msb[9] msb_n[0] msb_n[10] msb_n[11] msb_n[12] msb_n[13] msb_n[14]
+ msb_n[15]  msb_n[1] msb_n[2] msb_n[3] msb_n[4] msb_n[5] msb_n[6] msb_n[7] msb_n[8] msb_n[9]  rst_n test_mode
+ vccd1 vssd1
C0 _040_ vccd1 2.89fF
C1 _019_ vccd1 2.21fF
C2 _049_ vccd1 3.09fF
C3 cnt_r\[8\] vccd1 2.02fF
C4 _082_ vccd1 5.33fF
C5 _089_ vccd1 6.65fF
C6 clknet_2_2__leaf_clk vccd1 3.82fF
C7 _053_ vccd1 2.88fF
C8 clknet_2_0__leaf_clk vccd1 5.31fF
C9 vccd1 _045_ 3.19fF
C10 dac_in[5] vccd1 2.91fF
C11 _044_ vccd1 5.54fF
C12 _038_ vccd1 3.29fF
C13 net29 vccd1 2.36fF
C14 vccd1 _065_ 4.79fF
C15 vccd1 net28 2.20fF
C16 _041_ vccd1 11.19fF
C17 net12 vccd1 3.23fF
C18 net34 vccd1 2.13fF
C19 vccd1 clknet_2_3__leaf_clk 5.25fF
C20 _085_ vccd1 2.40fF
C21 vccd1 _063_ 5.70fF
C22 dac_in[3] vccd1 2.38fF
C23 net13 vccd1 2.15fF
C24 net37 vccd1 2.60fF
C25 clknet_2_1__leaf_clk vccd1 4.14fF
C26 net33 vccd1 2.21fF
C27 vccd1 _034_ 8.79fF
C28 cnt_r\[9\] _055_ 2.07fF
C29 _085_ _082_ 2.25fF
C30 net30 vccd1 3.63fF
C31 vccd1 net16 2.26fF
C32 _078_ vccd1 2.57fF
C33 clknet_2_2__leaf_clk _063_ 2.39fF
C34 _087_ vccd1 4.40fF
C35 _052_ vccd1 2.32fF
C36 clk vccd1 4.57fF
C37 _064_ vccd1 4.30fF
C38 vccd1 net19 2.25fF
C39 _037_ vccd1 3.80fF
C40 net3 vccd1 2.94fF
C41 vccd1 net18 2.57fF
C42 clknet_0_clk vccd1 2.98fF
X_131_ _044_ cnt_r\[2\] cnt_r\[0\] cnt_r\[1\] cnt_r\[3\] vssd1 vccd1 sky130_fd_sc_hd__and4_1
X_200_ vccd1 vssd1 _041_ _091_ sky130_fd_sc_hd__dlymetal6s2s_1
X_114_ net26 net20 vccd1 vssd1 sky130_fd_sc_hd__clkinv_2
Xoutput20 vccd1 vssd1 lsb[4] net20 sky130_fd_sc_hd__buf_2
Xoutput53 vccd1 vssd1 msb_n[3] net53 sky130_fd_sc_hd__buf_2
Xoutput42 vccd1 vssd1 msb[8] net42 sky130_fd_sc_hd__buf_2
Xoutput31 vccd1 vssd1 msb[12] net31 sky130_fd_sc_hd__buf_2
X_130_ vssd1 vccd1 _003_ _043_ sky130_fd_sc_hd__clkbuf_1
X_113_ net25 net19 vccd1 vssd1 sky130_fd_sc_hd__clkinv_2
Xoutput54 vccd1 vssd1 msb_n[4] net54 sky130_fd_sc_hd__buf_2
Xoutput43 vccd1 vssd1 msb[9] net43 sky130_fd_sc_hd__buf_2
Xoutput32 vccd1 vssd1 msb[13] net32 sky130_fd_sc_hd__buf_2
Xoutput21 vccd1 vssd1 lsb[5] net21 sky130_fd_sc_hd__buf_2
X_189_ vccd1 vssd1 _081_ _085_ sky130_fd_sc_hd__dlymetal6s2s_1
X_112_ net24 net18 vccd1 vssd1 sky130_fd_sc_hd__clkinv_2
Xoutput55 vccd1 vssd1 msb_n[5] net55 sky130_fd_sc_hd__buf_2
Xoutput33 vccd1 vssd1 msb[14] net33 sky130_fd_sc_hd__buf_2
Xoutput22 vccd1 vssd1 lsb_n[0] net22 sky130_fd_sc_hd__buf_2
Xoutput44 vccd1 vssd1 msb_n[0] net44 sky130_fd_sc_hd__buf_2
X_188_ _082_ _032_ _021_ _018_ vccd1 vssd1 sky130_fd_sc_hd__a21o_1
X_111_ net23 net17 vccd1 vssd1 sky130_fd_sc_hd__clkinv_2
Xoutput23 vccd1 vssd1 lsb_n[1] net23 sky130_fd_sc_hd__buf_2
Xoutput56 vccd1 vssd1 msb_n[6] net56 sky130_fd_sc_hd__buf_2
Xoutput45 vccd1 vssd1 msb_n[10] net45 sky130_fd_sc_hd__buf_2
Xoutput34 vccd1 vssd1 msb[15] net34 sky130_fd_sc_hd__buf_2
X_187_ vccd1 vssd1 _084_ _021_ sky130_fd_sc_hd__dlymetal6s2s_1
X_110_ net22 net16 vccd1 vssd1 sky130_fd_sc_hd__clkinv_2
X_239_ net40 clknet_2_1__leaf_clk _030_ vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1
Xoutput24 vccd1 vssd1 lsb_n[2] net24 sky130_fd_sc_hd__buf_2
Xoutput35 vccd1 vssd1 msb[1] net35 sky130_fd_sc_hd__buf_2
Xoutput57 vccd1 vssd1 msb_n[7] net57 sky130_fd_sc_hd__buf_2
Xoutput46 vccd1 vssd1 msb_n[11] net46 sky130_fd_sc_hd__buf_2
X_186_ vssd1 vccd1 _084_ _078_ net12 _083_ sky130_fd_sc_hd__and3_1
X_169_ vssd1 vccd1 _014_ _071_ sky130_fd_sc_hd__clkbuf_1
X_238_ net39 clknet_2_1__leaf_clk _029_ vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1
Xoutput36 vccd1 vssd1 msb[2] net36 sky130_fd_sc_hd__buf_2
Xoutput25 vccd1 vssd1 lsb_n[3] net25 sky130_fd_sc_hd__buf_2
Xoutput58 vccd1 vssd1 msb_n[8] net58 sky130_fd_sc_hd__buf_2
Xoutput47 vccd1 vssd1 msb_n[12] net47 sky130_fd_sc_hd__buf_2
Xoutput14 vccd1 vssd1 llsb net14 sky130_fd_sc_hd__buf_2
XPHY_0 vccd1 vssd1 sky130_fd_sc_hd__decap_3
X_185_ vssd1 vccd1 _064_ cnt_r\[8\] net9 _083_ sky130_fd_sc_hd__mux2_1
X_099_ net55 net39 vccd1 vssd1 sky130_fd_sc_hd__clkinv_2
X_237_ net38 clknet_2_3__leaf_clk _028_ vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1
X_168_ vccd1 vssd1 _071_ _070_ _063_ sky130_fd_sc_hd__and2_1
Xoutput26 vccd1 vssd1 lsb_n[4] net26 sky130_fd_sc_hd__buf_2
Xoutput37 vccd1 vssd1 msb[3] net37 sky130_fd_sc_hd__buf_2
Xoutput59 vccd1 vssd1 msb_n[9] net59 sky130_fd_sc_hd__buf_2
Xoutput48 vccd1 vssd1 msb_n[13] net48 sky130_fd_sc_hd__buf_2
Xoutput15 vccd1 vssd1 llsb_n net15 sky130_fd_sc_hd__buf_2
XPHY_1 vccd1 vssd1 sky130_fd_sc_hd__decap_3
X_184_ _080_ _082_ _081_ vssd1 vccd1 sky130_fd_sc_hd__or2_1
X_098_ net54 net38 vccd1 vssd1 sky130_fd_sc_hd__clkinv_2
X_167_ vssd1 vccd1 _065_ cnt_r\[2\] net3 _070_ sky130_fd_sc_hd__mux2_1
X_236_ net37 clknet_2_2__leaf_clk _027_ vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1
X_219_ cnt_r\[9\] clknet_2_0__leaf_clk _010_ vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1
Xoutput16 vccd1 vssd1 lsb[0] net16 sky130_fd_sc_hd__buf_2
Xoutput27 vccd1 vssd1 lsb_n[5] net27 sky130_fd_sc_hd__buf_2
Xoutput38 vccd1 vssd1 msb[4] net38 sky130_fd_sc_hd__buf_2
Xoutput49 vccd1 vssd1 msb_n[14] net49 sky130_fd_sc_hd__buf_2
XPHY_2 vccd1 vssd1 sky130_fd_sc_hd__decap_3
Xclkbuf_0_clk clknet_0_clk clk vssd1 vccd1 sky130_fd_sc_hd__clkbuf_16
X_183_ vssd1 vccd1 _064_ cnt_r\[7\] net8 _081_ sky130_fd_sc_hd__mux2_1
X_235_ net36 clknet_2_3__leaf_clk _026_ vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1
X_097_ net53 net37 vccd1 vssd1 sky130_fd_sc_hd__clkinv_2
X_166_ vssd1 vccd1 _013_ _069_ sky130_fd_sc_hd__clkbuf_1
X_218_ cnt_r\[8\] clknet_2_0__leaf_clk _009_ vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1
X_149_ _052_ _055_ cnt_r\[8\] _057_ vccd1 vssd1 sky130_fd_sc_hd__a21o_1
Xoutput17 vccd1 vssd1 lsb[1] net17 sky130_fd_sc_hd__buf_2
Xoutput28 vccd1 vssd1 msb[0] net28 sky130_fd_sc_hd__buf_2
Xoutput39 vccd1 vssd1 msb[5] net39 sky130_fd_sc_hd__buf_2
XPHY_3 vccd1 vssd1 sky130_fd_sc_hd__decap_3
Xclkbuf_2_0__f_clk clknet_2_0__leaf_clk clknet_0_clk vssd1 vccd1 sky130_fd_sc_hd__clkbuf_16
X_182_ vssd1 vccd1 _064_ cnt_r\[6\] net7 _080_ sky130_fd_sc_hd__mux2_1
X_096_ net52 net36 vccd1 vssd1 sky130_fd_sc_hd__clkinv_2
X_234_ net35 clknet_2_3__leaf_clk _025_ vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1
X_165_ vccd1 vssd1 _069_ _068_ _063_ sky130_fd_sc_hd__and2_1
X_217_ cnt_r\[7\] clknet_2_0__leaf_clk _008_ vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1
X_148_ _008_ _055_ _056_ _053_ vssd1 vccd1 sky130_fd_sc_hd__o21a_1
Xoutput18 vccd1 vssd1 lsb[2] net18 sky130_fd_sc_hd__buf_2
Xoutput29 vccd1 vssd1 msb[10] net29 sky130_fd_sc_hd__buf_2
XPHY_4 vccd1 vssd1 sky130_fd_sc_hd__decap_3
X_181_ vccd1 vssd1 _079_ _032_ sky130_fd_sc_hd__dlymetal6s2s_1
X_095_ net35 net51 vccd1 vssd1 sky130_fd_sc_hd__inv_2
X_164_ vssd1 vccd1 _065_ _038_ net2 _068_ sky130_fd_sc_hd__mux2_1
X_233_ net34 clknet_2_0__leaf_clk _024_ vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1
X_216_ cnt_r\[6\] clknet_2_0__leaf_clk _007_ vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1
X_147_ _055_ _037_ _056_ _053_ vccd1 vssd1 sky130_fd_sc_hd__a21oi_1
Xoutput19 vccd1 vssd1 lsb[3] net19 sky130_fd_sc_hd__buf_2
XPHY_5 vccd1 vssd1 sky130_fd_sc_hd__decap_3
X_180_ vccd1 vssd1 _079_ _078_ _033_ sky130_fd_sc_hd__and2_1
X_094_ net28 net44 vccd1 vssd1 sky130_fd_sc_hd__inv_2
X_232_ net33 clknet_2_1__leaf_clk _023_ vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1
X_163_ vssd1 vccd1 _012_ _067_ sky130_fd_sc_hd__clkbuf_1
X_146_ vccd1 vssd1 cnt_r\[7\] _055_ sky130_fd_sc_hd__dlymetal6s2s_1
X_215_ cnt_r\[5\] clknet_2_2__leaf_clk _006_ vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1
XPHY_6 vccd1 vssd1 sky130_fd_sc_hd__decap_3
X_129_ _040_ _041_ _043_ _042_ vssd1 vccd1 sky130_fd_sc_hd__and3b_1
X_093_ net15 net14 vccd1 vssd1 sky130_fd_sc_hd__clkinv_2
X_231_ net32 clknet_2_1__leaf_clk _022_ vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1
X_162_ vccd1 vssd1 _067_ _066_ _063_ sky130_fd_sc_hd__and2_1
Xinput1 vssd1 vccd1 net1 dac_in[0] sky130_fd_sc_hd__clkbuf_1
X_214_ cnt_r\[4\] clknet_2_2__leaf_clk _005_ vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1
X_145_ _054_ _007_ _053_ vssd1 vccd1 sky130_fd_sc_hd__nor2_1
XPHY_7 vccd1 vssd1 sky130_fd_sc_hd__decap_3
X_128_ _038_ _036_ cnt_r\[2\] _042_ vccd1 vssd1 sky130_fd_sc_hd__a21o_1
X_161_ vssd1 vccd1 _065_ _036_ net1 _066_ sky130_fd_sc_hd__mux2_1
X_230_ net31 clknet_2_1__leaf_clk _021_ vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1
Xinput2 vssd1 vccd1 net2 dac_in[1] sky130_fd_sc_hd__clkbuf_1
X_144_ vssd1 vccd1 _049_ cnt_r\[6\] _034_ _054_ sky130_fd_sc_hd__o21ai_1
X_213_ cnt_r\[3\] clknet_2_2__leaf_clk _004_ vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1
X_127_ vccd1 vssd1 _033_ _041_ sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_8 vccd1 vssd1 sky130_fd_sc_hd__decap_3
X_160_ _064_ _065_ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_2
Xinput3 vssd1 vccd1 net3 dac_in[2] sky130_fd_sc_hd__clkbuf_1
X_143_ vccd1 vssd1 _052_ _053_ sky130_fd_sc_hd__dlymetal6s2s_1
X_212_ cnt_r\[2\] clknet_2_2__leaf_clk _003_ vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1
XPHY_9 vccd1 vssd1 sky130_fd_sc_hd__decap_3
X_126_ vssd1 vccd1 _040_ _038_ cnt_r\[0\] cnt_r\[2\] sky130_fd_sc_hd__and3_1
X_109_ net34 net50 vccd1 vssd1 sky130_fd_sc_hd__inv_2
Xinput4 vssd1 vccd1 net4 dac_in[3] sky130_fd_sc_hd__clkbuf_1
Xclkbuf_2_1__f_clk clknet_2_1__leaf_clk clknet_0_clk vssd1 vccd1 sky130_fd_sc_hd__clkbuf_16
X_142_ _052_ cnt_r\[6\] cnt_r\[4\] cnt_r\[5\] _044_ vssd1 vccd1 sky130_fd_sc_hd__and4_1
X_211_ cnt_r\[1\] clknet_2_2__leaf_clk _002_ vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1
X_125_ _036_ _039_ _002_ _038_ vccd1 vssd1 sky130_fd_sc_hd__a21oi_1
X_108_ net49 net33 vccd1 vssd1 sky130_fd_sc_hd__clkinv_2
Xinput5 vssd1 vccd1 net5 dac_in[4] sky130_fd_sc_hd__clkbuf_1
X_141_ vssd1 vccd1 _006_ _051_ sky130_fd_sc_hd__clkbuf_1
X_210_ cnt_r\[0\] clknet_2_2__leaf_clk _001_ vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1
X_124_ vssd1 vccd1 _038_ _036_ _034_ _039_ sky130_fd_sc_hd__o21ai_1
X_107_ net48 net32 vccd1 vssd1 sky130_fd_sc_hd__clkinv_2
Xinput6 vssd1 vccd1 net6 dac_in[5] sky130_fd_sc_hd__clkbuf_1
X_140_ _049_ _041_ _051_ _050_ vssd1 vccd1 sky130_fd_sc_hd__and3b_1
X_123_ vccd1 vssd1 cnt_r\[1\] _038_ sky130_fd_sc_hd__dlymetal6s2s_1
X_106_ net47 net31 vccd1 vssd1 sky130_fd_sc_hd__clkinv_2
Xinput7 vssd1 vccd1 net7 dac_in[6] sky130_fd_sc_hd__clkbuf_1
X_199_ vssd1 vccd1 _024_ _090_ sky130_fd_sc_hd__clkbuf_1
X_122_ _037_ _001_ _036_ vssd1 vccd1 sky130_fd_sc_hd__nor2_1
Xinput10 vssd1 vccd1 net10 dac_in[9] sky130_fd_sc_hd__clkbuf_1
X_105_ net46 net30 vccd1 vssd1 sky130_fd_sc_hd__clkinv_2
Xinput8 vssd1 vccd1 net8 dac_in[7] sky130_fd_sc_hd__clkbuf_1
X_198_ vccd1 vssd1 _090_ _087_ _084_ sky130_fd_sc_hd__and2_1
X_121_ _037_ net12 vccd1 vssd1 sky130_fd_sc_hd__clkinv_2
Xinput11 vssd1 vccd1 net11 dummy sky130_fd_sc_hd__clkbuf_1
X_104_ net45 net29 vccd1 vssd1 sky130_fd_sc_hd__clkinv_2
Xinput9 vssd1 vccd1 net9 dac_in[8] sky130_fd_sc_hd__clkbuf_1
X_197_ vssd1 vccd1 _023_ _089_ sky130_fd_sc_hd__clkbuf_1
X_120_ vccd1 vssd1 cnt_r\[0\] _036_ sky130_fd_sc_hd__dlymetal6s2s_1
Xinput12 vssd1 vccd1 net12 rst_n sky130_fd_sc_hd__clkbuf_1
X_103_ net59 net43 vccd1 vssd1 sky130_fd_sc_hd__clkinv_2
X_196_ vccd1 vssd1 _089_ _085_ _021_ sky130_fd_sc_hd__and2_1
Xinput13 vssd1 vccd1 net13 test_mode sky130_fd_sc_hd__clkbuf_1
X_179_ vssd1 vccd1 net13 cnt_r\[9\] net10 _078_ sky130_fd_sc_hd__mux2_1
X_102_ net58 net42 vccd1 vssd1 sky130_fd_sc_hd__clkinv_2
Xclkbuf_2_2__f_clk clknet_2_2__leaf_clk clknet_0_clk vssd1 vccd1 sky130_fd_sc_hd__clkbuf_16
X_195_ vssd1 vccd1 _022_ _088_ sky130_fd_sc_hd__clkbuf_1
X_178_ vssd1 vccd1 _017_ _077_ sky130_fd_sc_hd__clkbuf_1
X_101_ net57 net41 vccd1 vssd1 sky130_fd_sc_hd__clkinv_2
X_194_ vccd1 vssd1 _088_ _082_ _021_ sky130_fd_sc_hd__and2_1
X_177_ vccd1 vssd1 _077_ _076_ _041_ sky130_fd_sc_hd__and2_1
X_100_ net56 net40 vccd1 vssd1 sky130_fd_sc_hd__clkinv_2
X_229_ net30 clknet_2_1__leaf_clk _020_ vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1
X_193_ _020_ _086_ _032_ _087_ vssd1 vccd1 sky130_fd_sc_hd__o21a_1
X_176_ vssd1 vccd1 _064_ cnt_r\[5\] net6 _076_ sky130_fd_sc_hd__mux2_1
X_228_ net29 clknet_2_0__leaf_clk _019_ vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1
X_159_ net13 _064_ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_2
X_192_ vccd1 vssd1 _087_ _085_ _080_ sky130_fd_sc_hd__and2_1
XPHY_10 vccd1 vssd1 sky130_fd_sc_hd__decap_3
X_175_ vssd1 vccd1 _016_ _075_ sky130_fd_sc_hd__clkbuf_1
X_158_ vccd1 vssd1 _033_ _063_ sky130_fd_sc_hd__dlymetal6s2s_1
X_227_ net43 clknet_2_1__leaf_clk _018_ vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1
XPHY_11 vccd1 vssd1 sky130_fd_sc_hd__decap_3
X_191_ vccd1 vssd1 _083_ _086_ sky130_fd_sc_hd__dlymetal6s2s_1
X_174_ vccd1 vssd1 _075_ _074_ _063_ sky130_fd_sc_hd__and2_1
X_226_ net21 clknet_2_3__leaf_clk _017_ vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1
X_157_ vssd1 vccd1 _011_ _062_ sky130_fd_sc_hd__clkbuf_1
X_209_ net28 clknet_2_3__leaf_clk _000_ vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1
XPHY_12 vccd1 vssd1 sky130_fd_sc_hd__decap_3
X_190_ _085_ _032_ _021_ _019_ vccd1 vssd1 sky130_fd_sc_hd__a21o_1
X_173_ vssd1 vccd1 _065_ _047_ net5 _074_ sky130_fd_sc_hd__mux2_1
X_225_ net20 clknet_2_3__leaf_clk _016_ vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1
X_156_ vccd1 vssd1 _062_ net11 _034_ sky130_fd_sc_hd__and2_1
X_139_ _045_ _047_ cnt_r\[5\] _050_ vccd1 vssd1 sky130_fd_sc_hd__a21o_1
X_208_ _086_ _079_ _034_ _087_ _031_ vssd1 vccd1 sky130_fd_sc_hd__a31o_1
Xclkbuf_2_3__f_clk clknet_2_3__leaf_clk clknet_0_clk vssd1 vccd1 sky130_fd_sc_hd__clkbuf_16
XPHY_13 vccd1 vssd1 sky130_fd_sc_hd__decap_3
X_241_ net42 clknet_2_1__leaf_clk _032_ vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1
X_172_ vssd1 vccd1 _015_ _073_ sky130_fd_sc_hd__clkbuf_1
X_224_ net19 clknet_2_3__leaf_clk _015_ vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1
X_155_ _060_ _061_ _010_ _058_ vccd1 vssd1 sky130_fd_sc_hd__a21oi_1
X_138_ vssd1 vccd1 _049_ cnt_r\[5\] _047_ _045_ sky130_fd_sc_hd__and3_1
X_207_ _086_ _079_ _091_ _085_ _030_ vssd1 vccd1 sky130_fd_sc_hd__a31o_1
XPHY_14 vccd1 vssd1 sky130_fd_sc_hd__decap_3
X_171_ vccd1 vssd1 _073_ _072_ _063_ sky130_fd_sc_hd__and2_1
X_240_ net41 clknet_2_1__leaf_clk _031_ vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1
X_223_ net18 clknet_2_3__leaf_clk _014_ vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1
X_154_ vssd1 vccd1 _055_ _053_ cnt_r\[8\] _061_ _037_ cnt_r\[9\] sky130_fd_sc_hd__a41o_1
X_137_ _005_ _047_ _048_ _045_ vssd1 vccd1 sky130_fd_sc_hd__o21a_1
X_206_ _086_ _032_ _091_ _082_ _029_ vssd1 vccd1 sky130_fd_sc_hd__a31o_1
XPHY_15 vccd1 vssd1 sky130_fd_sc_hd__decap_3
X_170_ vssd1 vccd1 _065_ cnt_r\[3\] net4 _072_ sky130_fd_sc_hd__mux2_1
X_153_ cnt_r\[9\] _060_ vccd1 vssd1 sky130_fd_sc_hd__inv_2
X_222_ net17 clknet_2_2__leaf_clk _013_ vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1
X_205_ _087_ _091_ _028_ _027_ vccd1 vssd1 sky130_fd_sc_hd__a21o_1
X_136_ _047_ _037_ _048_ _045_ vccd1 vssd1 sky130_fd_sc_hd__a21oi_1
X_119_ vssd1 vccd1 _000_ _035_ sky130_fd_sc_hd__clkbuf_1
XPHY_16 vccd1 vssd1 sky130_fd_sc_hd__decap_3
X_152_ vssd1 vccd1 _009_ _059_ sky130_fd_sc_hd__clkbuf_1
X_221_ net16 clknet_2_3__leaf_clk _012_ vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1
X_204_ _085_ _091_ _028_ _026_ vccd1 vssd1 sky130_fd_sc_hd__a21o_1
X_135_ vccd1 vssd1 cnt_r\[4\] _047_ sky130_fd_sc_hd__dlymetal6s2s_1
X_118_ vssd1 vccd1 _035_ _034_ sky130_fd_sc_hd__clkbuf_1
XPHY_17 vccd1 vssd1 sky130_fd_sc_hd__decap_3
X_220_ net14 clknet_2_3__leaf_clk _011_ vccd1 vssd1 sky130_fd_sc_hd__dfxtp_1
X_151_ vssd1 vccd1 _059_ _057_ _041_ _058_ sky130_fd_sc_hd__and3_1
X_203_ _082_ _091_ _028_ _025_ vccd1 vssd1 sky130_fd_sc_hd__a21o_1
X_134_ _004_ cnt_r\[3\] _046_ _040_ vssd1 vccd1 sky130_fd_sc_hd__o21a_1
X_117_ _033_ _034_ vssd1 vccd1 sky130_fd_sc_hd__clkbuf_2
XPHY_18 vccd1 vssd1 sky130_fd_sc_hd__decap_3
Xoutput50 vccd1 vssd1 msb_n[15] net50 sky130_fd_sc_hd__buf_2
X_150_ _058_ cnt_r\[8\] _053_ _055_ vssd1 vccd1 sky130_fd_sc_hd__nand3_1
X_133_ _045_ _046_ _037_ vssd1 vccd1 sky130_fd_sc_hd__nor2_1
X_202_ vssd1 vccd1 _028_ _092_ sky130_fd_sc_hd__clkbuf_1
X_116_ vccd1 vssd1 net12 _033_ sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_19 vccd1 vssd1 sky130_fd_sc_hd__decap_3
Xoutput51 vccd1 vssd1 msb_n[1] net51 sky130_fd_sc_hd__buf_2
Xoutput40 vccd1 vssd1 msb[6] net40 sky130_fd_sc_hd__buf_2
X_132_ vccd1 vssd1 _044_ _045_ sky130_fd_sc_hd__dlymetal6s2s_1
X_201_ _092_ _078_ _033_ _086_ vssd1 vccd1 sky130_fd_sc_hd__o21a_1
X_115_ net27 net21 vccd1 vssd1 sky130_fd_sc_hd__clkinv_2
Xoutput52 vccd1 vssd1 msb_n[2] net52 sky130_fd_sc_hd__buf_2
Xoutput41 vccd1 vssd1 msb[7] net41 sky130_fd_sc_hd__buf_2
Xoutput30 vccd1 vssd1 msb[11] net30 sky130_fd_sc_hd__buf_2
C43 _034_ vssd1 3.42fF
C44 _033_ vssd1 3.54fF
C45 _011_ vssd1 2.09fF
C46 _055_ vssd1 4.92fF
C47 clknet_2_3__leaf_clk vssd1 4.24fF
C48 clkbuf_2_3__f_clk/a_110_47# vssd1 2.12fF $ **FLOATING
C49 _065_ vssd1 4.34fF
C50 net28 vssd1 2.23fF
C51 vccd1 vssd1 824.63fF
C52 _020_ vssd1 3.56fF
C53 _041_ vssd1 4.07fF
C54 clkbuf_2_2__f_clk/a_110_47# vssd1 2.03fF $ **FLOATING
C55 net13 vssd1 2.50fF
C56 _023_ vssd1 2.24fF
C57 dac_in[8] vssd1 2.16fF
C58 _087_ vssd1 2.40fF
C59 _036_ vssd1 3.29fF
C60 net6 vssd1 2.30fF
C61 dac_in[5] vssd1 3.26fF
C62 cnt_r\[0\] vssd1 2.16fF
C63 cnt_r\[5\] vssd1 2.80fF
C64 clknet_2_1__leaf_clk vssd1 3.51fF
C65 clkbuf_2_1__f_clk/a_110_47# vssd1 2.09fF $ **FLOATING
C66 clknet_2_2__leaf_clk vssd1 2.40fF
C67 net34 vssd1 2.03fF
C68 _008_ vssd1 2.95fF
C69 cnt_r\[7\] vssd1 2.67fF
C70 _064_ vssd1 2.18fF
C71 clknet_0_clk vssd1 6.08fF
C72 clkbuf_2_0__f_clk/a_110_47# vssd1 2.06fF $ **FLOATING
C73 clkbuf_0_clk/a_110_47# vssd1 2.12fF $ **FLOATING
C74 cnt_r\[2\] vssd1 3.78fF
C75 _078_ vssd1 2.45fF
C76 clk vssd1 2.30fF
C77 _021_ vssd1 3.11fF
C78 _085_ vssd1 2.80fF
C79 _037_ vssd1 12.45fF
.ends



XDUT clk dac_in[0] dac_in[1] dac_in[2] dac_in[3] dac_in[4] dac_in[5] dac_in[6]  dac_in[7] dac_in[8]
+ dac_in[9] dummy llsb llsb_n lsb[0] lsb[1] lsb[2] lsb[3] lsb[4]  lsb[5] lsb_n[0] lsb_n[1] lsb_n[2] lsb_n[3]
+ lsb_n[4] lsb_n[5] msb[0] msb[10] msb[11]  msb[12] msb[13] msb[14] msb[15] msb[1] msb[2] msb[3] msb[4] msb[5]
+ msb[6] msb[7]  msb[8] msb[9] msb_n[0] msb_n[10] msb_n[11] msb_n[12] msb_n[13] msb_n[14] msb_n[15]
+  msb_n[1] msb_n[2] msb_n[3] msb_n[4] msb_n[5] msb_n[6] msb_n[7] msb_n[8] msb_n[9]  rst_n test_mode vccd1
+ vssd1 dac_con


**** end user architecture code
.ends

.GLOBAL GND
.end
