* NGSPICE file created from dac_con_flat.ext - technology: sky130A

.subckt dac_con_flat clk dac_in[0] dac_in[1] dac_in[2] dac_in[3] dac_in[4] dac_in[5]
+ dac_in[6] dac_in[7] dac_in[8] dac_in[9] dummy llsb llsb_n lsb[0] lsb[1] lsb[2] lsb[3]
+ lsb[4] lsb[5] lsb_n[0] lsb_n[1] lsb_n[2] lsb_n[3] lsb_n[4] lsb_n[5] msb[0] msb[10]
+ msb[11] msb[12] msb[13] msb[14] msb[15] msb[1] msb[2] msb[3] msb[4] msb[5] msb[6]
+ msb[7] msb[8] msb[9] msb_n[0] msb_n[10] msb_n[11] msb_n[12] msb_n[13] msb_n[14]
+ msb_n[15] msb_n[1] msb_n[2] msb_n[3] msb_n[4] msb_n[5] msb_n[6] msb_n[7] msb_n[8]
+ msb_n[9] rst_n test_mode vccd1 vssd1
X0 a_12627_4649# _196_.A a_12409_4373# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_4894_4373# a_4694_4673# a_5043_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2 vccd1 _133_.Y a_31480_3561# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=2.99018e+14p pd=2.87785e+09u as=0p ps=0u w=1e+06u l=150000u
X3 a_7624_7093# output46.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 a_31589_4221# _125_.A2 a_31517_4221# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 _094_.Y output28.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 _148_.B1 _133_.A a_3063_2473# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 vssd1 a_16180_3285# _208_.X vssd1 sky130_fd_pr__nfet_01v8 ad=1.91416e+14p pd=2.07373e+09u as=0p ps=0u w=650000u l=150000u
X8 a_22369_4943# _235_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X10 a_20131_2375# a_20227_2197# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 output23.A output17.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 output15.A _093_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X14 vccd1 a_5600_7093# msb[13] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X15 vssd1 a_13445_2375# _203_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_27422_4765# a_27149_4399# a_27337_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 vccd1 a_17911_4943# a_18079_4917# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_16507_4399# a_16378_4673# a_16087_4373# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X19 vssd1 output41.A a_15299_7127# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 a_8079_5309# a_7859_5321# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X22 vccd1 a_4687_4373# a_4694_4673# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X23 vccd1 _209_.CLK a_28547_3861# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X24 vccd1 a_14894_2335# a_14821_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 vssd1 a_15319_2491# a_15277_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 a_5967_5461# a_6251_5461# a_6186_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X27 a_36783_5162# _163_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X28 a_28389_3339# _162_.A a_28303_3339# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 vccd1 _177_.B a_25635_3105# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X31 _164_.A0 a_34159_2223# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X32 a_28423_2999# _171_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X33 a_2511_2767# _149_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X35 vssd1 _160_.X a_27684_3133# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X36 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X37 vccd1 output29.A a_10147_7127# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X38 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X39 a_35249_4399# _169_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X40 vccd1 _129_.X a_25787_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X41 a_33478_4511# a_33310_4765# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X42 a_5241_4399# a_4687_4373# a_4894_4373# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X43 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X44 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X45 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X46 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X47 a_16087_4373# a_16378_4673# a_16329_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X48 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X49 a_10483_5175# _196_.A a_10657_5281# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X50 a_21454_4373# a_21247_4373# a_21630_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X51 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X52 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X53 a_17995_4943# a_17213_4949# a_17911_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X54 vssd1 a_13327_4373# _193_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X55 a_14821_2589# a_14287_2223# a_14726_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X56 a_15098_3677# a_14851_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X57 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X58 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X59 a_35437_4175# ANTENNA__118__A.DIODE _125_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X60 a_33386_3829# a_33218_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X61 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X62 msb[13] a_5600_7093# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X63 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X64 a_22069_2741# _215_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X65 a_14851_3311# a_14722_3585# a_14431_3285# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X66 vccd1 _180_.B a_15147_4427# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X67 vssd1 _159_.X a_20769_2806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X68 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X69 a_6725_2223# a_6559_2223# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X70 a_7534_2741# a_7366_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X71 vssd1 a_23478_3855# _209_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X72 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X73 vccd1 dac_in[0] a_36091_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X74 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X75 _160_.X a_19623_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X76 output23.A output17.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X77 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X78 a_33037_4399# a_32871_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X79 _128_.B1 a_27463_3579# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X80 _155_.B1 a_2869_3087# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X81 _232_.CLK a_13069_3829# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X82 a_26300_6549# _094_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X83 vccd1 a_34944_2375# _168_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X84 _183_.A1 a_9799_2741# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X85 _133_.A _121_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X86 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X87 a_21630_4765# a_21383_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X88 a_35334_4765# a_34895_4399# a_35249_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X89 vccd1 ANTENNA__177__A.DIODE a_19106_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X90 a_35307_2223# input3.X a_34944_2375# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X91 vccd1 output19.A output25.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X92 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X93 vccd1 a_29154_3829# a_29081_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X94 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X95 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X96 a_10936_7093# output59.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X97 a_14115_5321# a_13979_5161# a_13695_5175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X98 vccd1 a_4307_4551# output30.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X99 a_17965_4649# _205_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X100 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X101 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X102 vssd1 a_10943_4373# a_10950_4673# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X103 vccd1 a_27590_4511# a_27517_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X104 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X105 msb[10] a_10147_7127# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X106 vccd1 output41.A output57.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X107 a_25030_2589# a_24591_2223# a_24945_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X108 clkbuf_2_3__f_clk.A a_20442_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X109 vccd1 a_22983_2375# _140_.A_N vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X110 vssd1 a_23478_2767# _222_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X111 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X112 a_17486_4943# a_17047_4949# a_17401_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X113 a_4894_4373# a_4687_4373# a_5070_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X114 a_30550_3311# a_30373_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X115 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X116 a_25539_2589# a_24757_2223# a_25455_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X117 _209_.CLK a_23478_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X118 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X119 a_33309_3145# a_32319_2773# a_33183_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X120 a_36417_2806# input1.X a_36203_2806# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X121 vccd1 a_16911_2986# _183_.A0 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X122 _233_.CLK a_13069_2741# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X123 clkbuf_2_3__f_clk.A a_20442_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X124 a_26300_6549# _094_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X125 vccd1 a_15151_2589# a_15319_2491# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X126 a_29081_3855# a_28547_3861# a_28986_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X127 a_23005_5321# a_22015_4949# a_22879_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X128 vssd1 _134_.X a_31369_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X129 a_15398_3894# _159_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X130 a_35460_4399# a_35061_4399# a_35334_4765# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X131 vccd1 output20.A a_31215_7127# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X132 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X133 a_15269_3311# a_14715_3285# a_14922_3285# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X134 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X135 vssd1 _149_.A2 a_8296_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X136 a_15269_3311# a_14722_3585# a_14922_3285# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X137 vssd1 a_28142_4917# a_28100_5321# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X138 a_28107_2550# input4.X a_28107_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X139 _232_.CLK a_13069_3829# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X140 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X141 a_21801_4399# a_21254_4673# a_21454_4373# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X142 a_21182_4399# a_20867_4551# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X143 a_18015_2806# _144_.A1 a_17556_2999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X144 a_4772_7093# output48.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X145 a_5070_4765# a_4823_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X146 vssd1 a_20867_4551# output38.A vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X147 a_25156_2223# a_24757_2223# a_25030_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X148 vssd1 a_8307_7127# msb[11] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X149 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X150 vccd1 a_9631_2767# a_9799_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X151 a_16403_3311# _206_.A2 a_16309_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X152 vccd1 a_22069_2741# _140_.C vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X153 vccd1 a_7539_4073# a_7546_3977# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X154 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X155 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X156 a_17612_5321# a_17213_4949# a_17486_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X157 a_22983_2375# _135_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X158 _222_.CLK a_23478_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X159 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X160 vccd1 _121_.A _133_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X161 a_7675_4233# a_7546_3977# a_7255_4087# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X162 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
D0 vssd1 _133_.A sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
X163 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X164 vccd1 a_29801_2999# a_29614_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X165 _159_.A a_1591_2223# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X166 vssd1 a_14563_7127# msb_n[7] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X167 vccd1 a_15991_4551# output40.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X168 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X169 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X170 _114_.Y output20.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X171 a_11762_4087# a_11858_3829# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X172 a_37703_4564# _157_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X173 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X174 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X175 vccd1 a_22067_2197# _137_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
D1 vssd1 dac_in[5] sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
X176 a_21023_2806# input6.X a_21023_3133# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X177 vccd1 clkbuf_2_3__f_clk.A a_13069_3829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X178 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X179 vccd1 a_29796_7093# lsb_n[4] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X180 vccd1 a_13069_2741# _233_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X181 a_16180_3285# _180_.X a_16309_3561# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X182 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X183 vssd1 a_36236_6549# lsb_n[0] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X184 _136_.Y _133_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X185 vssd1 a_25198_2335# a_25156_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X186 output50.A output34.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X187 a_7791_2767# a_6927_2773# a_7534_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X188 vssd1 a_13979_5161# a_13986_5065# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X189 a_31022_2197# a_30815_2197# a_31198_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X190 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X191 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X192 _235_.D a_20070_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X193 a_35007_2806# _125_.A2 a_34935_2806# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X194 vssd1 a_7534_2741# a_7492_3145# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X195 a_23431_3677# a_22733_3311# a_23174_3423# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X196 vssd1 _172_.A a_26431_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X197 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X198 a_7331_3677# a_6633_3311# a_7074_3423# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X199 vssd1 _196_.B a_12160_5263# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X200 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X201 msb[3] a_22804_7093# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X202 lsb[4] a_31215_7127# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
D2 vssd1 rst_n sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
X203 vssd1 a_26063_7127# msb[1] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X204 vccd1 _133_.A a_30469_4649# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X205 _205_.A1 a_19106_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X206 lsb_n[4] a_29796_7093# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X207 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X208 vssd1 _196_.A a_7081_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X209 vccd1 _135_.A a_17743_2197# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X210 a_33225_4399# _157_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X211 vccd1 a_14186_5220# a_14115_5321# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X212 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X213 a_31171_2223# a_30951_2223# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X214 vssd1 a_13069_3829# _232_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X215 vccd1 _203_.A2 a_19257_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X216 vccd1 ANTENNA__177__A.DIODE a_27215_4087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X217 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X218 vssd1 a_33108_7093# lsb_n[2] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X219 output48.A output32.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X220 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X221 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X222 vccd1 a_32747_5161# a_32754_5065# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X223 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X224 a_20446_2223# a_20131_2375# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X225 vssd1 a_38023_6039# llsb vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X226 a_7166_2335# a_6998_2589# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X227 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X228 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X229 a_16911_2986# dac_in[7] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X230 vssd1 a_15151_2589# a_15319_2491# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X231 vssd1 _209_.CLK a_27535_4949# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X232 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X233 a_13069_3829# clkbuf_2_3__f_clk.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X234 msb[7] a_15299_7127# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X235 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X236 a_5687_3463# ANTENNA__177__A.DIODE a_5921_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X237 output53.A output37.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X238 vccd1 _162_.B a_36399_4193# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X239 a_27956_7093# _115_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X240 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X241 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X242 a_29801_2999# _133_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X243 vssd1 _159_.X a_10465_3894# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X244 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X245 a_36783_5162# _163_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X246 a_33643_3855# a_32945_3861# a_33386_3829# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X247 a_31022_2197# a_30822_2497# a_31171_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X248 vccd1 output17.A output23.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X249 vccd1 _093_.A output15.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X250 vccd1 _201_.X a_19439_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X251 vssd1 a_17192_7093# msb[6] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X252 clkbuf_2_3__f_clk.A a_20442_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X253 vssd1 a_35631_7127# lsb[1] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X254 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X255 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X256 a_26870_3677# a_26431_3311# a_26785_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X257 vccd1 a_33844_7093# lsb[2] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X258 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X259 vssd1 a_25226_3285# a_25155_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X260 a_22921_3311# _141_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X261 a_6821_3311# _190_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X262 _209_.CLK a_23478_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X263 _209_.CLK a_23478_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X264 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X265 a_20442_3311# clk vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X266 a_35843_4765# a_35061_4399# a_35759_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X267 a_24757_2223# a_24591_2223# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X268 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X269 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X270 vssd1 _152_.A a_5823_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X271 vssd1 a_23478_2767# _222_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X272 vssd1 a_10839_2999# _198_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X273 a_7281_2767# _152_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X274 a_27463_2806# _173_.A0 a_27463_3133# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X275 a_32942_3677# a_32669_3311# a_32857_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X276 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X277 vssd1 _222_.CLK a_24591_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X278 msb[0] a_27220_7093# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X279 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X280 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X281 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X282 vssd1 a_9799_2741# a_9757_3145# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X283 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X284 a_31463_3133# _134_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X285 vccd1 output30.A a_8307_7127# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X286 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X287 vccd1 a_30435_2375# _134_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X288 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X289 a_17213_4949# a_17047_4949# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X290 a_8999_4074# _199_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X291 a_19885_3855# a_19708_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X292 a_31665_3133# _211_.Q a_31559_3133# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X293 vssd1 a_15991_4551# output40.A vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X294 a_27295_3677# a_26431_3311# a_27038_3423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X295 output19.A a_28015_4667# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X296 _211_.Q a_33351_2741# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X297 vccd1 a_13069_3829# _232_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X298 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X299 a_26996_3311# a_26597_3311# a_26870_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X300 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X301 vssd1 a_17192_3285# _239_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X302 vccd1 a_10483_5175# _195_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X303 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X304 a_8933_2773# a_8767_2773# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X305 vccd1 clkbuf_2_3__f_clk.A a_23478_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X306 vssd1 dac_in[0] a_36091_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X307 _155_.A1 _179_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X308 a_27391_2806# a_27209_2806# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X309 vssd1 a_14335_3463# output41.A vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X310 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X311 a_24735_3285# a_25019_3285# a_24954_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X312 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X313 a_28901_3855# _225_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X314 vccd1 _233_.CLK a_6559_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X315 vssd1 a_30815_2197# a_30822_2497# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X316 vssd1 _121_.A _133_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X317 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X318 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X319 _125_.A1 a_30054_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X320 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X321 a_20227_2197# a_20511_2197# a_20446_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X322 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X323 a_36599_3476# _166_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X324 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X325 vccd1 a_1644_6549# msb_n[15] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X326 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X327 _149_.B1 a_7959_2741# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X328 vssd1 a_33535_3579# a_33493_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X329 lsb[5] a_28784_6549# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X330 vssd1 a_22067_2197# _137_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X331 vccd1 a_13069_2741# _233_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X332 vssd1 a_37839_6575# llsb_n vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X333 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X334 _165_.B a_35007_2806# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X335 a_2585_3311# _149_.A1 a_2501_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X336 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X337 _222_.CLK a_23478_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X338 vccd1 _162_.A a_19793_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X339 a_28525_5321# a_27535_4949# a_28399_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X340 a_31307_3311# _126_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X341 a_10933_3894# _185_.A0 a_10719_3894# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X342 vccd1 _196_.A a_10483_5175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X343 a_17321_3311# _196_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X344 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X345 vssd1 a_20442_3311# clkbuf_2_3__f_clk.A vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X346 a_6251_5461# _232_.CLK vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X347 a_10003_3638# a_9821_3638# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X348 vccd1 a_6527_4373# a_6534_4673# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X349 vccd1 dac_in[2] a_29743_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X350 _180_.A a_11746_2223# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X351 msb[11] a_8307_7127# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X352 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X353 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X354 vssd1 _232_.D a_6805_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X355 a_34948_7093# output23.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X356 a_27847_4765# a_27149_4399# a_27590_4511# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X357 a_24639_3463# a_24735_3285# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X358 a_22454_4943# a_22181_4949# a_22369_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X359 _196_.B a_15242_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X360 vccd1 a_13599_5175# output42.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X361 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X362 a_25155_3311# a_25019_3285# a_24735_3285# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X363 a_7081_4399# a_6527_4373# a_6734_4373# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X364 vssd1 _159_.A a_14287_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X365 vccd1 a_26479_2388# input6.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X366 vssd1 a_32922_2375# a_32871_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X367 a_23006_3677# a_22567_3311# a_22921_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X368 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X369 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X370 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X371 vccd1 a_27463_3579# a_27379_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X372 _125_.Y _125_.A1 a_34702_4175# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X373 vccd1 a_7723_5161# a_7730_5065# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X374 a_25030_4765# a_24757_4399# a_24945_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X375 a_2511_2767# _179_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X376 a_23478_3855# clkbuf_2_3__f_clk.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X377 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X378 a_27038_3423# a_26870_3677# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X379 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X380 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X381 output20.A a_29579_3829# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X382 a_15398_4221# _159_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X383 a_20253_2767# a_20076_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X384 output35.A a_25623_4667# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X385 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X386 vssd1 _205_.B1 a_19426_5263# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
D3 vssd1 _133_.A sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
X387 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X388 msb_n[2] a_23540_7093# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X389 _133_.A _121_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X390 vccd1 a_4036_7093# msb[14] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X391 a_28871_4564# _178_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X392 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X393 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X394 a_25019_3285# _222_.CLK vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X395 vccd1 a_5687_3463# _152_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X396 vccd1 output17.A a_35631_7127# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X397 a_12242_2223# a_12065_2223# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X398 a_3697_2767# _149_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X399 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X400 vccd1 a_11863_5639# _196_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X401 vccd1 output41.A output57.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X402 a_23132_3311# a_22733_3311# a_23006_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X403 clkbuf_2_3__f_clk.A a_20442_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X404 a_18416_3561# _180_.A a_18243_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X405 a_7032_3311# a_6633_3311# a_6906_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X406 vssd1 output36.A a_24591_7127# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X407 vccd1 output20.A _114_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X408 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X409 vccd1 a_14922_3285# a_14851_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X410 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X411 a_30833_3311# a_30656_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X412 msb[14] a_4036_7093# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X413 _233_.CLK a_13069_2741# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X414 a_2593_3087# _145_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X415 vccd1 a_6147_4551# output31.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X416 a_10839_2999# _121_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X417 a_23935_2223# _135_.X _136_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X418 vccd1 a_25198_4511# a_25125_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X419 a_26785_3311# _130_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X420 clkbuf_2_3__f_clk.A a_20442_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X421 a_33218_3855# a_32779_3861# a_33133_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X422 llsb a_38023_6039# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X423 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
D4 vssd1 dac_in[0] sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
X424 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X425 a_19257_4943# _205_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X426 vccd1 a_31267_2741# _131_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X427 vccd1 _126_.X a_27488_4087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X428 vssd1 _129_.X a_25787_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X429 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X430 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X431 output35.A a_25623_4667# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X432 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X433 vccd1 a_22622_4917# a_22549_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X434 a_9374_2741# a_9206_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X435 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X436 a_17415_3311# _206_.A2 a_17321_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X437 _232_.CLK a_13069_3829# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X438 a_18785_2767# _144_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X439 vccd1 a_8999_4074# _199_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X440 vssd1 a_10936_7093# msb_n[9] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X441 a_6607_5487# a_6387_5487# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X442 vssd1 a_23174_3423# a_23132_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X443 vssd1 a_7074_3423# a_7032_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X444 vccd1 _126_.A a_31267_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X445 a_19970_2767# a_19793_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X446 a_15738_2767# a_15561_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X447 vccd1 _193_.X a_5241_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X448 vssd1 _159_.A a_10296_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X449 _157_.A a_37503_4193# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X450 vccd1 _222_.CLK a_26431_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X451 a_13630_4649# _205_.A2 a_13327_4373# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X452 _222_.CLK a_23478_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X453 msb_n[0] a_26300_6549# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
D5 vssd1 dummy sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
X454 vssd1 output32.A output48.A vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X455 a_25125_4765# a_24591_4399# a_25030_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X456 a_34944_2375# _128_.B1 a_35086_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X457 vssd1 a_7159_4087# output34.A vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X458 msb[6] a_17192_7093# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X459 a_21237_2806# input6.X a_21023_2806# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X460 _122_.Y _133_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X461 a_33344_4233# a_32945_3861# a_33218_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X462 a_10563_4551# a_10659_4373# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X463 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X464 a_12627_4649# _203_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X465 vssd1 a_9655_4087# _199_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X466 a_17192_3285# _180_.X a_17321_3561# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X467 vccd1 clkbuf_2_3__f_clk.A a_13069_3829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X468 vssd1 a_20504_7093# msb[4] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X469 a_32945_3861# a_32779_3861# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X470 a_6458_5461# a_6258_5761# a_6607_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X471 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X472 a_20260_5263# _205_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X473 vccd1 clk a_20442_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X474 vccd1 _125_.A2 a_34619_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X475 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X476 vssd1 _201_.X a_19439_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X477 vccd1 a_33735_4765# a_33903_4667# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X478 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X479 vccd1 _209_.CLK a_22015_4949# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X480 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X481 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X482 vccd1 a_30441_3829# _128_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X483 vssd1 _160_.X a_35228_3133# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X484 a_9655_4087# _198_.A a_9829_4193# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X485 vssd1 ANTENNA__118__A.DIODE a_37011_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X486 _171_.B a_28107_2550# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X487 vssd1 a_23478_3855# _209_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X488 a_33844_7093# output18.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X489 vccd1 a_33478_4511# a_33405_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X490 vssd1 a_16911_2986# _183_.A0 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X491 a_7681_4943# a_7343_5175# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X492 vccd1 _141_.A a_22659_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X493 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X494 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X495 _222_.CLK a_23478_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X496 a_36203_3133# a_35949_2806# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X497 a_6805_5487# a_6251_5461# a_6458_5461# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X498 _115_.A a_28567_4917# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X499 vccd1 _239_.D a_16925_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X500 a_33451_3677# a_32669_3311# a_33367_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X501 vssd1 a_16915_2197# ANTENNA__118__A.DIODE vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
D6 vssd1 ANTENNA__118__A.DIODE sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
X502 vccd1 _134_.X a_31369_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X503 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X504 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X505 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X506 a_27422_4765# a_26983_4399# a_27337_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X507 _174_.X a_28303_3339# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X508 a_22733_3311# a_22567_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X509 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X510 a_23217_2223# _215_.Q a_23145_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X511 vssd1 _133_.B a_22372_3087# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X512 vssd1 a_33367_3677# a_33535_3579# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X513 vccd1 _174_.B a_28303_3339# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X514 a_6633_3311# a_6467_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X515 _232_.CLK a_13069_3829# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X516 a_33405_4765# a_32871_4399# a_33310_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X517 llsb_n a_37839_6575# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X518 vssd1 a_33735_4765# a_33903_4667# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X519 vssd1 a_13069_2741# _233_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X520 vccd1 a_29579_3829# a_29495_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X521 a_17928_7093# output55.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X522 vccd1 a_29055_2388# input4.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X523 vccd1 _180_.A a_19474_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X524 output48.A output32.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X525 vssd1 output39.A output55.A vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X526 clkbuf_2_3__f_clk.A a_20442_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X527 a_18751_2388# dac_in[6] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X528 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X529 a_36599_3476# _166_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X530 a_21247_4373# _209_.CLK vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X531 _222_.CLK a_23478_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X532 vssd1 a_32926_2741# a_32884_3145# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X533 _233_.CLK a_13069_2741# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X534 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X535 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X536 a_27548_4399# a_27149_4399# a_27422_4765# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X537 vssd1 _209_.CLK a_28547_3861# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X538 msb_n[3] a_22068_7093# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X539 vccd1 a_5871_5639# output33.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X540 a_20070_4399# _205_.A1 a_19984_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X541 vssd1 a_23478_2767# _222_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X542 a_35885_4399# a_34895_4399# a_35759_4765# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X543 _203_.X a_19426_5263# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X544 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X545 vssd1 _205_.B1 a_21801_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X546 a_12794_3311# a_12617_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X547 vccd1 a_11150_4373# a_11079_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X548 _133_.Y _133_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X549 _215_.Q a_23599_3579# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X550 output29.A a_7499_3579# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X551 vssd1 output39.A a_18611_7127# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X552 msb_n[14] a_3116_6549# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X553 vccd1 a_12242_2767# a_12348_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X554 a_21023_3133# a_20769_2806# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X555 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X556 a_9121_2767# _217_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X557 _162_.B a_36203_2806# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X558 vccd1 a_15727_5175# _205_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X559 a_14453_2223# a_14287_2223# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X560 vssd1 a_26479_2388# input6.X vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X561 msb_n[8] a_12999_6575# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X562 _201_.X a_18416_3561# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X563 vccd1 a_33524_2375# _125_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X564 vccd1 _206_.A2 a_13630_4649# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X565 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X566 a_7439_5175# a_7723_5161# a_7658_5309# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X567 a_17401_4943# _238_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X568 a_20131_2375# a_20227_2197# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X569 a_12364_4087# _180_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X570 a_11506_3311# a_11329_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X571 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X572 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X573 vccd1 clkbuf_2_3__f_clk.A a_23478_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X574 vssd1 a_27590_4511# a_27548_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X575 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X576 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X577 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X578 msb[2] a_24591_7127# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X579 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X580 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X581 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X582 _232_.D a_2695_4399# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X583 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X584 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X585 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X586 a_9631_2767# a_8933_2773# a_9374_2741# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X587 a_33037_3677# a_32503_3311# a_32942_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X588 vccd1 output42.A a_13459_7127# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X589 vccd1 a_30120_2999# _133_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X590 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X591 a_35502_4511# a_35334_4765# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X592 vssd1 _183_.X a_15242_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X593 output46.A output30.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X594 a_13069_2741# clkbuf_2_3__f_clk.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X595 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X596 vssd1 _160_.X a_34753_2806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X597 vccd1 a_17762_3855# a_17868_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X598 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X599 _102_.Y output42.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X600 _115_.Y _115_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X601 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X602 vssd1 a_32367_5175# output28.A vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X603 a_20511_2197# _222_.CLK vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X604 output57.A output41.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X605 vccd1 a_20442_3311# clkbuf_2_3__f_clk.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X606 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X607 a_30744_4175# _125_.A1 a_30441_3829# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X608 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X609 _145_.Y _145_.B a_13649_3561# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X610 vccd1 a_28142_4917# a_28069_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X611 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X612 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X613 vccd1 _149_.X a_5687_3463# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X614 msb_n[9] a_10936_7093# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X615 _173_.A0 a_26431_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X616 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X617 msb_n[11] a_7624_7093# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X618 a_32673_2767# _125_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X619 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X620 _162_.A a_19474_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X621 a_22921_3311# _141_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X622 vccd1 a_20442_3311# clkbuf_2_3__f_clk.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X623 a_6821_3311# _190_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X624 a_21603_4399# a_21383_4399# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X625 vccd1 a_38163_2388# _156_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X626 vccd1 a_11987_7127# msb[9] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X627 a_37519_5162# _119_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X628 a_10878_4399# a_10563_4551# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X629 vccd1 a_23478_2767# _222_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X630 a_12525_2767# a_12348_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X631 vssd1 a_7993_4373# _149_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X632 output51.A output35.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X633 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X634 vssd1 a_13069_3829# _232_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X635 msb[15] a_2288_7093# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X636 a_17192_7093# output40.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X637 vssd1 a_35927_4667# a_35885_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X638 lsb_n[2] a_33108_7093# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X639 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X640 vssd1 a_14287_4399# _159_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X641 _133_.A _121_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X642 a_30659_3855# _128_.B1 a_30441_3829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X643 vssd1 a_7539_4073# a_7546_3977# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X644 a_27684_3133# _135_.X a_27463_2806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X645 a_6387_5487# a_6258_5761# a_5967_5461# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X646 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X647 a_27337_4399# _224_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X648 vssd1 a_13069_2741# _233_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X649 a_31389_3561# _134_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X650 a_7255_4087# a_7546_3977# a_7497_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X651 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X652 vssd1 a_5871_5639# output33.A vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X653 a_21454_4373# a_21254_4673# a_21603_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X654 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X655 vssd1 a_25623_2491# a_25581_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X656 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X657 _179_.A1 a_7591_2491# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X658 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X659 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X660 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X661 msb_n[1] a_25380_7093# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X662 _211_.Q a_33351_2741# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X663 vssd1 a_7959_2741# a_7917_3145# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X664 vccd1 _144_.A1 a_17743_2197# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X665 a_20718_2197# a_20511_2197# a_20894_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X666 a_32922_2375# a_33018_2197# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X667 vssd1 a_37703_4564# _157_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X668 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X669 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
D7 vssd1 ANTENNA__177__A.DIODE sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
X670 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X671 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X672 a_20442_3311# clk vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X673 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X674 vssd1 a_15738_2767# a_15844_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X675 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X676 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X677 a_25198_4511# a_25030_4765# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X678 vccd1 a_13069_3829# _232_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X679 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X680 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X681 a_12160_5263# _241_.D a_11857_4917# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X682 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X683 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X684 vssd1 a_11857_4917# _190_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X685 a_29518_2999# a_29614_2741# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X686 _233_.CLK a_13069_2741# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X687 a_21801_4399# a_21247_4373# a_21454_4373# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X688 a_20867_2223# a_20647_2223# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X689 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X690 a_27463_2806# _135_.X a_27391_2806# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X691 _163_.A a_36399_4193# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X692 vssd1 a_22804_7093# msb[3] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X693 vccd1 a_15319_2491# a_15235_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X694 _128_.B1 a_27463_3579# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
D8 vssd1 dac_in[4] sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
X695 a_20894_2589# a_20647_2223# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X696 a_14894_2335# a_14726_2589# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X697 vssd1 _208_.X a_15269_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X698 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X699 a_14894_2335# a_14726_2589# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X700 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X701 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X702 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X703 msb_n[6] a_16088_7093# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X704 a_27365_4215# _128_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X705 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X706 vccd1 _206_.A2 a_17965_4649# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X707 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X708 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X709 vssd1 a_32747_5161# a_32754_5065# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X710 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X711 vccd1 a_23478_3855# _209_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X712 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X713 _180_.X a_15147_4427# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X714 vccd1 _196_.A a_7081_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X715 vssd1 output38.A _098_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X716 a_16915_2197# _180_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X717 a_24945_4399# _203_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X718 a_20718_2197# a_20518_2497# a_20867_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X719 vccd1 ANTENNA__118__A.DIODE _145_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X720 a_10659_4373# a_10943_4373# a_10878_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X721 a_12075_4943# _196_.A a_11857_4917# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X722 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X723 _233_.CLK a_13069_2741# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X724 vccd1 _198_.A a_9655_4087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X725 vssd1 a_29055_2388# input4.X vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X726 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X727 a_28107_2550# _134_.A1 a_28035_2550# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X728 a_33108_7093# output24.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X729 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X730 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X731 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X732 _232_.CLK a_13069_3829# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X733 vssd1 a_26300_6549# msb_n[0] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X734 msb_n[13] a_4772_7093# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X735 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X736 vccd1 a_20867_4551# output38.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X737 _206_.A2 a_12298_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X738 a_18751_2388# dac_in[6] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X739 vssd1 a_20442_3311# clkbuf_2_3__f_clk.A vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X740 msb[5] a_18611_7127# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X741 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X742 a_28107_2223# a_27853_2550# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X743 a_9206_2767# a_8767_2773# a_9121_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X744 a_22068_7093# output53.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X745 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X746 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X747 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X748 vssd1 _205_.B1 a_20070_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X749 a_5357_2767# _151_.C vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X750 vccd1 a_31022_2197# a_30951_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X751 a_14922_3285# a_14715_3285# a_15098_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X752 vssd1 a_23478_3855# _209_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X753 vssd1 a_15299_7127# msb[7] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X754 a_6428_6549# _106_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X755 vccd1 a_13069_2741# _233_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X756 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X757 a_22879_4943# a_22015_4949# a_22622_4917# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X758 _222_.CLK a_23478_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X759 vccd1 a_28015_4667# a_27931_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X760 a_33478_4511# a_33310_4765# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X761 a_13445_2375# _192_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X762 a_26785_3311# _130_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X763 vccd1 a_33205_2375# a_33018_2197# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
D9 vssd1 dac_in[1] sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
X764 a_12045_4087# ANTENNA__177__A.DIODE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X765 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X766 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X767 a_25455_4765# a_24591_4399# a_25198_4511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X768 vccd1 _233_.CLK a_14287_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X769 _196_.A a_11010_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X770 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X771 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X772 vssd1 a_23478_3855# _209_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X773 a_37703_4564# _157_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X774 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X775 vccd1 a_20890_3855# a_20996_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X776 vssd1 a_8999_4074# _199_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X777 a_15071_3311# a_14851_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X778 _108_.Y output33.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X779 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X780 a_17486_4943# a_17213_4949# a_17401_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X781 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X782 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X783 vssd1 _159_.X a_19623_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X784 a_9332_3145# a_8933_2773# a_9206_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X785 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X786 a_16309_3561# ANTENNA__118__A.DIODE vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X787 vccd1 a_11762_4087# a_11711_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X788 vssd1 a_9738_2375# a_9687_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X789 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X790 vssd1 a_13599_5175# output42.A vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X791 vccd1 _135_.X a_22370_2473# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X792 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X793 a_6428_6549# _106_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X794 vccd1 output30.A output46.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X795 a_23478_3855# clkbuf_2_3__f_clk.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X796 vccd1 a_16371_4373# a_16378_4673# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X797 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X798 a_5849_3311# _151_.C vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X799 vccd1 output25.A a_31767_6575# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X800 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X801 a_8933_2773# a_8767_2773# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X802 vssd1 a_4687_4373# a_4694_4673# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X803 a_23557_3311# a_22567_3311# a_23431_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X804 a_7457_3311# a_6467_3311# a_7331_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X805 a_18037_5321# a_17047_4949# a_17911_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X806 vccd1 _160_.X a_36417_2806# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X807 _222_.CLK a_23478_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X808 a_35841_3339# _162_.A a_35755_3339# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X809 a_7534_2741# a_7366_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X810 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X811 _145_.B _140_.A_N a_18785_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X812 vccd1 a_27956_7093# lsb_n[5] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X813 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X814 vccd1 a_36599_3476# _166_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X815 vssd1 _125_.A1 a_30373_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X816 a_14922_3285# a_14722_3585# a_15071_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X817 a_31355_4087# _126_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X818 a_15256_4087# _183_.A0 a_15398_3894# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X819 vssd1 clkbuf_2_3__f_clk.A a_13069_2741# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X820 a_31480_3561# _126_.X a_31389_3561# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X821 vssd1 _133_.A _148_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X822 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X823 vccd1 output42.A _102_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X824 a_32463_5175# a_32754_5065# a_32705_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X825 _125_.Y _125_.B1 a_34619_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X826 vssd1 _125_.A2 a_30744_4175# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X827 a_6998_2589# a_6559_2223# a_6913_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X828 a_37589_4193# ANTENNA__118__A.DIODE a_37503_4193# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X829 a_37519_5162# _119_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X830 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X831 a_23006_3677# a_22733_3311# a_22921_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X832 a_6906_3677# a_6633_3311# a_6821_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X833 vssd1 output25.A a_31767_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X834 msb[12] a_6835_7127# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X835 vssd1 a_17928_7093# msb_n[5] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X836 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X837 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X838 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X839 vssd1 a_12364_4087# ANTENNA__177__A.DIODE vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X840 a_4645_4765# a_4307_4551# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X841 vccd1 _209_.CLK a_26983_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X842 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X843 vccd1 a_25623_4667# a_25539_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X844 vccd1 a_32319_7127# lsb[3] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X845 vssd1 a_38163_2388# _156_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X846 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X847 ANTENNA__118__A.DIODE a_16915_2197# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X848 a_32669_3311# a_32503_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X849 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X850 vccd1 _196_.A a_11863_5639# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X851 a_33037_4399# a_32871_4399# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X852 a_20504_7093# output38.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X853 a_33735_4765# a_32871_4399# a_33478_4511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X854 vccd1 a_14335_3463# output41.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X855 a_2288_7093# output34.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X856 vssd1 a_25455_2589# a_25623_2491# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X857 vccd1 a_17654_4917# a_17581_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X858 a_11789_3311# a_11612_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X859 a_33769_4233# a_32779_3861# a_33643_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X860 vssd1 a_7723_5161# a_7730_5065# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X861 a_20963_4373# a_21254_4673# a_21205_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X862 a_21383_4399# a_21254_4673# a_20963_4373# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X863 a_7423_2589# a_6559_2223# a_7166_2335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X864 a_33133_3855# _163_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X865 a_10901_4765# a_10563_4551# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X866 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X867 lsb[3] a_32319_7127# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X868 msb_n[15] a_1644_6549# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X869 vccd1 _232_.D a_6805_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X870 vccd1 a_29791_2388# _225_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X871 vccd1 a_17743_2197# _149_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X872 a_17985_3065# _159_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X873 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X874 _115_.A a_28567_4917# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X875 a_17743_2197# _215_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X876 a_13069_2741# clkbuf_2_3__f_clk.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X877 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X878 a_8093_4233# a_7546_3977# a_7746_4132# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X879 vccd1 a_32367_5175# output28.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X880 _177_.B a_21023_2806# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X881 _115_.Y _115_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X882 vssd1 a_32954_5220# a_32883_5321# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X883 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X884 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X885 a_21173_3855# a_20996_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X886 a_17581_4943# a_17047_4949# a_17486_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X887 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X888 vssd1 a_14715_3285# a_14722_3585# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X889 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X890 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X891 _160_.X a_19623_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X892 vccd1 output41.A a_15299_7127# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X893 a_9738_2375# a_9834_2197# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X894 vssd1 _205_.B1 a_20346_5263# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X895 vccd1 output38.A _098_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X896 vssd1 a_3116_6549# msb_n[14] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X897 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X898 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X899 output52.A output36.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X900 vssd1 a_34944_2375# _168_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X901 vssd1 a_23478_3855# _209_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X902 vccd1 a_19602_3855# a_19708_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X903 vccd1 clk a_20442_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X904 vssd1 a_12999_6575# msb_n[8] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X905 a_22983_2375# _135_.X a_23217_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X906 vssd1 a_23599_3579# a_23557_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X907 vssd1 a_7499_3579# a_7457_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X908 _222_.CLK a_23478_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X909 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X910 _232_.CLK a_13069_3829# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X911 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X912 vccd1 _232_.CLK a_17047_4949# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X913 a_30773_2589# a_30435_2375# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X914 a_7159_4087# a_7255_4087# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X915 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X916 vccd1 _160_.X a_27209_2806# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X917 a_4823_4399# a_4687_4373# a_4403_4373# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X918 a_7423_2589# a_6725_2223# a_7166_2335# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X919 vssd1 a_22983_2375# _140_.A_N vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X920 vccd1 _209_.CLK a_24591_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X921 a_16088_7093# output56.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X922 a_30550_3311# a_30373_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X923 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X924 vccd1 a_34948_7093# lsb_n[1] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X925 vccd1 a_33903_4667# a_33819_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X926 a_18045_3855# a_17868_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X927 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X928 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X929 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X930 a_11001_3133# _185_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X931 clkbuf_2_3__f_clk.A a_20442_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X932 a_20647_2223# a_20518_2497# a_20227_2197# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X933 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X934 msb_n[4] a_19676_7093# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X935 vccd1 a_7591_2491# a_7507_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X936 a_18243_3311# _206_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X937 a_8093_4233# a_7539_4073# a_7746_4132# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X938 vssd1 a_13069_2741# _233_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X939 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X940 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X941 a_20177_4943# _205_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X942 a_33493_3311# a_32503_3311# a_33367_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X943 a_7001_3677# a_6467_3311# a_6906_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X944 a_3116_6549# _108_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X945 lsb_n[3] a_31767_6575# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X946 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X947 _209_.CLK a_23478_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X948 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X949 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X950 vccd1 output28.A _094_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X951 a_30531_2197# a_30815_2197# a_30750_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X952 vccd1 _159_.A a_9821_3638# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X953 vccd1 _241_.D a_12627_4649# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X954 vssd1 _149_.A2 a_11746_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X955 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X956 vssd1 clkbuf_2_3__f_clk.A a_23478_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X957 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X958 a_10936_7093# output59.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X959 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X960 vssd1 a_29579_3829# a_29537_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X961 a_28399_4943# a_27535_4949# a_28142_4917# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X962 a_35545_3855# _125_.A2 _125_.B1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X963 vssd1 a_6734_4373# a_6663_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X964 vssd1 a_29518_2999# a_29467_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X965 vccd1 a_11023_2388# _185_.A0 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X966 vccd1 a_37471_7127# lsb[0] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X967 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X968 vssd1 _241_.D a_17836_4373# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X969 vssd1 a_28871_4564# _226_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X970 vccd1 a_13069_3829# _232_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X971 a_13545_4399# _241_.D a_13327_4373# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X972 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X973 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X974 a_23540_7093# output52.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X975 a_3116_6549# _108_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X976 _233_.CLK a_13069_2741# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X977 vssd1 _209_.CLK a_22015_4949# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
D10 vssd1 dac_in[3] sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
X978 a_32954_5220# a_32747_5161# a_33130_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X979 vssd1 output35.A output51.A vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X980 _173_.A0 a_26431_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X981 a_10943_4373# _232_.CLK vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X982 a_35334_4765# a_35061_4399# a_35249_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X983 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X984 a_6913_2223# _219_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X985 a_30951_2223# a_30815_2197# a_30531_2197# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X986 vccd1 output33.A _108_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X987 vssd1 a_17556_2999# _192_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X988 a_33110_3423# a_32942_3677# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X989 vssd1 _180_.X a_16180_3285# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X990 a_27446_4215# ANTENNA__177__A.DIODE a_27365_4215# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X991 vccd1 a_9411_7127# msb_n[10] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X992 vccd1 a_34955_3463# _169_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X993 vssd1 output20.A _114_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X994 lsb[0] a_37471_7127# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X995 a_7791_2767# a_7093_2773# a_7534_2741# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X996 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X997 vssd1 _145_.A a_12065_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X998 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X999 vccd1 a_23431_3677# a_23599_3579# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1000 vccd1 a_7331_3677# a_7499_3579# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1001 vssd1 _135_.X a_20713_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1002 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1003 lsb[2] a_33844_7093# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X1004 vccd1 _209_.CLK a_32871_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1005 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1006 vccd1 _196_.B a_19901_4649# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1007 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1008 a_34944_2375# input3.X a_35086_2550# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1009 a_23478_2767# clkbuf_2_3__f_clk.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1010 a_33130_4943# a_32883_5321# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1011 vccd1 a_19623_3311# _160_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1012 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X1013 a_22372_3087# _135_.X a_22069_2741# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1014 msb_n[10] a_9411_7127# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X1015 vccd1 a_35759_4765# a_35927_4667# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1016 a_8211_4649# _149_.B1 a_7993_4373# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1017 a_6243_4373# a_6527_4373# a_6462_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1018 vccd1 _145_.A a_3063_2473# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1019 lsb_n[5] a_27956_7093# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1020 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1021 vssd1 _126_.A a_30054_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1022 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1023 vccd1 a_7343_5175# output32.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1024 a_4307_4551# a_4403_4373# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1025 a_30815_2197# _222_.CLK vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1026 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1027 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1028 _195_.X a_7663_5487# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1029 vccd1 a_28567_4917# a_28483_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1030 vccd1 a_10147_7127# msb[10] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1031 a_35086_2550# _160_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1032 a_27295_3677# a_26597_3311# a_27038_3423# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1033 msb_n[5] a_17928_7093# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1034 _159_.X a_14287_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1035 vssd1 _241_.D a_17585_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1036 vssd1 output31.A a_6835_7127# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1037 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1038 vccd1 a_23478_2767# _222_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1039 a_10296_3311# _179_.A1 a_10075_3638# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1040 vccd1 a_6835_7127# msb[12] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1041 vssd1 a_36599_3476# _166_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1042 a_32922_2375# a_33018_2197# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1043 vssd1 _121_.A a_11746_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1044 a_34955_3463# _168_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1045 vssd1 a_12045_4087# a_11858_3829# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1046 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1047 a_35086_2223# _160_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1048 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1049 vssd1 a_17985_3065# a_17919_3133# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1050 vccd1 _196_.B a_15561_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1051 vccd1 a_33643_3855# a_33811_3829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1052 _185_.X a_10719_3894# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1053 a_10563_4551# a_10659_4373# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1054 _125_.B1 ANTENNA__118__A.DIODE vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X1055 _102_.Y output42.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1056 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1057 a_32883_5321# a_32754_5065# a_32463_5175# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1058 a_3615_3087# _145_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1059 vccd1 dac_in[1] a_34159_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1060 a_22287_2767# _215_.Q a_22069_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1061 vccd1 a_35502_4511# a_35429_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1062 a_33301_5321# a_32754_5065# a_32954_5220# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1063 a_33727_3855# a_32945_3861# a_33643_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1064 vssd1 a_23478_3855# _209_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1065 a_18141_2223# _215_.Q a_18035_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1066 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1067 a_35429_4765# a_34895_4399# a_35334_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1068 output19.A a_28015_4667# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1069 a_23515_3677# a_22733_3311# a_23431_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1070 a_7415_3677# a_6633_3311# a_7331_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1071 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X1072 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1073 vssd1 a_35759_4765# a_35927_4667# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1074 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1075 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1076 _155_.B1 a_2869_3087# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1077 a_29154_3829# a_28986_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X1078 vccd1 _222_.CLK a_32319_2773# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1079 a_20442_3311# clk vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1080 vccd1 a_7791_2767# a_7959_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1081 a_7539_4073# _233_.CLK vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1082 vccd1 _208_.X a_15269_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1083 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X1084 vssd1 a_22068_7093# msb_n[3] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X1085 vccd1 a_16578_4373# a_16507_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X1086 vccd1 _205_.B1 a_21801_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1087 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1088 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X1089 msb_n[12] a_6428_6549# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1090 a_34955_3463# _162_.A a_35129_3339# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1091 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1092 a_13445_2375# _183_.X a_13608_2473# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1093 a_35437_4175# _125_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1094 vccd1 output16.A _110_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1095 a_35228_3133# _125_.A2 a_35007_2806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1096 a_26965_3677# a_26431_3311# a_26870_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1097 vccd1 a_31767_6575# lsb_n[3] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1098 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1099 vssd1 _180_.A a_12065_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1100 vccd1 ANTENNA__118__A.DIODE a_37011_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1101 a_35007_3133# a_34753_2806# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1102 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1103 vssd1 a_29791_2388# _225_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1104 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1105 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X1106 vccd1 _199_.X a_8093_4233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1107 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1108 vssd1 a_23431_3677# a_23599_3579# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1109 vccd1 output15.A a_37839_6575# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1110 a_31267_2741# _211_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1111 vssd1 clkbuf_2_3__f_clk.A a_13069_2741# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1112 vssd1 a_7331_3677# a_7499_3579# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1113 a_37503_4193# ANTENNA__118__A.DIODE vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1114 a_22804_7093# output37.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1115 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X1116 vssd1 a_6527_4373# a_6534_4673# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1117 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1118 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1119 _205_.B1 a_19439_2223# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1120 vssd1 a_30550_3311# a_30656_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1121 a_29154_3829# a_28986_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1122 vccd1 _115_.A _115_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1123 vssd1 output34.A output50.A vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1124 vssd1 a_17654_4917# a_17612_5321# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1125 a_7875_2767# a_7093_2773# a_7791_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1126 _155_.A1 _179_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1127 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1128 vccd1 a_13069_3829# _232_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1129 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1130 _209_.CLK a_23478_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1131 vssd1 a_24591_7127# msb[2] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X1132 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1133 vccd1 a_29411_3855# a_29579_3829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1134 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1135 vccd1 a_31215_7127# lsb[4] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1136 vccd1 output36.A output52.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1137 vssd1 a_17836_4373# _238_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1138 lsb_n[1] a_34948_7093# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1139 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1140 vccd1 _128_.B1 a_31267_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1141 _125_.A1 a_30054_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1142 vccd1 a_33367_3677# a_33535_3579# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1143 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1144 vccd1 _159_.X a_21237_2806# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
D11 vssd1 _133_.A sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
X1145 a_33310_4765# a_33037_4399# a_33225_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1146 a_31355_4087# _126_.A a_31589_4221# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1147 vssd1 output15.A a_37839_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1148 a_32747_5161# _209_.CLK vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1149 vssd1 a_17911_4943# a_18079_4917# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1150 a_14186_5220# a_13979_5161# a_14362_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1151 a_15685_4153# _159_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1152 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1153 a_4307_4551# a_4403_4373# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1154 a_6485_4765# a_6147_4551# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1155 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1156 _180_.A a_11746_2223# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1157 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1158 a_19676_7093# _098_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1159 a_22197_3971# ANTENNA__177__A.DIODE vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1160 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1161 a_10075_3638# _179_.A1 a_10003_3638# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1162 vccd1 test_mode a_1591_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1163 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1164 a_16021_2767# a_15844_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1165 _144_.A1 a_15319_2491# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1166 a_7366_2767# a_6927_2773# a_7281_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1167 a_17965_4399# _203_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1168 a_31355_4087# _128_.B1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1169 a_11079_4399# a_10943_4373# a_10659_4373# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1170 _233_.CLK a_13069_2741# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1171 vssd1 a_13459_7127# msb[8] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X1172 a_23849_2473# _133_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1173 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1174 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1175 a_29411_3855# a_28547_3861# a_29154_3829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1176 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1177 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1178 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1179 a_12075_4943# _196_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1180 a_14362_4943# a_14115_5321# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1181 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1182 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X1183 vssd1 a_29154_3829# a_29112_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1184 vccd1 output38.A _098_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1185 _178_.A a_25635_3105# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1186 vssd1 a_2288_7093# msb[15] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X1187 vccd1 a_21454_4373# a_21383_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X1188 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1189 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1190 a_17401_4943# _238_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1191 a_7474_4221# a_7159_4087# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1192 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X1193 a_27337_4399# _224_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1194 vssd1 a_11023_2388# _185_.A0 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1195 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1196 vccd1 _125_.A1 a_30373_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1197 vssd1 a_5687_3463# _152_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1198 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1199 a_12242_2223# a_12065_2223# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1200 a_7492_3145# a_7093_2773# a_7366_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1201 _232_.CLK a_13069_3829# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1202 msb[13] a_5600_7093# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1203 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1204 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1205 a_7859_5321# a_7730_5065# a_7439_5175# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1206 vccd1 a_12409_4373# _188_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1207 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1208 a_24757_2223# a_24591_2223# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1209 vssd1 _135_.A a_20394_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1210 vssd1 a_27220_7093# msb[0] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1211 a_28986_3855# a_28547_3861# a_28901_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1212 vccd1 a_13069_2741# _233_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1213 _232_.D a_2695_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1214 a_10657_5281# _203_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1215 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1216 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1217 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1218 a_30833_3311# a_30656_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1219 _108_.Y output33.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1220 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1221 a_22983_2375# _133_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1222 a_9757_3145# a_8767_2773# a_9631_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1223 a_27379_3677# a_26597_3311# a_27295_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1224 vccd1 a_10340_2375# _149_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1225 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1226 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1227 clkbuf_2_3__f_clk.A a_20442_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1228 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1229 a_13327_4373# _241_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1230 a_6663_4399# a_6527_4373# a_6243_4373# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1231 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1232 _209_.CLK a_23478_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1233 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1234 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X1235 vccd1 _149_.A1 a_8211_4649# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1236 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1237 a_22285_2223# _136_.Y a_22067_2197# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1238 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1239 vssd1 output36.A output52.A vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1240 vccd1 _179_.A1 _155_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1241 vssd1 clkbuf_2_3__f_clk.A a_23478_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1242 _098_.Y output38.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1243 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1244 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X1245 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1246 a_27677_2806# _173_.A0 a_27463_2806# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1247 vssd1 _180_.X a_17266_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1248 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1249 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1250 a_15147_4427# _180_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1251 vccd1 a_19970_2767# a_20076_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1252 a_2785_3087# _149_.B1 a_2689_3087# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1253 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X1254 output36.A a_23047_4917# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1255 vssd1 _233_.CLK a_6559_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1256 vccd1 _159_.X a_10933_3894# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1257 vssd1 a_16088_7093# msb_n[6] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X1258 a_14533_5321# a_13986_5065# a_14186_5220# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1259 vccd1 a_36783_5162# _163_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1260 vssd1 a_28784_6549# lsb[5] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1261 vccd1 output36.A a_24591_7127# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1262 vccd1 a_10839_2999# _198_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1263 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1264 a_32682_5309# a_32367_5175# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1265 _195_.X a_7663_5487# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1266 vssd1 a_9631_2767# a_9799_2741# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1267 vssd1 _180_.B a_15233_4427# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1268 vssd1 _206_.A2 a_12617_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1269 a_14186_5220# a_13986_5065# a_14335_5309# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1270 a_6527_4373# _232_.CLK vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1271 a_9738_2375# a_9834_2197# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1272 vssd1 _180_.X a_17192_3285# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1273 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1274 vccd1 a_8307_7127# msb[11] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1275 a_24945_4399# _203_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1276 vccd1 _165_.B a_35755_3339# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1277 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1278 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1279 vssd1 clk a_20442_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1280 vssd1 dac_in[1] a_34159_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1281 vssd1 a_27038_3423# a_26996_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1282 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1283 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1284 a_25380_7093# output51.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1285 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1286 output24.A output18.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1287 a_36131_2806# a_35949_2806# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1288 a_29411_3855# a_28713_3861# a_29154_3829# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1289 _209_.CLK a_23478_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1290 vccd1 a_14563_7127# msb_n[7] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1291 vssd1 a_18611_7127# msb[5] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X1292 _179_.A1 a_7591_2491# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1293 _134_.X a_31480_3561# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1294 vccd1 a_33110_3423# a_33037_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1295 vccd1 a_37703_4564# _157_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1296 a_25581_2223# a_24591_2223# a_25455_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1297 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1298 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1299 vccd1 a_20442_3311# clkbuf_2_3__f_clk.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1300 a_11863_5639# _196_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1301 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1302 a_14533_5321# a_13979_5161# a_14186_5220# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1303 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1304 vssd1 a_23540_7093# msb_n[2] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
D12 vssd1 clk sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
X1305 a_13979_5161# _232_.CLK vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1306 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1307 input3.X a_29743_4399# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1308 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1309 vssd1 a_13069_3829# _232_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1310 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1311 _169_.X a_34527_4943# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1312 a_28784_6549# _115_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1313 vccd1 a_25019_3285# a_25026_3585# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1314 a_16309_3561# _205_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1315 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1316 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1317 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1318 vccd1 a_26063_7127# msb[1] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1319 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1320 lsb_n[4] a_29796_7093# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1321 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X1322 a_35502_4511# a_35334_4765# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X1323 _174_.X a_28303_3339# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1324 vccd1 a_23478_2767# _222_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1325 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1326 output52.A output36.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1327 lsb_n[0] a_36236_6549# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1328 vccd1 dac_in[9] a_8399_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
D13 vssd1 dac_in[8] sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
X1329 a_14726_2589# a_14287_2223# a_14641_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1330 _205_.B1 a_19439_2223# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1331 _196_.B a_15242_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1332 a_6147_4551# a_6243_4373# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1333 vccd1 a_33108_7093# lsb_n[2] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1334 msb_n[7] a_14563_7127# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1335 _209_.CLK a_23478_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1336 vccd1 a_38023_6039# llsb vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1337 a_34619_3855# _125_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1338 _232_.CLK a_13069_3829# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1339 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1340 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1341 vssd1 _205_.X a_25573_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1342 a_25198_2335# a_25030_2589# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1343 vccd1 a_23478_2767# _222_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1344 vssd1 _205_.A1 a_19425_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1345 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1346 vssd1 a_23478_3855# _209_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1347 a_20253_2767# a_20076_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1348 vssd1 a_13069_2741# _233_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1349 a_33844_7093# output18.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1350 a_19426_5263# _205_.B1 a_19257_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1351 a_28784_6549# _115_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1352 vssd1 a_28567_4917# a_28525_5321# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
D14 vssd1 ANTENNA__118__A.DIODE sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
X1353 vssd1 a_28423_2999# _172_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1354 vccd1 _180_.A a_18416_3561# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1355 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1356 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1357 a_20951_2806# a_20769_2806# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1358 a_6913_2223# _219_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1359 a_15151_2589# a_14287_2223# a_14894_2335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1360 a_22370_2473# _133_.B a_22067_2197# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1361 a_35061_4399# a_34895_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1362 a_26597_3311# a_26431_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
D15 vssd1 _133_.A sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
X1363 a_15715_3894# _183_.A1 a_15256_4087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1364 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1365 msb[1] a_26063_7127# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1366 a_14852_2223# a_14453_2223# a_14726_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1367 a_12794_3311# a_12617_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1368 vssd1 _222_.CLK a_26431_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1369 a_7159_4087# a_7255_4087# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1370 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1371 vccd1 a_17192_7093# msb[6] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1372 vssd1 a_4894_4373# a_4823_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1373 a_25455_4765# a_24757_4399# a_25198_4511# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1374 a_12525_2223# a_12348_2223# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1375 vssd1 test_mode a_1591_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1376 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X1377 vccd1 a_35631_7127# lsb[1] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1378 vssd1 a_23478_2767# _222_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1379 vssd1 output29.A output45.A vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1380 a_27701_4949# a_27535_4949# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1381 a_30435_2375# a_30531_2197# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1382 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1383 a_15685_4153# _159_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1384 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1385 a_10075_3638# _179_.A0 a_10075_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1386 vccd1 _145_.A a_2511_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1387 _151_.C _145_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1388 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1389 a_5600_7093# output32.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1390 a_17928_7093# output55.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1391 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1392 a_32926_2741# a_32758_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X1393 msb[9] a_11987_7127# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X1394 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X1395 a_5967_5461# a_6258_5761# a_6209_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1396 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1397 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1398 vssd1 a_33524_2375# _125_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1399 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1400 a_11506_3311# a_11329_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1401 _108_.Y output33.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1402 a_22097_3855# _140_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1403 a_22622_4917# a_22454_4943# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X1404 msb[0] a_27220_7093# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1405 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1406 vccd1 _126_.A a_30054_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1407 a_25226_3285# a_25019_3285# a_25402_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1408 lsb[1] a_35631_7127# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1409 a_13069_3829# clkbuf_2_3__f_clk.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1410 a_7658_5309# a_7343_5175# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1411 vssd1 a_14894_2335# a_14852_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1412 a_10340_2375# _183_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1413 _233_.CLK a_13069_2741# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1414 _098_.Y output38.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1415 a_27931_4765# a_27149_4399# a_27847_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1416 _141_.A a_22197_3971# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1417 a_22622_4917# a_22454_4943# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1418 a_35759_4765# a_34895_4399# a_35502_4511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1419 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1420 a_9715_2767# a_8933_2773# a_9631_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1421 _157_.A a_37503_4193# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1422 output46.A output30.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1423 _224_.D a_26431_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1424 vccd1 a_10021_2375# a_9834_2197# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1425 vccd1 _121_.A a_11746_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1426 a_30120_2999# _131_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1427 a_25375_3311# a_25155_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1428 vccd1 output39.A a_18611_7127# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1429 a_13914_5309# a_13599_5175# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1430 a_4403_4373# a_4687_4373# a_4622_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1431 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1432 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1433 vssd1 _232_.CLK a_17047_4949# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1434 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X1435 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1436 _145_.A a_11746_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1437 a_25402_3677# a_25155_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1438 vssd1 a_20442_3311# clkbuf_2_3__f_clk.A vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1439 vssd1 a_6428_6549# msb_n[12] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X1440 vssd1 _145_.B _145_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1441 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1442 a_35007_2806# _164_.A0 a_35007_3133# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1443 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1444 vccd1 a_6251_5461# a_6258_5761# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1445 a_28423_2999# _162_.A a_28597_3105# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1446 vccd1 a_23478_3855# _209_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1447 vccd1 a_9655_4087# _199_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1448 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X1449 vssd1 a_16578_4373# a_16507_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1450 vssd1 a_33643_3855# a_33811_3829# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1451 a_18416_3561# _206_.A2 a_18325_3561# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1452 _141_.X a_22659_4399# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1453 vssd1 a_20442_3311# clkbuf_2_3__f_clk.A vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1454 vccd1 a_20442_3311# clkbuf_2_3__f_clk.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1455 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1456 vccd1 _233_.CLK a_8767_2773# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1457 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1458 a_22067_2197# _136_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1459 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1460 vccd1 _205_.A2 a_20177_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1461 a_22733_3311# a_22567_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1462 a_6633_3311# a_6467_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1463 a_6147_4551# a_6243_4373# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1464 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1465 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1466 vssd1 _093_.A a_38023_6039# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1467 vssd1 a_36783_5162# _163_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1468 a_33735_4765# a_33037_4399# a_33478_4511# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1469 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1470 a_8211_4649# _149_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1471 a_25226_3285# a_25026_3585# a_25375_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1472 vssd1 a_13069_3829# _232_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1473 a_23478_2767# clkbuf_2_3__f_clk.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1474 a_27889_4943# _226_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1475 vccd1 _125_.A1 a_27249_2473# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1476 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1477 vccd1 _241_.D a_14533_5321# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1478 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1479 vccd1 _180_.A a_12065_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1480 vccd1 a_23478_2767# _222_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1481 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1482 a_10647_3894# a_10465_3894# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1483 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1484 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X1485 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1486 a_12242_2767# a_12065_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1487 vssd1 _134_.A1 a_31307_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1488 vssd1 a_19676_7093# msb_n[4] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X1489 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1490 a_20890_3855# a_20713_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1491 a_10483_5175# _203_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1492 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1493 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X1494 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1495 a_5871_5639# a_5967_5461# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1496 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X1497 a_14641_2223# _145_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1498 vccd1 a_30550_3311# a_30656_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1499 vssd1 a_14922_3285# a_14851_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1500 vssd1 a_7343_5175# output32.A vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1501 vccd1 a_35927_4667# a_35843_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1502 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1503 a_15901_5281# _196_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1504 vccd1 a_25455_2589# a_25623_2491# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1505 vssd1 _159_.X a_10940_4221# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1506 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1507 _219_.D _155_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1508 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1509 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X1510 a_33183_2767# a_32319_2773# a_32926_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1511 a_33524_2375# _211_.Q vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1512 a_25573_3311# a_25019_3285# a_25226_3285# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1513 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1514 _152_.X a_5823_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1515 a_22287_2767# _133_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1516 vccd1 a_17985_3065# a_18015_2806# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1517 _232_.CLK a_13069_3829# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1518 msb_n[2] a_23540_7093# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1519 vccd1 a_36236_6549# lsb_n[0] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1520 a_12409_4373# _196_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1521 a_25573_3311# a_25026_3585# a_25226_3285# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1522 a_20442_3311# clk vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1523 a_14673_3677# a_14335_3463# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1524 _114_.Y output20.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1525 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1526 output50.A output34.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1527 _094_.Y output28.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1528 a_20227_2197# a_20518_2497# a_20469_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1529 vccd1 _140_.C a_22197_3971# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1530 vccd1 output18.A output24.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1531 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1532 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1533 a_17192_7093# output40.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1534 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1535 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1536 vssd1 a_27215_4087# _129_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1537 a_17762_3855# a_17585_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1538 a_32758_2767# a_32319_2773# a_32673_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1539 _166_.A a_35755_3339# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1540 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1541 _169_.X a_34527_4943# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1542 a_7497_3855# a_7159_4087# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1543 clkbuf_2_3__f_clk.A a_20442_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1544 msb[14] a_4036_7093# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1545 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1546 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1547 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1548 a_14431_3285# a_14715_3285# a_14650_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1549 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X1550 a_29796_7093# _114_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1551 _203_.X a_19426_5263# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1552 vssd1 output57.A a_14563_7127# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1553 a_25030_4765# a_24591_4399# a_24945_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1554 vssd1 a_15256_4087# _183_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1555 _232_.CLK a_13069_3829# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1556 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1557 a_7549_2223# a_6559_2223# a_7423_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1558 vssd1 ANTENNA__177__A.DIODE a_19106_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1559 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1560 vccd1 a_10936_7093# msb_n[9] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1561 a_16915_2197# _180_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1562 vccd1 a_20511_2197# a_20518_2497# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1563 output59.A output43.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1564 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1565 vssd1 dac_in[9] a_8399_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1566 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1567 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1568 _162_.B a_36203_2806# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1569 a_32884_3145# a_32485_2773# a_32758_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1570 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1571 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1572 vssd1 a_7624_7093# msb_n[11] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1573 vccd1 _209_.CLK a_34895_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1574 vccd1 a_33351_2741# a_33267_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1575 vccd1 a_13069_3829# _232_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1576 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1577 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X1578 vssd1 output35.A a_26063_7127# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1579 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1580 _206_.A2 a_12298_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1581 _209_.CLK a_23478_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1582 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1583 a_25030_2589# a_24757_2223# a_24945_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1584 _233_.CLK a_13069_2741# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1585 a_14851_3311# a_14715_3285# a_14431_3285# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1586 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1587 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X1588 a_30750_2223# a_30435_2375# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1589 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1590 a_25156_4399# a_24757_4399# a_25030_4765# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1591 a_6998_2589# a_6725_2223# a_6913_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1592 vssd1 _137_.X a_21065_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1593 vccd1 a_20504_7093# msb[4] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1594 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1595 vssd1 a_16371_4373# a_16378_4673# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1596 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1597 a_27220_7093# output28.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1598 a_22879_4943# a_22181_4949# a_22622_4917# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1599 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1600 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1601 vssd1 _222_.CLK a_32319_2773# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1602 a_23174_3423# a_23006_3677# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X1603 a_7074_3423# a_6906_3677# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X1604 vssd1 output43.A a_11987_7127# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1605 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X1606 vssd1 a_33205_2375# a_33018_2197# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1607 a_23174_3423# a_23006_3677# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1608 a_13649_3561# _145_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1609 a_7074_3423# a_6906_3677# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1610 a_7539_4073# _233_.CLK vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1611 a_17836_4373# _205_.A1 a_18059_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1612 vccd1 a_28871_4564# _226_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1613 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1614 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1615 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1616 _196_.A a_11010_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1617 a_7675_4233# a_7539_4073# a_7255_4087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1618 a_28142_4917# a_27974_4943# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X1619 _110_.Y output16.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1620 a_5871_5639# a_5967_5461# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1621 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X1622 vssd1 a_15685_4153# a_15619_4221# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1623 vccd1 _125_.A1 a_30659_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1624 _222_.CLK a_23478_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
D16 vssd1 test_mode sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
X1625 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1626 a_10021_2375# _149_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1627 vssd1 a_25380_7093# msb_n[1] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1628 a_16180_3285# ANTENNA__118__A.DIODE a_16403_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1629 a_28142_4917# a_27974_4943# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1630 vssd1 a_25198_4511# a_25156_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1631 a_7255_4087# a_7539_4073# a_7474_4221# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1632 msb[8] a_13459_7127# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1633 a_27463_3133# a_27209_2806# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1634 a_32942_3677# a_32503_3311# a_32857_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1635 a_22285_2223# _135_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1636 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1637 vssd1 output18.A output24.A vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1638 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1639 a_14715_3285# _232_.CLK vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1640 _180_.B a_10075_3638# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1641 _209_.CLK a_23478_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1642 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X1643 a_16329_4765# a_15991_4551# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1644 a_7917_3145# a_6927_2773# a_7791_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1645 a_22068_7093# output53.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1646 a_33310_4765# a_32871_4399# a_33225_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1647 vccd1 a_25198_2335# a_25125_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1648 a_11762_4087# a_11858_3829# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1649 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1650 vccd1 output40.A output56.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1651 vssd1 clkbuf_2_3__f_clk.A a_13069_3829# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1652 a_9829_4193# _205_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1653 vssd1 _209_.CLK a_26983_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1654 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1655 vccd1 a_23478_2767# _222_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1656 a_7281_2767# _152_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1657 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1658 msb[4] a_20504_7093# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1659 a_18703_3087# _140_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1660 vssd1 a_13069_2741# _233_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1661 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1662 a_31267_2741# _134_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1663 output36.A a_23047_4917# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1664 vccd1 _206_.A2 a_12617_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1665 lsb[5] a_28784_6549# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1666 vccd1 a_21247_4373# a_21254_4673# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1667 vssd1 output30.A output46.A vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1668 vssd1 a_11150_4373# a_11079_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1669 _130_.X a_25787_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1670 vccd1 a_37839_6575# llsb_n vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1671 vccd1 a_28399_4943# a_28567_4917# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1672 _217_.D a_3788_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1673 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X1674 a_33367_3677# a_32503_3311# a_33110_3423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1675 a_6462_4399# a_6147_4551# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1676 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1677 vssd1 a_7591_2491# a_7549_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1678 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1679 a_25721_3105# ANTENNA__177__A.DIODE a_25635_3105# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1680 a_25125_2589# a_24591_2223# a_25030_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1681 a_7093_2773# a_6927_2773# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1682 a_32747_5161# _209_.CLK vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1683 a_33436_4399# a_33037_4399# a_33310_4765# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1684 vccd1 _222_.CLK a_22567_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1685 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1686 a_28303_3339# _162_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1687 a_25155_3311# a_25026_3585# a_24735_3285# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1688 vccd1 _233_.CLK a_6467_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1689 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X1690 vssd1 a_24639_3463# output37.A vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1691 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X1692 ANTENNA__118__A.DIODE a_16915_2197# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1693 a_28901_3855# _225_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1694 a_17919_3133# input7.X a_17556_2999# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1695 vccd1 _159_.A a_14287_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1696 a_4687_4373# _232_.CLK vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1697 _235_.D a_20070_4399# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1698 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X1699 input1.X a_36091_2223# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1700 _135_.X a_20394_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1701 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X1702 a_11789_3311# a_11612_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1703 a_7895_4221# a_7675_4233# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1704 a_13069_3829# clkbuf_2_3__f_clk.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1705 vccd1 _241_.D a_12075_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1706 _222_.CLK a_23478_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1707 vccd1 a_11857_4917# _190_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1708 vssd1 a_4772_7093# msb_n[13] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1709 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1710 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1711 a_20867_4551# a_20963_4373# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1712 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1713 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1714 _163_.A a_36399_4193# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1715 a_29801_2999# _133_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1716 _174_.B a_27463_2806# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1717 a_16507_4399# a_16371_4373# a_16087_4373# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1718 vssd1 a_33478_4511# a_33436_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1719 a_33205_2375# _125_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1720 a_10289_3638# _179_.A0 a_10075_3638# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1721 output39.A a_18079_4917# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1722 vssd1 a_17743_2197# _149_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1723 a_28713_3861# a_28547_3861# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1724 vccd1 a_7746_4132# a_7675_4233# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X1725 a_27973_4399# a_26983_4399# a_27847_4765# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1726 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1727 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1728 vssd1 _174_.B a_28389_3339# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1729 _151_.C _149_.B1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1730 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
D17 vssd1 ANTENNA__177__A.DIODE sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
X1731 vssd1 _209_.CLK a_24591_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1732 vccd1 _162_.A a_28423_2999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1733 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X1734 a_7439_5175# a_7730_5065# a_7681_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1735 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X1736 vssd1 a_5600_7093# msb[13] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1737 vccd1 a_6458_5461# a_6387_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X1738 a_5443_3087# _155_.A1 _219_.D vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1739 a_25539_4765# a_24757_4399# a_25455_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1740 _209_.CLK a_23478_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1741 vccd1 _205_.X a_25573_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1742 a_22284_4215# a_22097_3855# a_22197_3971# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1743 a_17698_2806# _159_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1744 vccd1 a_33535_3579# a_33451_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1745 vssd1 _115_.A _115_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1746 a_26870_3677# a_26597_3311# a_26785_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1747 vssd1 _233_.CLK a_14287_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1748 a_33110_3423# a_32942_3677# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X1749 _241_.D a_17266_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1750 a_2288_7093# output34.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1751 a_20504_7093# output38.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1752 vssd1 clk a_20442_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1753 vccd1 a_20442_3311# clkbuf_2_3__f_clk.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1754 a_27974_4943# a_27535_4949# a_27889_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1755 a_21065_2223# a_20511_2197# a_20718_2197# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1756 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1757 vssd1 _160_.X a_36424_3133# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1758 a_21065_2223# a_20518_2497# a_20718_2197# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1759 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1760 a_4036_7093# output33.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1761 a_16371_4373# _232_.CLK vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1762 a_31559_3133# _128_.B1 a_31463_3133# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1763 vssd1 a_13069_3829# _232_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1764 output52.A output36.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1765 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1766 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1767 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X1768 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1769 msb_n[9] a_10936_7093# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1770 a_27590_4511# a_27422_4765# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1771 vccd1 a_18751_2388# input7.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1772 msb_n[11] a_7624_7093# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1773 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1774 vssd1 a_31355_4087# _126_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1775 vssd1 clkbuf_2_3__f_clk.A a_23478_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1776 a_15727_5175# _196_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1777 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1778 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X1779 vssd1 a_7930_5220# a_7859_5321# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1780 a_10943_4373# _232_.CLK vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1781 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1782 a_32857_3311# _166_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1783 vccd1 a_15685_4153# a_15715_3894# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1784 vssd1 a_27463_3579# a_27421_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1785 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1786 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X1787 vssd1 a_13069_2741# _233_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1788 vccd1 output43.A output59.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1789 a_10340_2375# _183_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1790 vssd1 _162_.A a_19793_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1791 _232_.CLK a_13069_3829# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1792 lsb_n[2] a_33108_7093# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1793 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1794 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1795 a_27149_4399# a_26983_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1796 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1797 vssd1 _209_.CLK a_32871_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1798 _224_.D a_26431_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1799 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1800 a_28399_4943# a_27701_4949# a_28142_4917# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1801 _144_.A1 a_15319_2491# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1802 a_17985_3065# _159_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1803 a_33218_3855# a_32945_3861# a_33133_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1804 a_16088_7093# output56.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1805 _205_.X a_20346_5263# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1806 vccd1 _222_.CLK a_32503_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1807 msb[10] a_10147_7127# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X1808 a_13077_3311# a_12900_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1809 vccd1 a_23047_4917# a_22963_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1810 _126_.A a_25623_2491# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1811 vssd1 _159_.A a_9821_3638# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1812 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1813 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1814 _121_.A a_4351_2223# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1815 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1816 a_17321_3561# _205_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1817 msb_n[1] a_25380_7093# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1818 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X1819 a_7507_2589# a_6725_2223# a_7423_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1820 vssd1 output19.A a_32319_7127# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1821 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1822 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1823 vssd1 _196_.X a_2695_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1824 a_15991_4551# a_16087_4373# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1825 a_20867_4551# a_20963_4373# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1826 vssd1 a_1644_6549# msb_n[15] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1827 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1828 a_32954_5220# a_32754_5065# a_33103_5309# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1829 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1830 a_23478_3855# clkbuf_2_3__f_clk.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1831 vssd1 a_34955_3463# _169_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1832 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X1833 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1834 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1835 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
D18 vssd1 dac_in[2] sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
X1836 a_27215_4087# _128_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1837 a_19602_3855# a_19425_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1838 a_13979_5161# _232_.CLK vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1839 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X1840 a_32367_5175# a_32463_5175# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1841 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1842 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1843 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1844 vccd1 _209_.CLK a_32779_3861# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1845 a_30659_3855# _125_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1846 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1847 a_7124_2223# a_6725_2223# a_6998_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1848 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1849 vssd1 a_19623_3311# _160_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1850 vssd1 _160_.X a_27209_2806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1851 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1852 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1853 vccd1 a_22804_7093# msb[3] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1854 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1855 a_7930_5220# a_7723_5161# a_8106_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1856 vccd1 dac_in[4] a_26431_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1857 vccd1 a_12364_4087# ANTENNA__177__A.DIODE vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1858 a_3146_2223# _145_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1859 llsb_n a_37839_6575# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1860 a_7366_2767# a_7093_2773# a_7281_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1861 a_17654_4917# a_17486_4943# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X1862 vssd1 a_7423_2589# a_7591_2491# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1863 vccd1 a_23478_3855# _209_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1864 a_33301_5321# a_32747_5161# a_32954_5220# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1865 a_36485_4193# _162_.A a_36399_4193# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1866 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1867 a_23540_7093# output52.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1868 output56.A output40.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1869 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1870 vssd1 a_18079_4917# a_18037_5321# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1871 _222_.CLK a_23478_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1872 vccd1 _233_.CLK a_6927_2773# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1873 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1874 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1875 vccd1 a_37519_5162# _119_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1876 vssd1 a_31022_2197# a_30951_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1877 _233_.CLK a_13069_2741# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1878 a_14641_2223# _145_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1879 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1880 a_31480_3561# _133_.Y a_31307_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1881 vssd1 a_29796_7093# lsb_n[4] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1882 a_24757_4399# a_24591_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1883 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1884 a_33524_2375# _211_.Q vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1885 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1886 vccd1 a_33386_3829# a_33313_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1887 _152_.X a_5823_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1888 a_8106_4943# a_7859_5321# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1889 vssd1 a_7166_2335# a_7124_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1890 a_2689_3087# _149_.A1 a_2593_3087# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1891 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1892 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1893 vccd1 a_23174_3423# a_23101_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1894 vccd1 a_7074_3423# a_7001_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1895 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1896 a_19901_4649# _205_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1897 vccd1 a_32954_5220# a_32883_5321# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X1898 a_1644_6549# output50.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1899 _145_.Y _145_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1900 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1901 _177_.B a_21023_2806# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1902 a_30469_4649# _133_.B _133_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1903 vssd1 a_11863_5639# _196_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1904 vccd1 a_13069_2741# _233_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1905 msb[3] a_22804_7093# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1906 lsb[4] a_31215_7127# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X1907 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1908 a_31267_2741# _126_.A a_31665_3133# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1909 a_10940_4221# _149_.B1 a_10719_3894# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1910 msb_n[13] a_4772_7093# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1911 a_17654_4917# a_17486_4943# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1912 vccd1 a_20442_3311# clkbuf_2_3__f_clk.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1913 a_28986_3855# a_28713_3861# a_28901_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1914 _222_.CLK a_23478_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1915 _106_.Y output31.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1916 output45.A output29.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1917 a_13937_4943# a_13599_5175# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1918 a_20346_5263# _205_.B1 a_20177_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1919 a_34935_2806# a_34753_2806# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1920 a_33313_3855# a_32779_3861# a_33218_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1921 a_27701_4949# a_27535_4949# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1922 a_9655_4087# _205_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1923 vccd1 a_15299_7127# msb[7] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1924 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1925 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X1926 input1.X a_36091_2223# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1927 a_23101_3677# a_22567_3311# a_23006_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
D19 vssd1 dac_in[7] sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
X1928 a_3063_2473# _149_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1929 vssd1 a_20131_2375# _135_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1930 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1931 vccd1 _160_.X a_35949_2806# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1932 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1933 vssd1 clkbuf_2_3__f_clk.A a_13069_3829# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1934 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1935 vccd1 a_23478_2767# _222_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1936 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1937 vccd1 output31.A a_6835_7127# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1938 a_1644_6549# output50.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1939 a_29537_4233# a_28547_3861# a_29411_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1940 vccd1 a_7534_2741# a_7461_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1941 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1942 msb[7] a_15299_7127# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1943 a_25635_3105# ANTENNA__177__A.DIODE vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1944 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X1945 a_15991_4551# a_16087_4373# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1946 msb_n[0] a_26300_6549# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1947 vssd1 output16.A a_37471_7127# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1948 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1949 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1950 a_9121_2767# _217_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1951 output53.A output37.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1952 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1953 input3.X a_29743_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1954 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1955 a_8277_5321# a_7730_5065# a_7930_5220# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1956 a_12364_4087# _180_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1957 vssd1 _203_.A2 a_12712_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1958 a_30435_2375# a_30531_2197# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1959 vssd1 a_33844_7093# lsb[2] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1960 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1961 vccd1 _160_.X a_27677_2806# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1962 a_7461_2767# a_6927_2773# a_7366_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1963 _102_.Y output42.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1964 a_17911_4943# a_17047_4949# a_17654_4917# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1965 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1966 vccd1 _137_.X a_21065_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1967 vssd1 output45.A a_9411_7127# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1968 a_26479_2388# dac_in[5] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1969 clkbuf_2_3__f_clk.A a_20442_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1970 a_6725_2223# a_6559_2223# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1971 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1972 a_7930_5220# a_7730_5065# a_8079_5309# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1973 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1974 vccd1 a_29518_2999# a_29467_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1975 vssd1 _233_.CLK a_8767_2773# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1976 output24.A output18.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1977 a_36203_2806# input1.X a_36203_3133# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1978 vccd1 _183_.X a_15242_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1979 vssd1 a_27295_3677# a_27463_3579# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1980 a_7624_7093# output46.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1981 a_13069_2741# clkbuf_2_3__f_clk.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1982 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1983 _232_.CLK a_13069_3829# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1984 vccd1 a_7993_4373# _149_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1985 a_14335_3463# a_14431_3285# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1986 _217_.D a_3788_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1987 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1988 vssd1 a_18751_2388# input7.X vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X1989 vssd1 a_22069_2741# _140_.C vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1990 msb[12] a_6835_7127# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1991 a_30815_2197# _222_.CLK vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1992 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1993 vccd1 a_17928_7093# msb_n[5] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1994 a_22804_7093# output37.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1995 vccd1 _125_.A2 a_31355_4087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1996 output59.A output43.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1997 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1998 vccd1 _159_.X a_20769_2806# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1999 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X2000 a_13695_5175# a_13986_5065# a_13937_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2001 vccd1 a_14287_4399# _159_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2002 a_10021_2375# _149_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2003 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
D20 vssd1 ANTENNA__177__A.DIODE sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
X2004 vssd1 _180_.A a_19474_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2005 vccd1 a_17556_2999# _192_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2006 output46.A output30.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2007 a_32673_2767# _125_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2008 vccd1 _160_.X a_28321_2550# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2009 vssd1 _133_.B a_23935_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2010 vssd1 a_33351_2741# a_33309_3145# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2011 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2012 a_13599_5175# a_13695_5175# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2013 vssd1 a_29801_2999# a_29614_2741# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2014 output16.A a_33811_3829# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2015 a_8277_5321# a_7723_5161# a_7930_5220# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2016 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2017 vccd1 a_20718_2197# a_20647_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X2018 _222_.CLK a_23478_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2019 vssd1 output29.A a_10147_7127# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2020 vssd1 _160_.X a_28328_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2021 a_25455_2589# a_24591_2223# a_25198_2335# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2022 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2023 _233_.CLK a_13069_2741# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2024 vssd1 _188_.X a_11497_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2025 lsb[3] a_32319_7127# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2026 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X2027 vccd1 _135_.X a_22287_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2028 a_10075_3311# a_9821_3638# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2029 vccd1 a_13069_3829# _232_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2030 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2031 a_18325_3561# _180_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2032 vccd1 _119_.X a_33301_5321# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2033 vssd1 a_14186_5220# a_14115_5321# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2034 a_35759_4765# a_35061_4399# a_35502_4511# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2035 a_17556_2999# _144_.A1 a_17698_3133# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2036 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X2037 _130_.X a_25787_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2038 a_32485_2773# a_32319_2773# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2039 vccd1 a_16180_3285# _208_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2040 a_28321_2550# input4.X a_28107_2550# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2041 vccd1 a_27038_3423# a_26965_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2042 a_19676_7093# _098_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2043 vssd1 a_12242_2767# a_12348_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2044 output25.A output19.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2045 a_7723_5161# _232_.CLK vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2046 a_2869_3087# _133_.A a_2511_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2047 vccd1 a_13069_2741# _233_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2048 _205_.A1 a_19106_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2049 _110_.Y output16.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2050 _121_.A a_4351_2223# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2051 vssd1 _196_.A a_11329_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2052 msb[11] a_8307_7127# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2053 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2054 vssd1 a_28015_4667# a_27973_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2055 vccd1 a_13445_2375# _203_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2056 vccd1 _215_.Q a_22983_2375# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2057 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2058 vssd1 a_28399_4943# a_28567_4917# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2059 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2060 vssd1 a_10340_2375# _149_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2061 vssd1 clkbuf_2_3__f_clk.A a_23478_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2062 a_19340_5263# _203_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2063 vccd1 a_12045_4087# a_11858_3829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2064 a_16578_4373# a_16371_4373# a_16754_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2065 _185_.X a_10719_3894# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2066 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X2067 a_6527_4373# _232_.CLK vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2068 vccd1 a_15738_2767# a_15844_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2069 a_11863_5639# _196_.A a_12037_5515# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2070 vccd1 output29.A output45.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2071 _180_.X a_15147_4427# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2072 vccd1 a_13327_4373# _193_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2073 vssd1 _179_.A1 _155_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2074 vssd1 _159_.X a_21244_3133# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2075 a_4622_4399# a_4307_4551# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2076 msb_n[14] a_3116_6549# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2077 output55.A output39.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2078 a_17911_4943# a_17213_4949# a_17654_4917# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2079 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2080 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X2081 vssd1 a_37519_5162# _119_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2082 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X2083 vssd1 a_17762_3855# a_17868_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2084 a_29518_2999# a_29614_2741# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2085 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2086 vssd1 a_4036_7093# msb[14] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2087 _141_.X a_22659_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2088 msb_n[8] a_12999_6575# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2089 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X2090 a_35373_2197# _160_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2091 a_33205_2375# _125_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2092 a_13545_4399# _206_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2093 a_16754_4765# a_16507_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2094 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2095 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2096 vccd1 a_25623_2491# a_25539_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2097 output17.A a_33535_3579# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2098 vssd1 a_6458_5461# a_6387_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2099 a_4403_4373# a_4694_4673# a_4645_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2100 a_25198_2335# a_25030_2589# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X2101 vccd1 a_26300_6549# msb_n[0] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2102 a_35373_2197# _160_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2103 _119_.A a_37011_4399# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2104 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2105 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X2106 a_27889_4943# _226_.D vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2107 vccd1 _125_.A1 a_35545_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2108 vssd1 output20.A a_31215_7127# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2109 a_11299_4399# a_11079_4399# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2110 vssd1 _241_.D a_14533_5321# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2111 output39.A a_18079_4917# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2112 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2113 a_20070_4399# _205_.B1 a_19901_4649# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2114 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2115 a_4772_7093# output48.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2116 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X2117 a_10659_4373# a_10950_4673# a_10901_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2118 vssd1 a_23478_2767# _222_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2119 llsb a_38023_6039# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2120 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2121 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2122 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X2123 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2124 vssd1 a_25623_4667# a_25581_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2125 _233_.CLK a_13069_2741# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2126 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2127 a_27215_4087# a_27488_4087# a_27446_4215# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2128 _093_.A a_33903_4667# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2129 vssd1 _125_.A1 _122_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2130 clkbuf_2_3__f_clk.A a_20442_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2131 a_19885_3855# a_19708_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2132 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2133 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2134 vssd1 output31.A _106_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2135 a_29495_3855# a_28713_3861# a_29411_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2136 vssd1 a_23047_4917# a_23005_5321# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2137 vssd1 a_12242_2223# a_12348_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2138 a_36399_4193# _162_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2139 a_11150_4373# a_10950_4673# a_11299_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2140 vssd1 a_20442_3311# clkbuf_2_3__f_clk.A vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2141 vccd1 _160_.X a_27853_2550# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2142 a_22356_4215# ANTENNA__177__A.DIODE a_22284_4215# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2143 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2144 a_16306_4399# a_15991_4551# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2145 a_24945_2223# _122_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2146 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X2147 vssd1 a_10483_5175# _195_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2148 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2149 a_15151_2589# a_14453_2223# a_14894_2335# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2150 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2151 a_29055_2388# dac_in[3] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2152 lsb[0] a_37471_7127# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2153 msb[6] a_17192_7093# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2154 output24.A output18.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2155 vccd1 a_23478_3855# _209_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2156 vssd1 _160_.X a_27853_2550# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2157 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
D21 vssd1 dac_in[9] sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
X2158 output56.A output40.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2159 _222_.CLK a_23478_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2160 a_32926_2741# a_32758_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2161 lsb[2] a_33844_7093# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2162 a_33386_3829# a_33218_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X2163 output51.A output35.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2164 a_22181_4949# a_22015_4949# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2165 a_6883_4399# a_6663_4399# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2166 a_24977_3677# a_24639_3463# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2167 a_16309_3311# _205_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2168 vccd1 a_10943_4373# a_10950_4673# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
D22 vssd1 _133_.A sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
X2169 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2170 a_32857_3311# _166_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2171 a_12045_4087# ANTENNA__177__A.DIODE vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2172 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2173 a_16925_4399# a_16378_4673# a_16578_4373# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2174 a_35061_4399# a_34895_4399# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2175 a_30531_2197# a_30822_2497# a_30773_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2176 a_9206_2767# a_8933_2773# a_9121_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2177 vccd1 _206_.A2 a_16309_3561# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2178 vccd1 a_23478_3855# _209_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2179 vccd1 _222_.CLK a_24591_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2180 msb_n[10] a_9411_7127# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2181 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X2182 vssd1 a_13069_3829# _232_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2183 a_25380_7093# output51.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2184 _165_.B a_35007_2806# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2185 a_16021_2767# a_15844_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2186 vccd1 _195_.X a_8277_5321# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2187 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2188 a_11497_4399# a_10943_4373# a_11150_4373# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2189 _233_.CLK a_13069_2741# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2190 _093_.A a_33903_4667# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2191 a_14650_3311# a_14335_3463# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2192 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2193 output55.A output39.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2194 a_14335_5309# a_14115_5321# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2195 output15.A _093_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2196 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2197 a_7093_2773# a_6927_2773# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2198 vccd1 a_27847_4765# a_28015_4667# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2199 vccd1 a_33183_2767# a_33351_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2200 vssd1 output42.A _102_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2201 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2202 a_26479_2388# dac_in[5] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2203 msb_n[5] a_17928_7093# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2204 _178_.A a_25635_3105# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2205 a_6734_4373# a_6534_4673# a_6883_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2206 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X2207 output17.A a_33535_3579# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2208 a_14115_5321# a_13986_5065# a_13695_5175# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2209 a_23849_2473# _133_.A _136_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2210 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2211 vssd1 a_23478_3855# _209_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2212 a_2869_3087# _179_.A1 a_2785_3087# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2213 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X2214 vssd1 a_33903_4667# a_33861_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2215 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2216 vccd1 a_30815_2197# a_30822_2497# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2217 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X2218 output48.A output32.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2219 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X2220 a_27956_7093# _115_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2221 vccd1 clkbuf_2_3__f_clk.A a_13069_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2222 a_12525_2223# a_12348_2223# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2223 a_17939_2223# _131_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2224 a_29112_4233# a_28713_3861# a_28986_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2225 a_10719_3894# _185_.A0 a_10719_4221# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2226 msb_n[15] a_1644_6549# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2227 a_32758_2767# a_32485_2773# a_32673_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2228 vssd1 a_7791_2767# a_7959_2741# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
D23 vssd1 ANTENNA__118__A.DIODE sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
X2229 vssd1 _185_.X a_12298_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2230 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X2231 _179_.A0 a_8399_2223# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2232 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2233 vssd1 dac_in[4] a_26431_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2234 a_2501_3311# _145_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2235 _110_.Y output16.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2236 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2237 _232_.CLK a_13069_3829# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2238 vccd1 a_10563_4551# output43.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2239 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X2240 vssd1 _149_.A1 a_3615_3087# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
D24 vssd1 ANTENNA__177__A.DIODE sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
X2241 a_18059_4399# _206_.A2 a_17965_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2242 a_28713_3861# a_28547_3861# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2243 vccd1 a_22068_7093# msb_n[3] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2244 output53.A output37.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2245 vssd1 a_6251_5461# a_6258_5761# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2246 a_6906_3677# a_6467_3311# a_6821_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2247 vccd1 a_9374_2741# a_9301_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2248 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X2249 a_22369_4943# _235_.D vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2250 a_23145_2223# _133_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2251 a_11150_4373# a_10943_4373# a_11326_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2252 a_27517_4765# a_26983_4399# a_27422_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2253 vssd1 _133_.A _133_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2254 a_15619_4221# _183_.A0 a_15256_4087# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2255 vssd1 a_27847_4765# a_28015_4667# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2256 a_16087_4373# a_16371_4373# a_16306_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2257 vssd1 a_13069_2741# _233_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2258 vssd1 _198_.A a_11010_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2259 vssd1 output30.A a_8307_7127# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2260 _115_.Y _115_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2261 vccd1 a_24639_3463# output37.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2262 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2263 vccd1 a_3116_6549# msb_n[14] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2264 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X2265 a_24735_3285# a_25026_3585# a_24977_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2266 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X2267 a_38163_2388# dummy vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2268 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2269 msb_n[3] a_22068_7093# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2270 vssd1 a_10021_2375# a_9834_2197# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2271 vccd1 _149_.B1 a_2511_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2272 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X2273 vccd1 a_12999_6575# msb_n[8] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2274 a_19426_5263# _205_.A1 a_19340_5263# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2275 vssd1 a_31267_2741# _131_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2276 a_33643_3855# a_32779_3861# a_33386_3829# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2277 output56.A output40.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2278 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2279 a_35129_3339# _168_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2280 vssd1 a_29411_3855# a_29579_3829# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2281 vssd1 _126_.X a_27488_4087# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2282 vccd1 a_18079_4917# a_17995_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2283 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2284 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2285 vssd1 output19.A output25.A vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2286 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2287 a_23431_3677# a_22567_3311# a_23174_3423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2288 a_7331_3677# a_6467_3311# a_7074_3423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2289 a_9301_2767# a_8767_2773# a_9206_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2290 vssd1 a_20890_3855# a_20996_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2291 vccd1 a_25455_4765# a_25623_4667# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2292 a_13069_2741# clkbuf_2_3__f_clk.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2293 vssd1 a_33386_3829# a_33344_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2294 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2295 vssd1 a_35502_4511# a_35460_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2296 a_11326_4765# a_11079_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2297 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2298 vssd1 _144_.A1 a_18703_3087# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2299 clkbuf_2_3__f_clk.A a_20442_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2300 a_6209_5853# a_5871_5639# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2301 a_5600_7093# output32.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2302 vccd1 a_24591_7127# msb[2] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2303 vssd1 output41.A output57.A vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2304 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X2305 a_19970_2767# a_19793_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2306 a_15738_2767# a_15561_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2307 a_25019_3285# _222_.CLK vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2308 vccd1 _195_.A a_7663_5487# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2309 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2310 a_23478_3855# clkbuf_2_3__f_clk.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2311 vssd1 a_25019_3285# a_25026_3585# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2312 vssd1 a_20442_3311# clkbuf_2_3__f_clk.A vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2313 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2314 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2315 lsb_n[3] a_31767_6575# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2316 vccd1 a_23478_3855# _209_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2317 vccd1 a_32926_2741# a_32853_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2318 msb[2] a_24591_7127# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2319 a_32367_5175# a_32463_5175# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2320 a_6734_4373# a_6527_4373# a_6910_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2321 _222_.CLK a_23478_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2322 _222_.CLK a_23478_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2323 vssd1 a_21454_4373# a_21383_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
D25 vssd1 ANTENNA__118__A.DIODE sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
X2324 a_35403_2550# _128_.B1 a_34944_2375# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2325 vccd1 _180_.B a_10839_2999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2326 a_5687_3463# ANTENNA__177__A.DIODE vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2327 vssd1 a_12794_3311# a_12900_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2328 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2329 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X2330 vssd1 a_35373_2197# a_35307_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2331 vccd1 a_17192_3285# _239_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2332 a_34702_4175# _125_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2333 vccd1 a_23599_3579# a_23515_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2334 vccd1 a_7499_3579# a_7415_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2335 a_34948_7093# output23.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2336 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X2337 a_31198_2589# a_30951_2223# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2338 a_11073_3133# _180_.B a_11001_3133# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2339 a_17836_4373# _241_.D a_17965_4649# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2340 vssd1 a_25455_4765# a_25623_4667# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2341 a_15235_2589# a_14453_2223# a_15151_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2342 vccd1 a_13459_7127# msb[8] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X2343 a_5241_4399# a_4694_4673# a_4894_4373# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2344 a_32853_2767# a_32319_2773# a_32758_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2345 vssd1 a_30441_3829# _128_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2346 vssd1 a_4307_4551# output30.A vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2347 a_30951_2223# a_30822_2497# a_30531_2197# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2348 vccd1 a_13069_2741# _233_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2349 vccd1 a_22097_3855# a_22197_3971# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2350 a_6910_4765# a_6663_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2351 a_26597_3311# a_26431_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2352 vccd1 output35.A output51.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2353 a_33183_2767# a_32485_2773# a_32926_2741# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2354 vssd1 a_11506_3311# a_11612_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2355 vccd1 a_33811_3829# a_33727_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2356 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X2357 vccd1 rst_n a_4351_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2358 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2359 vccd1 a_2288_7093# msb[15] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2360 vccd1 clkbuf_2_3__f_clk.A a_23478_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2361 vccd1 _149_.A2 a_11746_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2362 a_11079_4399# a_10950_4673# a_10659_4373# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2363 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2364 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X2365 a_11497_4399# a_10950_4673# a_11150_4373# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2366 vccd1 _093_.A a_38023_6039# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2367 vccd1 _149_.A1 _151_.C vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2368 vssd1 a_11987_7127# msb[9] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2369 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2370 a_6387_5487# a_6251_5461# a_5967_5461# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2371 vssd1 a_10563_4551# output43.A vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2372 a_33133_3855# _163_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2373 vssd1 output33.A _108_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2374 a_35249_4399# _169_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2375 a_7166_2335# a_6998_2589# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2376 a_17321_3561# _196_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2377 a_36236_6549# _110_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2378 a_20963_4373# a_21247_4373# a_21182_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2379 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X2380 vssd1 _133_.A a_2869_3087# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2381 vccd1 output31.A _106_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2382 vccd1 output29.A output45.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2383 vccd1 a_20442_3311# clkbuf_2_3__f_clk.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2384 vssd1 output17.A a_35631_7127# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2385 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2386 vccd1 a_27220_7093# msb[0] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2387 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X2388 msb[15] a_2288_7093# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2389 vccd1 a_7959_2741# a_7875_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2390 _166_.A a_35755_3339# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2391 vssd1 _209_.CLK a_32779_3861# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2392 vssd1 _209_.CLK a_34895_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2393 clkbuf_2_3__f_clk.A a_20442_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2394 a_29055_2388# dac_in[3] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2395 vccd1 a_28423_2999# _172_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2396 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X2397 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X2398 a_36424_3133# _125_.A1 a_36203_2806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2399 vssd1 a_20718_2197# a_20647_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2400 vccd1 a_32922_2375# a_32871_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2401 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X2402 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2403 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2404 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X2405 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2406 vccd1 _145_.A a_12065_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2407 a_31369_2223# a_30815_2197# a_31022_2197# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2408 vssd1 _233_.CLK a_6927_2773# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2409 vssd1 a_19602_3855# a_19708_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2410 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X2411 vccd1 _135_.X a_20713_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2412 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2413 a_36236_6549# _110_.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2414 a_31369_2223# a_30822_2497# a_31022_2197# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2415 a_6251_5461# _232_.CLK vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2416 a_20469_2589# a_20131_2375# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2417 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X2418 a_23478_2767# clkbuf_2_3__f_clk.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2419 _232_.CLK a_13069_3829# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2420 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X2421 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X2422 a_6243_4373# a_6534_4673# a_6485_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2423 a_6663_4399# a_6534_4673# a_6243_4373# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2424 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X2425 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2426 output16.A a_33811_3829# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2427 vccd1 _160_.X a_35221_2806# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2428 vccd1 a_16088_7093# msb_n[6] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2429 a_22097_3855# _140_.A_N vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2430 vccd1 output17.A output23.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2431 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2432 clkbuf_2_3__f_clk.A a_20442_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2433 output59.A output43.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2434 vssd1 output17.A output23.A vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2435 vssd1 _093_.A output15.A vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2436 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2437 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2438 vccd1 _196_.A a_11329_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2439 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X2440 vccd1 a_4894_4373# a_4823_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X2441 a_36203_2806# _125_.A1 a_36131_2806# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2442 a_27421_3311# a_26431_3311# a_27295_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2443 vccd1 _159_.A a_10289_3638# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2444 vssd1 a_15727_5175# _205_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2445 _141_.A a_22197_3971# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2446 vssd1 _140_.C a_22356_4215# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2447 a_29796_7093# _114_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2448 vccd1 a_22879_4943# a_23047_4917# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2449 vccd1 _135_.X a_23849_2473# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2450 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X2451 msb_n[6] a_16088_7093# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2452 _209_.CLK a_23478_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2453 vccd1 _241_.D a_17585_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2454 vccd1 output57.A a_14563_7127# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2455 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X2456 a_33367_3677# a_32669_3311# a_33110_3423# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2457 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X2458 a_27974_4943# a_27701_4949# a_27889_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2459 a_35221_2806# _164_.A0 a_35007_2806# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2460 vccd1 output32.A output48.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2461 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2462 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X2463 _145_.A a_11746_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2464 a_17556_2999# input7.X a_17698_2806# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2465 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X2466 vssd1 a_21247_4373# a_21254_4673# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2467 vccd1 _206_.A2 a_17321_3561# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2468 a_7343_5175# a_7439_5175# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2469 vccd1 a_18611_7127# msb[5] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2470 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2471 a_15727_5175# _192_.A a_15901_5281# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2472 _179_.A0 a_8399_2223# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2473 _126_.A a_25623_2491# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2474 vssd1 a_30120_2999# _133_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2475 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2476 vccd1 _196_.X a_2695_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
D26 vssd1 dac_in[6] sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
X2477 a_33267_2767# a_32485_2773# a_33183_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2478 a_31517_4221# _128_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2479 vccd1 a_23478_3855# _209_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2480 vssd1 output16.A _110_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2481 a_32705_4943# a_32367_5175# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2482 vssd1 a_13069_3829# _232_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2483 vccd1 output35.A a_26063_7127# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2484 a_22963_4943# a_22181_4949# a_22879_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2485 vccd1 a_23540_7093# msb_n[2] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2486 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X2487 vccd1 output37.A output53.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2488 a_15233_4427# _180_.A a_15147_4427# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2489 _233_.CLK a_13069_2741# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2490 _180_.B a_10075_3638# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2491 vccd1 output34.A output50.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2492 vssd1 _125_.A2 a_35437_4175# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2493 vssd1 _183_.X a_13445_2375# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2494 a_13599_5175# a_13695_5175# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2495 vssd1 output28.A _094_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2496 a_20647_2223# a_20511_2197# a_20227_2197# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2497 a_27249_2473# _133_.A _122_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2498 msb[5] a_18611_7127# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2499 a_12712_4399# _241_.D a_12409_4373# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2500 a_14453_2223# a_14287_2223# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2501 a_27038_3423# a_26870_3677# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2502 a_35755_3339# _162_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2503 vccd1 a_17836_4373# _238_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2504 a_38163_2388# dummy vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2505 a_27220_7093# output28.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2506 a_4687_4373# _232_.CLK vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2507 a_28035_2550# a_27853_2550# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2508 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2509 _162_.A a_19474_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2510 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2511 vccd1 output43.A a_11987_7127# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2512 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2513 vccd1 a_20131_2375# _135_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2514 a_21205_4765# a_20867_4551# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2515 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2516 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2517 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X2518 vssd1 output40.A output56.A vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2519 vccd1 output19.A output25.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2520 a_12242_2767# a_12065_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2521 vssd1 _165_.B a_35841_3339# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2522 a_20890_3855# a_20713_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2523 msb_n[7] a_14563_7127# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2524 vccd1 a_7423_2589# a_7591_2491# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2525 a_21023_2806# _215_.Q a_20951_2806# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2526 a_12525_2767# a_12348_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2527 vccd1 clkbuf_2_3__f_clk.A a_13069_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2528 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2529 a_27590_4511# a_27422_4765# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X2530 a_5357_2767# _155_.B1 _219_.D vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2531 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2532 a_29791_2388# _174_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2533 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2534 vssd1 _195_.A a_7663_5487# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2535 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X2536 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X2537 a_33225_4399# _157_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2538 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2539 a_22454_4943# a_22015_4949# a_22369_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2540 _171_.B a_28107_2550# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2541 vccd1 a_12242_2223# a_12348_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2542 _209_.CLK a_23478_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2543 vccd1 a_13979_5161# a_13986_5065# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2544 a_30441_3829# _128_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2545 a_17965_4649# _203_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2546 a_20511_2197# _222_.CLK vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2547 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2548 a_9374_2741# a_9206_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X2549 a_24945_2223# _122_.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2550 a_12037_5515# _196_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2551 vssd1 a_20511_2197# a_20518_2497# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2552 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2553 vccd1 a_16915_2197# ANTENNA__118__A.DIODE vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2554 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2555 msb[1] a_26063_7127# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2556 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2557 a_32883_5321# a_32747_5161# a_32463_5175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2558 vssd1 a_23478_2767# _222_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2559 a_33819_4765# a_33037_4399# a_33735_4765# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2560 vccd1 output39.A output55.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2561 a_19984_4399# _196_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2562 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X2563 vssd1 _156_.B a_37589_4193# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2564 vccd1 a_27215_4087# _129_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2565 a_17762_3855# a_17585_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2566 vssd1 _196_.B a_15561_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2567 vccd1 _160_.X a_34753_2806# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2568 vssd1 _205_.A2 a_13545_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2569 a_7993_4373# _149_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2570 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2571 vssd1 a_27956_7093# lsb_n[5] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X2572 _183_.A1 a_9799_2741# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2573 msb[9] a_11987_7127# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2574 a_22580_5321# a_22181_4949# a_22454_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2575 a_32463_5175# a_32747_5161# a_32682_5309# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2576 a_16371_4373# _232_.CLK vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2577 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2578 _151_.C _149_.B1 a_2585_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2579 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X2580 a_32485_2773# a_32319_2773# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2581 a_14335_3463# a_14431_3285# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2582 a_18035_2223# _144_.A1 a_17939_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2583 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2584 _233_.CLK a_13069_2741# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2585 vccd1 a_15256_4087# _183_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2586 lsb[1] a_35631_7127# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2587 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X2588 a_7723_5161# _232_.CLK vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2589 vccd1 _209_.CLK a_27535_4949# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2590 a_21383_4399# a_21247_4373# a_20963_4373# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2591 clkbuf_2_3__f_clk.A a_20442_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2592 a_22549_4943# a_22015_4949# a_22454_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2593 vssd1 dac_in[2] a_29743_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2594 vssd1 rst_n a_4351_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2595 vssd1 a_30435_2375# _134_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2596 vccd1 _169_.A a_34527_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2597 vccd1 _188_.X a_11497_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2598 _159_.X a_14287_4399# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2599 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2600 vssd1 a_32319_7127# lsb[3] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2601 vssd1 a_20442_3311# clkbuf_2_3__f_clk.A vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2602 vssd1 output37.A output53.A vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2603 vssd1 output42.A a_13459_7127# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2604 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X2605 vccd1 _148_.B1 a_3788_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2606 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X2607 _106_.Y output31.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2608 output45.A output29.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2609 vssd1 a_33183_2767# a_33351_2741# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2610 a_15256_4087# _183_.A1 a_15398_4221# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2611 vssd1 _199_.X a_8093_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2612 a_14715_3285# _232_.CLK vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2613 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X2614 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2615 a_27149_4399# a_26983_4399# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2616 a_27847_4765# a_26983_4399# a_27590_4511# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2617 a_17743_2197# _131_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2618 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X2619 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X2620 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X2621 vccd1 _135_.A a_20394_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2622 _145_.B ANTENNA__118__A.DIODE a_18703_3087# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2623 a_11857_4917# _196_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2624 vccd1 _185_.X a_12298_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2625 a_11023_2388# dac_in[8] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2626 a_28871_4564# _178_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2627 vssd1 a_13069_3829# _232_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2628 vccd1 a_28784_6549# lsb[5] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2629 a_21247_4373# _209_.CLK vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2630 a_27215_4087# a_27488_4087# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2631 a_10719_3894# _149_.B1 a_10647_3894# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2632 msb_n[12] a_6428_6549# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2633 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X2634 a_17213_4949# a_17047_4949# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2635 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X2636 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X2637 vssd1 _177_.B a_25721_3105# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2638 vssd1 a_31767_6575# lsb_n[3] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2639 a_28597_3105# _171_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2640 vccd1 a_27295_3677# a_27463_3579# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2641 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X2642 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X2643 a_9631_2767# a_8767_2773# a_9374_2741# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2644 vssd1 output43.A output59.A vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2645 vssd1 _151_.C a_5443_3087# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2646 a_3788_2767# _148_.B1 a_3615_3087# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2647 vccd1 _198_.A a_11010_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2648 vccd1 clkbuf_2_3__f_clk.A a_23478_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2649 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2650 vssd1 a_9374_2741# a_9332_3145# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2651 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2652 a_10839_2999# _185_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2653 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X2654 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2655 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X2656 a_24639_3463# a_24735_3285# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2657 vssd1 _222_.CLK a_22567_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2658 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2659 a_7081_4399# a_6534_4673# a_6734_4373# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2660 vssd1 _233_.CLK a_6467_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2661 a_4036_7093# output33.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2662 vccd1 a_7166_2335# a_7093_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2663 vssd1 a_6147_4551# output31.A vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2664 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X2665 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2666 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X2667 vccd1 a_19676_7093# msb_n[4] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2668 a_33068_3311# a_32669_3311# a_32942_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2669 vccd1 _180_.X a_17266_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2670 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X2671 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2672 a_16727_4399# a_16507_4399# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2673 a_13077_3311# a_12900_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2674 vccd1 _093_.A output15.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2675 a_28328_2223# _134_.A1 a_28107_2550# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2676 a_17192_3285# _205_.A1 a_17415_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2677 vssd1 a_34948_7093# lsb_n[1] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X2678 a_5687_3463# _151_.C vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2679 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2680 vssd1 _119_.X a_33301_5321# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2681 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2682 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2683 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2684 vssd1 a_11762_4087# a_11711_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2685 msb_n[4] a_19676_7093# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2686 a_17698_3133# _159_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2687 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X2688 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2689 a_28483_4943# a_27701_4949# a_28399_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2690 a_7093_2589# a_6559_2223# a_6998_2589# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2691 _164_.A0 a_34159_2223# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2692 a_3788_2767# _145_.A a_3697_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2693 vccd1 _172_.A a_26431_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2694 _201_.X a_18416_3561# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2695 a_24757_4399# a_24591_4399# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2696 vccd1 a_9799_2741# a_9715_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2697 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2698 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X2699 a_17743_2197# _135_.A a_18141_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2700 vssd1 a_33110_3423# a_33068_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2701 a_7859_5321# a_7723_5161# a_7439_5175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2702 a_16578_4373# a_16378_4673# a_16727_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2703 a_5921_3311# _149_.X a_5849_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2704 a_7746_4132# a_7539_4073# a_7922_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2705 a_22181_4949# a_22015_4949# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2706 _209_.CLK a_23478_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2707 lsb_n[0] a_36236_6549# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2708 _232_.CLK a_13069_3829# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2709 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X2710 vccd1 _102_.Y a_12999_6575# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2711 vccd1 a_12794_3311# a_12900_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2712 vssd1 a_37471_7127# lsb[0] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2713 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2714 vssd1 a_13069_2741# _233_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2715 vssd1 _125_.B1 _125_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2716 _135_.X a_20394_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2717 a_6458_5461# a_6251_5461# a_6634_5853# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2718 vccd1 output19.A a_32319_7127# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2719 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X2720 a_21244_3133# _215_.Q a_21023_2806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2721 a_16911_2986# dac_in[7] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2722 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2723 a_7922_3855# a_7675_4233# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2724 vccd1 a_13069_3829# _232_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2725 a_16925_4399# a_16371_4373# a_16578_4373# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2726 _174_.B a_27463_2806# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2727 vccd1 a_11506_3311# a_11612_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2728 vssd1 a_9411_7127# msb_n[10] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2729 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2730 a_13695_5175# a_13979_5161# a_13914_5309# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2731 vccd1 a_35373_2197# a_35403_2550# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2732 output18.A a_35927_4667# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2733 vssd1 _141_.A a_22659_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2734 _209_.CLK a_23478_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2735 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X2736 vccd1 a_7624_7093# msb_n[11] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2737 output25.A output19.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2738 vccd1 _192_.A a_15727_5175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2739 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X2740 vssd1 _102_.Y a_12999_6575# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2741 _119_.A a_37011_4399# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2742 vssd1 a_12409_4373# _188_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2743 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X2744 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X2745 vccd1 a_6734_4373# a_6663_4399# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X2746 a_29791_2388# _174_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2747 a_10839_2999# _121_.A a_11073_3133# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2748 a_6634_5853# a_6387_5487# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2749 a_7343_5175# a_7439_5175# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2750 vssd1 a_20442_3311# clkbuf_2_3__f_clk.A vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2751 a_33108_7093# output24.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2752 vccd1 _155_.A1 a_5357_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2753 _114_.Y output20.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2754 vssd1 a_19970_2767# a_20076_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2755 a_33103_5309# a_32883_5321# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2756 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X2757 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2758 vccd1 _205_.A1 a_19425_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2759 vccd1 a_23478_3855# _209_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2760 _241_.D a_17266_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2761 lsb_n[5] a_27956_7093# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2762 vssd1 _193_.X a_5241_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2763 vccd1 a_13069_2741# _233_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2764 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X2765 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2766 vccd1 a_25226_3285# a_25155_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X2767 vccd1 _152_.A a_5823_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2768 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2769 vccd1 _162_.A a_34955_3463# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2770 _148_.B1 _149_.A1 a_3146_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2771 a_28100_5321# a_27701_4949# a_27974_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2772 a_21173_3855# a_20996_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2773 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2774 a_14431_3285# a_14722_3585# a_14673_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2775 output55.A output39.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2776 a_8296_4399# _149_.A1 a_7993_4373# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2777 a_8999_4074# _199_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X2778 a_32669_3311# a_32503_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2779 vssd1 a_10147_7127# msb[10] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2780 a_25581_4399# a_24591_4399# a_25455_4765# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2781 a_28069_4943# a_27535_4949# a_27974_4943# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2782 vssd1 a_6835_7127# msb[12] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2783 vssd1 _222_.CLK a_32503_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2784 vssd1 a_33811_3829# a_33769_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2785 output18.A a_35927_4667# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2786 vccd1 a_25380_7093# msb_n[1] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2787 vssd1 _169_.A a_34527_4943# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2788 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2789 vccd1 a_23478_2767# _222_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2790 vccd1 a_31355_4087# _126_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2791 msb[8] a_13459_7127# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2792 _149_.B1 a_7959_2741# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2793 vccd1 a_7930_5220# a_7859_5321# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X2794 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X2795 a_15277_2223# a_14287_2223# a_15151_2589# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2796 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X2797 a_6186_5487# a_5871_5639# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2798 _215_.Q a_23599_3579# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2799 output29.A a_7499_3579# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2800 vccd1 a_6428_6549# msb_n[12] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2801 vssd1 a_22622_4917# a_22580_5321# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2802 a_25455_2589# a_24757_2223# a_25198_2335# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2803 vccd1 a_20442_3311# clkbuf_2_3__f_clk.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2804 msb[4] a_20504_7093# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2805 _159_.A a_1591_2223# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
D27 vssd1 ANTENNA__118__A.DIODE sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
X2806 output57.A output41.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2807 a_32945_3861# a_32779_3861# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2808 a_18045_3855# a_17868_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2809 a_13069_3829# clkbuf_2_3__f_clk.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2810 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X2811 clkbuf_2_3__f_clk.A a_20442_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2812 _233_.CLK a_13069_2741# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2813 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2814 a_7746_4132# a_7546_3977# a_7895_4221# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2815 vssd1 _195_.X a_8277_5321# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2816 vssd1 _133_.B a_22285_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2817 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X2818 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X2819 a_6805_5487# a_6258_5761# a_6458_5461# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2820 a_20346_5263# _205_.A1 a_20260_5263# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2821 vccd1 a_14715_3285# a_14722_3585# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2822 a_13608_2473# _192_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2823 _134_.X a_31480_3561# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2824 vccd1 _156_.B a_37503_4193# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2825 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X2826 vssd1 _239_.D a_16925_4399# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2827 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X2828 a_14726_2589# a_14453_2223# a_14641_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2829 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X2830 vccd1 output31.A _106_.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2831 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X2832 _205_.X a_20346_5263# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2833 a_4823_4399# a_4694_4673# a_4403_4373# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2834 a_25198_4511# a_25030_4765# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2835 vssd1 a_23478_2767# _222_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2836 vssd1 _162_.B a_36485_4193# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2837 a_30120_2999# _131_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2838 vssd1 a_22879_4943# a_23047_4917# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2839 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X2840 output20.A a_29579_3829# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2841 a_5043_4399# a_4823_4399# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2842 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X2843 vccd1 output16.A a_37471_7127# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2844 a_11023_2388# dac_in[8] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2845 vccd1 _159_.X a_19623_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2846 _209_.CLK a_23478_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2847 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2848 vccd1 a_9738_2375# a_9687_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2849 a_24954_3311# a_24639_3463# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2850 _232_.CLK a_13069_3829# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2851 vssd1 a_23478_2767# _222_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2852 vssd1 a_7746_4132# a_7675_4233# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2853 vccd1 a_7159_4087# output34.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2854 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
D28 vssd1 ANTENNA__177__A.DIODE sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
X2855 a_19602_3855# a_19425_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2856 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X2857 a_33861_4399# a_32871_4399# a_33735_4765# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2858 vccd1 output45.A a_9411_7127# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2859 vssd1 a_31215_7127# lsb[4] vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2860 a_10719_4221# a_10465_3894# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2861 vccd1 a_4772_7093# msb_n[13] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2862 lsb_n[1] a_34948_7093# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2863 vssd1 _160_.X a_35949_2806# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2864 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2865 vccd1 vssd1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X2866 vssd1 vccd1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X2867 vccd1 _159_.X a_10465_3894# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2868 a_23478_2767# clkbuf_2_3__f_clk.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2869 vccd1 a_13069_3829# _232_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2870 vssd1 _180_.B a_18243_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
C0 vccd1 _196_.X 6.62fF
C1 vccd1 _133_.A 3.83fF
C2 vccd1 _203_.A2 5.41fF
C3 vccd1 _121_.A 3.29fF
C4 vccd1 _190_.X 2.19fF
C5 vccd1 _196_.B 2.39fF
C6 vccd1 _131_.X 5.60fF
C7 vccd1 _145_.A 2.90fF
C8 vccd1 ANTENNA__177__A.DIODE 11.31fF
C9 vccd1 output33.A 2.21fF
C10 vccd1 output18.A 2.58fF
C11 vccd1 dac_in[5] 2.88fF
C12 vccd1 output37.A 2.59fF
C13 vccd1 dac_in[3] 2.38fF
C14 vccd1 output30.A 3.48fF
C15 vccd1 output28.A 2.21fF
C16 vccd1 _160_.X 4.90fF
C17 vccd1 input3.X 2.97fF
C18 vccd1 output19.A 2.18fF
C19 vccd1 _209_.CLK 5.33fF
C20 vccd1 clk 3.53fF
C21 vccd1 _222_.CLK 3.92fF
C22 vccd1 _206_.A2 2.02fF
C23 _149_.A1 _179_.A1 2.07fF
C24 vccd1 _232_.CLK 4.34fF
C25 vccd1 output29.A 2.33fF
C26 vccd1 output16.A 2.33fF
C27 vccd1 _162_.A 4.77fF
C28 vccd1 _133_.B 3.22fF
C29 vccd1 _233_.CLK 5.38fF
C30 vccd1 _159_.X 4.39fF
C31 vccd1 _149_.A2 2.39fF
C32 vccd1 _125_.A2 3.33fF
C33 vccd1 clkbuf_2_3__f_clk.A 3.09fF
C34 vccd1 ANTENNA__118__A.DIODE 8.79fF
C35 vccd1 _205_.A2 4.46fF
C36 _162_.A _222_.CLK 2.35fF
C37 _196_.B _203_.A2 2.25fF
C38 vccd1 _140_.A_N 3.06fF
C39 vccd1 _180_.B 2.61fF
C40 vccd1 _126_.X 2.89fF
C41 dac_in[8] vssd1 2.19fF
C42 input6.X vssd1 2.35fF $ **FLOATING
C43 _217_.D vssd1 2.93fF $ **FLOATING
C44 dac_in[5] vssd1 3.30fF
C45 _215_.Q vssd1 2.76fF $ **FLOATING
C46 _222_.CLK vssd1 2.59fF $ **FLOATING
C47 _160_.X vssd1 4.32fF $ **FLOATING
C48 _126_.A vssd1 2.20fF $ **FLOATING
C49 _125_.A1 vssd1 3.32fF $ **FLOATING
C50 _128_.B1 vssd1 3.78fF $ **FLOATING
C51 _183_.A1 vssd1 2.73fF $ **FLOATING
C52 clkbuf_2_3__f_clk.A vssd1 6.28fF $ **FLOATING
C53 _233_.CLK vssd1 2.05fF $ **FLOATING
C54 _157_.X vssd1 2.09fF $ **FLOATING
C55 _133_.A vssd1 15.42fF $ **FLOATING
C56 _180_.B vssd1 2.44fF $ **FLOATING
C57 _180_.A vssd1 3.56fF $ **FLOATING
C58 _159_.X vssd1 2.30fF $ **FLOATING
C59 _159_.A vssd1 4.09fF $ **FLOATING
C60 _149_.A1 vssd1 4.90fF $ **FLOATING
C61 _193_.X vssd1 3.55fF $ **FLOATING
C62 ANTENNA__177__A.DIODE vssd1 4.23fF $ **FLOATING
C63 _209_.CLK vssd1 4.48fF $ **FLOATING
C64 _205_.A2 vssd1 2.48fF $ **FLOATING
C65 ANTENNA__118__A.DIODE vssd1 2.87fF $ **FLOATING
C66 _196_.A vssd1 3.13fF $ **FLOATING
C67 _196_.B vssd1 2.93fF $ **FLOATING
C68 _232_.CLK vssd1 3.63fF $ **FLOATING
C69 _232_.D vssd1 2.24fF $ **FLOATING
C70 output28.A vssd1 2.24fF $ **FLOATING
C71 output34.A vssd1 2.13fF $ **FLOATING
C72 vccd1 vssd1 858.36fF
.ends
