magic
tech sky130A
magscale 1 2
timestamp 1672468680
<< pwell >>
rect 1063 558 2009 3120
<< psubdiff >>
rect 1099 3050 1223 3084
rect 1429 3050 1643 3084
rect 1849 3050 1973 3084
rect 1099 2960 1133 3050
rect 1519 2960 1553 3050
rect 1099 628 1133 718
rect 1519 628 1553 718
rect 1939 628 1973 3050
rect 1099 594 1195 628
rect 1457 594 1615 628
rect 1877 594 1973 628
<< psubdiffcont >>
rect 1223 3050 1429 3084
rect 1643 3050 1849 3084
rect 1099 718 1133 2960
rect 1519 718 1553 2960
rect 1195 594 1457 628
rect 1615 594 1877 628
<< xpolycontact >>
rect 1257 2522 1395 2954
rect 1257 1990 1395 2422
rect 1677 2522 1815 2954
rect 1677 1990 1815 2422
<< ppolyres >>
rect 1257 2422 1395 2522
rect 1677 2422 1815 2522
<< locali >>
rect 1099 3050 1223 3084
rect 1429 3050 1445 3084
rect 1519 3050 1643 3084
rect 1849 3050 1865 3084
rect 1099 2960 1133 3050
rect 1519 2960 1553 3050
rect 1133 2954 1167 2960
rect 1553 2954 1587 2960
rect 1155 724 1167 2954
rect 1133 718 1167 724
rect 1575 724 1587 2954
rect 1553 718 1587 724
rect 1099 628 1133 718
rect 1519 628 1553 718
rect 1099 594 1195 628
rect 1457 594 1473 628
rect 1519 594 1615 628
rect 1877 594 1893 628
<< viali >>
rect 1111 724 1133 2954
rect 1133 724 1155 2954
rect 1273 2539 1379 2936
rect 1273 2008 1379 2405
rect 1531 724 1553 2954
rect 1553 724 1575 2954
rect 1693 2539 1799 2936
rect 1693 2008 1799 2405
<< metal1 >>
rect 1099 2954 1220 2960
rect 1519 2954 1640 2960
rect 1099 724 1111 2954
rect 1155 2950 1220 2954
rect 1155 2810 1160 2950
rect 1155 2800 1220 2810
rect 1257 2936 1395 2954
rect 1155 1868 1167 2800
rect 1257 2539 1273 2936
rect 1379 2539 1395 2936
rect 1257 2527 1395 2539
rect 1250 2410 1400 2420
rect 1250 2000 1260 2410
rect 1390 2000 1400 2410
rect 1250 1990 1400 2000
rect 1303 1980 1349 1990
rect 1155 724 1170 1868
rect 1099 718 1170 724
rect 1519 724 1531 2954
rect 1575 2950 1640 2954
rect 1575 2810 1580 2950
rect 1575 2800 1640 2810
rect 1677 2936 1815 2954
rect 1575 1868 1587 2800
rect 1677 2610 1693 2936
rect 1677 2550 1690 2610
rect 1677 2539 1693 2550
rect 1799 2610 1815 2936
rect 1800 2550 1815 2610
rect 1799 2539 1815 2550
rect 1677 2527 1815 2539
rect 1670 2410 1820 2420
rect 1670 2000 1680 2410
rect 1810 2000 1820 2410
rect 1670 1990 1820 2000
rect 1723 1980 1769 1990
rect 1575 724 1590 1868
rect 1519 718 1590 724
<< via1 >>
rect 1160 2810 1220 2950
rect 1273 2539 1379 2936
rect 1260 2405 1390 2410
rect 1260 2008 1273 2405
rect 1273 2008 1379 2405
rect 1379 2008 1390 2405
rect 1260 2000 1390 2008
rect 1580 2810 1640 2950
rect 1690 2550 1693 2610
rect 1693 2539 1799 2936
rect 1799 2550 1800 2610
rect 1680 2405 1810 2410
rect 1680 2008 1693 2405
rect 1693 2008 1799 2405
rect 1799 2008 1810 2405
rect 1680 2000 1810 2008
<< metal2 >>
rect 1150 3190 1230 3200
rect 1150 3130 1160 3190
rect 1220 3130 1230 3190
rect 1150 3120 1230 3130
rect 1570 3190 1650 3200
rect 1570 3130 1580 3190
rect 1640 3130 1650 3190
rect 1570 3120 1650 3130
rect 1160 2950 1220 3120
rect 1160 2800 1220 2810
rect 1257 2936 1395 2954
rect 1257 2610 1273 2936
rect 1379 2620 1395 2936
rect 1580 2950 1640 3120
rect 1580 2800 1640 2810
rect 1677 2936 1815 2954
rect 1677 2620 1693 2936
rect 1379 2610 1693 2620
rect 1799 2610 1815 2936
rect 1257 2550 1270 2610
rect 1380 2550 1690 2610
rect 1800 2550 1815 2610
rect 1257 2539 1273 2550
rect 1379 2539 1693 2550
rect 1799 2539 1815 2550
rect 1257 2530 1815 2539
rect 1257 2527 1395 2530
rect 1677 2527 1815 2530
rect 1250 2410 1400 2420
rect 1670 2410 1820 2420
rect 1250 2000 1260 2410
rect 1390 2320 1680 2410
rect 1390 2000 1400 2320
rect 1250 1990 1400 2000
rect 1670 2000 1680 2320
rect 1810 2000 1820 2410
rect 1670 1990 1820 2000
<< via2 >>
rect 1160 3130 1220 3190
rect 1580 3130 1640 3190
rect 1270 2550 1273 2610
rect 1273 2550 1379 2610
rect 1379 2550 1380 2610
rect 1690 2340 1800 2400
<< metal3 >>
rect 1060 3290 2010 3370
rect 1060 3190 2010 3200
rect 1060 3130 1160 3190
rect 1220 3130 1580 3190
rect 1640 3130 2010 3190
rect 1060 3120 2010 3130
rect 1060 2610 1390 2620
rect 1060 2550 1270 2610
rect 1380 2550 1390 2610
rect 1060 2540 1390 2550
rect 1830 2540 2010 2620
rect 1830 2410 1910 2540
rect 1680 2400 1910 2410
rect 1680 2340 1690 2400
rect 1800 2340 1910 2400
rect 1680 2330 1910 2340
<< comment >>
rect 1099 2960 1133 3084
rect 1519 2960 1553 3084
rect 1099 594 1133 718
rect 1519 594 1553 718
<< labels >>
rlabel metal3 1520 3120 1560 3200 1 VSUB
port 4 n
rlabel metal3 1940 3120 1980 3200 1 VSUB
port 4 n
rlabel metal3 1990 2540 2010 2620 1 IN
port 5 n
rlabel metal3 1060 2540 1080 2620 1 IO1
port 6 n
<< end >>
