magic
tech sky130A
magscale 1 2
timestamp 1670808485
<< nwell >>
rect 1066 6789 18898 7355
rect 1066 5701 18898 6267
rect 1066 4613 18898 5179
rect 1066 3525 18898 4091
rect 1066 2437 18898 3003
<< pwell >>
rect 1133 7595 1167 7633
rect 1411 7604 1443 7626
rect 1869 7595 1903 7633
rect 1961 7595 1995 7633
rect 3065 7595 3099 7633
rect 3616 7605 3640 7627
rect 3803 7604 3835 7626
rect 4261 7595 4295 7633
rect 4353 7595 4387 7633
rect 5459 7604 5491 7626
rect 5917 7595 5951 7633
rect 6009 7595 6043 7633
rect 6377 7595 6411 7633
rect 7481 7595 7515 7633
rect 7849 7595 7883 7633
rect 8217 7595 8251 7633
rect 8768 7605 8792 7627
rect 8953 7595 8987 7633
rect 9597 7603 9631 7633
rect 1105 7433 1379 7595
rect 1565 7459 1931 7595
rect 1565 7413 1834 7459
rect 1933 7433 3035 7595
rect 3037 7433 3587 7595
rect 3683 7421 3769 7578
rect 3957 7459 4323 7595
rect 3957 7413 4226 7459
rect 4325 7433 5427 7595
rect 5613 7459 5979 7595
rect 5613 7413 5882 7459
rect 5981 7433 6255 7595
rect 6259 7421 6345 7578
rect 6349 7433 7451 7595
rect 7453 7433 7819 7595
rect 7821 7459 8187 7595
rect 7918 7413 8187 7459
rect 8189 7433 8739 7595
rect 8835 7421 8921 7578
rect 8925 7433 9475 7595
rect 9477 7413 9655 7603
rect 9689 7595 9723 7633
rect 10057 7595 10091 7633
rect 10425 7595 10459 7633
rect 11161 7595 11195 7633
rect 11529 7595 11563 7633
rect 12265 7595 12299 7633
rect 12633 7595 12667 7633
rect 13737 7595 13771 7633
rect 14105 7595 14139 7633
rect 14473 7595 14507 7633
rect 14841 7595 14875 7633
rect 15945 7595 15979 7633
rect 16496 7605 16520 7627
rect 16683 7604 16715 7626
rect 16865 7595 16899 7633
rect 17233 7595 17267 7633
rect 17968 7605 17992 7627
rect 18061 7595 18095 7633
rect 18431 7604 18463 7626
rect 18797 7595 18831 7633
rect 9661 7433 10027 7595
rect 10029 7459 10395 7595
rect 10397 7433 11131 7595
rect 11133 7433 11407 7595
rect 11411 7421 11497 7578
rect 11501 7433 12235 7595
rect 12237 7459 12603 7595
rect 12334 7413 12603 7459
rect 12605 7433 13707 7595
rect 13709 7433 13983 7595
rect 13987 7421 14073 7578
rect 14077 7433 14443 7595
rect 14445 7459 14811 7595
rect 14542 7413 14811 7459
rect 14813 7433 15915 7595
rect 15917 7433 16467 7595
rect 16563 7421 16649 7578
rect 16837 7459 17203 7595
rect 16934 7413 17203 7459
rect 17205 7433 17939 7595
rect 18033 7459 18399 7595
rect 18130 7413 18399 7459
rect 18585 7433 18859 7595
rect 1105 6549 1379 6711
rect 1381 6549 2483 6711
rect 2485 6549 3587 6711
rect 3683 6566 3769 6723
rect 3773 6549 4875 6711
rect 4877 6549 5979 6711
rect 5981 6549 7083 6711
rect 7085 6549 8187 6711
rect 8189 6549 8739 6711
rect 8835 6566 8921 6723
rect 8925 6549 10027 6711
rect 10029 6549 11131 6711
rect 11133 6549 12235 6711
rect 12237 6549 13339 6711
rect 13341 6549 13891 6711
rect 13987 6566 14073 6723
rect 14077 6549 15179 6711
rect 15181 6549 16283 6711
rect 16285 6549 17387 6711
rect 17389 6549 18491 6711
rect 18585 6549 18859 6711
rect 1133 6507 1167 6549
rect 1409 6507 1443 6549
rect 2513 6507 2547 6549
rect 3617 6539 3651 6545
rect 3616 6517 3651 6539
rect 3617 6507 3651 6517
rect 3801 6511 3835 6549
rect 4721 6507 4755 6545
rect 4905 6511 4939 6549
rect 5825 6507 5859 6545
rect 6009 6511 6043 6549
rect 6192 6517 6216 6539
rect 6377 6507 6411 6545
rect 7113 6511 7147 6549
rect 7481 6507 7515 6545
rect 8217 6511 8251 6549
rect 8585 6507 8619 6545
rect 8768 6517 8792 6539
rect 8953 6511 8987 6549
rect 9689 6507 9723 6545
rect 10057 6511 10091 6549
rect 10793 6507 10827 6545
rect 11161 6511 11195 6549
rect 11344 6517 11368 6539
rect 11529 6507 11563 6545
rect 12265 6511 12299 6549
rect 12633 6507 12667 6545
rect 13369 6511 13403 6549
rect 13737 6507 13771 6545
rect 13920 6517 13944 6539
rect 14105 6511 14139 6549
rect 14841 6507 14875 6545
rect 15209 6511 15243 6549
rect 15945 6507 15979 6545
rect 16313 6511 16347 6549
rect 16496 6517 16520 6539
rect 16681 6507 16715 6545
rect 17417 6511 17451 6549
rect 17785 6507 17819 6545
rect 18520 6517 18544 6539
rect 18797 6507 18831 6549
rect 1105 6345 1379 6507
rect 1381 6345 2483 6507
rect 2485 6345 3587 6507
rect 3589 6345 4691 6507
rect 4693 6345 5795 6507
rect 5797 6345 6163 6507
rect 6259 6333 6345 6490
rect 6349 6345 7451 6507
rect 7453 6345 8555 6507
rect 8557 6345 9659 6507
rect 9661 6345 10763 6507
rect 10765 6345 11315 6507
rect 11411 6333 11497 6490
rect 11501 6345 12603 6507
rect 12605 6345 13707 6507
rect 13709 6345 14811 6507
rect 14813 6345 15915 6507
rect 15917 6345 16467 6507
rect 16563 6333 16649 6490
rect 16653 6345 17755 6507
rect 17757 6345 18491 6507
rect 18585 6345 18859 6507
rect 1105 5461 1379 5623
rect 1381 5461 2115 5623
rect 2209 5461 2483 5617
rect 2485 5461 3035 5623
rect 3037 5461 3311 5617
rect 3313 5461 3679 5623
rect 3683 5478 3769 5635
rect 3773 5461 4875 5623
rect 4877 5461 5979 5623
rect 5981 5461 6715 5623
rect 6717 5597 6903 5643
rect 6717 5461 7497 5597
rect 7545 5461 8647 5623
rect 8835 5478 8921 5635
rect 8925 5461 9659 5623
rect 9845 5597 10031 5643
rect 11081 5625 11271 5643
rect 9845 5461 10625 5597
rect 10673 5461 11039 5623
rect 11081 5461 11467 5625
rect 11501 5461 12235 5623
rect 12237 5597 12423 5643
rect 12237 5461 13017 5597
rect 13065 5461 13799 5623
rect 13987 5478 14073 5635
rect 14261 5597 14447 5643
rect 14261 5461 15041 5597
rect 15089 5461 16191 5623
rect 16193 5461 17295 5623
rect 17297 5461 18399 5623
rect 18585 5461 18859 5623
rect 1133 5419 1167 5461
rect 1409 5419 1443 5461
rect 2144 5429 2168 5451
rect 2237 5423 2271 5461
rect 2329 5423 2363 5457
rect 2329 5419 2359 5423
rect 2421 5419 2455 5457
rect 2513 5423 2547 5461
rect 2788 5429 2812 5451
rect 3249 5423 3283 5461
rect 3249 5419 3279 5423
rect 3341 5419 3375 5461
rect 3709 5419 3743 5457
rect 3801 5423 3835 5461
rect 4077 5419 4111 5457
rect 4445 5419 4479 5457
rect 4721 5419 4755 5457
rect 4905 5423 4939 5461
rect 6009 5419 6043 5461
rect 6103 5428 6135 5450
rect 6377 5419 6411 5457
rect 6708 5419 6742 5457
rect 6800 5423 6834 5461
rect 7481 5419 7515 5457
rect 7573 5423 7607 5461
rect 7904 5419 7938 5457
rect 8677 5419 8711 5457
rect 8953 5423 8987 5461
rect 9044 5429 9068 5451
rect 9137 5419 9171 5457
rect 9689 5419 9723 5457
rect 9928 5423 9962 5461
rect 10480 5419 10514 5457
rect 10701 5423 10735 5461
rect 11437 5457 11467 5461
rect 11255 5428 11287 5450
rect 11437 5423 11471 5457
rect 11529 5419 11563 5461
rect 12320 5423 12354 5461
rect 12633 5419 12667 5457
rect 13000 5429 13024 5451
rect 13093 5423 13127 5461
rect 13148 5419 13182 5457
rect 13831 5430 13863 5452
rect 13921 5419 13955 5457
rect 14107 5430 14139 5452
rect 14344 5423 14378 5461
rect 15025 5419 15059 5457
rect 15117 5423 15151 5461
rect 16129 5419 16163 5457
rect 16221 5423 16255 5461
rect 16496 5429 16520 5451
rect 16681 5419 16715 5457
rect 17325 5423 17359 5461
rect 17785 5419 17819 5457
rect 18431 5430 18463 5452
rect 18520 5429 18544 5451
rect 18797 5419 18831 5461
rect 1105 5257 1379 5419
rect 1381 5257 1931 5419
rect 1973 5255 2359 5419
rect 2393 5257 2759 5419
rect 2893 5255 3279 5419
rect 3313 5257 3679 5419
rect 3681 5283 4047 5419
rect 1973 5237 2163 5255
rect 2893 5237 3083 5255
rect 3778 5237 4047 5283
rect 4049 5257 4415 5419
rect 4419 5237 4689 5419
rect 4693 5257 5795 5419
rect 5797 5263 6071 5419
rect 6259 5245 6345 5402
rect 6349 5257 6623 5419
rect 6625 5283 7405 5419
rect 6625 5237 6811 5283
rect 7453 5257 7819 5419
rect 7821 5283 8601 5419
rect 7821 5237 8007 5283
rect 8649 5257 9015 5419
rect 9109 5237 9659 5419
rect 9661 5257 10395 5419
rect 10397 5283 11177 5419
rect 10397 5237 10583 5283
rect 11411 5245 11497 5402
rect 11501 5257 12603 5419
rect 12605 5257 12971 5419
rect 13065 5283 13845 5419
rect 13065 5237 13251 5283
rect 13893 5257 14995 5419
rect 14997 5257 16099 5419
rect 16101 5257 16467 5419
rect 16563 5245 16649 5402
rect 16653 5257 17755 5419
rect 17757 5257 18491 5419
rect 18585 5257 18859 5419
rect 1105 4373 1379 4535
rect 1381 4373 1931 4535
rect 2728 4509 2910 4553
rect 3217 4509 3487 4555
rect 2025 4373 3487 4509
rect 3683 4390 3769 4547
rect 3997 4537 4187 4555
rect 3997 4373 4383 4537
rect 4417 4373 4783 4535
rect 4877 4373 5427 4555
rect 5429 4373 5795 4535
rect 5797 4373 6347 4555
rect 6349 4373 6715 4535
rect 7420 4509 7602 4553
rect 7909 4509 8179 4555
rect 6717 4373 8179 4509
rect 8189 4373 8739 4535
rect 8835 4390 8921 4547
rect 8925 4373 9659 4535
rect 9661 4373 9935 4535
rect 9945 4509 10215 4555
rect 10522 4509 10704 4553
rect 9945 4373 11407 4509
rect 11409 4373 11775 4535
rect 11777 4373 12327 4555
rect 12329 4373 12695 4535
rect 12697 4373 13247 4555
rect 13249 4373 13983 4535
rect 13987 4390 14073 4547
rect 14581 4537 14771 4555
rect 14077 4373 14351 4535
rect 14385 4373 14771 4537
rect 14813 4373 15915 4535
rect 15917 4373 17019 4535
rect 17021 4373 18123 4535
rect 18125 4373 18491 4535
rect 18585 4373 18859 4535
rect 1133 4331 1167 4373
rect 1409 4331 1443 4373
rect 1961 4363 1995 4369
rect 1960 4341 1995 4363
rect 1961 4331 1995 4341
rect 2053 4335 2087 4373
rect 4353 4369 4383 4373
rect 2237 4331 2271 4369
rect 3527 4342 3559 4364
rect 3803 4342 3835 4364
rect 3985 4331 4019 4369
rect 4077 4331 4111 4369
rect 4353 4335 4387 4369
rect 4445 4335 4479 4373
rect 4812 4341 4836 4363
rect 4905 4335 4939 4373
rect 5457 4335 5491 4373
rect 5825 4335 5859 4373
rect 6009 4331 6043 4369
rect 6103 4340 6135 4362
rect 6377 4331 6411 4373
rect 6745 4335 6779 4373
rect 6929 4331 6963 4369
rect 7481 4331 7515 4369
rect 7849 4331 7883 4369
rect 8217 4335 8251 4373
rect 8768 4341 8792 4363
rect 8953 4335 8987 4373
rect 9689 4331 9723 4373
rect 10424 4341 10448 4363
rect 10517 4331 10551 4369
rect 11069 4331 11103 4369
rect 11345 4335 11379 4373
rect 11437 4335 11471 4373
rect 11531 4340 11563 4362
rect 11713 4331 11747 4369
rect 11805 4335 11839 4373
rect 12357 4335 12391 4373
rect 12725 4335 12759 4373
rect 13185 4331 13219 4369
rect 13277 4335 13311 4373
rect 14105 4335 14139 4373
rect 14385 4369 14415 4373
rect 14289 4331 14323 4369
rect 14381 4335 14415 4369
rect 14841 4335 14875 4373
rect 15392 4341 15416 4363
rect 15669 4331 15703 4369
rect 15761 4331 15795 4369
rect 15945 4335 15979 4373
rect 16496 4341 16520 4363
rect 16683 4340 16715 4362
rect 16865 4335 16899 4369
rect 17049 4335 17083 4373
rect 16869 4331 16899 4335
rect 17325 4331 17359 4369
rect 18153 4335 18187 4373
rect 18431 4340 18463 4362
rect 18520 4341 18544 4363
rect 18797 4331 18831 4373
rect 1105 4169 1379 4331
rect 1381 4169 1931 4331
rect 1933 4175 2207 4331
rect 2209 4169 2575 4331
rect 2585 4195 4047 4331
rect 2585 4149 2855 4195
rect 3162 4151 3344 4195
rect 4049 4169 4599 4331
rect 4609 4195 6071 4331
rect 4609 4149 4879 4195
rect 5186 4151 5368 4195
rect 6259 4157 6345 4314
rect 6349 4169 6899 4331
rect 6901 4149 7451 4331
rect 7453 4169 7819 4331
rect 7821 4195 9642 4331
rect 9661 4169 10395 4331
rect 10489 4149 11039 4331
rect 11041 4169 11407 4331
rect 11411 4157 11497 4314
rect 11685 4195 13147 4331
rect 12388 4151 12570 4195
rect 12877 4149 13147 4195
rect 13157 4169 14259 4331
rect 14261 4169 15363 4331
rect 15457 4175 15731 4331
rect 15733 4169 16467 4331
rect 16563 4157 16649 4314
rect 16869 4167 17255 4331
rect 17297 4169 18399 4331
rect 18585 4169 18859 4331
rect 17065 4149 17255 4167
rect 1105 3285 1379 3447
rect 1381 3285 1931 3447
rect 2728 3421 2910 3465
rect 3217 3421 3487 3467
rect 2025 3285 3487 3421
rect 3683 3302 3769 3459
rect 4660 3421 4842 3465
rect 5149 3421 5419 3467
rect 3957 3285 5419 3421
rect 5429 3285 6163 3447
rect 6257 3285 6807 3467
rect 6809 3285 7175 3447
rect 7880 3421 8062 3465
rect 8369 3421 8639 3467
rect 7177 3285 8639 3421
rect 8835 3302 8921 3459
rect 8925 3285 9659 3447
rect 10456 3421 10638 3465
rect 10945 3421 11215 3467
rect 9753 3285 11215 3421
rect 11225 3285 11775 3447
rect 12480 3421 12662 3465
rect 12969 3421 13239 3467
rect 11777 3285 13239 3421
rect 13249 3285 13983 3447
rect 13987 3302 14073 3459
rect 16417 3449 16607 3467
rect 17245 3449 17435 3467
rect 14077 3285 15179 3447
rect 15181 3285 15731 3447
rect 15733 3285 16007 3441
rect 16009 3285 16375 3447
rect 16417 3285 16803 3449
rect 16837 3285 17203 3447
rect 17245 3285 17631 3449
rect 17665 3285 18399 3447
rect 18585 3285 18859 3447
rect 1133 3243 1167 3285
rect 1409 3243 1443 3285
rect 1776 3253 1800 3275
rect 1869 3243 1903 3281
rect 1960 3253 1984 3275
rect 2053 3247 2087 3285
rect 2237 3243 2271 3281
rect 3527 3254 3559 3276
rect 3803 3254 3835 3276
rect 3985 3247 4019 3285
rect 4353 3243 4387 3281
rect 4445 3243 4479 3281
rect 5457 3247 5491 3285
rect 5549 3243 5583 3281
rect 6192 3253 6216 3275
rect 6285 3247 6319 3285
rect 6377 3243 6411 3281
rect 6837 3247 6871 3285
rect 7112 3253 7136 3275
rect 7205 3251 7239 3285
rect 7297 3251 7331 3281
rect 1105 3081 1379 3243
rect 1381 3081 1747 3243
rect 1841 3107 2207 3243
rect 2209 3081 2575 3243
rect 2594 3107 4415 3243
rect 4417 3081 5519 3243
rect 5521 3081 6255 3243
rect 6259 3069 6345 3226
rect 6349 3081 7083 3243
rect 7177 3061 7355 3251
rect 7389 3243 7423 3281
rect 7757 3243 7791 3281
rect 8679 3254 8711 3276
rect 8953 3247 8987 3285
rect 9597 3243 9631 3281
rect 9688 3253 9712 3275
rect 9781 3247 9815 3285
rect 10701 3243 10735 3281
rect 11253 3247 11287 3285
rect 11531 3252 11563 3274
rect 11713 3243 11747 3281
rect 11805 3247 11839 3285
rect 13185 3243 13219 3281
rect 13277 3247 13311 3285
rect 14105 3247 14139 3285
rect 14289 3243 14323 3281
rect 15209 3247 15243 3285
rect 15393 3243 15427 3281
rect 15945 3247 15979 3285
rect 16037 3247 16071 3285
rect 16773 3281 16803 3285
rect 16496 3253 16520 3275
rect 16683 3252 16715 3274
rect 16773 3247 16807 3281
rect 16865 3247 16899 3285
rect 17601 3281 17631 3285
rect 17049 3243 17083 3281
rect 17141 3243 17175 3281
rect 17601 3247 17635 3281
rect 17693 3247 17727 3285
rect 18245 3243 18279 3281
rect 18431 3254 18463 3276
rect 18797 3243 18831 3285
rect 7361 3081 7727 3243
rect 7729 3107 9550 3243
rect 9569 3081 10671 3243
rect 10673 3081 11407 3243
rect 11411 3069 11497 3226
rect 11685 3107 13147 3243
rect 12388 3063 12570 3107
rect 12877 3061 13147 3107
rect 13157 3081 14259 3243
rect 14261 3081 15363 3243
rect 15365 3081 16467 3243
rect 16563 3069 16649 3226
rect 16837 3087 17111 3243
rect 17113 3081 18215 3243
rect 18217 3081 18583 3243
rect 18585 3081 18859 3243
rect 1105 2197 1379 2359
rect 1381 2197 1931 2359
rect 2033 2333 2303 2379
rect 2610 2333 2792 2377
rect 2033 2197 3495 2333
rect 3683 2214 3769 2371
rect 1133 2159 1167 2197
rect 1409 2159 1443 2197
rect 1960 2165 1984 2187
rect 3433 2159 3467 2197
rect 3957 2189 4135 2379
rect 4141 2197 4507 2359
rect 5304 2333 5486 2377
rect 5793 2333 6063 2379
rect 4601 2197 6063 2333
rect 6259 2214 6345 2371
rect 6349 2197 7083 2359
rect 7185 2333 7455 2379
rect 7762 2333 7944 2377
rect 7185 2197 8647 2333
rect 8835 2214 8921 2371
rect 8925 2197 9659 2359
rect 10456 2333 10638 2377
rect 10945 2333 11215 2379
rect 9753 2197 11215 2333
rect 11411 2214 11497 2371
rect 11501 2197 11867 2359
rect 11877 2333 12147 2379
rect 12454 2333 12636 2377
rect 11877 2197 13339 2333
rect 13341 2197 13891 2359
rect 13987 2214 14073 2371
rect 14537 2197 15639 2359
rect 15641 2197 16375 2359
rect 16563 2214 16649 2371
rect 16837 2197 17111 2353
rect 17113 2197 17479 2359
rect 17578 2333 17847 2379
rect 17481 2197 17847 2333
rect 17849 2197 18583 2359
rect 18585 2197 18859 2359
rect 3527 2166 3559 2188
rect 3803 2166 3835 2188
rect 4077 2159 4111 2189
rect 4169 2159 4203 2197
rect 4536 2165 4560 2187
rect 4629 2159 4663 2197
rect 6103 2166 6135 2188
rect 6377 2159 6411 2197
rect 7112 2165 7136 2187
rect 8585 2159 8619 2197
rect 8679 2166 8711 2188
rect 8953 2159 8987 2197
rect 9688 2165 9712 2187
rect 9781 2159 9815 2197
rect 11255 2166 11287 2188
rect 11529 2159 11563 2197
rect 13277 2159 13311 2197
rect 13369 2159 13403 2197
rect 13920 2165 13944 2187
rect 14107 2166 14139 2188
rect 14473 2159 14507 2193
rect 14565 2159 14599 2197
rect 15669 2159 15703 2197
rect 16407 2166 16439 2188
rect 16683 2166 16715 2188
rect 17049 2159 17083 2197
rect 17141 2159 17175 2197
rect 17509 2159 17543 2197
rect 17877 2159 17911 2197
rect 18797 2159 18831 2197
<< scnmos >>
rect 1183 7459 1301 7569
rect 1644 7439 1674 7569
rect 1728 7439 1758 7569
rect 1823 7485 1853 7569
rect 2011 7459 2957 7569
rect 3115 7459 3509 7569
rect 4036 7439 4066 7569
rect 4120 7439 4150 7569
rect 4215 7485 4245 7569
rect 4403 7459 5349 7569
rect 5692 7439 5722 7569
rect 5776 7439 5806 7569
rect 5871 7485 5901 7569
rect 6059 7459 6177 7569
rect 6427 7459 7373 7569
rect 7531 7459 7741 7569
rect 7899 7485 7929 7569
rect 7994 7439 8024 7569
rect 8078 7439 8108 7569
rect 8267 7459 8661 7569
rect 9003 7459 9397 7569
rect 9739 7459 9949 7569
rect 10108 7485 10138 7569
rect 10203 7485 10233 7569
rect 10287 7485 10317 7569
rect 10475 7459 11053 7569
rect 11211 7459 11329 7569
rect 11579 7459 12157 7569
rect 12315 7485 12345 7569
rect 12410 7439 12440 7569
rect 12494 7439 12524 7569
rect 12683 7459 13629 7569
rect 13787 7459 13905 7569
rect 14155 7459 14365 7569
rect 14523 7485 14553 7569
rect 14618 7439 14648 7569
rect 14702 7439 14732 7569
rect 14891 7459 15837 7569
rect 15995 7459 16389 7569
rect 16915 7485 16945 7569
rect 17010 7439 17040 7569
rect 17094 7439 17124 7569
rect 17283 7459 17861 7569
rect 18111 7485 18141 7569
rect 18206 7439 18236 7569
rect 18290 7439 18320 7569
rect 18663 7459 18781 7569
rect 1183 6575 1301 6685
rect 1459 6575 2405 6685
rect 2563 6575 3509 6685
rect 3851 6575 4797 6685
rect 4955 6575 5901 6685
rect 6059 6575 7005 6685
rect 7163 6575 8109 6685
rect 8267 6575 8661 6685
rect 9003 6575 9949 6685
rect 10107 6575 11053 6685
rect 11211 6575 12157 6685
rect 12315 6575 13261 6685
rect 13419 6575 13813 6685
rect 14155 6575 15101 6685
rect 15259 6575 16205 6685
rect 16363 6575 17309 6685
rect 17467 6575 18413 6685
rect 18663 6575 18781 6685
rect 1183 6371 1301 6481
rect 1459 6371 2405 6481
rect 2563 6371 3509 6481
rect 3667 6371 4613 6481
rect 4771 6371 5717 6481
rect 5875 6371 6085 6481
rect 6427 6371 7373 6481
rect 7531 6371 8477 6481
rect 8635 6371 9581 6481
rect 9739 6371 10685 6481
rect 10843 6371 11237 6481
rect 11579 6371 12525 6481
rect 12683 6371 13629 6481
rect 13787 6371 14733 6481
rect 14891 6371 15837 6481
rect 15995 6371 16389 6481
rect 16731 6371 17677 6481
rect 17835 6371 18413 6481
rect 18663 6371 18781 6481
rect 1183 5487 1301 5597
rect 1459 5487 2037 5597
rect 2287 5487 2317 5591
rect 2375 5487 2405 5591
rect 2563 5487 2957 5597
rect 3115 5487 3145 5591
rect 3203 5487 3233 5591
rect 3391 5487 3601 5597
rect 3851 5487 4797 5597
rect 4955 5487 5901 5597
rect 6059 5487 6637 5597
rect 6795 5487 6825 5617
rect 6904 5487 6934 5571
rect 7000 5487 7030 5571
rect 7125 5487 7155 5571
rect 7221 5487 7251 5571
rect 7389 5487 7419 5571
rect 7623 5487 8569 5597
rect 9003 5487 9581 5597
rect 9923 5487 9953 5617
rect 10032 5487 10062 5571
rect 10128 5487 10158 5571
rect 10253 5487 10283 5571
rect 10349 5487 10379 5571
rect 10517 5487 10547 5571
rect 10751 5487 10961 5597
rect 11163 5487 11193 5617
rect 11271 5515 11301 5599
rect 11355 5515 11385 5599
rect 11579 5487 12157 5597
rect 12315 5487 12345 5617
rect 12424 5487 12454 5571
rect 12520 5487 12550 5571
rect 12645 5487 12675 5571
rect 12741 5487 12771 5571
rect 12909 5487 12939 5571
rect 13143 5487 13721 5597
rect 14339 5487 14369 5617
rect 14448 5487 14478 5571
rect 14544 5487 14574 5571
rect 14669 5487 14699 5571
rect 14765 5487 14795 5571
rect 14933 5487 14963 5571
rect 15167 5487 16113 5597
rect 16271 5487 17217 5597
rect 17375 5487 18321 5597
rect 18663 5487 18781 5597
rect 1183 5283 1301 5393
rect 1459 5283 1853 5393
rect 2055 5263 2085 5393
rect 2163 5281 2193 5365
rect 2247 5281 2277 5365
rect 2471 5283 2681 5393
rect 2975 5263 3005 5393
rect 3083 5281 3113 5365
rect 3167 5281 3197 5365
rect 3391 5283 3601 5393
rect 3759 5309 3789 5393
rect 3854 5263 3884 5393
rect 3938 5263 3968 5393
rect 4127 5283 4337 5393
rect 4497 5263 4527 5393
rect 4581 5263 4611 5393
rect 4771 5283 5717 5393
rect 5875 5289 5905 5393
rect 5963 5289 5993 5393
rect 6427 5283 6545 5393
rect 6703 5263 6733 5393
rect 6812 5309 6842 5393
rect 6908 5309 6938 5393
rect 7033 5309 7063 5393
rect 7129 5309 7159 5393
rect 7297 5309 7327 5393
rect 7531 5283 7741 5393
rect 7899 5263 7929 5393
rect 8008 5309 8038 5393
rect 8104 5309 8134 5393
rect 8229 5309 8259 5393
rect 8325 5309 8355 5393
rect 8493 5309 8523 5393
rect 8727 5283 8937 5393
rect 9187 5263 9217 5393
rect 9375 5263 9405 5393
rect 9467 5263 9497 5393
rect 9551 5263 9581 5393
rect 9739 5283 10317 5393
rect 10475 5263 10505 5393
rect 10584 5309 10614 5393
rect 10680 5309 10710 5393
rect 10805 5309 10835 5393
rect 10901 5309 10931 5393
rect 11069 5309 11099 5393
rect 11579 5283 12525 5393
rect 12683 5283 12893 5393
rect 13143 5263 13173 5393
rect 13252 5309 13282 5393
rect 13348 5309 13378 5393
rect 13473 5309 13503 5393
rect 13569 5309 13599 5393
rect 13737 5309 13767 5393
rect 13971 5283 14917 5393
rect 15075 5283 16021 5393
rect 16179 5283 16389 5393
rect 16731 5283 17677 5393
rect 17835 5283 18413 5393
rect 18663 5283 18781 5393
rect 1183 4399 1301 4509
rect 1459 4399 1853 4509
rect 2103 4399 2133 4483
rect 2187 4399 2217 4483
rect 2375 4399 2405 4483
rect 2487 4399 2517 4471
rect 2586 4399 2616 4471
rect 2685 4399 2715 4483
rect 2804 4399 2834 4527
rect 2905 4399 2935 4471
rect 3011 4399 3041 4471
rect 3106 4399 3136 4483
rect 3295 4399 3325 4529
rect 3379 4399 3409 4529
rect 4079 4399 4109 4529
rect 4187 4427 4217 4511
rect 4271 4427 4301 4511
rect 4495 4399 4705 4509
rect 4955 4399 4985 4529
rect 5143 4399 5173 4529
rect 5235 4399 5265 4529
rect 5319 4399 5349 4529
rect 5507 4399 5717 4509
rect 5875 4399 5905 4529
rect 6063 4399 6093 4529
rect 6155 4399 6185 4529
rect 6239 4399 6269 4529
rect 6427 4399 6637 4509
rect 6795 4399 6825 4483
rect 6879 4399 6909 4483
rect 7067 4399 7097 4483
rect 7179 4399 7209 4471
rect 7278 4399 7308 4471
rect 7377 4399 7407 4483
rect 7496 4399 7526 4527
rect 7597 4399 7627 4471
rect 7703 4399 7733 4471
rect 7798 4399 7828 4483
rect 7987 4399 8017 4529
rect 8071 4399 8101 4529
rect 8267 4399 8661 4509
rect 9003 4399 9581 4509
rect 9739 4399 9857 4509
rect 10023 4399 10053 4529
rect 10107 4399 10137 4529
rect 10296 4399 10326 4483
rect 10391 4399 10421 4471
rect 10497 4399 10527 4471
rect 10598 4399 10628 4527
rect 10717 4399 10747 4483
rect 10816 4399 10846 4471
rect 10915 4399 10945 4471
rect 11027 4399 11057 4483
rect 11215 4399 11245 4483
rect 11299 4399 11329 4483
rect 11487 4399 11697 4509
rect 11855 4399 11885 4529
rect 12043 4399 12073 4529
rect 12135 4399 12165 4529
rect 12219 4399 12249 4529
rect 12407 4399 12617 4509
rect 12775 4399 12805 4529
rect 12963 4399 12993 4529
rect 13055 4399 13085 4529
rect 13139 4399 13169 4529
rect 13327 4399 13905 4509
rect 14155 4399 14273 4509
rect 14467 4427 14497 4511
rect 14551 4427 14581 4511
rect 14659 4399 14689 4529
rect 14891 4399 15837 4509
rect 15995 4399 16941 4509
rect 17099 4399 18045 4509
rect 18203 4399 18413 4509
rect 18663 4399 18781 4509
rect 1183 4195 1301 4305
rect 1459 4195 1853 4305
rect 2011 4201 2041 4305
rect 2099 4201 2129 4305
rect 2287 4195 2497 4305
rect 2663 4175 2693 4305
rect 2747 4175 2777 4305
rect 2936 4221 2966 4305
rect 3031 4233 3061 4305
rect 3137 4233 3167 4305
rect 3238 4177 3268 4305
rect 3357 4221 3387 4305
rect 3456 4233 3486 4305
rect 3555 4233 3585 4305
rect 3667 4221 3697 4305
rect 3855 4221 3885 4305
rect 3939 4221 3969 4305
rect 4127 4195 4521 4305
rect 4687 4175 4717 4305
rect 4771 4175 4801 4305
rect 4960 4221 4990 4305
rect 5055 4233 5085 4305
rect 5161 4233 5191 4305
rect 5262 4177 5292 4305
rect 5381 4221 5411 4305
rect 5480 4233 5510 4305
rect 5579 4233 5609 4305
rect 5691 4221 5721 4305
rect 5879 4221 5909 4305
rect 5963 4221 5993 4305
rect 6427 4195 6821 4305
rect 6979 4175 7009 4305
rect 7167 4175 7197 4305
rect 7259 4175 7289 4305
rect 7343 4175 7373 4305
rect 7531 4195 7741 4305
rect 7900 4221 7930 4305
rect 7986 4221 8016 4305
rect 8072 4221 8102 4305
rect 8158 4221 8188 4305
rect 8244 4221 8274 4305
rect 8330 4221 8360 4305
rect 8416 4221 8446 4305
rect 8502 4221 8532 4305
rect 8588 4221 8618 4305
rect 8674 4221 8704 4305
rect 8760 4221 8790 4305
rect 8846 4221 8876 4305
rect 8931 4221 8961 4305
rect 9017 4221 9047 4305
rect 9103 4221 9133 4305
rect 9189 4221 9219 4305
rect 9275 4221 9305 4305
rect 9361 4221 9391 4305
rect 9447 4221 9477 4305
rect 9533 4221 9563 4305
rect 9739 4195 10317 4305
rect 10567 4175 10597 4305
rect 10755 4175 10785 4305
rect 10847 4175 10877 4305
rect 10931 4175 10961 4305
rect 11119 4195 11329 4305
rect 11763 4221 11793 4305
rect 11847 4221 11877 4305
rect 12035 4221 12065 4305
rect 12147 4233 12177 4305
rect 12246 4233 12276 4305
rect 12345 4221 12375 4305
rect 12464 4177 12494 4305
rect 12565 4233 12595 4305
rect 12671 4233 12701 4305
rect 12766 4221 12796 4305
rect 12955 4175 12985 4305
rect 13039 4175 13069 4305
rect 13235 4195 14181 4305
rect 14339 4195 15285 4305
rect 15535 4201 15565 4305
rect 15623 4201 15653 4305
rect 15811 4195 16389 4305
rect 16951 4193 16981 4277
rect 17035 4193 17065 4277
rect 17143 4175 17173 4305
rect 17375 4195 18321 4305
rect 18663 4195 18781 4305
rect 1183 3311 1301 3421
rect 1459 3311 1853 3421
rect 2103 3311 2133 3395
rect 2187 3311 2217 3395
rect 2375 3311 2405 3395
rect 2487 3311 2517 3383
rect 2586 3311 2616 3383
rect 2685 3311 2715 3395
rect 2804 3311 2834 3439
rect 2905 3311 2935 3383
rect 3011 3311 3041 3383
rect 3106 3311 3136 3395
rect 3295 3311 3325 3441
rect 3379 3311 3409 3441
rect 4035 3311 4065 3395
rect 4119 3311 4149 3395
rect 4307 3311 4337 3395
rect 4419 3311 4449 3383
rect 4518 3311 4548 3383
rect 4617 3311 4647 3395
rect 4736 3311 4766 3439
rect 4837 3311 4867 3383
rect 4943 3311 4973 3383
rect 5038 3311 5068 3395
rect 5227 3311 5257 3441
rect 5311 3311 5341 3441
rect 5507 3311 6085 3421
rect 6335 3311 6365 3441
rect 6523 3311 6553 3441
rect 6615 3311 6645 3441
rect 6699 3311 6729 3441
rect 6887 3311 7097 3421
rect 7255 3311 7285 3395
rect 7339 3311 7369 3395
rect 7527 3311 7557 3395
rect 7639 3311 7669 3383
rect 7738 3311 7768 3383
rect 7837 3311 7867 3395
rect 7956 3311 7986 3439
rect 8057 3311 8087 3383
rect 8163 3311 8193 3383
rect 8258 3311 8288 3395
rect 8447 3311 8477 3441
rect 8531 3311 8561 3441
rect 9003 3311 9581 3421
rect 9831 3311 9861 3395
rect 9915 3311 9945 3395
rect 10103 3311 10133 3395
rect 10215 3311 10245 3383
rect 10314 3311 10344 3383
rect 10413 3311 10443 3395
rect 10532 3311 10562 3439
rect 10633 3311 10663 3383
rect 10739 3311 10769 3383
rect 10834 3311 10864 3395
rect 11023 3311 11053 3441
rect 11107 3311 11137 3441
rect 11303 3311 11697 3421
rect 11855 3311 11885 3395
rect 11939 3311 11969 3395
rect 12127 3311 12157 3395
rect 12239 3311 12269 3383
rect 12338 3311 12368 3383
rect 12437 3311 12467 3395
rect 12556 3311 12586 3439
rect 12657 3311 12687 3383
rect 12763 3311 12793 3383
rect 12858 3311 12888 3395
rect 13047 3311 13077 3441
rect 13131 3311 13161 3441
rect 13327 3311 13905 3421
rect 14155 3311 15101 3421
rect 15259 3311 15653 3421
rect 15811 3311 15841 3415
rect 15899 3311 15929 3415
rect 16087 3311 16297 3421
rect 16499 3311 16529 3441
rect 16607 3339 16637 3423
rect 16691 3339 16721 3423
rect 16915 3311 17125 3421
rect 17327 3311 17357 3441
rect 17435 3339 17465 3423
rect 17519 3339 17549 3423
rect 17743 3311 18321 3421
rect 18663 3311 18781 3421
rect 1183 3107 1301 3217
rect 1459 3107 1669 3217
rect 1920 3133 1950 3217
rect 2015 3133 2045 3217
rect 2099 3133 2129 3217
rect 2287 3107 2497 3217
rect 2673 3133 2703 3217
rect 2759 3133 2789 3217
rect 2845 3133 2875 3217
rect 2931 3133 2961 3217
rect 3017 3133 3047 3217
rect 3103 3133 3133 3217
rect 3189 3133 3219 3217
rect 3275 3133 3305 3217
rect 3360 3133 3390 3217
rect 3446 3133 3476 3217
rect 3532 3133 3562 3217
rect 3618 3133 3648 3217
rect 3704 3133 3734 3217
rect 3790 3133 3820 3217
rect 3876 3133 3906 3217
rect 3962 3133 3992 3217
rect 4048 3133 4078 3217
rect 4134 3133 4164 3217
rect 4220 3133 4250 3217
rect 4306 3133 4336 3217
rect 4495 3107 5441 3217
rect 5599 3107 6177 3217
rect 6427 3107 7005 3217
rect 7439 3107 7649 3217
rect 7808 3133 7838 3217
rect 7894 3133 7924 3217
rect 7980 3133 8010 3217
rect 8066 3133 8096 3217
rect 8152 3133 8182 3217
rect 8238 3133 8268 3217
rect 8324 3133 8354 3217
rect 8410 3133 8440 3217
rect 8496 3133 8526 3217
rect 8582 3133 8612 3217
rect 8668 3133 8698 3217
rect 8754 3133 8784 3217
rect 8839 3133 8869 3217
rect 8925 3133 8955 3217
rect 9011 3133 9041 3217
rect 9097 3133 9127 3217
rect 9183 3133 9213 3217
rect 9269 3133 9299 3217
rect 9355 3133 9385 3217
rect 9441 3133 9471 3217
rect 9647 3107 10593 3217
rect 10751 3107 11329 3217
rect 11763 3133 11793 3217
rect 11847 3133 11877 3217
rect 12035 3133 12065 3217
rect 12147 3145 12177 3217
rect 12246 3145 12276 3217
rect 12345 3133 12375 3217
rect 12464 3089 12494 3217
rect 12565 3145 12595 3217
rect 12671 3145 12701 3217
rect 12766 3133 12796 3217
rect 12955 3087 12985 3217
rect 13039 3087 13069 3217
rect 13235 3107 14181 3217
rect 14339 3107 15285 3217
rect 15443 3107 16389 3217
rect 16915 3113 16945 3217
rect 17003 3113 17033 3217
rect 17191 3107 18137 3217
rect 18295 3107 18505 3217
rect 18663 3107 18781 3217
rect 1183 2223 1301 2333
rect 1459 2223 1853 2333
rect 2111 2223 2141 2353
rect 2195 2223 2225 2353
rect 2384 2223 2414 2307
rect 2479 2223 2509 2295
rect 2585 2223 2615 2295
rect 2686 2223 2716 2351
rect 2805 2223 2835 2307
rect 2904 2223 2934 2295
rect 3003 2223 3033 2295
rect 3115 2223 3145 2307
rect 3303 2223 3333 2307
rect 3387 2223 3417 2307
rect 4219 2223 4429 2333
rect 4679 2223 4709 2307
rect 4763 2223 4793 2307
rect 4951 2223 4981 2307
rect 5063 2223 5093 2295
rect 5162 2223 5192 2295
rect 5261 2223 5291 2307
rect 5380 2223 5410 2351
rect 5481 2223 5511 2295
rect 5587 2223 5617 2295
rect 5682 2223 5712 2307
rect 5871 2223 5901 2353
rect 5955 2223 5985 2353
rect 6427 2223 7005 2333
rect 7263 2223 7293 2353
rect 7347 2223 7377 2353
rect 7536 2223 7566 2307
rect 7631 2223 7661 2295
rect 7737 2223 7767 2295
rect 7838 2223 7868 2351
rect 7957 2223 7987 2307
rect 8056 2223 8086 2295
rect 8155 2223 8185 2295
rect 8267 2223 8297 2307
rect 8455 2223 8485 2307
rect 8539 2223 8569 2307
rect 9003 2223 9581 2333
rect 9831 2223 9861 2307
rect 9915 2223 9945 2307
rect 10103 2223 10133 2307
rect 10215 2223 10245 2295
rect 10314 2223 10344 2295
rect 10413 2223 10443 2307
rect 10532 2223 10562 2351
rect 10633 2223 10663 2295
rect 10739 2223 10769 2295
rect 10834 2223 10864 2307
rect 11023 2223 11053 2353
rect 11107 2223 11137 2353
rect 11579 2223 11789 2333
rect 11955 2223 11985 2353
rect 12039 2223 12069 2353
rect 12228 2223 12258 2307
rect 12323 2223 12353 2295
rect 12429 2223 12459 2295
rect 12530 2223 12560 2351
rect 12649 2223 12679 2307
rect 12748 2223 12778 2295
rect 12847 2223 12877 2295
rect 12959 2223 12989 2307
rect 13147 2223 13177 2307
rect 13231 2223 13261 2307
rect 13419 2223 13813 2333
rect 14615 2223 15561 2333
rect 15719 2223 16297 2333
rect 16915 2223 16945 2327
rect 17003 2223 17033 2327
rect 17191 2223 17401 2333
rect 17559 2223 17589 2307
rect 17654 2223 17684 2353
rect 17738 2223 17768 2353
rect 17927 2223 18505 2333
rect 18663 2223 18781 2333
<< scpmoshvt >>
rect 1183 7119 1301 7293
rect 1644 7119 1674 7319
rect 1728 7119 1758 7319
rect 1823 7127 1853 7255
rect 2011 7119 2957 7293
rect 3115 7119 3509 7293
rect 4036 7119 4066 7319
rect 4120 7119 4150 7319
rect 4215 7127 4245 7255
rect 4403 7119 5349 7293
rect 5692 7119 5722 7319
rect 5776 7119 5806 7319
rect 5871 7127 5901 7255
rect 6059 7119 6177 7293
rect 6427 7119 7373 7293
rect 7531 7119 7741 7293
rect 7899 7127 7929 7255
rect 7994 7119 8024 7319
rect 8078 7119 8108 7319
rect 8267 7119 8661 7293
rect 9003 7119 9397 7293
rect 9739 7119 9949 7293
rect 10108 7119 10138 7319
rect 10203 7119 10233 7319
rect 10287 7119 10317 7319
rect 10475 7119 11053 7293
rect 11211 7119 11329 7293
rect 11579 7119 12157 7293
rect 12315 7127 12345 7255
rect 12410 7119 12440 7319
rect 12494 7119 12524 7319
rect 12683 7119 13629 7293
rect 13787 7119 13905 7293
rect 14155 7119 14365 7293
rect 14523 7127 14553 7255
rect 14618 7119 14648 7319
rect 14702 7119 14732 7319
rect 14891 7119 15837 7293
rect 15995 7119 16389 7293
rect 16915 7127 16945 7255
rect 17010 7119 17040 7319
rect 17094 7119 17124 7319
rect 17283 7119 17861 7293
rect 18111 7127 18141 7255
rect 18206 7119 18236 7319
rect 18290 7119 18320 7319
rect 18663 7119 18781 7293
rect 1183 6851 1301 7025
rect 1459 6851 2405 7025
rect 2563 6851 3509 7025
rect 3851 6851 4797 7025
rect 4955 6851 5901 7025
rect 6059 6851 7005 7025
rect 7163 6851 8109 7025
rect 8267 6851 8661 7025
rect 9003 6851 9949 7025
rect 10107 6851 11053 7025
rect 11211 6851 12157 7025
rect 12315 6851 13261 7025
rect 13419 6851 13813 7025
rect 14155 6851 15101 7025
rect 15259 6851 16205 7025
rect 16363 6851 17309 7025
rect 17467 6851 18413 7025
rect 18663 6851 18781 7025
rect 1183 6031 1301 6205
rect 1459 6031 2405 6205
rect 2563 6031 3509 6205
rect 3667 6031 4613 6205
rect 4771 6031 5717 6205
rect 5875 6031 6085 6205
rect 6427 6031 7373 6205
rect 7531 6031 8477 6205
rect 8635 6031 9581 6205
rect 9739 6031 10685 6205
rect 10843 6031 11237 6205
rect 11579 6031 12525 6205
rect 12683 6031 13629 6205
rect 13787 6031 14733 6205
rect 14891 6031 15837 6205
rect 15995 6031 16389 6205
rect 16731 6031 17677 6205
rect 17835 6031 18413 6205
rect 18663 6031 18781 6205
rect 1183 5763 1301 5937
rect 1459 5763 2037 5937
rect 2287 5779 2317 5937
rect 2375 5779 2405 5937
rect 2563 5763 2957 5937
rect 3115 5779 3145 5937
rect 3203 5779 3233 5937
rect 3391 5763 3601 5937
rect 3851 5763 4797 5937
rect 4955 5763 5901 5937
rect 6059 5763 6637 5937
rect 6795 5737 6825 5937
rect 6904 5814 6934 5898
rect 7007 5814 7037 5898
rect 7221 5814 7251 5898
rect 7293 5814 7323 5898
rect 7389 5814 7419 5898
rect 7623 5763 8569 5937
rect 9003 5763 9581 5937
rect 9923 5737 9953 5937
rect 10032 5814 10062 5898
rect 10135 5814 10165 5898
rect 10349 5814 10379 5898
rect 10421 5814 10451 5898
rect 10517 5814 10547 5898
rect 10751 5763 10961 5937
rect 11163 5737 11193 5937
rect 11271 5811 11301 5895
rect 11355 5811 11385 5895
rect 11579 5763 12157 5937
rect 12315 5737 12345 5937
rect 12424 5814 12454 5898
rect 12527 5814 12557 5898
rect 12741 5814 12771 5898
rect 12813 5814 12843 5898
rect 12909 5814 12939 5898
rect 13143 5763 13721 5937
rect 14339 5737 14369 5937
rect 14448 5814 14478 5898
rect 14551 5814 14581 5898
rect 14765 5814 14795 5898
rect 14837 5814 14867 5898
rect 14933 5814 14963 5898
rect 15167 5763 16113 5937
rect 16271 5763 17217 5937
rect 17375 5763 18321 5937
rect 18663 5763 18781 5937
rect 1183 4943 1301 5117
rect 1459 4943 1853 5117
rect 2055 4943 2085 5143
rect 2163 4985 2193 5069
rect 2247 4985 2277 5069
rect 2471 4943 2681 5117
rect 2975 4943 3005 5143
rect 3083 4985 3113 5069
rect 3167 4985 3197 5069
rect 3391 4943 3601 5117
rect 3759 4951 3789 5079
rect 3854 4943 3884 5143
rect 3938 4943 3968 5143
rect 4127 4943 4337 5117
rect 4497 4943 4527 5143
rect 4581 4943 4611 5143
rect 4771 4943 5717 5117
rect 5875 4943 5905 5101
rect 5963 4943 5993 5101
rect 6427 4943 6545 5117
rect 6703 4943 6733 5143
rect 6812 4982 6842 5066
rect 6915 4982 6945 5066
rect 7129 4982 7159 5066
rect 7201 4982 7231 5066
rect 7297 4982 7327 5066
rect 7531 4943 7741 5117
rect 7899 4943 7929 5143
rect 8008 4982 8038 5066
rect 8111 4982 8141 5066
rect 8325 4982 8355 5066
rect 8397 4982 8427 5066
rect 8493 4982 8523 5066
rect 8727 4943 8937 5117
rect 9191 4943 9221 5143
rect 9352 4943 9382 5143
rect 9460 4943 9490 5143
rect 9551 4943 9581 5143
rect 9739 4943 10317 5117
rect 10475 4943 10505 5143
rect 10584 4982 10614 5066
rect 10687 4982 10717 5066
rect 10901 4982 10931 5066
rect 10973 4982 11003 5066
rect 11069 4982 11099 5066
rect 11579 4943 12525 5117
rect 12683 4943 12893 5117
rect 13143 4943 13173 5143
rect 13252 4982 13282 5066
rect 13355 4982 13385 5066
rect 13569 4982 13599 5066
rect 13641 4982 13671 5066
rect 13737 4982 13767 5066
rect 13971 4943 14917 5117
rect 15075 4943 16021 5117
rect 16179 4943 16389 5117
rect 16731 4943 17677 5117
rect 17835 4943 18413 5117
rect 18663 4943 18781 5117
rect 1183 4675 1301 4849
rect 1459 4675 1853 4849
rect 2103 4715 2133 4843
rect 2187 4715 2217 4843
rect 2375 4765 2405 4849
rect 2460 4765 2490 4849
rect 2555 4765 2585 4849
rect 2658 4765 2688 4849
rect 2790 4699 2820 4849
rect 2885 4765 2915 4849
rect 2969 4765 2999 4849
rect 3083 4765 3113 4849
rect 3293 4649 3323 4849
rect 3377 4649 3407 4849
rect 4079 4649 4109 4849
rect 4187 4723 4217 4807
rect 4271 4723 4301 4807
rect 4495 4675 4705 4849
rect 4959 4649 4989 4849
rect 5120 4649 5150 4849
rect 5228 4649 5258 4849
rect 5319 4649 5349 4849
rect 5507 4675 5717 4849
rect 5879 4649 5909 4849
rect 6040 4649 6070 4849
rect 6148 4649 6178 4849
rect 6239 4649 6269 4849
rect 6427 4675 6637 4849
rect 6795 4715 6825 4843
rect 6879 4715 6909 4843
rect 7067 4765 7097 4849
rect 7152 4765 7182 4849
rect 7247 4765 7277 4849
rect 7350 4765 7380 4849
rect 7482 4699 7512 4849
rect 7577 4765 7607 4849
rect 7661 4765 7691 4849
rect 7775 4765 7805 4849
rect 7985 4649 8015 4849
rect 8069 4649 8099 4849
rect 8267 4675 8661 4849
rect 9003 4675 9581 4849
rect 9739 4675 9857 4849
rect 10025 4649 10055 4849
rect 10109 4649 10139 4849
rect 10319 4765 10349 4849
rect 10433 4765 10463 4849
rect 10517 4765 10547 4849
rect 10612 4699 10642 4849
rect 10744 4765 10774 4849
rect 10847 4765 10877 4849
rect 10942 4765 10972 4849
rect 11027 4765 11057 4849
rect 11215 4715 11245 4843
rect 11299 4715 11329 4843
rect 11487 4675 11697 4849
rect 11859 4649 11889 4849
rect 12020 4649 12050 4849
rect 12128 4649 12158 4849
rect 12219 4649 12249 4849
rect 12407 4675 12617 4849
rect 12779 4649 12809 4849
rect 12940 4649 12970 4849
rect 13048 4649 13078 4849
rect 13139 4649 13169 4849
rect 13327 4675 13905 4849
rect 14155 4675 14273 4849
rect 14467 4723 14497 4807
rect 14551 4723 14581 4807
rect 14659 4649 14689 4849
rect 14891 4675 15837 4849
rect 15995 4675 16941 4849
rect 17099 4675 18045 4849
rect 18203 4675 18413 4849
rect 18663 4675 18781 4849
rect 1183 3855 1301 4029
rect 1459 3855 1853 4029
rect 2011 3855 2041 4013
rect 2099 3855 2129 4013
rect 2287 3855 2497 4029
rect 2665 3855 2695 4055
rect 2749 3855 2779 4055
rect 2959 3855 2989 3939
rect 3073 3855 3103 3939
rect 3157 3855 3187 3939
rect 3252 3855 3282 4005
rect 3384 3855 3414 3939
rect 3487 3855 3517 3939
rect 3582 3855 3612 3939
rect 3667 3855 3697 3939
rect 3855 3861 3885 3989
rect 3939 3861 3969 3989
rect 4127 3855 4521 4029
rect 4689 3855 4719 4055
rect 4773 3855 4803 4055
rect 4983 3855 5013 3939
rect 5097 3855 5127 3939
rect 5181 3855 5211 3939
rect 5276 3855 5306 4005
rect 5408 3855 5438 3939
rect 5511 3855 5541 3939
rect 5606 3855 5636 3939
rect 5691 3855 5721 3939
rect 5879 3861 5909 3989
rect 5963 3861 5993 3989
rect 6427 3855 6821 4029
rect 6983 3855 7013 4055
rect 7144 3855 7174 4055
rect 7252 3855 7282 4055
rect 7343 3855 7373 4055
rect 7531 3855 7741 4029
rect 7900 3855 7930 4055
rect 7986 3855 8016 4055
rect 8072 3855 8102 4055
rect 8158 3855 8188 4055
rect 8244 3855 8274 4055
rect 8330 3855 8360 4055
rect 8416 3855 8446 4055
rect 8502 3855 8532 4055
rect 8588 3855 8618 4055
rect 8674 3855 8704 4055
rect 8760 3855 8790 4055
rect 8846 3855 8876 4055
rect 8931 3855 8961 4055
rect 9017 3855 9047 4055
rect 9103 3855 9133 4055
rect 9189 3855 9219 4055
rect 9275 3855 9305 4055
rect 9361 3855 9391 4055
rect 9447 3855 9477 4055
rect 9533 3855 9563 4055
rect 9739 3855 10317 4029
rect 10571 3855 10601 4055
rect 10732 3855 10762 4055
rect 10840 3855 10870 4055
rect 10931 3855 10961 4055
rect 11119 3855 11329 4029
rect 11763 3861 11793 3989
rect 11847 3861 11877 3989
rect 12035 3855 12065 3939
rect 12120 3855 12150 3939
rect 12215 3855 12245 3939
rect 12318 3855 12348 3939
rect 12450 3855 12480 4005
rect 12545 3855 12575 3939
rect 12629 3855 12659 3939
rect 12743 3855 12773 3939
rect 12953 3855 12983 4055
rect 13037 3855 13067 4055
rect 13235 3855 14181 4029
rect 14339 3855 15285 4029
rect 15535 3855 15565 4013
rect 15623 3855 15653 4013
rect 15811 3855 16389 4029
rect 16951 3897 16981 3981
rect 17035 3897 17065 3981
rect 17143 3855 17173 4055
rect 17375 3855 18321 4029
rect 18663 3855 18781 4029
rect 1183 3587 1301 3761
rect 1459 3587 1853 3761
rect 2103 3627 2133 3755
rect 2187 3627 2217 3755
rect 2375 3677 2405 3761
rect 2460 3677 2490 3761
rect 2555 3677 2585 3761
rect 2658 3677 2688 3761
rect 2790 3611 2820 3761
rect 2885 3677 2915 3761
rect 2969 3677 2999 3761
rect 3083 3677 3113 3761
rect 3293 3561 3323 3761
rect 3377 3561 3407 3761
rect 4035 3627 4065 3755
rect 4119 3627 4149 3755
rect 4307 3677 4337 3761
rect 4392 3677 4422 3761
rect 4487 3677 4517 3761
rect 4590 3677 4620 3761
rect 4722 3611 4752 3761
rect 4817 3677 4847 3761
rect 4901 3677 4931 3761
rect 5015 3677 5045 3761
rect 5225 3561 5255 3761
rect 5309 3561 5339 3761
rect 5507 3587 6085 3761
rect 6339 3561 6369 3761
rect 6500 3561 6530 3761
rect 6608 3561 6638 3761
rect 6699 3561 6729 3761
rect 6887 3587 7097 3761
rect 7255 3627 7285 3755
rect 7339 3627 7369 3755
rect 7527 3677 7557 3761
rect 7612 3677 7642 3761
rect 7707 3677 7737 3761
rect 7810 3677 7840 3761
rect 7942 3611 7972 3761
rect 8037 3677 8067 3761
rect 8121 3677 8151 3761
rect 8235 3677 8265 3761
rect 8445 3561 8475 3761
rect 8529 3561 8559 3761
rect 9003 3587 9581 3761
rect 9831 3627 9861 3755
rect 9915 3627 9945 3755
rect 10103 3677 10133 3761
rect 10188 3677 10218 3761
rect 10283 3677 10313 3761
rect 10386 3677 10416 3761
rect 10518 3611 10548 3761
rect 10613 3677 10643 3761
rect 10697 3677 10727 3761
rect 10811 3677 10841 3761
rect 11021 3561 11051 3761
rect 11105 3561 11135 3761
rect 11303 3587 11697 3761
rect 11855 3627 11885 3755
rect 11939 3627 11969 3755
rect 12127 3677 12157 3761
rect 12212 3677 12242 3761
rect 12307 3677 12337 3761
rect 12410 3677 12440 3761
rect 12542 3611 12572 3761
rect 12637 3677 12667 3761
rect 12721 3677 12751 3761
rect 12835 3677 12865 3761
rect 13045 3561 13075 3761
rect 13129 3561 13159 3761
rect 13327 3587 13905 3761
rect 14155 3587 15101 3761
rect 15259 3587 15653 3761
rect 15811 3603 15841 3761
rect 15899 3603 15929 3761
rect 16087 3587 16297 3761
rect 16499 3561 16529 3761
rect 16607 3635 16637 3719
rect 16691 3635 16721 3719
rect 16915 3587 17125 3761
rect 17327 3561 17357 3761
rect 17435 3635 17465 3719
rect 17519 3635 17549 3719
rect 17743 3587 18321 3761
rect 18663 3587 18781 3761
rect 1183 2767 1301 2941
rect 1459 2767 1669 2941
rect 1920 2767 1950 2967
rect 2015 2767 2045 2967
rect 2099 2767 2129 2967
rect 2287 2767 2497 2941
rect 2673 2767 2703 2967
rect 2759 2767 2789 2967
rect 2845 2767 2875 2967
rect 2931 2767 2961 2967
rect 3017 2767 3047 2967
rect 3103 2767 3133 2967
rect 3189 2767 3219 2967
rect 3275 2767 3305 2967
rect 3360 2767 3390 2967
rect 3446 2767 3476 2967
rect 3532 2767 3562 2967
rect 3618 2767 3648 2967
rect 3704 2767 3734 2967
rect 3790 2767 3820 2967
rect 3876 2767 3906 2967
rect 3962 2767 3992 2967
rect 4048 2767 4078 2967
rect 4134 2767 4164 2967
rect 4220 2767 4250 2967
rect 4306 2767 4336 2967
rect 4495 2767 5441 2941
rect 5599 2767 6177 2941
rect 6427 2767 7005 2941
rect 7439 2767 7649 2941
rect 7808 2767 7838 2967
rect 7894 2767 7924 2967
rect 7980 2767 8010 2967
rect 8066 2767 8096 2967
rect 8152 2767 8182 2967
rect 8238 2767 8268 2967
rect 8324 2767 8354 2967
rect 8410 2767 8440 2967
rect 8496 2767 8526 2967
rect 8582 2767 8612 2967
rect 8668 2767 8698 2967
rect 8754 2767 8784 2967
rect 8839 2767 8869 2967
rect 8925 2767 8955 2967
rect 9011 2767 9041 2967
rect 9097 2767 9127 2967
rect 9183 2767 9213 2967
rect 9269 2767 9299 2967
rect 9355 2767 9385 2967
rect 9441 2767 9471 2967
rect 9647 2767 10593 2941
rect 10751 2767 11329 2941
rect 11763 2773 11793 2901
rect 11847 2773 11877 2901
rect 12035 2767 12065 2851
rect 12120 2767 12150 2851
rect 12215 2767 12245 2851
rect 12318 2767 12348 2851
rect 12450 2767 12480 2917
rect 12545 2767 12575 2851
rect 12629 2767 12659 2851
rect 12743 2767 12773 2851
rect 12953 2767 12983 2967
rect 13037 2767 13067 2967
rect 13235 2767 14181 2941
rect 14339 2767 15285 2941
rect 15443 2767 16389 2941
rect 16915 2767 16945 2925
rect 17003 2767 17033 2925
rect 17191 2767 18137 2941
rect 18295 2767 18505 2941
rect 18663 2767 18781 2941
rect 1183 2499 1301 2673
rect 1459 2499 1853 2673
rect 2113 2473 2143 2673
rect 2197 2473 2227 2673
rect 2407 2589 2437 2673
rect 2521 2589 2551 2673
rect 2605 2589 2635 2673
rect 2700 2523 2730 2673
rect 2832 2589 2862 2673
rect 2935 2589 2965 2673
rect 3030 2589 3060 2673
rect 3115 2589 3145 2673
rect 3303 2539 3333 2667
rect 3387 2539 3417 2667
rect 4219 2499 4429 2673
rect 4679 2539 4709 2667
rect 4763 2539 4793 2667
rect 4951 2589 4981 2673
rect 5036 2589 5066 2673
rect 5131 2589 5161 2673
rect 5234 2589 5264 2673
rect 5366 2523 5396 2673
rect 5461 2589 5491 2673
rect 5545 2589 5575 2673
rect 5659 2589 5689 2673
rect 5869 2473 5899 2673
rect 5953 2473 5983 2673
rect 6427 2499 7005 2673
rect 7265 2473 7295 2673
rect 7349 2473 7379 2673
rect 7559 2589 7589 2673
rect 7673 2589 7703 2673
rect 7757 2589 7787 2673
rect 7852 2523 7882 2673
rect 7984 2589 8014 2673
rect 8087 2589 8117 2673
rect 8182 2589 8212 2673
rect 8267 2589 8297 2673
rect 8455 2539 8485 2667
rect 8539 2539 8569 2667
rect 9003 2499 9581 2673
rect 9831 2539 9861 2667
rect 9915 2539 9945 2667
rect 10103 2589 10133 2673
rect 10188 2589 10218 2673
rect 10283 2589 10313 2673
rect 10386 2589 10416 2673
rect 10518 2523 10548 2673
rect 10613 2589 10643 2673
rect 10697 2589 10727 2673
rect 10811 2589 10841 2673
rect 11021 2473 11051 2673
rect 11105 2473 11135 2673
rect 11579 2499 11789 2673
rect 11957 2473 11987 2673
rect 12041 2473 12071 2673
rect 12251 2589 12281 2673
rect 12365 2589 12395 2673
rect 12449 2589 12479 2673
rect 12544 2523 12574 2673
rect 12676 2589 12706 2673
rect 12779 2589 12809 2673
rect 12874 2589 12904 2673
rect 12959 2589 12989 2673
rect 13147 2539 13177 2667
rect 13231 2539 13261 2667
rect 13419 2499 13813 2673
rect 14615 2499 15561 2673
rect 15719 2499 16297 2673
rect 16915 2515 16945 2673
rect 17003 2515 17033 2673
rect 17191 2499 17401 2673
rect 17559 2537 17589 2665
rect 17654 2473 17684 2673
rect 17738 2473 17768 2673
rect 17927 2499 18505 2673
rect 18663 2499 18781 2673
<< ndiff >>
rect 1131 7536 1183 7569
rect 1131 7502 1139 7536
rect 1173 7502 1183 7536
rect 1131 7459 1183 7502
rect 1301 7536 1353 7569
rect 1301 7502 1311 7536
rect 1345 7502 1353 7536
rect 1301 7459 1353 7502
rect 1591 7553 1644 7569
rect 1591 7519 1600 7553
rect 1634 7519 1644 7553
rect 1591 7485 1644 7519
rect 1591 7451 1600 7485
rect 1634 7451 1644 7485
rect 1591 7439 1644 7451
rect 1674 7527 1728 7569
rect 1674 7493 1684 7527
rect 1718 7493 1728 7527
rect 1674 7439 1728 7493
rect 1758 7557 1823 7569
rect 1758 7523 1770 7557
rect 1804 7523 1823 7557
rect 1758 7485 1823 7523
rect 1853 7544 1905 7569
rect 1853 7510 1863 7544
rect 1897 7510 1905 7544
rect 1853 7485 1905 7510
rect 1959 7538 2011 7569
rect 1959 7504 1967 7538
rect 2001 7504 2011 7538
rect 1758 7439 1808 7485
rect 1959 7459 2011 7504
rect 2957 7538 3009 7569
rect 2957 7504 2967 7538
rect 3001 7504 3009 7538
rect 2957 7459 3009 7504
rect 3063 7538 3115 7569
rect 3063 7504 3071 7538
rect 3105 7504 3115 7538
rect 3063 7459 3115 7504
rect 3509 7538 3561 7569
rect 3983 7553 4036 7569
rect 3509 7504 3519 7538
rect 3553 7504 3561 7538
rect 3509 7459 3561 7504
rect 3983 7519 3992 7553
rect 4026 7519 4036 7553
rect 3983 7485 4036 7519
rect 3983 7451 3992 7485
rect 4026 7451 4036 7485
rect 3983 7439 4036 7451
rect 4066 7527 4120 7569
rect 4066 7493 4076 7527
rect 4110 7493 4120 7527
rect 4066 7439 4120 7493
rect 4150 7557 4215 7569
rect 4150 7523 4162 7557
rect 4196 7523 4215 7557
rect 4150 7485 4215 7523
rect 4245 7544 4297 7569
rect 4245 7510 4255 7544
rect 4289 7510 4297 7544
rect 4245 7485 4297 7510
rect 4351 7538 4403 7569
rect 4351 7504 4359 7538
rect 4393 7504 4403 7538
rect 4150 7439 4200 7485
rect 4351 7459 4403 7504
rect 5349 7538 5401 7569
rect 5349 7504 5359 7538
rect 5393 7504 5401 7538
rect 5349 7459 5401 7504
rect 5639 7553 5692 7569
rect 5639 7519 5648 7553
rect 5682 7519 5692 7553
rect 5639 7485 5692 7519
rect 5639 7451 5648 7485
rect 5682 7451 5692 7485
rect 5639 7439 5692 7451
rect 5722 7527 5776 7569
rect 5722 7493 5732 7527
rect 5766 7493 5776 7527
rect 5722 7439 5776 7493
rect 5806 7557 5871 7569
rect 5806 7523 5818 7557
rect 5852 7523 5871 7557
rect 5806 7485 5871 7523
rect 5901 7544 5953 7569
rect 5901 7510 5911 7544
rect 5945 7510 5953 7544
rect 5901 7485 5953 7510
rect 6007 7536 6059 7569
rect 6007 7502 6015 7536
rect 6049 7502 6059 7536
rect 5806 7439 5856 7485
rect 6007 7459 6059 7502
rect 6177 7536 6229 7569
rect 6177 7502 6187 7536
rect 6221 7502 6229 7536
rect 6177 7459 6229 7502
rect 6375 7538 6427 7569
rect 6375 7504 6383 7538
rect 6417 7504 6427 7538
rect 6375 7459 6427 7504
rect 7373 7538 7425 7569
rect 7373 7504 7383 7538
rect 7417 7504 7425 7538
rect 7373 7459 7425 7504
rect 7479 7531 7531 7569
rect 7479 7497 7487 7531
rect 7521 7497 7531 7531
rect 7479 7459 7531 7497
rect 7741 7531 7793 7569
rect 7741 7497 7751 7531
rect 7785 7497 7793 7531
rect 7741 7459 7793 7497
rect 7847 7544 7899 7569
rect 7847 7510 7855 7544
rect 7889 7510 7899 7544
rect 7847 7485 7899 7510
rect 7929 7557 7994 7569
rect 7929 7523 7948 7557
rect 7982 7523 7994 7557
rect 7929 7485 7994 7523
rect 7944 7439 7994 7485
rect 8024 7527 8078 7569
rect 8024 7493 8034 7527
rect 8068 7493 8078 7527
rect 8024 7439 8078 7493
rect 8108 7553 8161 7569
rect 8108 7519 8118 7553
rect 8152 7519 8161 7553
rect 8108 7485 8161 7519
rect 8108 7451 8118 7485
rect 8152 7451 8161 7485
rect 8215 7538 8267 7569
rect 8215 7504 8223 7538
rect 8257 7504 8267 7538
rect 8215 7459 8267 7504
rect 8661 7538 8713 7569
rect 8661 7504 8671 7538
rect 8705 7504 8713 7538
rect 8661 7459 8713 7504
rect 8108 7439 8161 7451
rect 8951 7538 9003 7569
rect 8951 7504 8959 7538
rect 8993 7504 9003 7538
rect 8951 7459 9003 7504
rect 9397 7538 9449 7569
rect 9397 7504 9407 7538
rect 9441 7504 9449 7538
rect 9397 7459 9449 7504
rect 9687 7531 9739 7569
rect 9687 7497 9695 7531
rect 9729 7497 9739 7531
rect 9687 7459 9739 7497
rect 9949 7531 10001 7569
rect 9949 7497 9959 7531
rect 9993 7497 10001 7531
rect 9949 7459 10001 7497
rect 10055 7549 10108 7569
rect 10055 7515 10063 7549
rect 10097 7515 10108 7549
rect 10055 7485 10108 7515
rect 10138 7553 10203 7569
rect 10138 7519 10149 7553
rect 10183 7519 10203 7553
rect 10138 7485 10203 7519
rect 10233 7549 10287 7569
rect 10233 7515 10243 7549
rect 10277 7515 10287 7549
rect 10233 7485 10287 7515
rect 10317 7553 10369 7569
rect 10317 7519 10327 7553
rect 10361 7519 10369 7553
rect 10317 7485 10369 7519
rect 10423 7538 10475 7569
rect 10423 7504 10431 7538
rect 10465 7504 10475 7538
rect 10423 7459 10475 7504
rect 11053 7538 11105 7569
rect 11053 7504 11063 7538
rect 11097 7504 11105 7538
rect 11053 7459 11105 7504
rect 11159 7536 11211 7569
rect 11159 7502 11167 7536
rect 11201 7502 11211 7536
rect 11159 7459 11211 7502
rect 11329 7536 11381 7569
rect 11329 7502 11339 7536
rect 11373 7502 11381 7536
rect 11329 7459 11381 7502
rect 11527 7538 11579 7569
rect 11527 7504 11535 7538
rect 11569 7504 11579 7538
rect 11527 7459 11579 7504
rect 12157 7538 12209 7569
rect 12157 7504 12167 7538
rect 12201 7504 12209 7538
rect 12157 7459 12209 7504
rect 12263 7544 12315 7569
rect 12263 7510 12271 7544
rect 12305 7510 12315 7544
rect 12263 7485 12315 7510
rect 12345 7557 12410 7569
rect 12345 7523 12364 7557
rect 12398 7523 12410 7557
rect 12345 7485 12410 7523
rect 12360 7439 12410 7485
rect 12440 7527 12494 7569
rect 12440 7493 12450 7527
rect 12484 7493 12494 7527
rect 12440 7439 12494 7493
rect 12524 7553 12577 7569
rect 12524 7519 12534 7553
rect 12568 7519 12577 7553
rect 12524 7485 12577 7519
rect 12524 7451 12534 7485
rect 12568 7451 12577 7485
rect 12631 7538 12683 7569
rect 12631 7504 12639 7538
rect 12673 7504 12683 7538
rect 12631 7459 12683 7504
rect 13629 7538 13681 7569
rect 13629 7504 13639 7538
rect 13673 7504 13681 7538
rect 13629 7459 13681 7504
rect 13735 7536 13787 7569
rect 13735 7502 13743 7536
rect 13777 7502 13787 7536
rect 13735 7459 13787 7502
rect 13905 7536 13957 7569
rect 13905 7502 13915 7536
rect 13949 7502 13957 7536
rect 13905 7459 13957 7502
rect 12524 7439 12577 7451
rect 14103 7531 14155 7569
rect 14103 7497 14111 7531
rect 14145 7497 14155 7531
rect 14103 7459 14155 7497
rect 14365 7531 14417 7569
rect 14365 7497 14375 7531
rect 14409 7497 14417 7531
rect 14365 7459 14417 7497
rect 14471 7544 14523 7569
rect 14471 7510 14479 7544
rect 14513 7510 14523 7544
rect 14471 7485 14523 7510
rect 14553 7557 14618 7569
rect 14553 7523 14572 7557
rect 14606 7523 14618 7557
rect 14553 7485 14618 7523
rect 14568 7439 14618 7485
rect 14648 7527 14702 7569
rect 14648 7493 14658 7527
rect 14692 7493 14702 7527
rect 14648 7439 14702 7493
rect 14732 7553 14785 7569
rect 14732 7519 14742 7553
rect 14776 7519 14785 7553
rect 14732 7485 14785 7519
rect 14732 7451 14742 7485
rect 14776 7451 14785 7485
rect 14839 7538 14891 7569
rect 14839 7504 14847 7538
rect 14881 7504 14891 7538
rect 14839 7459 14891 7504
rect 15837 7538 15889 7569
rect 15837 7504 15847 7538
rect 15881 7504 15889 7538
rect 15837 7459 15889 7504
rect 15943 7538 15995 7569
rect 15943 7504 15951 7538
rect 15985 7504 15995 7538
rect 15943 7459 15995 7504
rect 16389 7538 16441 7569
rect 16389 7504 16399 7538
rect 16433 7504 16441 7538
rect 16389 7459 16441 7504
rect 16863 7544 16915 7569
rect 16863 7510 16871 7544
rect 16905 7510 16915 7544
rect 16863 7485 16915 7510
rect 16945 7557 17010 7569
rect 16945 7523 16964 7557
rect 16998 7523 17010 7557
rect 16945 7485 17010 7523
rect 14732 7439 14785 7451
rect 16960 7439 17010 7485
rect 17040 7527 17094 7569
rect 17040 7493 17050 7527
rect 17084 7493 17094 7527
rect 17040 7439 17094 7493
rect 17124 7553 17177 7569
rect 17124 7519 17134 7553
rect 17168 7519 17177 7553
rect 17124 7485 17177 7519
rect 17124 7451 17134 7485
rect 17168 7451 17177 7485
rect 17231 7538 17283 7569
rect 17231 7504 17239 7538
rect 17273 7504 17283 7538
rect 17231 7459 17283 7504
rect 17861 7538 17913 7569
rect 17861 7504 17871 7538
rect 17905 7504 17913 7538
rect 17861 7459 17913 7504
rect 18059 7544 18111 7569
rect 18059 7510 18067 7544
rect 18101 7510 18111 7544
rect 18059 7485 18111 7510
rect 18141 7557 18206 7569
rect 18141 7523 18160 7557
rect 18194 7523 18206 7557
rect 18141 7485 18206 7523
rect 17124 7439 17177 7451
rect 18156 7439 18206 7485
rect 18236 7527 18290 7569
rect 18236 7493 18246 7527
rect 18280 7493 18290 7527
rect 18236 7439 18290 7493
rect 18320 7553 18373 7569
rect 18320 7519 18330 7553
rect 18364 7519 18373 7553
rect 18320 7485 18373 7519
rect 18320 7451 18330 7485
rect 18364 7451 18373 7485
rect 18611 7536 18663 7569
rect 18611 7502 18619 7536
rect 18653 7502 18663 7536
rect 18611 7459 18663 7502
rect 18781 7536 18833 7569
rect 18781 7502 18791 7536
rect 18825 7502 18833 7536
rect 18781 7459 18833 7502
rect 18320 7439 18373 7451
rect 1131 6642 1183 6685
rect 1131 6608 1139 6642
rect 1173 6608 1183 6642
rect 1131 6575 1183 6608
rect 1301 6642 1353 6685
rect 1301 6608 1311 6642
rect 1345 6608 1353 6642
rect 1301 6575 1353 6608
rect 1407 6640 1459 6685
rect 1407 6606 1415 6640
rect 1449 6606 1459 6640
rect 1407 6575 1459 6606
rect 2405 6640 2457 6685
rect 2405 6606 2415 6640
rect 2449 6606 2457 6640
rect 2405 6575 2457 6606
rect 2511 6640 2563 6685
rect 2511 6606 2519 6640
rect 2553 6606 2563 6640
rect 2511 6575 2563 6606
rect 3509 6640 3561 6685
rect 3509 6606 3519 6640
rect 3553 6606 3561 6640
rect 3509 6575 3561 6606
rect 3799 6640 3851 6685
rect 3799 6606 3807 6640
rect 3841 6606 3851 6640
rect 3799 6575 3851 6606
rect 4797 6640 4849 6685
rect 4797 6606 4807 6640
rect 4841 6606 4849 6640
rect 4797 6575 4849 6606
rect 4903 6640 4955 6685
rect 4903 6606 4911 6640
rect 4945 6606 4955 6640
rect 4903 6575 4955 6606
rect 5901 6640 5953 6685
rect 5901 6606 5911 6640
rect 5945 6606 5953 6640
rect 5901 6575 5953 6606
rect 6007 6640 6059 6685
rect 6007 6606 6015 6640
rect 6049 6606 6059 6640
rect 6007 6575 6059 6606
rect 7005 6640 7057 6685
rect 7005 6606 7015 6640
rect 7049 6606 7057 6640
rect 7005 6575 7057 6606
rect 7111 6640 7163 6685
rect 7111 6606 7119 6640
rect 7153 6606 7163 6640
rect 7111 6575 7163 6606
rect 8109 6640 8161 6685
rect 8109 6606 8119 6640
rect 8153 6606 8161 6640
rect 8109 6575 8161 6606
rect 8215 6640 8267 6685
rect 8215 6606 8223 6640
rect 8257 6606 8267 6640
rect 8215 6575 8267 6606
rect 8661 6640 8713 6685
rect 8661 6606 8671 6640
rect 8705 6606 8713 6640
rect 8661 6575 8713 6606
rect 8951 6640 9003 6685
rect 8951 6606 8959 6640
rect 8993 6606 9003 6640
rect 8951 6575 9003 6606
rect 9949 6640 10001 6685
rect 9949 6606 9959 6640
rect 9993 6606 10001 6640
rect 9949 6575 10001 6606
rect 10055 6640 10107 6685
rect 10055 6606 10063 6640
rect 10097 6606 10107 6640
rect 10055 6575 10107 6606
rect 11053 6640 11105 6685
rect 11053 6606 11063 6640
rect 11097 6606 11105 6640
rect 11053 6575 11105 6606
rect 11159 6640 11211 6685
rect 11159 6606 11167 6640
rect 11201 6606 11211 6640
rect 11159 6575 11211 6606
rect 12157 6640 12209 6685
rect 12157 6606 12167 6640
rect 12201 6606 12209 6640
rect 12157 6575 12209 6606
rect 12263 6640 12315 6685
rect 12263 6606 12271 6640
rect 12305 6606 12315 6640
rect 12263 6575 12315 6606
rect 13261 6640 13313 6685
rect 13261 6606 13271 6640
rect 13305 6606 13313 6640
rect 13261 6575 13313 6606
rect 13367 6640 13419 6685
rect 13367 6606 13375 6640
rect 13409 6606 13419 6640
rect 13367 6575 13419 6606
rect 13813 6640 13865 6685
rect 13813 6606 13823 6640
rect 13857 6606 13865 6640
rect 13813 6575 13865 6606
rect 14103 6640 14155 6685
rect 14103 6606 14111 6640
rect 14145 6606 14155 6640
rect 14103 6575 14155 6606
rect 15101 6640 15153 6685
rect 15101 6606 15111 6640
rect 15145 6606 15153 6640
rect 15101 6575 15153 6606
rect 15207 6640 15259 6685
rect 15207 6606 15215 6640
rect 15249 6606 15259 6640
rect 15207 6575 15259 6606
rect 16205 6640 16257 6685
rect 16205 6606 16215 6640
rect 16249 6606 16257 6640
rect 16205 6575 16257 6606
rect 16311 6640 16363 6685
rect 16311 6606 16319 6640
rect 16353 6606 16363 6640
rect 16311 6575 16363 6606
rect 17309 6640 17361 6685
rect 17309 6606 17319 6640
rect 17353 6606 17361 6640
rect 17309 6575 17361 6606
rect 17415 6640 17467 6685
rect 17415 6606 17423 6640
rect 17457 6606 17467 6640
rect 17415 6575 17467 6606
rect 18413 6640 18465 6685
rect 18413 6606 18423 6640
rect 18457 6606 18465 6640
rect 18413 6575 18465 6606
rect 18611 6642 18663 6685
rect 18611 6608 18619 6642
rect 18653 6608 18663 6642
rect 18611 6575 18663 6608
rect 18781 6642 18833 6685
rect 18781 6608 18791 6642
rect 18825 6608 18833 6642
rect 18781 6575 18833 6608
rect 1131 6448 1183 6481
rect 1131 6414 1139 6448
rect 1173 6414 1183 6448
rect 1131 6371 1183 6414
rect 1301 6448 1353 6481
rect 1301 6414 1311 6448
rect 1345 6414 1353 6448
rect 1301 6371 1353 6414
rect 1407 6450 1459 6481
rect 1407 6416 1415 6450
rect 1449 6416 1459 6450
rect 1407 6371 1459 6416
rect 2405 6450 2457 6481
rect 2405 6416 2415 6450
rect 2449 6416 2457 6450
rect 2405 6371 2457 6416
rect 2511 6450 2563 6481
rect 2511 6416 2519 6450
rect 2553 6416 2563 6450
rect 2511 6371 2563 6416
rect 3509 6450 3561 6481
rect 3509 6416 3519 6450
rect 3553 6416 3561 6450
rect 3509 6371 3561 6416
rect 3615 6450 3667 6481
rect 3615 6416 3623 6450
rect 3657 6416 3667 6450
rect 3615 6371 3667 6416
rect 4613 6450 4665 6481
rect 4613 6416 4623 6450
rect 4657 6416 4665 6450
rect 4613 6371 4665 6416
rect 4719 6450 4771 6481
rect 4719 6416 4727 6450
rect 4761 6416 4771 6450
rect 4719 6371 4771 6416
rect 5717 6450 5769 6481
rect 5717 6416 5727 6450
rect 5761 6416 5769 6450
rect 5717 6371 5769 6416
rect 5823 6443 5875 6481
rect 5823 6409 5831 6443
rect 5865 6409 5875 6443
rect 5823 6371 5875 6409
rect 6085 6443 6137 6481
rect 6085 6409 6095 6443
rect 6129 6409 6137 6443
rect 6085 6371 6137 6409
rect 6375 6450 6427 6481
rect 6375 6416 6383 6450
rect 6417 6416 6427 6450
rect 6375 6371 6427 6416
rect 7373 6450 7425 6481
rect 7373 6416 7383 6450
rect 7417 6416 7425 6450
rect 7373 6371 7425 6416
rect 7479 6450 7531 6481
rect 7479 6416 7487 6450
rect 7521 6416 7531 6450
rect 7479 6371 7531 6416
rect 8477 6450 8529 6481
rect 8477 6416 8487 6450
rect 8521 6416 8529 6450
rect 8477 6371 8529 6416
rect 8583 6450 8635 6481
rect 8583 6416 8591 6450
rect 8625 6416 8635 6450
rect 8583 6371 8635 6416
rect 9581 6450 9633 6481
rect 9581 6416 9591 6450
rect 9625 6416 9633 6450
rect 9581 6371 9633 6416
rect 9687 6450 9739 6481
rect 9687 6416 9695 6450
rect 9729 6416 9739 6450
rect 9687 6371 9739 6416
rect 10685 6450 10737 6481
rect 10685 6416 10695 6450
rect 10729 6416 10737 6450
rect 10685 6371 10737 6416
rect 10791 6450 10843 6481
rect 10791 6416 10799 6450
rect 10833 6416 10843 6450
rect 10791 6371 10843 6416
rect 11237 6450 11289 6481
rect 11237 6416 11247 6450
rect 11281 6416 11289 6450
rect 11237 6371 11289 6416
rect 11527 6450 11579 6481
rect 11527 6416 11535 6450
rect 11569 6416 11579 6450
rect 11527 6371 11579 6416
rect 12525 6450 12577 6481
rect 12525 6416 12535 6450
rect 12569 6416 12577 6450
rect 12525 6371 12577 6416
rect 12631 6450 12683 6481
rect 12631 6416 12639 6450
rect 12673 6416 12683 6450
rect 12631 6371 12683 6416
rect 13629 6450 13681 6481
rect 13629 6416 13639 6450
rect 13673 6416 13681 6450
rect 13629 6371 13681 6416
rect 13735 6450 13787 6481
rect 13735 6416 13743 6450
rect 13777 6416 13787 6450
rect 13735 6371 13787 6416
rect 14733 6450 14785 6481
rect 14733 6416 14743 6450
rect 14777 6416 14785 6450
rect 14733 6371 14785 6416
rect 14839 6450 14891 6481
rect 14839 6416 14847 6450
rect 14881 6416 14891 6450
rect 14839 6371 14891 6416
rect 15837 6450 15889 6481
rect 15837 6416 15847 6450
rect 15881 6416 15889 6450
rect 15837 6371 15889 6416
rect 15943 6450 15995 6481
rect 15943 6416 15951 6450
rect 15985 6416 15995 6450
rect 15943 6371 15995 6416
rect 16389 6450 16441 6481
rect 16389 6416 16399 6450
rect 16433 6416 16441 6450
rect 16389 6371 16441 6416
rect 16679 6450 16731 6481
rect 16679 6416 16687 6450
rect 16721 6416 16731 6450
rect 16679 6371 16731 6416
rect 17677 6450 17729 6481
rect 17677 6416 17687 6450
rect 17721 6416 17729 6450
rect 17677 6371 17729 6416
rect 17783 6450 17835 6481
rect 17783 6416 17791 6450
rect 17825 6416 17835 6450
rect 17783 6371 17835 6416
rect 18413 6450 18465 6481
rect 18413 6416 18423 6450
rect 18457 6416 18465 6450
rect 18413 6371 18465 6416
rect 18611 6448 18663 6481
rect 18611 6414 18619 6448
rect 18653 6414 18663 6448
rect 18611 6371 18663 6414
rect 18781 6448 18833 6481
rect 18781 6414 18791 6448
rect 18825 6414 18833 6448
rect 18781 6371 18833 6414
rect 1131 5554 1183 5597
rect 1131 5520 1139 5554
rect 1173 5520 1183 5554
rect 1131 5487 1183 5520
rect 1301 5554 1353 5597
rect 1301 5520 1311 5554
rect 1345 5520 1353 5554
rect 1301 5487 1353 5520
rect 1407 5552 1459 5597
rect 1407 5518 1415 5552
rect 1449 5518 1459 5552
rect 1407 5487 1459 5518
rect 2037 5552 2089 5597
rect 2037 5518 2047 5552
rect 2081 5518 2089 5552
rect 2037 5487 2089 5518
rect 2235 5546 2287 5591
rect 2235 5512 2243 5546
rect 2277 5512 2287 5546
rect 2235 5487 2287 5512
rect 2317 5533 2375 5591
rect 2317 5499 2329 5533
rect 2363 5499 2375 5533
rect 2317 5487 2375 5499
rect 2405 5563 2457 5591
rect 2405 5529 2415 5563
rect 2449 5529 2457 5563
rect 2405 5487 2457 5529
rect 2511 5552 2563 5597
rect 2511 5518 2519 5552
rect 2553 5518 2563 5552
rect 2511 5487 2563 5518
rect 2957 5552 3009 5597
rect 2957 5518 2967 5552
rect 3001 5518 3009 5552
rect 2957 5487 3009 5518
rect 3063 5563 3115 5591
rect 3063 5529 3071 5563
rect 3105 5529 3115 5563
rect 3063 5487 3115 5529
rect 3145 5533 3203 5591
rect 3145 5499 3157 5533
rect 3191 5499 3203 5533
rect 3145 5487 3203 5499
rect 3233 5546 3285 5591
rect 3233 5512 3243 5546
rect 3277 5512 3285 5546
rect 3233 5487 3285 5512
rect 3339 5559 3391 5597
rect 3339 5525 3347 5559
rect 3381 5525 3391 5559
rect 3339 5487 3391 5525
rect 3601 5559 3653 5597
rect 3601 5525 3611 5559
rect 3645 5525 3653 5559
rect 3601 5487 3653 5525
rect 3799 5552 3851 5597
rect 3799 5518 3807 5552
rect 3841 5518 3851 5552
rect 3799 5487 3851 5518
rect 4797 5552 4849 5597
rect 4797 5518 4807 5552
rect 4841 5518 4849 5552
rect 4797 5487 4849 5518
rect 4903 5552 4955 5597
rect 4903 5518 4911 5552
rect 4945 5518 4955 5552
rect 4903 5487 4955 5518
rect 5901 5552 5953 5597
rect 5901 5518 5911 5552
rect 5945 5518 5953 5552
rect 5901 5487 5953 5518
rect 6007 5552 6059 5597
rect 6007 5518 6015 5552
rect 6049 5518 6059 5552
rect 6007 5487 6059 5518
rect 6637 5552 6689 5597
rect 6637 5518 6647 5552
rect 6681 5518 6689 5552
rect 6637 5487 6689 5518
rect 6743 5552 6795 5617
rect 6743 5518 6751 5552
rect 6785 5518 6795 5552
rect 6743 5487 6795 5518
rect 6825 5571 6877 5617
rect 6825 5533 6904 5571
rect 6825 5499 6835 5533
rect 6869 5499 6904 5533
rect 6825 5487 6904 5499
rect 6934 5487 7000 5571
rect 7030 5548 7125 5571
rect 7030 5514 7042 5548
rect 7076 5514 7125 5548
rect 7030 5487 7125 5514
rect 7155 5487 7221 5571
rect 7251 5548 7389 5571
rect 7251 5514 7277 5548
rect 7311 5514 7345 5548
rect 7379 5514 7389 5548
rect 7251 5487 7389 5514
rect 7419 5548 7471 5571
rect 7419 5514 7429 5548
rect 7463 5514 7471 5548
rect 7419 5487 7471 5514
rect 7571 5552 7623 5597
rect 7571 5518 7579 5552
rect 7613 5518 7623 5552
rect 7571 5487 7623 5518
rect 8569 5552 8621 5597
rect 8569 5518 8579 5552
rect 8613 5518 8621 5552
rect 8569 5487 8621 5518
rect 8951 5552 9003 5597
rect 8951 5518 8959 5552
rect 8993 5518 9003 5552
rect 8951 5487 9003 5518
rect 9581 5552 9633 5597
rect 9581 5518 9591 5552
rect 9625 5518 9633 5552
rect 9581 5487 9633 5518
rect 9871 5552 9923 5617
rect 9871 5518 9879 5552
rect 9913 5518 9923 5552
rect 9871 5487 9923 5518
rect 9953 5571 10005 5617
rect 9953 5533 10032 5571
rect 9953 5499 9963 5533
rect 9997 5499 10032 5533
rect 9953 5487 10032 5499
rect 10062 5487 10128 5571
rect 10158 5548 10253 5571
rect 10158 5514 10170 5548
rect 10204 5514 10253 5548
rect 10158 5487 10253 5514
rect 10283 5487 10349 5571
rect 10379 5548 10517 5571
rect 10379 5514 10405 5548
rect 10439 5514 10473 5548
rect 10507 5514 10517 5548
rect 10379 5487 10517 5514
rect 10547 5548 10599 5571
rect 10547 5514 10557 5548
rect 10591 5514 10599 5548
rect 10547 5487 10599 5514
rect 10699 5559 10751 5597
rect 10699 5525 10707 5559
rect 10741 5525 10751 5559
rect 10699 5487 10751 5525
rect 10961 5559 11013 5597
rect 10961 5525 10971 5559
rect 11005 5525 11013 5559
rect 10961 5487 11013 5525
rect 11107 5533 11163 5617
rect 11107 5499 11119 5533
rect 11153 5499 11163 5533
rect 11107 5487 11163 5499
rect 11193 5599 11245 5617
rect 11193 5533 11271 5599
rect 11193 5499 11203 5533
rect 11237 5515 11271 5533
rect 11301 5515 11355 5599
rect 11385 5561 11441 5599
rect 11385 5527 11395 5561
rect 11429 5527 11441 5561
rect 11385 5515 11441 5527
rect 11527 5552 11579 5597
rect 11527 5518 11535 5552
rect 11569 5518 11579 5552
rect 11237 5499 11245 5515
rect 11193 5487 11245 5499
rect 11527 5487 11579 5518
rect 12157 5552 12209 5597
rect 12157 5518 12167 5552
rect 12201 5518 12209 5552
rect 12157 5487 12209 5518
rect 12263 5552 12315 5617
rect 12263 5518 12271 5552
rect 12305 5518 12315 5552
rect 12263 5487 12315 5518
rect 12345 5571 12397 5617
rect 12345 5533 12424 5571
rect 12345 5499 12355 5533
rect 12389 5499 12424 5533
rect 12345 5487 12424 5499
rect 12454 5487 12520 5571
rect 12550 5548 12645 5571
rect 12550 5514 12562 5548
rect 12596 5514 12645 5548
rect 12550 5487 12645 5514
rect 12675 5487 12741 5571
rect 12771 5548 12909 5571
rect 12771 5514 12797 5548
rect 12831 5514 12865 5548
rect 12899 5514 12909 5548
rect 12771 5487 12909 5514
rect 12939 5548 12991 5571
rect 12939 5514 12949 5548
rect 12983 5514 12991 5548
rect 12939 5487 12991 5514
rect 13091 5552 13143 5597
rect 13091 5518 13099 5552
rect 13133 5518 13143 5552
rect 13091 5487 13143 5518
rect 13721 5552 13773 5597
rect 13721 5518 13731 5552
rect 13765 5518 13773 5552
rect 13721 5487 13773 5518
rect 14287 5552 14339 5617
rect 14287 5518 14295 5552
rect 14329 5518 14339 5552
rect 14287 5487 14339 5518
rect 14369 5571 14421 5617
rect 14369 5533 14448 5571
rect 14369 5499 14379 5533
rect 14413 5499 14448 5533
rect 14369 5487 14448 5499
rect 14478 5487 14544 5571
rect 14574 5548 14669 5571
rect 14574 5514 14586 5548
rect 14620 5514 14669 5548
rect 14574 5487 14669 5514
rect 14699 5487 14765 5571
rect 14795 5548 14933 5571
rect 14795 5514 14821 5548
rect 14855 5514 14889 5548
rect 14923 5514 14933 5548
rect 14795 5487 14933 5514
rect 14963 5548 15015 5571
rect 14963 5514 14973 5548
rect 15007 5514 15015 5548
rect 14963 5487 15015 5514
rect 15115 5552 15167 5597
rect 15115 5518 15123 5552
rect 15157 5518 15167 5552
rect 15115 5487 15167 5518
rect 16113 5552 16165 5597
rect 16113 5518 16123 5552
rect 16157 5518 16165 5552
rect 16113 5487 16165 5518
rect 16219 5552 16271 5597
rect 16219 5518 16227 5552
rect 16261 5518 16271 5552
rect 16219 5487 16271 5518
rect 17217 5552 17269 5597
rect 17217 5518 17227 5552
rect 17261 5518 17269 5552
rect 17217 5487 17269 5518
rect 17323 5552 17375 5597
rect 17323 5518 17331 5552
rect 17365 5518 17375 5552
rect 17323 5487 17375 5518
rect 18321 5552 18373 5597
rect 18321 5518 18331 5552
rect 18365 5518 18373 5552
rect 18321 5487 18373 5518
rect 18611 5554 18663 5597
rect 18611 5520 18619 5554
rect 18653 5520 18663 5554
rect 18611 5487 18663 5520
rect 18781 5554 18833 5597
rect 18781 5520 18791 5554
rect 18825 5520 18833 5554
rect 18781 5487 18833 5520
rect 1131 5360 1183 5393
rect 1131 5326 1139 5360
rect 1173 5326 1183 5360
rect 1131 5283 1183 5326
rect 1301 5360 1353 5393
rect 1301 5326 1311 5360
rect 1345 5326 1353 5360
rect 1301 5283 1353 5326
rect 1407 5362 1459 5393
rect 1407 5328 1415 5362
rect 1449 5328 1459 5362
rect 1407 5283 1459 5328
rect 1853 5362 1905 5393
rect 1853 5328 1863 5362
rect 1897 5328 1905 5362
rect 1853 5283 1905 5328
rect 1999 5381 2055 5393
rect 1999 5347 2011 5381
rect 2045 5347 2055 5381
rect 1999 5263 2055 5347
rect 2085 5381 2137 5393
rect 2085 5347 2095 5381
rect 2129 5365 2137 5381
rect 2129 5347 2163 5365
rect 2085 5281 2163 5347
rect 2193 5281 2247 5365
rect 2277 5353 2333 5365
rect 2277 5319 2287 5353
rect 2321 5319 2333 5353
rect 2277 5281 2333 5319
rect 2419 5355 2471 5393
rect 2419 5321 2427 5355
rect 2461 5321 2471 5355
rect 2419 5283 2471 5321
rect 2681 5355 2733 5393
rect 2681 5321 2691 5355
rect 2725 5321 2733 5355
rect 2681 5283 2733 5321
rect 2919 5381 2975 5393
rect 2919 5347 2931 5381
rect 2965 5347 2975 5381
rect 2085 5263 2137 5281
rect 2919 5263 2975 5347
rect 3005 5381 3057 5393
rect 3005 5347 3015 5381
rect 3049 5365 3057 5381
rect 3049 5347 3083 5365
rect 3005 5281 3083 5347
rect 3113 5281 3167 5365
rect 3197 5353 3253 5365
rect 3197 5319 3207 5353
rect 3241 5319 3253 5353
rect 3197 5281 3253 5319
rect 3339 5355 3391 5393
rect 3339 5321 3347 5355
rect 3381 5321 3391 5355
rect 3339 5283 3391 5321
rect 3601 5355 3653 5393
rect 3601 5321 3611 5355
rect 3645 5321 3653 5355
rect 3601 5283 3653 5321
rect 3707 5368 3759 5393
rect 3707 5334 3715 5368
rect 3749 5334 3759 5368
rect 3707 5309 3759 5334
rect 3789 5381 3854 5393
rect 3789 5347 3808 5381
rect 3842 5347 3854 5381
rect 3789 5309 3854 5347
rect 3005 5263 3057 5281
rect 3804 5263 3854 5309
rect 3884 5351 3938 5393
rect 3884 5317 3894 5351
rect 3928 5317 3938 5351
rect 3884 5263 3938 5317
rect 3968 5377 4021 5393
rect 3968 5343 3978 5377
rect 4012 5343 4021 5377
rect 3968 5309 4021 5343
rect 3968 5275 3978 5309
rect 4012 5275 4021 5309
rect 4075 5355 4127 5393
rect 4075 5321 4083 5355
rect 4117 5321 4127 5355
rect 4075 5283 4127 5321
rect 4337 5355 4389 5393
rect 4337 5321 4347 5355
rect 4381 5321 4389 5355
rect 4337 5283 4389 5321
rect 4445 5381 4497 5393
rect 4445 5347 4453 5381
rect 4487 5347 4497 5381
rect 4445 5309 4497 5347
rect 3968 5263 4021 5275
rect 4445 5275 4453 5309
rect 4487 5275 4497 5309
rect 4445 5263 4497 5275
rect 4527 5381 4581 5393
rect 4527 5347 4537 5381
rect 4571 5347 4581 5381
rect 4527 5309 4581 5347
rect 4527 5275 4537 5309
rect 4571 5275 4581 5309
rect 4527 5263 4581 5275
rect 4611 5381 4663 5393
rect 4611 5347 4621 5381
rect 4655 5347 4663 5381
rect 4611 5309 4663 5347
rect 4611 5275 4621 5309
rect 4655 5275 4663 5309
rect 4719 5362 4771 5393
rect 4719 5328 4727 5362
rect 4761 5328 4771 5362
rect 4719 5283 4771 5328
rect 5717 5362 5769 5393
rect 5717 5328 5727 5362
rect 5761 5328 5769 5362
rect 5717 5283 5769 5328
rect 5823 5351 5875 5393
rect 5823 5317 5831 5351
rect 5865 5317 5875 5351
rect 5823 5289 5875 5317
rect 5905 5381 5963 5393
rect 5905 5347 5917 5381
rect 5951 5347 5963 5381
rect 5905 5289 5963 5347
rect 5993 5368 6045 5393
rect 5993 5334 6003 5368
rect 6037 5334 6045 5368
rect 5993 5289 6045 5334
rect 4611 5263 4663 5275
rect 6375 5360 6427 5393
rect 6375 5326 6383 5360
rect 6417 5326 6427 5360
rect 6375 5283 6427 5326
rect 6545 5360 6597 5393
rect 6545 5326 6555 5360
rect 6589 5326 6597 5360
rect 6545 5283 6597 5326
rect 6651 5362 6703 5393
rect 6651 5328 6659 5362
rect 6693 5328 6703 5362
rect 6651 5263 6703 5328
rect 6733 5381 6812 5393
rect 6733 5347 6743 5381
rect 6777 5347 6812 5381
rect 6733 5309 6812 5347
rect 6842 5309 6908 5393
rect 6938 5366 7033 5393
rect 6938 5332 6950 5366
rect 6984 5332 7033 5366
rect 6938 5309 7033 5332
rect 7063 5309 7129 5393
rect 7159 5366 7297 5393
rect 7159 5332 7185 5366
rect 7219 5332 7253 5366
rect 7287 5332 7297 5366
rect 7159 5309 7297 5332
rect 7327 5366 7379 5393
rect 7327 5332 7337 5366
rect 7371 5332 7379 5366
rect 7327 5309 7379 5332
rect 7479 5355 7531 5393
rect 7479 5321 7487 5355
rect 7521 5321 7531 5355
rect 6733 5263 6785 5309
rect 7479 5283 7531 5321
rect 7741 5355 7793 5393
rect 7741 5321 7751 5355
rect 7785 5321 7793 5355
rect 7741 5283 7793 5321
rect 7847 5362 7899 5393
rect 7847 5328 7855 5362
rect 7889 5328 7899 5362
rect 7847 5263 7899 5328
rect 7929 5381 8008 5393
rect 7929 5347 7939 5381
rect 7973 5347 8008 5381
rect 7929 5309 8008 5347
rect 8038 5309 8104 5393
rect 8134 5366 8229 5393
rect 8134 5332 8146 5366
rect 8180 5332 8229 5366
rect 8134 5309 8229 5332
rect 8259 5309 8325 5393
rect 8355 5366 8493 5393
rect 8355 5332 8381 5366
rect 8415 5332 8449 5366
rect 8483 5332 8493 5366
rect 8355 5309 8493 5332
rect 8523 5366 8575 5393
rect 8523 5332 8533 5366
rect 8567 5332 8575 5366
rect 8523 5309 8575 5332
rect 8675 5355 8727 5393
rect 8675 5321 8683 5355
rect 8717 5321 8727 5355
rect 7929 5263 7981 5309
rect 8675 5283 8727 5321
rect 8937 5355 8989 5393
rect 8937 5321 8947 5355
rect 8981 5321 8989 5355
rect 8937 5283 8989 5321
rect 9135 5378 9187 5393
rect 9135 5344 9143 5378
rect 9177 5344 9187 5378
rect 9135 5310 9187 5344
rect 9135 5276 9143 5310
rect 9177 5276 9187 5310
rect 9135 5263 9187 5276
rect 9217 5381 9269 5393
rect 9217 5347 9227 5381
rect 9261 5347 9269 5381
rect 9217 5263 9269 5347
rect 9323 5377 9375 5393
rect 9323 5343 9331 5377
rect 9365 5343 9375 5377
rect 9323 5309 9375 5343
rect 9323 5275 9331 5309
rect 9365 5275 9375 5309
rect 9323 5263 9375 5275
rect 9405 5313 9467 5393
rect 9405 5279 9423 5313
rect 9457 5279 9467 5313
rect 9405 5263 9467 5279
rect 9497 5381 9551 5393
rect 9497 5347 9507 5381
rect 9541 5347 9551 5381
rect 9497 5263 9551 5347
rect 9581 5377 9633 5393
rect 9581 5343 9591 5377
rect 9625 5343 9633 5377
rect 9581 5309 9633 5343
rect 9581 5275 9591 5309
rect 9625 5275 9633 5309
rect 9687 5362 9739 5393
rect 9687 5328 9695 5362
rect 9729 5328 9739 5362
rect 9687 5283 9739 5328
rect 10317 5362 10369 5393
rect 10317 5328 10327 5362
rect 10361 5328 10369 5362
rect 10317 5283 10369 5328
rect 10423 5362 10475 5393
rect 10423 5328 10431 5362
rect 10465 5328 10475 5362
rect 9581 5263 9633 5275
rect 10423 5263 10475 5328
rect 10505 5381 10584 5393
rect 10505 5347 10515 5381
rect 10549 5347 10584 5381
rect 10505 5309 10584 5347
rect 10614 5309 10680 5393
rect 10710 5366 10805 5393
rect 10710 5332 10722 5366
rect 10756 5332 10805 5366
rect 10710 5309 10805 5332
rect 10835 5309 10901 5393
rect 10931 5366 11069 5393
rect 10931 5332 10957 5366
rect 10991 5332 11025 5366
rect 11059 5332 11069 5366
rect 10931 5309 11069 5332
rect 11099 5366 11151 5393
rect 11099 5332 11109 5366
rect 11143 5332 11151 5366
rect 11099 5309 11151 5332
rect 10505 5263 10557 5309
rect 11527 5362 11579 5393
rect 11527 5328 11535 5362
rect 11569 5328 11579 5362
rect 11527 5283 11579 5328
rect 12525 5362 12577 5393
rect 12525 5328 12535 5362
rect 12569 5328 12577 5362
rect 12525 5283 12577 5328
rect 12631 5355 12683 5393
rect 12631 5321 12639 5355
rect 12673 5321 12683 5355
rect 12631 5283 12683 5321
rect 12893 5355 12945 5393
rect 12893 5321 12903 5355
rect 12937 5321 12945 5355
rect 12893 5283 12945 5321
rect 13091 5362 13143 5393
rect 13091 5328 13099 5362
rect 13133 5328 13143 5362
rect 13091 5263 13143 5328
rect 13173 5381 13252 5393
rect 13173 5347 13183 5381
rect 13217 5347 13252 5381
rect 13173 5309 13252 5347
rect 13282 5309 13348 5393
rect 13378 5366 13473 5393
rect 13378 5332 13390 5366
rect 13424 5332 13473 5366
rect 13378 5309 13473 5332
rect 13503 5309 13569 5393
rect 13599 5366 13737 5393
rect 13599 5332 13625 5366
rect 13659 5332 13693 5366
rect 13727 5332 13737 5366
rect 13599 5309 13737 5332
rect 13767 5366 13819 5393
rect 13767 5332 13777 5366
rect 13811 5332 13819 5366
rect 13767 5309 13819 5332
rect 13919 5362 13971 5393
rect 13919 5328 13927 5362
rect 13961 5328 13971 5362
rect 13173 5263 13225 5309
rect 13919 5283 13971 5328
rect 14917 5362 14969 5393
rect 14917 5328 14927 5362
rect 14961 5328 14969 5362
rect 14917 5283 14969 5328
rect 15023 5362 15075 5393
rect 15023 5328 15031 5362
rect 15065 5328 15075 5362
rect 15023 5283 15075 5328
rect 16021 5362 16073 5393
rect 16021 5328 16031 5362
rect 16065 5328 16073 5362
rect 16021 5283 16073 5328
rect 16127 5355 16179 5393
rect 16127 5321 16135 5355
rect 16169 5321 16179 5355
rect 16127 5283 16179 5321
rect 16389 5355 16441 5393
rect 16389 5321 16399 5355
rect 16433 5321 16441 5355
rect 16389 5283 16441 5321
rect 16679 5362 16731 5393
rect 16679 5328 16687 5362
rect 16721 5328 16731 5362
rect 16679 5283 16731 5328
rect 17677 5362 17729 5393
rect 17677 5328 17687 5362
rect 17721 5328 17729 5362
rect 17677 5283 17729 5328
rect 17783 5362 17835 5393
rect 17783 5328 17791 5362
rect 17825 5328 17835 5362
rect 17783 5283 17835 5328
rect 18413 5362 18465 5393
rect 18413 5328 18423 5362
rect 18457 5328 18465 5362
rect 18413 5283 18465 5328
rect 18611 5360 18663 5393
rect 18611 5326 18619 5360
rect 18653 5326 18663 5360
rect 18611 5283 18663 5326
rect 18781 5360 18833 5393
rect 18781 5326 18791 5360
rect 18825 5326 18833 5360
rect 18781 5283 18833 5326
rect 1131 4466 1183 4509
rect 1131 4432 1139 4466
rect 1173 4432 1183 4466
rect 1131 4399 1183 4432
rect 1301 4466 1353 4509
rect 1301 4432 1311 4466
rect 1345 4432 1353 4466
rect 1301 4399 1353 4432
rect 1407 4464 1459 4509
rect 1407 4430 1415 4464
rect 1449 4430 1459 4464
rect 1407 4399 1459 4430
rect 1853 4464 1905 4509
rect 1853 4430 1863 4464
rect 1897 4430 1905 4464
rect 1853 4399 1905 4430
rect 2051 4471 2103 4483
rect 2051 4437 2059 4471
rect 2093 4437 2103 4471
rect 2051 4399 2103 4437
rect 2133 4445 2187 4483
rect 2133 4411 2143 4445
rect 2177 4411 2187 4445
rect 2133 4399 2187 4411
rect 2217 4471 2269 4483
rect 2217 4437 2227 4471
rect 2261 4437 2269 4471
rect 2217 4399 2269 4437
rect 2323 4445 2375 4483
rect 2323 4411 2331 4445
rect 2365 4411 2375 4445
rect 2323 4399 2375 4411
rect 2405 4471 2455 4483
rect 2754 4483 2804 4527
rect 2635 4471 2685 4483
rect 2405 4459 2487 4471
rect 2405 4425 2416 4459
rect 2450 4425 2487 4459
rect 2405 4399 2487 4425
rect 2517 4459 2586 4471
rect 2517 4425 2527 4459
rect 2561 4425 2586 4459
rect 2517 4399 2586 4425
rect 2616 4399 2685 4471
rect 2715 4453 2804 4483
rect 2715 4419 2726 4453
rect 2760 4419 2804 4453
rect 2715 4399 2804 4419
rect 2834 4471 2884 4527
rect 3243 4514 3295 4529
rect 3056 4471 3106 4483
rect 2834 4459 2905 4471
rect 2834 4425 2845 4459
rect 2879 4425 2905 4459
rect 2834 4399 2905 4425
rect 2935 4459 3011 4471
rect 2935 4425 2948 4459
rect 2982 4425 3011 4459
rect 2935 4399 3011 4425
rect 3041 4399 3106 4471
rect 3136 4459 3188 4483
rect 3136 4425 3146 4459
rect 3180 4425 3188 4459
rect 3136 4399 3188 4425
rect 3243 4480 3251 4514
rect 3285 4480 3295 4514
rect 3243 4446 3295 4480
rect 3243 4412 3251 4446
rect 3285 4412 3295 4446
rect 3243 4399 3295 4412
rect 3325 4475 3379 4529
rect 3325 4441 3335 4475
rect 3369 4441 3379 4475
rect 3325 4399 3379 4441
rect 3409 4516 3461 4529
rect 3409 4482 3419 4516
rect 3453 4482 3461 4516
rect 3409 4448 3461 4482
rect 3409 4414 3419 4448
rect 3453 4414 3461 4448
rect 4023 4445 4079 4529
rect 3409 4399 3461 4414
rect 4023 4411 4035 4445
rect 4069 4411 4079 4445
rect 4023 4399 4079 4411
rect 4109 4511 4161 4529
rect 4109 4445 4187 4511
rect 4109 4411 4119 4445
rect 4153 4427 4187 4445
rect 4217 4427 4271 4511
rect 4301 4473 4357 4511
rect 4903 4516 4955 4529
rect 4301 4439 4311 4473
rect 4345 4439 4357 4473
rect 4301 4427 4357 4439
rect 4443 4471 4495 4509
rect 4443 4437 4451 4471
rect 4485 4437 4495 4471
rect 4153 4411 4161 4427
rect 4109 4399 4161 4411
rect 4443 4399 4495 4437
rect 4705 4471 4757 4509
rect 4705 4437 4715 4471
rect 4749 4437 4757 4471
rect 4705 4399 4757 4437
rect 4903 4482 4911 4516
rect 4945 4482 4955 4516
rect 4903 4448 4955 4482
rect 4903 4414 4911 4448
rect 4945 4414 4955 4448
rect 4903 4399 4955 4414
rect 4985 4445 5037 4529
rect 4985 4411 4995 4445
rect 5029 4411 5037 4445
rect 4985 4399 5037 4411
rect 5091 4517 5143 4529
rect 5091 4483 5099 4517
rect 5133 4483 5143 4517
rect 5091 4449 5143 4483
rect 5091 4415 5099 4449
rect 5133 4415 5143 4449
rect 5091 4399 5143 4415
rect 5173 4513 5235 4529
rect 5173 4479 5191 4513
rect 5225 4479 5235 4513
rect 5173 4399 5235 4479
rect 5265 4445 5319 4529
rect 5265 4411 5275 4445
rect 5309 4411 5319 4445
rect 5265 4399 5319 4411
rect 5349 4517 5401 4529
rect 5349 4483 5359 4517
rect 5393 4483 5401 4517
rect 5823 4516 5875 4529
rect 5349 4449 5401 4483
rect 5349 4415 5359 4449
rect 5393 4415 5401 4449
rect 5349 4399 5401 4415
rect 5455 4471 5507 4509
rect 5455 4437 5463 4471
rect 5497 4437 5507 4471
rect 5455 4399 5507 4437
rect 5717 4471 5769 4509
rect 5717 4437 5727 4471
rect 5761 4437 5769 4471
rect 5717 4399 5769 4437
rect 5823 4482 5831 4516
rect 5865 4482 5875 4516
rect 5823 4448 5875 4482
rect 5823 4414 5831 4448
rect 5865 4414 5875 4448
rect 5823 4399 5875 4414
rect 5905 4445 5957 4529
rect 5905 4411 5915 4445
rect 5949 4411 5957 4445
rect 5905 4399 5957 4411
rect 6011 4517 6063 4529
rect 6011 4483 6019 4517
rect 6053 4483 6063 4517
rect 6011 4449 6063 4483
rect 6011 4415 6019 4449
rect 6053 4415 6063 4449
rect 6011 4399 6063 4415
rect 6093 4513 6155 4529
rect 6093 4479 6111 4513
rect 6145 4479 6155 4513
rect 6093 4399 6155 4479
rect 6185 4445 6239 4529
rect 6185 4411 6195 4445
rect 6229 4411 6239 4445
rect 6185 4399 6239 4411
rect 6269 4517 6321 4529
rect 6269 4483 6279 4517
rect 6313 4483 6321 4517
rect 6269 4449 6321 4483
rect 6269 4415 6279 4449
rect 6313 4415 6321 4449
rect 6269 4399 6321 4415
rect 6375 4471 6427 4509
rect 6375 4437 6383 4471
rect 6417 4437 6427 4471
rect 6375 4399 6427 4437
rect 6637 4471 6689 4509
rect 6637 4437 6647 4471
rect 6681 4437 6689 4471
rect 6637 4399 6689 4437
rect 6743 4471 6795 4483
rect 6743 4437 6751 4471
rect 6785 4437 6795 4471
rect 6743 4399 6795 4437
rect 6825 4445 6879 4483
rect 6825 4411 6835 4445
rect 6869 4411 6879 4445
rect 6825 4399 6879 4411
rect 6909 4471 6961 4483
rect 6909 4437 6919 4471
rect 6953 4437 6961 4471
rect 6909 4399 6961 4437
rect 7015 4445 7067 4483
rect 7015 4411 7023 4445
rect 7057 4411 7067 4445
rect 7015 4399 7067 4411
rect 7097 4471 7147 4483
rect 7446 4483 7496 4527
rect 7327 4471 7377 4483
rect 7097 4459 7179 4471
rect 7097 4425 7108 4459
rect 7142 4425 7179 4459
rect 7097 4399 7179 4425
rect 7209 4459 7278 4471
rect 7209 4425 7219 4459
rect 7253 4425 7278 4459
rect 7209 4399 7278 4425
rect 7308 4399 7377 4471
rect 7407 4453 7496 4483
rect 7407 4419 7418 4453
rect 7452 4419 7496 4453
rect 7407 4399 7496 4419
rect 7526 4471 7576 4527
rect 7935 4514 7987 4529
rect 7748 4471 7798 4483
rect 7526 4459 7597 4471
rect 7526 4425 7537 4459
rect 7571 4425 7597 4459
rect 7526 4399 7597 4425
rect 7627 4459 7703 4471
rect 7627 4425 7640 4459
rect 7674 4425 7703 4459
rect 7627 4399 7703 4425
rect 7733 4399 7798 4471
rect 7828 4459 7880 4483
rect 7828 4425 7838 4459
rect 7872 4425 7880 4459
rect 7828 4399 7880 4425
rect 7935 4480 7943 4514
rect 7977 4480 7987 4514
rect 7935 4446 7987 4480
rect 7935 4412 7943 4446
rect 7977 4412 7987 4446
rect 7935 4399 7987 4412
rect 8017 4475 8071 4529
rect 8017 4441 8027 4475
rect 8061 4441 8071 4475
rect 8017 4399 8071 4441
rect 8101 4516 8153 4529
rect 8101 4482 8111 4516
rect 8145 4482 8153 4516
rect 8101 4448 8153 4482
rect 8101 4414 8111 4448
rect 8145 4414 8153 4448
rect 8101 4399 8153 4414
rect 8215 4464 8267 4509
rect 8215 4430 8223 4464
rect 8257 4430 8267 4464
rect 8215 4399 8267 4430
rect 8661 4464 8713 4509
rect 8661 4430 8671 4464
rect 8705 4430 8713 4464
rect 8661 4399 8713 4430
rect 9971 4516 10023 4529
rect 8951 4464 9003 4509
rect 8951 4430 8959 4464
rect 8993 4430 9003 4464
rect 8951 4399 9003 4430
rect 9581 4464 9633 4509
rect 9581 4430 9591 4464
rect 9625 4430 9633 4464
rect 9581 4399 9633 4430
rect 9687 4466 9739 4509
rect 9687 4432 9695 4466
rect 9729 4432 9739 4466
rect 9687 4399 9739 4432
rect 9857 4466 9909 4509
rect 9857 4432 9867 4466
rect 9901 4432 9909 4466
rect 9857 4399 9909 4432
rect 9971 4482 9979 4516
rect 10013 4482 10023 4516
rect 9971 4448 10023 4482
rect 9971 4414 9979 4448
rect 10013 4414 10023 4448
rect 9971 4399 10023 4414
rect 10053 4475 10107 4529
rect 10053 4441 10063 4475
rect 10097 4441 10107 4475
rect 10053 4399 10107 4441
rect 10137 4514 10189 4529
rect 10137 4480 10147 4514
rect 10181 4480 10189 4514
rect 10137 4446 10189 4480
rect 10137 4412 10147 4446
rect 10181 4412 10189 4446
rect 10137 4399 10189 4412
rect 10244 4459 10296 4483
rect 10244 4425 10252 4459
rect 10286 4425 10296 4459
rect 10244 4399 10296 4425
rect 10326 4471 10376 4483
rect 10548 4471 10598 4527
rect 10326 4399 10391 4471
rect 10421 4459 10497 4471
rect 10421 4425 10450 4459
rect 10484 4425 10497 4459
rect 10421 4399 10497 4425
rect 10527 4459 10598 4471
rect 10527 4425 10553 4459
rect 10587 4425 10598 4459
rect 10527 4399 10598 4425
rect 10628 4483 10678 4527
rect 10628 4453 10717 4483
rect 10628 4419 10672 4453
rect 10706 4419 10717 4453
rect 10628 4399 10717 4419
rect 10747 4471 10797 4483
rect 11803 4516 11855 4529
rect 10977 4471 11027 4483
rect 10747 4399 10816 4471
rect 10846 4459 10915 4471
rect 10846 4425 10871 4459
rect 10905 4425 10915 4459
rect 10846 4399 10915 4425
rect 10945 4459 11027 4471
rect 10945 4425 10982 4459
rect 11016 4425 11027 4459
rect 10945 4399 11027 4425
rect 11057 4445 11109 4483
rect 11057 4411 11067 4445
rect 11101 4411 11109 4445
rect 11057 4399 11109 4411
rect 11163 4471 11215 4483
rect 11163 4437 11171 4471
rect 11205 4437 11215 4471
rect 11163 4399 11215 4437
rect 11245 4445 11299 4483
rect 11245 4411 11255 4445
rect 11289 4411 11299 4445
rect 11245 4399 11299 4411
rect 11329 4471 11381 4483
rect 11329 4437 11339 4471
rect 11373 4437 11381 4471
rect 11329 4399 11381 4437
rect 11435 4471 11487 4509
rect 11435 4437 11443 4471
rect 11477 4437 11487 4471
rect 11435 4399 11487 4437
rect 11697 4471 11749 4509
rect 11697 4437 11707 4471
rect 11741 4437 11749 4471
rect 11697 4399 11749 4437
rect 11803 4482 11811 4516
rect 11845 4482 11855 4516
rect 11803 4448 11855 4482
rect 11803 4414 11811 4448
rect 11845 4414 11855 4448
rect 11803 4399 11855 4414
rect 11885 4445 11937 4529
rect 11885 4411 11895 4445
rect 11929 4411 11937 4445
rect 11885 4399 11937 4411
rect 11991 4517 12043 4529
rect 11991 4483 11999 4517
rect 12033 4483 12043 4517
rect 11991 4449 12043 4483
rect 11991 4415 11999 4449
rect 12033 4415 12043 4449
rect 11991 4399 12043 4415
rect 12073 4513 12135 4529
rect 12073 4479 12091 4513
rect 12125 4479 12135 4513
rect 12073 4399 12135 4479
rect 12165 4445 12219 4529
rect 12165 4411 12175 4445
rect 12209 4411 12219 4445
rect 12165 4399 12219 4411
rect 12249 4517 12301 4529
rect 12249 4483 12259 4517
rect 12293 4483 12301 4517
rect 12723 4516 12775 4529
rect 12249 4449 12301 4483
rect 12249 4415 12259 4449
rect 12293 4415 12301 4449
rect 12249 4399 12301 4415
rect 12355 4471 12407 4509
rect 12355 4437 12363 4471
rect 12397 4437 12407 4471
rect 12355 4399 12407 4437
rect 12617 4471 12669 4509
rect 12617 4437 12627 4471
rect 12661 4437 12669 4471
rect 12617 4399 12669 4437
rect 12723 4482 12731 4516
rect 12765 4482 12775 4516
rect 12723 4448 12775 4482
rect 12723 4414 12731 4448
rect 12765 4414 12775 4448
rect 12723 4399 12775 4414
rect 12805 4445 12857 4529
rect 12805 4411 12815 4445
rect 12849 4411 12857 4445
rect 12805 4399 12857 4411
rect 12911 4517 12963 4529
rect 12911 4483 12919 4517
rect 12953 4483 12963 4517
rect 12911 4449 12963 4483
rect 12911 4415 12919 4449
rect 12953 4415 12963 4449
rect 12911 4399 12963 4415
rect 12993 4513 13055 4529
rect 12993 4479 13011 4513
rect 13045 4479 13055 4513
rect 12993 4399 13055 4479
rect 13085 4445 13139 4529
rect 13085 4411 13095 4445
rect 13129 4411 13139 4445
rect 13085 4399 13139 4411
rect 13169 4517 13221 4529
rect 13169 4483 13179 4517
rect 13213 4483 13221 4517
rect 13169 4449 13221 4483
rect 13169 4415 13179 4449
rect 13213 4415 13221 4449
rect 13169 4399 13221 4415
rect 13275 4464 13327 4509
rect 13275 4430 13283 4464
rect 13317 4430 13327 4464
rect 13275 4399 13327 4430
rect 13905 4464 13957 4509
rect 13905 4430 13915 4464
rect 13949 4430 13957 4464
rect 13905 4399 13957 4430
rect 14607 4511 14659 4529
rect 14103 4466 14155 4509
rect 14103 4432 14111 4466
rect 14145 4432 14155 4466
rect 14103 4399 14155 4432
rect 14273 4466 14325 4509
rect 14273 4432 14283 4466
rect 14317 4432 14325 4466
rect 14273 4399 14325 4432
rect 14411 4473 14467 4511
rect 14411 4439 14423 4473
rect 14457 4439 14467 4473
rect 14411 4427 14467 4439
rect 14497 4427 14551 4511
rect 14581 4445 14659 4511
rect 14581 4427 14615 4445
rect 14607 4411 14615 4427
rect 14649 4411 14659 4445
rect 14607 4399 14659 4411
rect 14689 4445 14745 4529
rect 14689 4411 14699 4445
rect 14733 4411 14745 4445
rect 14689 4399 14745 4411
rect 14839 4464 14891 4509
rect 14839 4430 14847 4464
rect 14881 4430 14891 4464
rect 14839 4399 14891 4430
rect 15837 4464 15889 4509
rect 15837 4430 15847 4464
rect 15881 4430 15889 4464
rect 15837 4399 15889 4430
rect 15943 4464 15995 4509
rect 15943 4430 15951 4464
rect 15985 4430 15995 4464
rect 15943 4399 15995 4430
rect 16941 4464 16993 4509
rect 16941 4430 16951 4464
rect 16985 4430 16993 4464
rect 16941 4399 16993 4430
rect 17047 4464 17099 4509
rect 17047 4430 17055 4464
rect 17089 4430 17099 4464
rect 17047 4399 17099 4430
rect 18045 4464 18097 4509
rect 18045 4430 18055 4464
rect 18089 4430 18097 4464
rect 18045 4399 18097 4430
rect 18151 4471 18203 4509
rect 18151 4437 18159 4471
rect 18193 4437 18203 4471
rect 18151 4399 18203 4437
rect 18413 4471 18465 4509
rect 18413 4437 18423 4471
rect 18457 4437 18465 4471
rect 18413 4399 18465 4437
rect 18611 4466 18663 4509
rect 18611 4432 18619 4466
rect 18653 4432 18663 4466
rect 18611 4399 18663 4432
rect 18781 4466 18833 4509
rect 18781 4432 18791 4466
rect 18825 4432 18833 4466
rect 18781 4399 18833 4432
rect 1131 4272 1183 4305
rect 1131 4238 1139 4272
rect 1173 4238 1183 4272
rect 1131 4195 1183 4238
rect 1301 4272 1353 4305
rect 1301 4238 1311 4272
rect 1345 4238 1353 4272
rect 1301 4195 1353 4238
rect 1407 4274 1459 4305
rect 1407 4240 1415 4274
rect 1449 4240 1459 4274
rect 1407 4195 1459 4240
rect 1853 4274 1905 4305
rect 1853 4240 1863 4274
rect 1897 4240 1905 4274
rect 1853 4195 1905 4240
rect 1959 4280 2011 4305
rect 1959 4246 1967 4280
rect 2001 4246 2011 4280
rect 1959 4201 2011 4246
rect 2041 4293 2099 4305
rect 2041 4259 2053 4293
rect 2087 4259 2099 4293
rect 2041 4201 2099 4259
rect 2129 4263 2181 4305
rect 2129 4229 2139 4263
rect 2173 4229 2181 4263
rect 2129 4201 2181 4229
rect 2235 4267 2287 4305
rect 2235 4233 2243 4267
rect 2277 4233 2287 4267
rect 2235 4195 2287 4233
rect 2497 4267 2549 4305
rect 2497 4233 2507 4267
rect 2541 4233 2549 4267
rect 2497 4195 2549 4233
rect 2611 4290 2663 4305
rect 2611 4256 2619 4290
rect 2653 4256 2663 4290
rect 2611 4222 2663 4256
rect 2611 4188 2619 4222
rect 2653 4188 2663 4222
rect 2611 4175 2663 4188
rect 2693 4263 2747 4305
rect 2693 4229 2703 4263
rect 2737 4229 2747 4263
rect 2693 4175 2747 4229
rect 2777 4292 2829 4305
rect 2777 4258 2787 4292
rect 2821 4258 2829 4292
rect 2777 4224 2829 4258
rect 2777 4190 2787 4224
rect 2821 4190 2829 4224
rect 2884 4279 2936 4305
rect 2884 4245 2892 4279
rect 2926 4245 2936 4279
rect 2884 4221 2936 4245
rect 2966 4233 3031 4305
rect 3061 4279 3137 4305
rect 3061 4245 3090 4279
rect 3124 4245 3137 4279
rect 3061 4233 3137 4245
rect 3167 4279 3238 4305
rect 3167 4245 3193 4279
rect 3227 4245 3238 4279
rect 3167 4233 3238 4245
rect 2966 4221 3016 4233
rect 2777 4175 2829 4190
rect 3188 4177 3238 4233
rect 3268 4285 3357 4305
rect 3268 4251 3312 4285
rect 3346 4251 3357 4285
rect 3268 4221 3357 4251
rect 3387 4233 3456 4305
rect 3486 4279 3555 4305
rect 3486 4245 3511 4279
rect 3545 4245 3555 4279
rect 3486 4233 3555 4245
rect 3585 4279 3667 4305
rect 3585 4245 3622 4279
rect 3656 4245 3667 4279
rect 3585 4233 3667 4245
rect 3387 4221 3437 4233
rect 3268 4177 3318 4221
rect 3617 4221 3667 4233
rect 3697 4293 3749 4305
rect 3697 4259 3707 4293
rect 3741 4259 3749 4293
rect 3697 4221 3749 4259
rect 3803 4267 3855 4305
rect 3803 4233 3811 4267
rect 3845 4233 3855 4267
rect 3803 4221 3855 4233
rect 3885 4293 3939 4305
rect 3885 4259 3895 4293
rect 3929 4259 3939 4293
rect 3885 4221 3939 4259
rect 3969 4267 4021 4305
rect 3969 4233 3979 4267
rect 4013 4233 4021 4267
rect 3969 4221 4021 4233
rect 4075 4274 4127 4305
rect 4075 4240 4083 4274
rect 4117 4240 4127 4274
rect 4075 4195 4127 4240
rect 4521 4274 4573 4305
rect 4521 4240 4531 4274
rect 4565 4240 4573 4274
rect 4521 4195 4573 4240
rect 4635 4290 4687 4305
rect 4635 4256 4643 4290
rect 4677 4256 4687 4290
rect 4635 4222 4687 4256
rect 4635 4188 4643 4222
rect 4677 4188 4687 4222
rect 4635 4175 4687 4188
rect 4717 4263 4771 4305
rect 4717 4229 4727 4263
rect 4761 4229 4771 4263
rect 4717 4175 4771 4229
rect 4801 4292 4853 4305
rect 4801 4258 4811 4292
rect 4845 4258 4853 4292
rect 4801 4224 4853 4258
rect 4801 4190 4811 4224
rect 4845 4190 4853 4224
rect 4908 4279 4960 4305
rect 4908 4245 4916 4279
rect 4950 4245 4960 4279
rect 4908 4221 4960 4245
rect 4990 4233 5055 4305
rect 5085 4279 5161 4305
rect 5085 4245 5114 4279
rect 5148 4245 5161 4279
rect 5085 4233 5161 4245
rect 5191 4279 5262 4305
rect 5191 4245 5217 4279
rect 5251 4245 5262 4279
rect 5191 4233 5262 4245
rect 4990 4221 5040 4233
rect 4801 4175 4853 4190
rect 5212 4177 5262 4233
rect 5292 4285 5381 4305
rect 5292 4251 5336 4285
rect 5370 4251 5381 4285
rect 5292 4221 5381 4251
rect 5411 4233 5480 4305
rect 5510 4279 5579 4305
rect 5510 4245 5535 4279
rect 5569 4245 5579 4279
rect 5510 4233 5579 4245
rect 5609 4279 5691 4305
rect 5609 4245 5646 4279
rect 5680 4245 5691 4279
rect 5609 4233 5691 4245
rect 5411 4221 5461 4233
rect 5292 4177 5342 4221
rect 5641 4221 5691 4233
rect 5721 4293 5773 4305
rect 5721 4259 5731 4293
rect 5765 4259 5773 4293
rect 5721 4221 5773 4259
rect 5827 4267 5879 4305
rect 5827 4233 5835 4267
rect 5869 4233 5879 4267
rect 5827 4221 5879 4233
rect 5909 4293 5963 4305
rect 5909 4259 5919 4293
rect 5953 4259 5963 4293
rect 5909 4221 5963 4259
rect 5993 4267 6045 4305
rect 5993 4233 6003 4267
rect 6037 4233 6045 4267
rect 5993 4221 6045 4233
rect 6375 4274 6427 4305
rect 6375 4240 6383 4274
rect 6417 4240 6427 4274
rect 6375 4195 6427 4240
rect 6821 4274 6873 4305
rect 6821 4240 6831 4274
rect 6865 4240 6873 4274
rect 6821 4195 6873 4240
rect 6927 4290 6979 4305
rect 6927 4256 6935 4290
rect 6969 4256 6979 4290
rect 6927 4222 6979 4256
rect 6927 4188 6935 4222
rect 6969 4188 6979 4222
rect 6927 4175 6979 4188
rect 7009 4293 7061 4305
rect 7009 4259 7019 4293
rect 7053 4259 7061 4293
rect 7009 4175 7061 4259
rect 7115 4289 7167 4305
rect 7115 4255 7123 4289
rect 7157 4255 7167 4289
rect 7115 4221 7167 4255
rect 7115 4187 7123 4221
rect 7157 4187 7167 4221
rect 7115 4175 7167 4187
rect 7197 4225 7259 4305
rect 7197 4191 7215 4225
rect 7249 4191 7259 4225
rect 7197 4175 7259 4191
rect 7289 4293 7343 4305
rect 7289 4259 7299 4293
rect 7333 4259 7343 4293
rect 7289 4175 7343 4259
rect 7373 4289 7425 4305
rect 7373 4255 7383 4289
rect 7417 4255 7425 4289
rect 7373 4221 7425 4255
rect 7373 4187 7383 4221
rect 7417 4187 7425 4221
rect 7479 4267 7531 4305
rect 7479 4233 7487 4267
rect 7521 4233 7531 4267
rect 7479 4195 7531 4233
rect 7741 4267 7793 4305
rect 7741 4233 7751 4267
rect 7785 4233 7793 4267
rect 7741 4195 7793 4233
rect 7847 4293 7900 4305
rect 7847 4259 7855 4293
rect 7889 4259 7900 4293
rect 7847 4221 7900 4259
rect 7930 4280 7986 4305
rect 7930 4246 7941 4280
rect 7975 4246 7986 4280
rect 7930 4221 7986 4246
rect 8016 4280 8072 4305
rect 8016 4246 8027 4280
rect 8061 4246 8072 4280
rect 8016 4221 8072 4246
rect 8102 4280 8158 4305
rect 8102 4246 8113 4280
rect 8147 4246 8158 4280
rect 8102 4221 8158 4246
rect 8188 4280 8244 4305
rect 8188 4246 8199 4280
rect 8233 4246 8244 4280
rect 8188 4221 8244 4246
rect 8274 4280 8330 4305
rect 8274 4246 8285 4280
rect 8319 4246 8330 4280
rect 8274 4221 8330 4246
rect 8360 4289 8416 4305
rect 8360 4255 8371 4289
rect 8405 4255 8416 4289
rect 8360 4221 8416 4255
rect 8446 4280 8502 4305
rect 8446 4246 8457 4280
rect 8491 4246 8502 4280
rect 8446 4221 8502 4246
rect 8532 4289 8588 4305
rect 8532 4255 8543 4289
rect 8577 4255 8588 4289
rect 8532 4221 8588 4255
rect 8618 4280 8674 4305
rect 8618 4246 8629 4280
rect 8663 4246 8674 4280
rect 8618 4221 8674 4246
rect 8704 4289 8760 4305
rect 8704 4255 8715 4289
rect 8749 4255 8760 4289
rect 8704 4221 8760 4255
rect 8790 4280 8846 4305
rect 8790 4246 8801 4280
rect 8835 4246 8846 4280
rect 8790 4221 8846 4246
rect 8876 4289 8931 4305
rect 8876 4255 8887 4289
rect 8921 4255 8931 4289
rect 8876 4221 8931 4255
rect 8961 4280 9017 4305
rect 8961 4246 8972 4280
rect 9006 4246 9017 4280
rect 8961 4221 9017 4246
rect 9047 4289 9103 4305
rect 9047 4255 9058 4289
rect 9092 4255 9103 4289
rect 9047 4221 9103 4255
rect 9133 4280 9189 4305
rect 9133 4246 9144 4280
rect 9178 4246 9189 4280
rect 9133 4221 9189 4246
rect 9219 4289 9275 4305
rect 9219 4255 9230 4289
rect 9264 4255 9275 4289
rect 9219 4221 9275 4255
rect 9305 4280 9361 4305
rect 9305 4246 9316 4280
rect 9350 4246 9361 4280
rect 9305 4221 9361 4246
rect 9391 4289 9447 4305
rect 9391 4255 9402 4289
rect 9436 4255 9447 4289
rect 9391 4221 9447 4255
rect 9477 4280 9533 4305
rect 9477 4246 9488 4280
rect 9522 4246 9533 4280
rect 9477 4221 9533 4246
rect 9563 4289 9616 4305
rect 9563 4255 9574 4289
rect 9608 4255 9616 4289
rect 9563 4221 9616 4255
rect 9687 4274 9739 4305
rect 9687 4240 9695 4274
rect 9729 4240 9739 4274
rect 7373 4175 7425 4187
rect 9687 4195 9739 4240
rect 10317 4274 10369 4305
rect 10317 4240 10327 4274
rect 10361 4240 10369 4274
rect 10317 4195 10369 4240
rect 10515 4290 10567 4305
rect 10515 4256 10523 4290
rect 10557 4256 10567 4290
rect 10515 4222 10567 4256
rect 10515 4188 10523 4222
rect 10557 4188 10567 4222
rect 10515 4175 10567 4188
rect 10597 4293 10649 4305
rect 10597 4259 10607 4293
rect 10641 4259 10649 4293
rect 10597 4175 10649 4259
rect 10703 4289 10755 4305
rect 10703 4255 10711 4289
rect 10745 4255 10755 4289
rect 10703 4221 10755 4255
rect 10703 4187 10711 4221
rect 10745 4187 10755 4221
rect 10703 4175 10755 4187
rect 10785 4225 10847 4305
rect 10785 4191 10803 4225
rect 10837 4191 10847 4225
rect 10785 4175 10847 4191
rect 10877 4293 10931 4305
rect 10877 4259 10887 4293
rect 10921 4259 10931 4293
rect 10877 4175 10931 4259
rect 10961 4289 11013 4305
rect 10961 4255 10971 4289
rect 11005 4255 11013 4289
rect 10961 4221 11013 4255
rect 10961 4187 10971 4221
rect 11005 4187 11013 4221
rect 11067 4267 11119 4305
rect 11067 4233 11075 4267
rect 11109 4233 11119 4267
rect 11067 4195 11119 4233
rect 11329 4267 11381 4305
rect 11329 4233 11339 4267
rect 11373 4233 11381 4267
rect 11329 4195 11381 4233
rect 11711 4267 11763 4305
rect 11711 4233 11719 4267
rect 11753 4233 11763 4267
rect 11711 4221 11763 4233
rect 11793 4293 11847 4305
rect 11793 4259 11803 4293
rect 11837 4259 11847 4293
rect 11793 4221 11847 4259
rect 11877 4267 11929 4305
rect 11877 4233 11887 4267
rect 11921 4233 11929 4267
rect 11877 4221 11929 4233
rect 11983 4293 12035 4305
rect 11983 4259 11991 4293
rect 12025 4259 12035 4293
rect 11983 4221 12035 4259
rect 12065 4279 12147 4305
rect 12065 4245 12076 4279
rect 12110 4245 12147 4279
rect 12065 4233 12147 4245
rect 12177 4279 12246 4305
rect 12177 4245 12187 4279
rect 12221 4245 12246 4279
rect 12177 4233 12246 4245
rect 12276 4233 12345 4305
rect 12065 4221 12115 4233
rect 10961 4175 11013 4187
rect 12295 4221 12345 4233
rect 12375 4285 12464 4305
rect 12375 4251 12386 4285
rect 12420 4251 12464 4285
rect 12375 4221 12464 4251
rect 12414 4177 12464 4221
rect 12494 4279 12565 4305
rect 12494 4245 12505 4279
rect 12539 4245 12565 4279
rect 12494 4233 12565 4245
rect 12595 4279 12671 4305
rect 12595 4245 12608 4279
rect 12642 4245 12671 4279
rect 12595 4233 12671 4245
rect 12701 4233 12766 4305
rect 12494 4177 12544 4233
rect 12716 4221 12766 4233
rect 12796 4279 12848 4305
rect 12796 4245 12806 4279
rect 12840 4245 12848 4279
rect 12796 4221 12848 4245
rect 12903 4292 12955 4305
rect 12903 4258 12911 4292
rect 12945 4258 12955 4292
rect 12903 4224 12955 4258
rect 12903 4190 12911 4224
rect 12945 4190 12955 4224
rect 12903 4175 12955 4190
rect 12985 4263 13039 4305
rect 12985 4229 12995 4263
rect 13029 4229 13039 4263
rect 12985 4175 13039 4229
rect 13069 4290 13121 4305
rect 13069 4256 13079 4290
rect 13113 4256 13121 4290
rect 13069 4222 13121 4256
rect 13069 4188 13079 4222
rect 13113 4188 13121 4222
rect 13183 4274 13235 4305
rect 13183 4240 13191 4274
rect 13225 4240 13235 4274
rect 13183 4195 13235 4240
rect 14181 4274 14233 4305
rect 14181 4240 14191 4274
rect 14225 4240 14233 4274
rect 14181 4195 14233 4240
rect 14287 4274 14339 4305
rect 14287 4240 14295 4274
rect 14329 4240 14339 4274
rect 14287 4195 14339 4240
rect 15285 4274 15337 4305
rect 15285 4240 15295 4274
rect 15329 4240 15337 4274
rect 15285 4195 15337 4240
rect 15483 4263 15535 4305
rect 15483 4229 15491 4263
rect 15525 4229 15535 4263
rect 15483 4201 15535 4229
rect 15565 4293 15623 4305
rect 15565 4259 15577 4293
rect 15611 4259 15623 4293
rect 15565 4201 15623 4259
rect 15653 4280 15705 4305
rect 15653 4246 15663 4280
rect 15697 4246 15705 4280
rect 15653 4201 15705 4246
rect 15759 4274 15811 4305
rect 15759 4240 15767 4274
rect 15801 4240 15811 4274
rect 13069 4175 13121 4188
rect 15759 4195 15811 4240
rect 16389 4274 16441 4305
rect 16389 4240 16399 4274
rect 16433 4240 16441 4274
rect 16389 4195 16441 4240
rect 17091 4293 17143 4305
rect 17091 4277 17099 4293
rect 16895 4265 16951 4277
rect 16895 4231 16907 4265
rect 16941 4231 16951 4265
rect 16895 4193 16951 4231
rect 16981 4193 17035 4277
rect 17065 4259 17099 4277
rect 17133 4259 17143 4293
rect 17065 4193 17143 4259
rect 17091 4175 17143 4193
rect 17173 4293 17229 4305
rect 17173 4259 17183 4293
rect 17217 4259 17229 4293
rect 17173 4175 17229 4259
rect 17323 4274 17375 4305
rect 17323 4240 17331 4274
rect 17365 4240 17375 4274
rect 17323 4195 17375 4240
rect 18321 4274 18373 4305
rect 18321 4240 18331 4274
rect 18365 4240 18373 4274
rect 18321 4195 18373 4240
rect 18611 4272 18663 4305
rect 18611 4238 18619 4272
rect 18653 4238 18663 4272
rect 18611 4195 18663 4238
rect 18781 4272 18833 4305
rect 18781 4238 18791 4272
rect 18825 4238 18833 4272
rect 18781 4195 18833 4238
rect 1131 3378 1183 3421
rect 1131 3344 1139 3378
rect 1173 3344 1183 3378
rect 1131 3311 1183 3344
rect 1301 3378 1353 3421
rect 1301 3344 1311 3378
rect 1345 3344 1353 3378
rect 1301 3311 1353 3344
rect 1407 3376 1459 3421
rect 1407 3342 1415 3376
rect 1449 3342 1459 3376
rect 1407 3311 1459 3342
rect 1853 3376 1905 3421
rect 1853 3342 1863 3376
rect 1897 3342 1905 3376
rect 1853 3311 1905 3342
rect 2051 3383 2103 3395
rect 2051 3349 2059 3383
rect 2093 3349 2103 3383
rect 2051 3311 2103 3349
rect 2133 3357 2187 3395
rect 2133 3323 2143 3357
rect 2177 3323 2187 3357
rect 2133 3311 2187 3323
rect 2217 3383 2269 3395
rect 2217 3349 2227 3383
rect 2261 3349 2269 3383
rect 2217 3311 2269 3349
rect 2323 3357 2375 3395
rect 2323 3323 2331 3357
rect 2365 3323 2375 3357
rect 2323 3311 2375 3323
rect 2405 3383 2455 3395
rect 2754 3395 2804 3439
rect 2635 3383 2685 3395
rect 2405 3371 2487 3383
rect 2405 3337 2416 3371
rect 2450 3337 2487 3371
rect 2405 3311 2487 3337
rect 2517 3371 2586 3383
rect 2517 3337 2527 3371
rect 2561 3337 2586 3371
rect 2517 3311 2586 3337
rect 2616 3311 2685 3383
rect 2715 3365 2804 3395
rect 2715 3331 2726 3365
rect 2760 3331 2804 3365
rect 2715 3311 2804 3331
rect 2834 3383 2884 3439
rect 3243 3426 3295 3441
rect 3056 3383 3106 3395
rect 2834 3371 2905 3383
rect 2834 3337 2845 3371
rect 2879 3337 2905 3371
rect 2834 3311 2905 3337
rect 2935 3371 3011 3383
rect 2935 3337 2948 3371
rect 2982 3337 3011 3371
rect 2935 3311 3011 3337
rect 3041 3311 3106 3383
rect 3136 3371 3188 3395
rect 3136 3337 3146 3371
rect 3180 3337 3188 3371
rect 3136 3311 3188 3337
rect 3243 3392 3251 3426
rect 3285 3392 3295 3426
rect 3243 3358 3295 3392
rect 3243 3324 3251 3358
rect 3285 3324 3295 3358
rect 3243 3311 3295 3324
rect 3325 3387 3379 3441
rect 3325 3353 3335 3387
rect 3369 3353 3379 3387
rect 3325 3311 3379 3353
rect 3409 3428 3461 3441
rect 3409 3394 3419 3428
rect 3453 3394 3461 3428
rect 3409 3360 3461 3394
rect 3409 3326 3419 3360
rect 3453 3326 3461 3360
rect 3983 3383 4035 3395
rect 3983 3349 3991 3383
rect 4025 3349 4035 3383
rect 3409 3311 3461 3326
rect 3983 3311 4035 3349
rect 4065 3357 4119 3395
rect 4065 3323 4075 3357
rect 4109 3323 4119 3357
rect 4065 3311 4119 3323
rect 4149 3383 4201 3395
rect 4149 3349 4159 3383
rect 4193 3349 4201 3383
rect 4149 3311 4201 3349
rect 4255 3357 4307 3395
rect 4255 3323 4263 3357
rect 4297 3323 4307 3357
rect 4255 3311 4307 3323
rect 4337 3383 4387 3395
rect 4686 3395 4736 3439
rect 4567 3383 4617 3395
rect 4337 3371 4419 3383
rect 4337 3337 4348 3371
rect 4382 3337 4419 3371
rect 4337 3311 4419 3337
rect 4449 3371 4518 3383
rect 4449 3337 4459 3371
rect 4493 3337 4518 3371
rect 4449 3311 4518 3337
rect 4548 3311 4617 3383
rect 4647 3365 4736 3395
rect 4647 3331 4658 3365
rect 4692 3331 4736 3365
rect 4647 3311 4736 3331
rect 4766 3383 4816 3439
rect 5175 3426 5227 3441
rect 4988 3383 5038 3395
rect 4766 3371 4837 3383
rect 4766 3337 4777 3371
rect 4811 3337 4837 3371
rect 4766 3311 4837 3337
rect 4867 3371 4943 3383
rect 4867 3337 4880 3371
rect 4914 3337 4943 3371
rect 4867 3311 4943 3337
rect 4973 3311 5038 3383
rect 5068 3371 5120 3395
rect 5068 3337 5078 3371
rect 5112 3337 5120 3371
rect 5068 3311 5120 3337
rect 5175 3392 5183 3426
rect 5217 3392 5227 3426
rect 5175 3358 5227 3392
rect 5175 3324 5183 3358
rect 5217 3324 5227 3358
rect 5175 3311 5227 3324
rect 5257 3387 5311 3441
rect 5257 3353 5267 3387
rect 5301 3353 5311 3387
rect 5257 3311 5311 3353
rect 5341 3428 5393 3441
rect 5341 3394 5351 3428
rect 5385 3394 5393 3428
rect 6283 3428 6335 3441
rect 5341 3360 5393 3394
rect 5341 3326 5351 3360
rect 5385 3326 5393 3360
rect 5341 3311 5393 3326
rect 5455 3376 5507 3421
rect 5455 3342 5463 3376
rect 5497 3342 5507 3376
rect 5455 3311 5507 3342
rect 6085 3376 6137 3421
rect 6085 3342 6095 3376
rect 6129 3342 6137 3376
rect 6085 3311 6137 3342
rect 6283 3394 6291 3428
rect 6325 3394 6335 3428
rect 6283 3360 6335 3394
rect 6283 3326 6291 3360
rect 6325 3326 6335 3360
rect 6283 3311 6335 3326
rect 6365 3357 6417 3441
rect 6365 3323 6375 3357
rect 6409 3323 6417 3357
rect 6365 3311 6417 3323
rect 6471 3429 6523 3441
rect 6471 3395 6479 3429
rect 6513 3395 6523 3429
rect 6471 3361 6523 3395
rect 6471 3327 6479 3361
rect 6513 3327 6523 3361
rect 6471 3311 6523 3327
rect 6553 3425 6615 3441
rect 6553 3391 6571 3425
rect 6605 3391 6615 3425
rect 6553 3311 6615 3391
rect 6645 3357 6699 3441
rect 6645 3323 6655 3357
rect 6689 3323 6699 3357
rect 6645 3311 6699 3323
rect 6729 3429 6781 3441
rect 6729 3395 6739 3429
rect 6773 3395 6781 3429
rect 6729 3361 6781 3395
rect 6729 3327 6739 3361
rect 6773 3327 6781 3361
rect 6729 3311 6781 3327
rect 6835 3383 6887 3421
rect 6835 3349 6843 3383
rect 6877 3349 6887 3383
rect 6835 3311 6887 3349
rect 7097 3383 7149 3421
rect 7097 3349 7107 3383
rect 7141 3349 7149 3383
rect 7097 3311 7149 3349
rect 7203 3383 7255 3395
rect 7203 3349 7211 3383
rect 7245 3349 7255 3383
rect 7203 3311 7255 3349
rect 7285 3357 7339 3395
rect 7285 3323 7295 3357
rect 7329 3323 7339 3357
rect 7285 3311 7339 3323
rect 7369 3383 7421 3395
rect 7369 3349 7379 3383
rect 7413 3349 7421 3383
rect 7369 3311 7421 3349
rect 7475 3357 7527 3395
rect 7475 3323 7483 3357
rect 7517 3323 7527 3357
rect 7475 3311 7527 3323
rect 7557 3383 7607 3395
rect 7906 3395 7956 3439
rect 7787 3383 7837 3395
rect 7557 3371 7639 3383
rect 7557 3337 7568 3371
rect 7602 3337 7639 3371
rect 7557 3311 7639 3337
rect 7669 3371 7738 3383
rect 7669 3337 7679 3371
rect 7713 3337 7738 3371
rect 7669 3311 7738 3337
rect 7768 3311 7837 3383
rect 7867 3365 7956 3395
rect 7867 3331 7878 3365
rect 7912 3331 7956 3365
rect 7867 3311 7956 3331
rect 7986 3383 8036 3439
rect 8395 3426 8447 3441
rect 8208 3383 8258 3395
rect 7986 3371 8057 3383
rect 7986 3337 7997 3371
rect 8031 3337 8057 3371
rect 7986 3311 8057 3337
rect 8087 3371 8163 3383
rect 8087 3337 8100 3371
rect 8134 3337 8163 3371
rect 8087 3311 8163 3337
rect 8193 3311 8258 3383
rect 8288 3371 8340 3395
rect 8288 3337 8298 3371
rect 8332 3337 8340 3371
rect 8288 3311 8340 3337
rect 8395 3392 8403 3426
rect 8437 3392 8447 3426
rect 8395 3358 8447 3392
rect 8395 3324 8403 3358
rect 8437 3324 8447 3358
rect 8395 3311 8447 3324
rect 8477 3387 8531 3441
rect 8477 3353 8487 3387
rect 8521 3353 8531 3387
rect 8477 3311 8531 3353
rect 8561 3428 8613 3441
rect 8561 3394 8571 3428
rect 8605 3394 8613 3428
rect 8561 3360 8613 3394
rect 8561 3326 8571 3360
rect 8605 3326 8613 3360
rect 8951 3376 9003 3421
rect 8951 3342 8959 3376
rect 8993 3342 9003 3376
rect 8561 3311 8613 3326
rect 8951 3311 9003 3342
rect 9581 3376 9633 3421
rect 9581 3342 9591 3376
rect 9625 3342 9633 3376
rect 9581 3311 9633 3342
rect 9779 3383 9831 3395
rect 9779 3349 9787 3383
rect 9821 3349 9831 3383
rect 9779 3311 9831 3349
rect 9861 3357 9915 3395
rect 9861 3323 9871 3357
rect 9905 3323 9915 3357
rect 9861 3311 9915 3323
rect 9945 3383 9997 3395
rect 9945 3349 9955 3383
rect 9989 3349 9997 3383
rect 9945 3311 9997 3349
rect 10051 3357 10103 3395
rect 10051 3323 10059 3357
rect 10093 3323 10103 3357
rect 10051 3311 10103 3323
rect 10133 3383 10183 3395
rect 10482 3395 10532 3439
rect 10363 3383 10413 3395
rect 10133 3371 10215 3383
rect 10133 3337 10144 3371
rect 10178 3337 10215 3371
rect 10133 3311 10215 3337
rect 10245 3371 10314 3383
rect 10245 3337 10255 3371
rect 10289 3337 10314 3371
rect 10245 3311 10314 3337
rect 10344 3311 10413 3383
rect 10443 3365 10532 3395
rect 10443 3331 10454 3365
rect 10488 3331 10532 3365
rect 10443 3311 10532 3331
rect 10562 3383 10612 3439
rect 10971 3426 11023 3441
rect 10784 3383 10834 3395
rect 10562 3371 10633 3383
rect 10562 3337 10573 3371
rect 10607 3337 10633 3371
rect 10562 3311 10633 3337
rect 10663 3371 10739 3383
rect 10663 3337 10676 3371
rect 10710 3337 10739 3371
rect 10663 3311 10739 3337
rect 10769 3311 10834 3383
rect 10864 3371 10916 3395
rect 10864 3337 10874 3371
rect 10908 3337 10916 3371
rect 10864 3311 10916 3337
rect 10971 3392 10979 3426
rect 11013 3392 11023 3426
rect 10971 3358 11023 3392
rect 10971 3324 10979 3358
rect 11013 3324 11023 3358
rect 10971 3311 11023 3324
rect 11053 3387 11107 3441
rect 11053 3353 11063 3387
rect 11097 3353 11107 3387
rect 11053 3311 11107 3353
rect 11137 3428 11189 3441
rect 11137 3394 11147 3428
rect 11181 3394 11189 3428
rect 11137 3360 11189 3394
rect 11137 3326 11147 3360
rect 11181 3326 11189 3360
rect 11137 3311 11189 3326
rect 11251 3376 11303 3421
rect 11251 3342 11259 3376
rect 11293 3342 11303 3376
rect 11251 3311 11303 3342
rect 11697 3376 11749 3421
rect 11697 3342 11707 3376
rect 11741 3342 11749 3376
rect 11697 3311 11749 3342
rect 11803 3383 11855 3395
rect 11803 3349 11811 3383
rect 11845 3349 11855 3383
rect 11803 3311 11855 3349
rect 11885 3357 11939 3395
rect 11885 3323 11895 3357
rect 11929 3323 11939 3357
rect 11885 3311 11939 3323
rect 11969 3383 12021 3395
rect 11969 3349 11979 3383
rect 12013 3349 12021 3383
rect 11969 3311 12021 3349
rect 12075 3357 12127 3395
rect 12075 3323 12083 3357
rect 12117 3323 12127 3357
rect 12075 3311 12127 3323
rect 12157 3383 12207 3395
rect 12506 3395 12556 3439
rect 12387 3383 12437 3395
rect 12157 3371 12239 3383
rect 12157 3337 12168 3371
rect 12202 3337 12239 3371
rect 12157 3311 12239 3337
rect 12269 3371 12338 3383
rect 12269 3337 12279 3371
rect 12313 3337 12338 3371
rect 12269 3311 12338 3337
rect 12368 3311 12437 3383
rect 12467 3365 12556 3395
rect 12467 3331 12478 3365
rect 12512 3331 12556 3365
rect 12467 3311 12556 3331
rect 12586 3383 12636 3439
rect 12995 3426 13047 3441
rect 12808 3383 12858 3395
rect 12586 3371 12657 3383
rect 12586 3337 12597 3371
rect 12631 3337 12657 3371
rect 12586 3311 12657 3337
rect 12687 3371 12763 3383
rect 12687 3337 12700 3371
rect 12734 3337 12763 3371
rect 12687 3311 12763 3337
rect 12793 3311 12858 3383
rect 12888 3371 12940 3395
rect 12888 3337 12898 3371
rect 12932 3337 12940 3371
rect 12888 3311 12940 3337
rect 12995 3392 13003 3426
rect 13037 3392 13047 3426
rect 12995 3358 13047 3392
rect 12995 3324 13003 3358
rect 13037 3324 13047 3358
rect 12995 3311 13047 3324
rect 13077 3387 13131 3441
rect 13077 3353 13087 3387
rect 13121 3353 13131 3387
rect 13077 3311 13131 3353
rect 13161 3428 13213 3441
rect 13161 3394 13171 3428
rect 13205 3394 13213 3428
rect 13161 3360 13213 3394
rect 13161 3326 13171 3360
rect 13205 3326 13213 3360
rect 13161 3311 13213 3326
rect 13275 3376 13327 3421
rect 13275 3342 13283 3376
rect 13317 3342 13327 3376
rect 13275 3311 13327 3342
rect 13905 3376 13957 3421
rect 13905 3342 13915 3376
rect 13949 3342 13957 3376
rect 13905 3311 13957 3342
rect 14103 3376 14155 3421
rect 14103 3342 14111 3376
rect 14145 3342 14155 3376
rect 14103 3311 14155 3342
rect 15101 3376 15153 3421
rect 15101 3342 15111 3376
rect 15145 3342 15153 3376
rect 15101 3311 15153 3342
rect 15207 3376 15259 3421
rect 15207 3342 15215 3376
rect 15249 3342 15259 3376
rect 15207 3311 15259 3342
rect 15653 3376 15705 3421
rect 15653 3342 15663 3376
rect 15697 3342 15705 3376
rect 15653 3311 15705 3342
rect 15759 3387 15811 3415
rect 15759 3353 15767 3387
rect 15801 3353 15811 3387
rect 15759 3311 15811 3353
rect 15841 3357 15899 3415
rect 15841 3323 15853 3357
rect 15887 3323 15899 3357
rect 15841 3311 15899 3323
rect 15929 3370 15981 3415
rect 15929 3336 15939 3370
rect 15973 3336 15981 3370
rect 15929 3311 15981 3336
rect 16035 3383 16087 3421
rect 16035 3349 16043 3383
rect 16077 3349 16087 3383
rect 16035 3311 16087 3349
rect 16297 3383 16349 3421
rect 16297 3349 16307 3383
rect 16341 3349 16349 3383
rect 16297 3311 16349 3349
rect 16443 3357 16499 3441
rect 16443 3323 16455 3357
rect 16489 3323 16499 3357
rect 16443 3311 16499 3323
rect 16529 3423 16581 3441
rect 16529 3357 16607 3423
rect 16529 3323 16539 3357
rect 16573 3339 16607 3357
rect 16637 3339 16691 3423
rect 16721 3385 16777 3423
rect 16721 3351 16731 3385
rect 16765 3351 16777 3385
rect 16721 3339 16777 3351
rect 16863 3383 16915 3421
rect 16863 3349 16871 3383
rect 16905 3349 16915 3383
rect 16573 3323 16581 3339
rect 16529 3311 16581 3323
rect 16863 3311 16915 3349
rect 17125 3383 17177 3421
rect 17125 3349 17135 3383
rect 17169 3349 17177 3383
rect 17125 3311 17177 3349
rect 17271 3357 17327 3441
rect 17271 3323 17283 3357
rect 17317 3323 17327 3357
rect 17271 3311 17327 3323
rect 17357 3423 17409 3441
rect 17357 3357 17435 3423
rect 17357 3323 17367 3357
rect 17401 3339 17435 3357
rect 17465 3339 17519 3423
rect 17549 3385 17605 3423
rect 17549 3351 17559 3385
rect 17593 3351 17605 3385
rect 17549 3339 17605 3351
rect 17691 3376 17743 3421
rect 17691 3342 17699 3376
rect 17733 3342 17743 3376
rect 17401 3323 17409 3339
rect 17357 3311 17409 3323
rect 17691 3311 17743 3342
rect 18321 3376 18373 3421
rect 18321 3342 18331 3376
rect 18365 3342 18373 3376
rect 18321 3311 18373 3342
rect 18611 3378 18663 3421
rect 18611 3344 18619 3378
rect 18653 3344 18663 3378
rect 18611 3311 18663 3344
rect 18781 3378 18833 3421
rect 18781 3344 18791 3378
rect 18825 3344 18833 3378
rect 18781 3311 18833 3344
rect 1131 3184 1183 3217
rect 1131 3150 1139 3184
rect 1173 3150 1183 3184
rect 1131 3107 1183 3150
rect 1301 3184 1353 3217
rect 1301 3150 1311 3184
rect 1345 3150 1353 3184
rect 1301 3107 1353 3150
rect 1407 3179 1459 3217
rect 1407 3145 1415 3179
rect 1449 3145 1459 3179
rect 1407 3107 1459 3145
rect 1669 3179 1721 3217
rect 1669 3145 1679 3179
rect 1713 3145 1721 3179
rect 1669 3107 1721 3145
rect 1867 3197 1920 3217
rect 1867 3163 1875 3197
rect 1909 3163 1920 3197
rect 1867 3133 1920 3163
rect 1950 3201 2015 3217
rect 1950 3167 1961 3201
rect 1995 3167 2015 3201
rect 1950 3133 2015 3167
rect 2045 3197 2099 3217
rect 2045 3163 2055 3197
rect 2089 3163 2099 3197
rect 2045 3133 2099 3163
rect 2129 3201 2181 3217
rect 2129 3167 2139 3201
rect 2173 3167 2181 3201
rect 2129 3133 2181 3167
rect 2235 3179 2287 3217
rect 2235 3145 2243 3179
rect 2277 3145 2287 3179
rect 2235 3107 2287 3145
rect 2497 3179 2549 3217
rect 2497 3145 2507 3179
rect 2541 3145 2549 3179
rect 2497 3107 2549 3145
rect 2620 3201 2673 3217
rect 2620 3167 2628 3201
rect 2662 3167 2673 3201
rect 2620 3133 2673 3167
rect 2703 3192 2759 3217
rect 2703 3158 2714 3192
rect 2748 3158 2759 3192
rect 2703 3133 2759 3158
rect 2789 3201 2845 3217
rect 2789 3167 2800 3201
rect 2834 3167 2845 3201
rect 2789 3133 2845 3167
rect 2875 3192 2931 3217
rect 2875 3158 2886 3192
rect 2920 3158 2931 3192
rect 2875 3133 2931 3158
rect 2961 3201 3017 3217
rect 2961 3167 2972 3201
rect 3006 3167 3017 3201
rect 2961 3133 3017 3167
rect 3047 3192 3103 3217
rect 3047 3158 3058 3192
rect 3092 3158 3103 3192
rect 3047 3133 3103 3158
rect 3133 3201 3189 3217
rect 3133 3167 3144 3201
rect 3178 3167 3189 3201
rect 3133 3133 3189 3167
rect 3219 3192 3275 3217
rect 3219 3158 3230 3192
rect 3264 3158 3275 3192
rect 3219 3133 3275 3158
rect 3305 3201 3360 3217
rect 3305 3167 3315 3201
rect 3349 3167 3360 3201
rect 3305 3133 3360 3167
rect 3390 3192 3446 3217
rect 3390 3158 3401 3192
rect 3435 3158 3446 3192
rect 3390 3133 3446 3158
rect 3476 3201 3532 3217
rect 3476 3167 3487 3201
rect 3521 3167 3532 3201
rect 3476 3133 3532 3167
rect 3562 3192 3618 3217
rect 3562 3158 3573 3192
rect 3607 3158 3618 3192
rect 3562 3133 3618 3158
rect 3648 3201 3704 3217
rect 3648 3167 3659 3201
rect 3693 3167 3704 3201
rect 3648 3133 3704 3167
rect 3734 3192 3790 3217
rect 3734 3158 3745 3192
rect 3779 3158 3790 3192
rect 3734 3133 3790 3158
rect 3820 3201 3876 3217
rect 3820 3167 3831 3201
rect 3865 3167 3876 3201
rect 3820 3133 3876 3167
rect 3906 3192 3962 3217
rect 3906 3158 3917 3192
rect 3951 3158 3962 3192
rect 3906 3133 3962 3158
rect 3992 3192 4048 3217
rect 3992 3158 4003 3192
rect 4037 3158 4048 3192
rect 3992 3133 4048 3158
rect 4078 3192 4134 3217
rect 4078 3158 4089 3192
rect 4123 3158 4134 3192
rect 4078 3133 4134 3158
rect 4164 3192 4220 3217
rect 4164 3158 4175 3192
rect 4209 3158 4220 3192
rect 4164 3133 4220 3158
rect 4250 3192 4306 3217
rect 4250 3158 4261 3192
rect 4295 3158 4306 3192
rect 4250 3133 4306 3158
rect 4336 3205 4389 3217
rect 4336 3171 4347 3205
rect 4381 3171 4389 3205
rect 4336 3133 4389 3171
rect 4443 3186 4495 3217
rect 4443 3152 4451 3186
rect 4485 3152 4495 3186
rect 4443 3107 4495 3152
rect 5441 3186 5493 3217
rect 5441 3152 5451 3186
rect 5485 3152 5493 3186
rect 5441 3107 5493 3152
rect 5547 3186 5599 3217
rect 5547 3152 5555 3186
rect 5589 3152 5599 3186
rect 5547 3107 5599 3152
rect 6177 3186 6229 3217
rect 6177 3152 6187 3186
rect 6221 3152 6229 3186
rect 6177 3107 6229 3152
rect 6375 3186 6427 3217
rect 6375 3152 6383 3186
rect 6417 3152 6427 3186
rect 6375 3107 6427 3152
rect 7005 3186 7057 3217
rect 7005 3152 7015 3186
rect 7049 3152 7057 3186
rect 7005 3107 7057 3152
rect 7387 3179 7439 3217
rect 7387 3145 7395 3179
rect 7429 3145 7439 3179
rect 7387 3107 7439 3145
rect 7649 3179 7701 3217
rect 7649 3145 7659 3179
rect 7693 3145 7701 3179
rect 7649 3107 7701 3145
rect 7755 3205 7808 3217
rect 7755 3171 7763 3205
rect 7797 3171 7808 3205
rect 7755 3133 7808 3171
rect 7838 3192 7894 3217
rect 7838 3158 7849 3192
rect 7883 3158 7894 3192
rect 7838 3133 7894 3158
rect 7924 3192 7980 3217
rect 7924 3158 7935 3192
rect 7969 3158 7980 3192
rect 7924 3133 7980 3158
rect 8010 3192 8066 3217
rect 8010 3158 8021 3192
rect 8055 3158 8066 3192
rect 8010 3133 8066 3158
rect 8096 3192 8152 3217
rect 8096 3158 8107 3192
rect 8141 3158 8152 3192
rect 8096 3133 8152 3158
rect 8182 3192 8238 3217
rect 8182 3158 8193 3192
rect 8227 3158 8238 3192
rect 8182 3133 8238 3158
rect 8268 3201 8324 3217
rect 8268 3167 8279 3201
rect 8313 3167 8324 3201
rect 8268 3133 8324 3167
rect 8354 3192 8410 3217
rect 8354 3158 8365 3192
rect 8399 3158 8410 3192
rect 8354 3133 8410 3158
rect 8440 3201 8496 3217
rect 8440 3167 8451 3201
rect 8485 3167 8496 3201
rect 8440 3133 8496 3167
rect 8526 3192 8582 3217
rect 8526 3158 8537 3192
rect 8571 3158 8582 3192
rect 8526 3133 8582 3158
rect 8612 3201 8668 3217
rect 8612 3167 8623 3201
rect 8657 3167 8668 3201
rect 8612 3133 8668 3167
rect 8698 3192 8754 3217
rect 8698 3158 8709 3192
rect 8743 3158 8754 3192
rect 8698 3133 8754 3158
rect 8784 3201 8839 3217
rect 8784 3167 8795 3201
rect 8829 3167 8839 3201
rect 8784 3133 8839 3167
rect 8869 3192 8925 3217
rect 8869 3158 8880 3192
rect 8914 3158 8925 3192
rect 8869 3133 8925 3158
rect 8955 3201 9011 3217
rect 8955 3167 8966 3201
rect 9000 3167 9011 3201
rect 8955 3133 9011 3167
rect 9041 3192 9097 3217
rect 9041 3158 9052 3192
rect 9086 3158 9097 3192
rect 9041 3133 9097 3158
rect 9127 3201 9183 3217
rect 9127 3167 9138 3201
rect 9172 3167 9183 3201
rect 9127 3133 9183 3167
rect 9213 3192 9269 3217
rect 9213 3158 9224 3192
rect 9258 3158 9269 3192
rect 9213 3133 9269 3158
rect 9299 3201 9355 3217
rect 9299 3167 9310 3201
rect 9344 3167 9355 3201
rect 9299 3133 9355 3167
rect 9385 3192 9441 3217
rect 9385 3158 9396 3192
rect 9430 3158 9441 3192
rect 9385 3133 9441 3158
rect 9471 3201 9524 3217
rect 9471 3167 9482 3201
rect 9516 3167 9524 3201
rect 9471 3133 9524 3167
rect 9595 3186 9647 3217
rect 9595 3152 9603 3186
rect 9637 3152 9647 3186
rect 9595 3107 9647 3152
rect 10593 3186 10645 3217
rect 10593 3152 10603 3186
rect 10637 3152 10645 3186
rect 10593 3107 10645 3152
rect 10699 3186 10751 3217
rect 10699 3152 10707 3186
rect 10741 3152 10751 3186
rect 10699 3107 10751 3152
rect 11329 3186 11381 3217
rect 11329 3152 11339 3186
rect 11373 3152 11381 3186
rect 11329 3107 11381 3152
rect 11711 3179 11763 3217
rect 11711 3145 11719 3179
rect 11753 3145 11763 3179
rect 11711 3133 11763 3145
rect 11793 3205 11847 3217
rect 11793 3171 11803 3205
rect 11837 3171 11847 3205
rect 11793 3133 11847 3171
rect 11877 3179 11929 3217
rect 11877 3145 11887 3179
rect 11921 3145 11929 3179
rect 11877 3133 11929 3145
rect 11983 3205 12035 3217
rect 11983 3171 11991 3205
rect 12025 3171 12035 3205
rect 11983 3133 12035 3171
rect 12065 3191 12147 3217
rect 12065 3157 12076 3191
rect 12110 3157 12147 3191
rect 12065 3145 12147 3157
rect 12177 3191 12246 3217
rect 12177 3157 12187 3191
rect 12221 3157 12246 3191
rect 12177 3145 12246 3157
rect 12276 3145 12345 3217
rect 12065 3133 12115 3145
rect 12295 3133 12345 3145
rect 12375 3197 12464 3217
rect 12375 3163 12386 3197
rect 12420 3163 12464 3197
rect 12375 3133 12464 3163
rect 12414 3089 12464 3133
rect 12494 3191 12565 3217
rect 12494 3157 12505 3191
rect 12539 3157 12565 3191
rect 12494 3145 12565 3157
rect 12595 3191 12671 3217
rect 12595 3157 12608 3191
rect 12642 3157 12671 3191
rect 12595 3145 12671 3157
rect 12701 3145 12766 3217
rect 12494 3089 12544 3145
rect 12716 3133 12766 3145
rect 12796 3191 12848 3217
rect 12796 3157 12806 3191
rect 12840 3157 12848 3191
rect 12796 3133 12848 3157
rect 12903 3204 12955 3217
rect 12903 3170 12911 3204
rect 12945 3170 12955 3204
rect 12903 3136 12955 3170
rect 12903 3102 12911 3136
rect 12945 3102 12955 3136
rect 12903 3087 12955 3102
rect 12985 3175 13039 3217
rect 12985 3141 12995 3175
rect 13029 3141 13039 3175
rect 12985 3087 13039 3141
rect 13069 3202 13121 3217
rect 13069 3168 13079 3202
rect 13113 3168 13121 3202
rect 13069 3134 13121 3168
rect 13069 3100 13079 3134
rect 13113 3100 13121 3134
rect 13183 3186 13235 3217
rect 13183 3152 13191 3186
rect 13225 3152 13235 3186
rect 13183 3107 13235 3152
rect 14181 3186 14233 3217
rect 14181 3152 14191 3186
rect 14225 3152 14233 3186
rect 14181 3107 14233 3152
rect 14287 3186 14339 3217
rect 14287 3152 14295 3186
rect 14329 3152 14339 3186
rect 14287 3107 14339 3152
rect 15285 3186 15337 3217
rect 15285 3152 15295 3186
rect 15329 3152 15337 3186
rect 15285 3107 15337 3152
rect 15391 3186 15443 3217
rect 15391 3152 15399 3186
rect 15433 3152 15443 3186
rect 15391 3107 15443 3152
rect 16389 3186 16441 3217
rect 16389 3152 16399 3186
rect 16433 3152 16441 3186
rect 16389 3107 16441 3152
rect 13069 3087 13121 3100
rect 16863 3175 16915 3217
rect 16863 3141 16871 3175
rect 16905 3141 16915 3175
rect 16863 3113 16915 3141
rect 16945 3205 17003 3217
rect 16945 3171 16957 3205
rect 16991 3171 17003 3205
rect 16945 3113 17003 3171
rect 17033 3192 17085 3217
rect 17033 3158 17043 3192
rect 17077 3158 17085 3192
rect 17033 3113 17085 3158
rect 17139 3186 17191 3217
rect 17139 3152 17147 3186
rect 17181 3152 17191 3186
rect 17139 3107 17191 3152
rect 18137 3186 18189 3217
rect 18137 3152 18147 3186
rect 18181 3152 18189 3186
rect 18137 3107 18189 3152
rect 18243 3179 18295 3217
rect 18243 3145 18251 3179
rect 18285 3145 18295 3179
rect 18243 3107 18295 3145
rect 18505 3179 18557 3217
rect 18505 3145 18515 3179
rect 18549 3145 18557 3179
rect 18505 3107 18557 3145
rect 18611 3184 18663 3217
rect 18611 3150 18619 3184
rect 18653 3150 18663 3184
rect 18611 3107 18663 3150
rect 18781 3184 18833 3217
rect 18781 3150 18791 3184
rect 18825 3150 18833 3184
rect 18781 3107 18833 3150
rect 2059 2340 2111 2353
rect 1131 2290 1183 2333
rect 1131 2256 1139 2290
rect 1173 2256 1183 2290
rect 1131 2223 1183 2256
rect 1301 2290 1353 2333
rect 1301 2256 1311 2290
rect 1345 2256 1353 2290
rect 1301 2223 1353 2256
rect 1407 2288 1459 2333
rect 1407 2254 1415 2288
rect 1449 2254 1459 2288
rect 1407 2223 1459 2254
rect 1853 2288 1905 2333
rect 1853 2254 1863 2288
rect 1897 2254 1905 2288
rect 1853 2223 1905 2254
rect 2059 2306 2067 2340
rect 2101 2306 2111 2340
rect 2059 2272 2111 2306
rect 2059 2238 2067 2272
rect 2101 2238 2111 2272
rect 2059 2223 2111 2238
rect 2141 2299 2195 2353
rect 2141 2265 2151 2299
rect 2185 2265 2195 2299
rect 2141 2223 2195 2265
rect 2225 2338 2277 2353
rect 2225 2304 2235 2338
rect 2269 2304 2277 2338
rect 2225 2270 2277 2304
rect 2225 2236 2235 2270
rect 2269 2236 2277 2270
rect 2225 2223 2277 2236
rect 2332 2283 2384 2307
rect 2332 2249 2340 2283
rect 2374 2249 2384 2283
rect 2332 2223 2384 2249
rect 2414 2295 2464 2307
rect 2636 2295 2686 2351
rect 2414 2223 2479 2295
rect 2509 2283 2585 2295
rect 2509 2249 2538 2283
rect 2572 2249 2585 2283
rect 2509 2223 2585 2249
rect 2615 2283 2686 2295
rect 2615 2249 2641 2283
rect 2675 2249 2686 2283
rect 2615 2223 2686 2249
rect 2716 2307 2766 2351
rect 2716 2277 2805 2307
rect 2716 2243 2760 2277
rect 2794 2243 2805 2277
rect 2716 2223 2805 2243
rect 2835 2295 2885 2307
rect 3065 2295 3115 2307
rect 2835 2223 2904 2295
rect 2934 2283 3003 2295
rect 2934 2249 2959 2283
rect 2993 2249 3003 2283
rect 2934 2223 3003 2249
rect 3033 2283 3115 2295
rect 3033 2249 3070 2283
rect 3104 2249 3115 2283
rect 3033 2223 3115 2249
rect 3145 2269 3197 2307
rect 3145 2235 3155 2269
rect 3189 2235 3197 2269
rect 3145 2223 3197 2235
rect 3251 2295 3303 2307
rect 3251 2261 3259 2295
rect 3293 2261 3303 2295
rect 3251 2223 3303 2261
rect 3333 2269 3387 2307
rect 3333 2235 3343 2269
rect 3377 2235 3387 2269
rect 3333 2223 3387 2235
rect 3417 2295 3469 2307
rect 3417 2261 3427 2295
rect 3461 2261 3469 2295
rect 3417 2223 3469 2261
rect 4167 2295 4219 2333
rect 4167 2261 4175 2295
rect 4209 2261 4219 2295
rect 4167 2223 4219 2261
rect 4429 2295 4481 2333
rect 4429 2261 4439 2295
rect 4473 2261 4481 2295
rect 4429 2223 4481 2261
rect 4627 2295 4679 2307
rect 4627 2261 4635 2295
rect 4669 2261 4679 2295
rect 4627 2223 4679 2261
rect 4709 2269 4763 2307
rect 4709 2235 4719 2269
rect 4753 2235 4763 2269
rect 4709 2223 4763 2235
rect 4793 2295 4845 2307
rect 4793 2261 4803 2295
rect 4837 2261 4845 2295
rect 4793 2223 4845 2261
rect 4899 2269 4951 2307
rect 4899 2235 4907 2269
rect 4941 2235 4951 2269
rect 4899 2223 4951 2235
rect 4981 2295 5031 2307
rect 5330 2307 5380 2351
rect 5211 2295 5261 2307
rect 4981 2283 5063 2295
rect 4981 2249 4992 2283
rect 5026 2249 5063 2283
rect 4981 2223 5063 2249
rect 5093 2283 5162 2295
rect 5093 2249 5103 2283
rect 5137 2249 5162 2283
rect 5093 2223 5162 2249
rect 5192 2223 5261 2295
rect 5291 2277 5380 2307
rect 5291 2243 5302 2277
rect 5336 2243 5380 2277
rect 5291 2223 5380 2243
rect 5410 2295 5460 2351
rect 5819 2338 5871 2353
rect 5632 2295 5682 2307
rect 5410 2283 5481 2295
rect 5410 2249 5421 2283
rect 5455 2249 5481 2283
rect 5410 2223 5481 2249
rect 5511 2283 5587 2295
rect 5511 2249 5524 2283
rect 5558 2249 5587 2283
rect 5511 2223 5587 2249
rect 5617 2223 5682 2295
rect 5712 2283 5764 2307
rect 5712 2249 5722 2283
rect 5756 2249 5764 2283
rect 5712 2223 5764 2249
rect 5819 2304 5827 2338
rect 5861 2304 5871 2338
rect 5819 2270 5871 2304
rect 5819 2236 5827 2270
rect 5861 2236 5871 2270
rect 5819 2223 5871 2236
rect 5901 2299 5955 2353
rect 5901 2265 5911 2299
rect 5945 2265 5955 2299
rect 5901 2223 5955 2265
rect 5985 2340 6037 2353
rect 5985 2306 5995 2340
rect 6029 2306 6037 2340
rect 5985 2272 6037 2306
rect 5985 2238 5995 2272
rect 6029 2238 6037 2272
rect 7211 2340 7263 2353
rect 6375 2288 6427 2333
rect 6375 2254 6383 2288
rect 6417 2254 6427 2288
rect 5985 2223 6037 2238
rect 6375 2223 6427 2254
rect 7005 2288 7057 2333
rect 7005 2254 7015 2288
rect 7049 2254 7057 2288
rect 7005 2223 7057 2254
rect 7211 2306 7219 2340
rect 7253 2306 7263 2340
rect 7211 2272 7263 2306
rect 7211 2238 7219 2272
rect 7253 2238 7263 2272
rect 7211 2223 7263 2238
rect 7293 2299 7347 2353
rect 7293 2265 7303 2299
rect 7337 2265 7347 2299
rect 7293 2223 7347 2265
rect 7377 2338 7429 2353
rect 7377 2304 7387 2338
rect 7421 2304 7429 2338
rect 7377 2270 7429 2304
rect 7377 2236 7387 2270
rect 7421 2236 7429 2270
rect 7377 2223 7429 2236
rect 7484 2283 7536 2307
rect 7484 2249 7492 2283
rect 7526 2249 7536 2283
rect 7484 2223 7536 2249
rect 7566 2295 7616 2307
rect 7788 2295 7838 2351
rect 7566 2223 7631 2295
rect 7661 2283 7737 2295
rect 7661 2249 7690 2283
rect 7724 2249 7737 2283
rect 7661 2223 7737 2249
rect 7767 2283 7838 2295
rect 7767 2249 7793 2283
rect 7827 2249 7838 2283
rect 7767 2223 7838 2249
rect 7868 2307 7918 2351
rect 7868 2277 7957 2307
rect 7868 2243 7912 2277
rect 7946 2243 7957 2277
rect 7868 2223 7957 2243
rect 7987 2295 8037 2307
rect 8217 2295 8267 2307
rect 7987 2223 8056 2295
rect 8086 2283 8155 2295
rect 8086 2249 8111 2283
rect 8145 2249 8155 2283
rect 8086 2223 8155 2249
rect 8185 2283 8267 2295
rect 8185 2249 8222 2283
rect 8256 2249 8267 2283
rect 8185 2223 8267 2249
rect 8297 2269 8349 2307
rect 8297 2235 8307 2269
rect 8341 2235 8349 2269
rect 8297 2223 8349 2235
rect 8403 2295 8455 2307
rect 8403 2261 8411 2295
rect 8445 2261 8455 2295
rect 8403 2223 8455 2261
rect 8485 2269 8539 2307
rect 8485 2235 8495 2269
rect 8529 2235 8539 2269
rect 8485 2223 8539 2235
rect 8569 2295 8621 2307
rect 8569 2261 8579 2295
rect 8613 2261 8621 2295
rect 8569 2223 8621 2261
rect 8951 2288 9003 2333
rect 8951 2254 8959 2288
rect 8993 2254 9003 2288
rect 8951 2223 9003 2254
rect 9581 2288 9633 2333
rect 9581 2254 9591 2288
rect 9625 2254 9633 2288
rect 9581 2223 9633 2254
rect 9779 2295 9831 2307
rect 9779 2261 9787 2295
rect 9821 2261 9831 2295
rect 9779 2223 9831 2261
rect 9861 2269 9915 2307
rect 9861 2235 9871 2269
rect 9905 2235 9915 2269
rect 9861 2223 9915 2235
rect 9945 2295 9997 2307
rect 9945 2261 9955 2295
rect 9989 2261 9997 2295
rect 9945 2223 9997 2261
rect 10051 2269 10103 2307
rect 10051 2235 10059 2269
rect 10093 2235 10103 2269
rect 10051 2223 10103 2235
rect 10133 2295 10183 2307
rect 10482 2307 10532 2351
rect 10363 2295 10413 2307
rect 10133 2283 10215 2295
rect 10133 2249 10144 2283
rect 10178 2249 10215 2283
rect 10133 2223 10215 2249
rect 10245 2283 10314 2295
rect 10245 2249 10255 2283
rect 10289 2249 10314 2283
rect 10245 2223 10314 2249
rect 10344 2223 10413 2295
rect 10443 2277 10532 2307
rect 10443 2243 10454 2277
rect 10488 2243 10532 2277
rect 10443 2223 10532 2243
rect 10562 2295 10612 2351
rect 10971 2338 11023 2353
rect 10784 2295 10834 2307
rect 10562 2283 10633 2295
rect 10562 2249 10573 2283
rect 10607 2249 10633 2283
rect 10562 2223 10633 2249
rect 10663 2283 10739 2295
rect 10663 2249 10676 2283
rect 10710 2249 10739 2283
rect 10663 2223 10739 2249
rect 10769 2223 10834 2295
rect 10864 2283 10916 2307
rect 10864 2249 10874 2283
rect 10908 2249 10916 2283
rect 10864 2223 10916 2249
rect 10971 2304 10979 2338
rect 11013 2304 11023 2338
rect 10971 2270 11023 2304
rect 10971 2236 10979 2270
rect 11013 2236 11023 2270
rect 10971 2223 11023 2236
rect 11053 2299 11107 2353
rect 11053 2265 11063 2299
rect 11097 2265 11107 2299
rect 11053 2223 11107 2265
rect 11137 2340 11189 2353
rect 11137 2306 11147 2340
rect 11181 2306 11189 2340
rect 11137 2272 11189 2306
rect 11137 2238 11147 2272
rect 11181 2238 11189 2272
rect 11903 2340 11955 2353
rect 11527 2295 11579 2333
rect 11527 2261 11535 2295
rect 11569 2261 11579 2295
rect 11137 2223 11189 2238
rect 11527 2223 11579 2261
rect 11789 2295 11841 2333
rect 11789 2261 11799 2295
rect 11833 2261 11841 2295
rect 11789 2223 11841 2261
rect 11903 2306 11911 2340
rect 11945 2306 11955 2340
rect 11903 2272 11955 2306
rect 11903 2238 11911 2272
rect 11945 2238 11955 2272
rect 11903 2223 11955 2238
rect 11985 2299 12039 2353
rect 11985 2265 11995 2299
rect 12029 2265 12039 2299
rect 11985 2223 12039 2265
rect 12069 2338 12121 2353
rect 12069 2304 12079 2338
rect 12113 2304 12121 2338
rect 12069 2270 12121 2304
rect 12069 2236 12079 2270
rect 12113 2236 12121 2270
rect 12069 2223 12121 2236
rect 12176 2283 12228 2307
rect 12176 2249 12184 2283
rect 12218 2249 12228 2283
rect 12176 2223 12228 2249
rect 12258 2295 12308 2307
rect 12480 2295 12530 2351
rect 12258 2223 12323 2295
rect 12353 2283 12429 2295
rect 12353 2249 12382 2283
rect 12416 2249 12429 2283
rect 12353 2223 12429 2249
rect 12459 2283 12530 2295
rect 12459 2249 12485 2283
rect 12519 2249 12530 2283
rect 12459 2223 12530 2249
rect 12560 2307 12610 2351
rect 12560 2277 12649 2307
rect 12560 2243 12604 2277
rect 12638 2243 12649 2277
rect 12560 2223 12649 2243
rect 12679 2295 12729 2307
rect 12909 2295 12959 2307
rect 12679 2223 12748 2295
rect 12778 2283 12847 2295
rect 12778 2249 12803 2283
rect 12837 2249 12847 2283
rect 12778 2223 12847 2249
rect 12877 2283 12959 2295
rect 12877 2249 12914 2283
rect 12948 2249 12959 2283
rect 12877 2223 12959 2249
rect 12989 2269 13041 2307
rect 12989 2235 12999 2269
rect 13033 2235 13041 2269
rect 12989 2223 13041 2235
rect 13095 2295 13147 2307
rect 13095 2261 13103 2295
rect 13137 2261 13147 2295
rect 13095 2223 13147 2261
rect 13177 2269 13231 2307
rect 13177 2235 13187 2269
rect 13221 2235 13231 2269
rect 13177 2223 13231 2235
rect 13261 2295 13313 2307
rect 13261 2261 13271 2295
rect 13305 2261 13313 2295
rect 13261 2223 13313 2261
rect 13367 2288 13419 2333
rect 13367 2254 13375 2288
rect 13409 2254 13419 2288
rect 13367 2223 13419 2254
rect 13813 2288 13865 2333
rect 13813 2254 13823 2288
rect 13857 2254 13865 2288
rect 13813 2223 13865 2254
rect 14563 2288 14615 2333
rect 14563 2254 14571 2288
rect 14605 2254 14615 2288
rect 14563 2223 14615 2254
rect 15561 2288 15613 2333
rect 15561 2254 15571 2288
rect 15605 2254 15613 2288
rect 15561 2223 15613 2254
rect 15667 2288 15719 2333
rect 15667 2254 15675 2288
rect 15709 2254 15719 2288
rect 15667 2223 15719 2254
rect 16297 2288 16349 2333
rect 16297 2254 16307 2288
rect 16341 2254 16349 2288
rect 16297 2223 16349 2254
rect 16863 2299 16915 2327
rect 16863 2265 16871 2299
rect 16905 2265 16915 2299
rect 16863 2223 16915 2265
rect 16945 2269 17003 2327
rect 16945 2235 16957 2269
rect 16991 2235 17003 2269
rect 16945 2223 17003 2235
rect 17033 2282 17085 2327
rect 17033 2248 17043 2282
rect 17077 2248 17085 2282
rect 17033 2223 17085 2248
rect 17139 2295 17191 2333
rect 17139 2261 17147 2295
rect 17181 2261 17191 2295
rect 17139 2223 17191 2261
rect 17401 2295 17453 2333
rect 17604 2307 17654 2353
rect 17401 2261 17411 2295
rect 17445 2261 17453 2295
rect 17401 2223 17453 2261
rect 17507 2282 17559 2307
rect 17507 2248 17515 2282
rect 17549 2248 17559 2282
rect 17507 2223 17559 2248
rect 17589 2269 17654 2307
rect 17589 2235 17608 2269
rect 17642 2235 17654 2269
rect 17589 2223 17654 2235
rect 17684 2299 17738 2353
rect 17684 2265 17694 2299
rect 17728 2265 17738 2299
rect 17684 2223 17738 2265
rect 17768 2341 17821 2353
rect 17768 2307 17778 2341
rect 17812 2307 17821 2341
rect 17768 2273 17821 2307
rect 17768 2239 17778 2273
rect 17812 2239 17821 2273
rect 17768 2223 17821 2239
rect 17875 2288 17927 2333
rect 17875 2254 17883 2288
rect 17917 2254 17927 2288
rect 17875 2223 17927 2254
rect 18505 2288 18557 2333
rect 18505 2254 18515 2288
rect 18549 2254 18557 2288
rect 18505 2223 18557 2254
rect 18611 2290 18663 2333
rect 18611 2256 18619 2290
rect 18653 2256 18663 2290
rect 18611 2223 18663 2256
rect 18781 2290 18833 2333
rect 18781 2256 18791 2290
rect 18825 2256 18833 2290
rect 18781 2223 18833 2256
<< pdiff >>
rect 1591 7301 1644 7319
rect 1131 7260 1183 7293
rect 1131 7226 1139 7260
rect 1173 7226 1183 7260
rect 1131 7165 1183 7226
rect 1131 7131 1139 7165
rect 1173 7131 1183 7165
rect 1131 7119 1183 7131
rect 1301 7260 1353 7293
rect 1301 7226 1311 7260
rect 1345 7226 1353 7260
rect 1301 7165 1353 7226
rect 1301 7131 1311 7165
rect 1345 7131 1353 7165
rect 1301 7119 1353 7131
rect 1591 7267 1600 7301
rect 1634 7267 1644 7301
rect 1591 7233 1644 7267
rect 1591 7199 1600 7233
rect 1634 7199 1644 7233
rect 1591 7165 1644 7199
rect 1591 7131 1600 7165
rect 1634 7131 1644 7165
rect 1591 7119 1644 7131
rect 1674 7270 1728 7319
rect 1674 7236 1684 7270
rect 1718 7236 1728 7270
rect 1674 7189 1728 7236
rect 1674 7155 1684 7189
rect 1718 7155 1728 7189
rect 1674 7119 1728 7155
rect 1758 7255 1808 7319
rect 1758 7241 1823 7255
rect 1758 7207 1770 7241
rect 1804 7207 1823 7241
rect 1758 7173 1823 7207
rect 1758 7139 1770 7173
rect 1804 7139 1823 7173
rect 1758 7127 1823 7139
rect 1853 7241 1905 7255
rect 1853 7207 1863 7241
rect 1897 7207 1905 7241
rect 1853 7173 1905 7207
rect 1853 7139 1863 7173
rect 1897 7139 1905 7173
rect 1853 7127 1905 7139
rect 1959 7165 2011 7293
rect 1959 7131 1967 7165
rect 2001 7131 2011 7165
rect 1758 7119 1808 7127
rect 1959 7119 2011 7131
rect 2957 7165 3009 7293
rect 2957 7131 2967 7165
rect 3001 7131 3009 7165
rect 2957 7119 3009 7131
rect 3063 7267 3115 7293
rect 3063 7233 3071 7267
rect 3105 7233 3115 7267
rect 3063 7165 3115 7233
rect 3063 7131 3071 7165
rect 3105 7131 3115 7165
rect 3063 7119 3115 7131
rect 3509 7267 3561 7293
rect 3509 7233 3519 7267
rect 3553 7233 3561 7267
rect 3509 7165 3561 7233
rect 3509 7131 3519 7165
rect 3553 7131 3561 7165
rect 3983 7301 4036 7319
rect 3983 7267 3992 7301
rect 4026 7267 4036 7301
rect 3983 7233 4036 7267
rect 3983 7199 3992 7233
rect 4026 7199 4036 7233
rect 3983 7165 4036 7199
rect 3509 7119 3561 7131
rect 3983 7131 3992 7165
rect 4026 7131 4036 7165
rect 3983 7119 4036 7131
rect 4066 7270 4120 7319
rect 4066 7236 4076 7270
rect 4110 7236 4120 7270
rect 4066 7189 4120 7236
rect 4066 7155 4076 7189
rect 4110 7155 4120 7189
rect 4066 7119 4120 7155
rect 4150 7255 4200 7319
rect 5639 7301 5692 7319
rect 4150 7241 4215 7255
rect 4150 7207 4162 7241
rect 4196 7207 4215 7241
rect 4150 7173 4215 7207
rect 4150 7139 4162 7173
rect 4196 7139 4215 7173
rect 4150 7127 4215 7139
rect 4245 7241 4297 7255
rect 4245 7207 4255 7241
rect 4289 7207 4297 7241
rect 4245 7173 4297 7207
rect 4245 7139 4255 7173
rect 4289 7139 4297 7173
rect 4245 7127 4297 7139
rect 4351 7165 4403 7293
rect 4351 7131 4359 7165
rect 4393 7131 4403 7165
rect 4150 7119 4200 7127
rect 4351 7119 4403 7131
rect 5349 7165 5401 7293
rect 5349 7131 5359 7165
rect 5393 7131 5401 7165
rect 5349 7119 5401 7131
rect 5639 7267 5648 7301
rect 5682 7267 5692 7301
rect 5639 7233 5692 7267
rect 5639 7199 5648 7233
rect 5682 7199 5692 7233
rect 5639 7165 5692 7199
rect 5639 7131 5648 7165
rect 5682 7131 5692 7165
rect 5639 7119 5692 7131
rect 5722 7270 5776 7319
rect 5722 7236 5732 7270
rect 5766 7236 5776 7270
rect 5722 7189 5776 7236
rect 5722 7155 5732 7189
rect 5766 7155 5776 7189
rect 5722 7119 5776 7155
rect 5806 7255 5856 7319
rect 6007 7260 6059 7293
rect 5806 7241 5871 7255
rect 5806 7207 5818 7241
rect 5852 7207 5871 7241
rect 5806 7173 5871 7207
rect 5806 7139 5818 7173
rect 5852 7139 5871 7173
rect 5806 7127 5871 7139
rect 5901 7241 5953 7255
rect 5901 7207 5911 7241
rect 5945 7207 5953 7241
rect 5901 7173 5953 7207
rect 5901 7139 5911 7173
rect 5945 7139 5953 7173
rect 5901 7127 5953 7139
rect 6007 7226 6015 7260
rect 6049 7226 6059 7260
rect 6007 7165 6059 7226
rect 6007 7131 6015 7165
rect 6049 7131 6059 7165
rect 5806 7119 5856 7127
rect 6007 7119 6059 7131
rect 6177 7260 6229 7293
rect 6177 7226 6187 7260
rect 6221 7226 6229 7260
rect 6177 7165 6229 7226
rect 6177 7131 6187 7165
rect 6221 7131 6229 7165
rect 6375 7165 6427 7293
rect 6177 7119 6229 7131
rect 6375 7131 6383 7165
rect 6417 7131 6427 7165
rect 6375 7119 6427 7131
rect 7373 7165 7425 7293
rect 7373 7131 7383 7165
rect 7417 7131 7425 7165
rect 7373 7119 7425 7131
rect 7479 7267 7531 7293
rect 7479 7233 7487 7267
rect 7521 7233 7531 7267
rect 7479 7165 7531 7233
rect 7479 7131 7487 7165
rect 7521 7131 7531 7165
rect 7479 7119 7531 7131
rect 7741 7267 7793 7293
rect 7741 7233 7751 7267
rect 7785 7233 7793 7267
rect 7944 7255 7994 7319
rect 7741 7165 7793 7233
rect 7741 7131 7751 7165
rect 7785 7131 7793 7165
rect 7741 7119 7793 7131
rect 7847 7241 7899 7255
rect 7847 7207 7855 7241
rect 7889 7207 7899 7241
rect 7847 7173 7899 7207
rect 7847 7139 7855 7173
rect 7889 7139 7899 7173
rect 7847 7127 7899 7139
rect 7929 7241 7994 7255
rect 7929 7207 7948 7241
rect 7982 7207 7994 7241
rect 7929 7173 7994 7207
rect 7929 7139 7948 7173
rect 7982 7139 7994 7173
rect 7929 7127 7994 7139
rect 7944 7119 7994 7127
rect 8024 7270 8078 7319
rect 8024 7236 8034 7270
rect 8068 7236 8078 7270
rect 8024 7189 8078 7236
rect 8024 7155 8034 7189
rect 8068 7155 8078 7189
rect 8024 7119 8078 7155
rect 8108 7301 8161 7319
rect 8108 7267 8118 7301
rect 8152 7267 8161 7301
rect 8108 7233 8161 7267
rect 8108 7199 8118 7233
rect 8152 7199 8161 7233
rect 8108 7165 8161 7199
rect 8108 7131 8118 7165
rect 8152 7131 8161 7165
rect 8108 7119 8161 7131
rect 8215 7267 8267 7293
rect 8215 7233 8223 7267
rect 8257 7233 8267 7267
rect 8215 7165 8267 7233
rect 8215 7131 8223 7165
rect 8257 7131 8267 7165
rect 8215 7119 8267 7131
rect 8661 7267 8713 7293
rect 8661 7233 8671 7267
rect 8705 7233 8713 7267
rect 8661 7165 8713 7233
rect 8661 7131 8671 7165
rect 8705 7131 8713 7165
rect 8951 7267 9003 7293
rect 8951 7233 8959 7267
rect 8993 7233 9003 7267
rect 8951 7165 9003 7233
rect 8661 7119 8713 7131
rect 8951 7131 8959 7165
rect 8993 7131 9003 7165
rect 8951 7119 9003 7131
rect 9397 7267 9449 7293
rect 9397 7233 9407 7267
rect 9441 7233 9449 7267
rect 9397 7165 9449 7233
rect 9397 7131 9407 7165
rect 9441 7131 9449 7165
rect 9397 7119 9449 7131
rect 9687 7267 9739 7293
rect 9687 7233 9695 7267
rect 9729 7233 9739 7267
rect 9687 7165 9739 7233
rect 9687 7131 9695 7165
rect 9729 7131 9739 7165
rect 9687 7119 9739 7131
rect 9949 7267 10001 7293
rect 9949 7233 9959 7267
rect 9993 7233 10001 7267
rect 9949 7165 10001 7233
rect 9949 7131 9959 7165
rect 9993 7131 10001 7165
rect 9949 7119 10001 7131
rect 10055 7284 10108 7319
rect 10055 7250 10063 7284
rect 10097 7250 10108 7284
rect 10055 7179 10108 7250
rect 10055 7145 10063 7179
rect 10097 7145 10108 7179
rect 10055 7119 10108 7145
rect 10138 7245 10203 7319
rect 10138 7211 10149 7245
rect 10183 7211 10203 7245
rect 10138 7177 10203 7211
rect 10138 7143 10149 7177
rect 10183 7143 10203 7177
rect 10138 7119 10203 7143
rect 10233 7179 10287 7319
rect 10233 7145 10243 7179
rect 10277 7145 10287 7179
rect 10233 7119 10287 7145
rect 10317 7174 10369 7319
rect 10317 7140 10327 7174
rect 10361 7140 10369 7174
rect 10317 7119 10369 7140
rect 10423 7267 10475 7293
rect 10423 7233 10431 7267
rect 10465 7233 10475 7267
rect 10423 7165 10475 7233
rect 10423 7131 10431 7165
rect 10465 7131 10475 7165
rect 10423 7119 10475 7131
rect 11053 7267 11105 7293
rect 11053 7233 11063 7267
rect 11097 7233 11105 7267
rect 11053 7165 11105 7233
rect 11053 7131 11063 7165
rect 11097 7131 11105 7165
rect 11053 7119 11105 7131
rect 11159 7260 11211 7293
rect 11159 7226 11167 7260
rect 11201 7226 11211 7260
rect 11159 7165 11211 7226
rect 11159 7131 11167 7165
rect 11201 7131 11211 7165
rect 11159 7119 11211 7131
rect 11329 7260 11381 7293
rect 11329 7226 11339 7260
rect 11373 7226 11381 7260
rect 11329 7165 11381 7226
rect 11329 7131 11339 7165
rect 11373 7131 11381 7165
rect 11527 7267 11579 7293
rect 11527 7233 11535 7267
rect 11569 7233 11579 7267
rect 11527 7165 11579 7233
rect 11329 7119 11381 7131
rect 11527 7131 11535 7165
rect 11569 7131 11579 7165
rect 11527 7119 11579 7131
rect 12157 7267 12209 7293
rect 12157 7233 12167 7267
rect 12201 7233 12209 7267
rect 12360 7255 12410 7319
rect 12157 7165 12209 7233
rect 12157 7131 12167 7165
rect 12201 7131 12209 7165
rect 12157 7119 12209 7131
rect 12263 7241 12315 7255
rect 12263 7207 12271 7241
rect 12305 7207 12315 7241
rect 12263 7173 12315 7207
rect 12263 7139 12271 7173
rect 12305 7139 12315 7173
rect 12263 7127 12315 7139
rect 12345 7241 12410 7255
rect 12345 7207 12364 7241
rect 12398 7207 12410 7241
rect 12345 7173 12410 7207
rect 12345 7139 12364 7173
rect 12398 7139 12410 7173
rect 12345 7127 12410 7139
rect 12360 7119 12410 7127
rect 12440 7270 12494 7319
rect 12440 7236 12450 7270
rect 12484 7236 12494 7270
rect 12440 7189 12494 7236
rect 12440 7155 12450 7189
rect 12484 7155 12494 7189
rect 12440 7119 12494 7155
rect 12524 7301 12577 7319
rect 12524 7267 12534 7301
rect 12568 7267 12577 7301
rect 12524 7233 12577 7267
rect 12524 7199 12534 7233
rect 12568 7199 12577 7233
rect 12524 7165 12577 7199
rect 12524 7131 12534 7165
rect 12568 7131 12577 7165
rect 12524 7119 12577 7131
rect 12631 7165 12683 7293
rect 12631 7131 12639 7165
rect 12673 7131 12683 7165
rect 12631 7119 12683 7131
rect 13629 7165 13681 7293
rect 13629 7131 13639 7165
rect 13673 7131 13681 7165
rect 13629 7119 13681 7131
rect 13735 7260 13787 7293
rect 13735 7226 13743 7260
rect 13777 7226 13787 7260
rect 13735 7165 13787 7226
rect 13735 7131 13743 7165
rect 13777 7131 13787 7165
rect 13735 7119 13787 7131
rect 13905 7260 13957 7293
rect 13905 7226 13915 7260
rect 13949 7226 13957 7260
rect 13905 7165 13957 7226
rect 13905 7131 13915 7165
rect 13949 7131 13957 7165
rect 14103 7267 14155 7293
rect 14103 7233 14111 7267
rect 14145 7233 14155 7267
rect 14103 7165 14155 7233
rect 13905 7119 13957 7131
rect 14103 7131 14111 7165
rect 14145 7131 14155 7165
rect 14103 7119 14155 7131
rect 14365 7267 14417 7293
rect 14365 7233 14375 7267
rect 14409 7233 14417 7267
rect 14568 7255 14618 7319
rect 14365 7165 14417 7233
rect 14365 7131 14375 7165
rect 14409 7131 14417 7165
rect 14365 7119 14417 7131
rect 14471 7241 14523 7255
rect 14471 7207 14479 7241
rect 14513 7207 14523 7241
rect 14471 7173 14523 7207
rect 14471 7139 14479 7173
rect 14513 7139 14523 7173
rect 14471 7127 14523 7139
rect 14553 7241 14618 7255
rect 14553 7207 14572 7241
rect 14606 7207 14618 7241
rect 14553 7173 14618 7207
rect 14553 7139 14572 7173
rect 14606 7139 14618 7173
rect 14553 7127 14618 7139
rect 14568 7119 14618 7127
rect 14648 7270 14702 7319
rect 14648 7236 14658 7270
rect 14692 7236 14702 7270
rect 14648 7189 14702 7236
rect 14648 7155 14658 7189
rect 14692 7155 14702 7189
rect 14648 7119 14702 7155
rect 14732 7301 14785 7319
rect 14732 7267 14742 7301
rect 14776 7267 14785 7301
rect 14732 7233 14785 7267
rect 14732 7199 14742 7233
rect 14776 7199 14785 7233
rect 14732 7165 14785 7199
rect 14732 7131 14742 7165
rect 14776 7131 14785 7165
rect 14732 7119 14785 7131
rect 14839 7165 14891 7293
rect 14839 7131 14847 7165
rect 14881 7131 14891 7165
rect 14839 7119 14891 7131
rect 15837 7165 15889 7293
rect 15837 7131 15847 7165
rect 15881 7131 15889 7165
rect 15837 7119 15889 7131
rect 15943 7267 15995 7293
rect 15943 7233 15951 7267
rect 15985 7233 15995 7267
rect 15943 7165 15995 7233
rect 15943 7131 15951 7165
rect 15985 7131 15995 7165
rect 15943 7119 15995 7131
rect 16389 7267 16441 7293
rect 16389 7233 16399 7267
rect 16433 7233 16441 7267
rect 16389 7165 16441 7233
rect 16389 7131 16399 7165
rect 16433 7131 16441 7165
rect 16960 7255 17010 7319
rect 16863 7241 16915 7255
rect 16863 7207 16871 7241
rect 16905 7207 16915 7241
rect 16863 7173 16915 7207
rect 16863 7139 16871 7173
rect 16905 7139 16915 7173
rect 16389 7119 16441 7131
rect 16863 7127 16915 7139
rect 16945 7241 17010 7255
rect 16945 7207 16964 7241
rect 16998 7207 17010 7241
rect 16945 7173 17010 7207
rect 16945 7139 16964 7173
rect 16998 7139 17010 7173
rect 16945 7127 17010 7139
rect 16960 7119 17010 7127
rect 17040 7270 17094 7319
rect 17040 7236 17050 7270
rect 17084 7236 17094 7270
rect 17040 7189 17094 7236
rect 17040 7155 17050 7189
rect 17084 7155 17094 7189
rect 17040 7119 17094 7155
rect 17124 7301 17177 7319
rect 17124 7267 17134 7301
rect 17168 7267 17177 7301
rect 17124 7233 17177 7267
rect 17124 7199 17134 7233
rect 17168 7199 17177 7233
rect 17124 7165 17177 7199
rect 17124 7131 17134 7165
rect 17168 7131 17177 7165
rect 17124 7119 17177 7131
rect 17231 7267 17283 7293
rect 17231 7233 17239 7267
rect 17273 7233 17283 7267
rect 17231 7165 17283 7233
rect 17231 7131 17239 7165
rect 17273 7131 17283 7165
rect 17231 7119 17283 7131
rect 17861 7267 17913 7293
rect 17861 7233 17871 7267
rect 17905 7233 17913 7267
rect 18156 7255 18206 7319
rect 17861 7165 17913 7233
rect 17861 7131 17871 7165
rect 17905 7131 17913 7165
rect 17861 7119 17913 7131
rect 18059 7241 18111 7255
rect 18059 7207 18067 7241
rect 18101 7207 18111 7241
rect 18059 7173 18111 7207
rect 18059 7139 18067 7173
rect 18101 7139 18111 7173
rect 18059 7127 18111 7139
rect 18141 7241 18206 7255
rect 18141 7207 18160 7241
rect 18194 7207 18206 7241
rect 18141 7173 18206 7207
rect 18141 7139 18160 7173
rect 18194 7139 18206 7173
rect 18141 7127 18206 7139
rect 18156 7119 18206 7127
rect 18236 7270 18290 7319
rect 18236 7236 18246 7270
rect 18280 7236 18290 7270
rect 18236 7189 18290 7236
rect 18236 7155 18246 7189
rect 18280 7155 18290 7189
rect 18236 7119 18290 7155
rect 18320 7301 18373 7319
rect 18320 7267 18330 7301
rect 18364 7267 18373 7301
rect 18320 7233 18373 7267
rect 18320 7199 18330 7233
rect 18364 7199 18373 7233
rect 18320 7165 18373 7199
rect 18320 7131 18330 7165
rect 18364 7131 18373 7165
rect 18320 7119 18373 7131
rect 18611 7260 18663 7293
rect 18611 7226 18619 7260
rect 18653 7226 18663 7260
rect 18611 7165 18663 7226
rect 18611 7131 18619 7165
rect 18653 7131 18663 7165
rect 18611 7119 18663 7131
rect 18781 7260 18833 7293
rect 18781 7226 18791 7260
rect 18825 7226 18833 7260
rect 18781 7165 18833 7226
rect 18781 7131 18791 7165
rect 18825 7131 18833 7165
rect 18781 7119 18833 7131
rect 1131 7013 1183 7025
rect 1131 6979 1139 7013
rect 1173 6979 1183 7013
rect 1131 6918 1183 6979
rect 1131 6884 1139 6918
rect 1173 6884 1183 6918
rect 1131 6851 1183 6884
rect 1301 7013 1353 7025
rect 1301 6979 1311 7013
rect 1345 6979 1353 7013
rect 1301 6918 1353 6979
rect 1301 6884 1311 6918
rect 1345 6884 1353 6918
rect 1301 6851 1353 6884
rect 1407 7013 1459 7025
rect 1407 6979 1415 7013
rect 1449 6979 1459 7013
rect 1407 6851 1459 6979
rect 2405 7013 2457 7025
rect 2405 6979 2415 7013
rect 2449 6979 2457 7013
rect 2405 6851 2457 6979
rect 2511 7013 2563 7025
rect 2511 6979 2519 7013
rect 2553 6979 2563 7013
rect 2511 6851 2563 6979
rect 3509 7013 3561 7025
rect 3509 6979 3519 7013
rect 3553 6979 3561 7013
rect 3799 7013 3851 7025
rect 3509 6851 3561 6979
rect 3799 6979 3807 7013
rect 3841 6979 3851 7013
rect 3799 6851 3851 6979
rect 4797 7013 4849 7025
rect 4797 6979 4807 7013
rect 4841 6979 4849 7013
rect 4797 6851 4849 6979
rect 4903 7013 4955 7025
rect 4903 6979 4911 7013
rect 4945 6979 4955 7013
rect 4903 6851 4955 6979
rect 5901 7013 5953 7025
rect 5901 6979 5911 7013
rect 5945 6979 5953 7013
rect 5901 6851 5953 6979
rect 6007 7013 6059 7025
rect 6007 6979 6015 7013
rect 6049 6979 6059 7013
rect 6007 6851 6059 6979
rect 7005 7013 7057 7025
rect 7005 6979 7015 7013
rect 7049 6979 7057 7013
rect 7005 6851 7057 6979
rect 7111 7013 7163 7025
rect 7111 6979 7119 7013
rect 7153 6979 7163 7013
rect 7111 6851 7163 6979
rect 8109 7013 8161 7025
rect 8109 6979 8119 7013
rect 8153 6979 8161 7013
rect 8109 6851 8161 6979
rect 8215 7013 8267 7025
rect 8215 6979 8223 7013
rect 8257 6979 8267 7013
rect 8215 6911 8267 6979
rect 8215 6877 8223 6911
rect 8257 6877 8267 6911
rect 8215 6851 8267 6877
rect 8661 7013 8713 7025
rect 8661 6979 8671 7013
rect 8705 6979 8713 7013
rect 8951 7013 9003 7025
rect 8661 6911 8713 6979
rect 8661 6877 8671 6911
rect 8705 6877 8713 6911
rect 8661 6851 8713 6877
rect 8951 6979 8959 7013
rect 8993 6979 9003 7013
rect 8951 6851 9003 6979
rect 9949 7013 10001 7025
rect 9949 6979 9959 7013
rect 9993 6979 10001 7013
rect 9949 6851 10001 6979
rect 10055 7013 10107 7025
rect 10055 6979 10063 7013
rect 10097 6979 10107 7013
rect 10055 6851 10107 6979
rect 11053 7013 11105 7025
rect 11053 6979 11063 7013
rect 11097 6979 11105 7013
rect 11053 6851 11105 6979
rect 11159 7013 11211 7025
rect 11159 6979 11167 7013
rect 11201 6979 11211 7013
rect 11159 6851 11211 6979
rect 12157 7013 12209 7025
rect 12157 6979 12167 7013
rect 12201 6979 12209 7013
rect 12157 6851 12209 6979
rect 12263 7013 12315 7025
rect 12263 6979 12271 7013
rect 12305 6979 12315 7013
rect 12263 6851 12315 6979
rect 13261 7013 13313 7025
rect 13261 6979 13271 7013
rect 13305 6979 13313 7013
rect 13261 6851 13313 6979
rect 13367 7013 13419 7025
rect 13367 6979 13375 7013
rect 13409 6979 13419 7013
rect 13367 6911 13419 6979
rect 13367 6877 13375 6911
rect 13409 6877 13419 6911
rect 13367 6851 13419 6877
rect 13813 7013 13865 7025
rect 13813 6979 13823 7013
rect 13857 6979 13865 7013
rect 14103 7013 14155 7025
rect 13813 6911 13865 6979
rect 13813 6877 13823 6911
rect 13857 6877 13865 6911
rect 13813 6851 13865 6877
rect 14103 6979 14111 7013
rect 14145 6979 14155 7013
rect 14103 6851 14155 6979
rect 15101 7013 15153 7025
rect 15101 6979 15111 7013
rect 15145 6979 15153 7013
rect 15101 6851 15153 6979
rect 15207 7013 15259 7025
rect 15207 6979 15215 7013
rect 15249 6979 15259 7013
rect 15207 6851 15259 6979
rect 16205 7013 16257 7025
rect 16205 6979 16215 7013
rect 16249 6979 16257 7013
rect 16205 6851 16257 6979
rect 16311 7013 16363 7025
rect 16311 6979 16319 7013
rect 16353 6979 16363 7013
rect 16311 6851 16363 6979
rect 17309 7013 17361 7025
rect 17309 6979 17319 7013
rect 17353 6979 17361 7013
rect 17309 6851 17361 6979
rect 17415 7013 17467 7025
rect 17415 6979 17423 7013
rect 17457 6979 17467 7013
rect 17415 6851 17467 6979
rect 18413 7013 18465 7025
rect 18413 6979 18423 7013
rect 18457 6979 18465 7013
rect 18413 6851 18465 6979
rect 18611 7013 18663 7025
rect 18611 6979 18619 7013
rect 18653 6979 18663 7013
rect 18611 6918 18663 6979
rect 18611 6884 18619 6918
rect 18653 6884 18663 6918
rect 18611 6851 18663 6884
rect 18781 7013 18833 7025
rect 18781 6979 18791 7013
rect 18825 6979 18833 7013
rect 18781 6918 18833 6979
rect 18781 6884 18791 6918
rect 18825 6884 18833 6918
rect 18781 6851 18833 6884
rect 1131 6172 1183 6205
rect 1131 6138 1139 6172
rect 1173 6138 1183 6172
rect 1131 6077 1183 6138
rect 1131 6043 1139 6077
rect 1173 6043 1183 6077
rect 1131 6031 1183 6043
rect 1301 6172 1353 6205
rect 1301 6138 1311 6172
rect 1345 6138 1353 6172
rect 1301 6077 1353 6138
rect 1301 6043 1311 6077
rect 1345 6043 1353 6077
rect 1301 6031 1353 6043
rect 1407 6077 1459 6205
rect 1407 6043 1415 6077
rect 1449 6043 1459 6077
rect 1407 6031 1459 6043
rect 2405 6077 2457 6205
rect 2405 6043 2415 6077
rect 2449 6043 2457 6077
rect 2405 6031 2457 6043
rect 2511 6077 2563 6205
rect 2511 6043 2519 6077
rect 2553 6043 2563 6077
rect 2511 6031 2563 6043
rect 3509 6077 3561 6205
rect 3509 6043 3519 6077
rect 3553 6043 3561 6077
rect 3509 6031 3561 6043
rect 3615 6077 3667 6205
rect 3615 6043 3623 6077
rect 3657 6043 3667 6077
rect 3615 6031 3667 6043
rect 4613 6077 4665 6205
rect 4613 6043 4623 6077
rect 4657 6043 4665 6077
rect 4613 6031 4665 6043
rect 4719 6077 4771 6205
rect 4719 6043 4727 6077
rect 4761 6043 4771 6077
rect 4719 6031 4771 6043
rect 5717 6077 5769 6205
rect 5717 6043 5727 6077
rect 5761 6043 5769 6077
rect 5717 6031 5769 6043
rect 5823 6179 5875 6205
rect 5823 6145 5831 6179
rect 5865 6145 5875 6179
rect 5823 6077 5875 6145
rect 5823 6043 5831 6077
rect 5865 6043 5875 6077
rect 5823 6031 5875 6043
rect 6085 6179 6137 6205
rect 6085 6145 6095 6179
rect 6129 6145 6137 6179
rect 6085 6077 6137 6145
rect 6085 6043 6095 6077
rect 6129 6043 6137 6077
rect 6375 6077 6427 6205
rect 6085 6031 6137 6043
rect 6375 6043 6383 6077
rect 6417 6043 6427 6077
rect 6375 6031 6427 6043
rect 7373 6077 7425 6205
rect 7373 6043 7383 6077
rect 7417 6043 7425 6077
rect 7373 6031 7425 6043
rect 7479 6077 7531 6205
rect 7479 6043 7487 6077
rect 7521 6043 7531 6077
rect 7479 6031 7531 6043
rect 8477 6077 8529 6205
rect 8477 6043 8487 6077
rect 8521 6043 8529 6077
rect 8477 6031 8529 6043
rect 8583 6077 8635 6205
rect 8583 6043 8591 6077
rect 8625 6043 8635 6077
rect 8583 6031 8635 6043
rect 9581 6077 9633 6205
rect 9581 6043 9591 6077
rect 9625 6043 9633 6077
rect 9581 6031 9633 6043
rect 9687 6077 9739 6205
rect 9687 6043 9695 6077
rect 9729 6043 9739 6077
rect 9687 6031 9739 6043
rect 10685 6077 10737 6205
rect 10685 6043 10695 6077
rect 10729 6043 10737 6077
rect 10685 6031 10737 6043
rect 10791 6179 10843 6205
rect 10791 6145 10799 6179
rect 10833 6145 10843 6179
rect 10791 6077 10843 6145
rect 10791 6043 10799 6077
rect 10833 6043 10843 6077
rect 10791 6031 10843 6043
rect 11237 6179 11289 6205
rect 11237 6145 11247 6179
rect 11281 6145 11289 6179
rect 11237 6077 11289 6145
rect 11237 6043 11247 6077
rect 11281 6043 11289 6077
rect 11527 6077 11579 6205
rect 11237 6031 11289 6043
rect 11527 6043 11535 6077
rect 11569 6043 11579 6077
rect 11527 6031 11579 6043
rect 12525 6077 12577 6205
rect 12525 6043 12535 6077
rect 12569 6043 12577 6077
rect 12525 6031 12577 6043
rect 12631 6077 12683 6205
rect 12631 6043 12639 6077
rect 12673 6043 12683 6077
rect 12631 6031 12683 6043
rect 13629 6077 13681 6205
rect 13629 6043 13639 6077
rect 13673 6043 13681 6077
rect 13629 6031 13681 6043
rect 13735 6077 13787 6205
rect 13735 6043 13743 6077
rect 13777 6043 13787 6077
rect 13735 6031 13787 6043
rect 14733 6077 14785 6205
rect 14733 6043 14743 6077
rect 14777 6043 14785 6077
rect 14733 6031 14785 6043
rect 14839 6077 14891 6205
rect 14839 6043 14847 6077
rect 14881 6043 14891 6077
rect 14839 6031 14891 6043
rect 15837 6077 15889 6205
rect 15837 6043 15847 6077
rect 15881 6043 15889 6077
rect 15837 6031 15889 6043
rect 15943 6179 15995 6205
rect 15943 6145 15951 6179
rect 15985 6145 15995 6179
rect 15943 6077 15995 6145
rect 15943 6043 15951 6077
rect 15985 6043 15995 6077
rect 15943 6031 15995 6043
rect 16389 6179 16441 6205
rect 16389 6145 16399 6179
rect 16433 6145 16441 6179
rect 16389 6077 16441 6145
rect 16389 6043 16399 6077
rect 16433 6043 16441 6077
rect 16679 6077 16731 6205
rect 16389 6031 16441 6043
rect 16679 6043 16687 6077
rect 16721 6043 16731 6077
rect 16679 6031 16731 6043
rect 17677 6077 17729 6205
rect 17677 6043 17687 6077
rect 17721 6043 17729 6077
rect 17677 6031 17729 6043
rect 17783 6179 17835 6205
rect 17783 6145 17791 6179
rect 17825 6145 17835 6179
rect 17783 6077 17835 6145
rect 17783 6043 17791 6077
rect 17825 6043 17835 6077
rect 17783 6031 17835 6043
rect 18413 6179 18465 6205
rect 18413 6145 18423 6179
rect 18457 6145 18465 6179
rect 18413 6077 18465 6145
rect 18413 6043 18423 6077
rect 18457 6043 18465 6077
rect 18413 6031 18465 6043
rect 18611 6172 18663 6205
rect 18611 6138 18619 6172
rect 18653 6138 18663 6172
rect 18611 6077 18663 6138
rect 18611 6043 18619 6077
rect 18653 6043 18663 6077
rect 18611 6031 18663 6043
rect 18781 6172 18833 6205
rect 18781 6138 18791 6172
rect 18825 6138 18833 6172
rect 18781 6077 18833 6138
rect 18781 6043 18791 6077
rect 18825 6043 18833 6077
rect 18781 6031 18833 6043
rect 1131 5925 1183 5937
rect 1131 5891 1139 5925
rect 1173 5891 1183 5925
rect 1131 5830 1183 5891
rect 1131 5796 1139 5830
rect 1173 5796 1183 5830
rect 1131 5763 1183 5796
rect 1301 5925 1353 5937
rect 1301 5891 1311 5925
rect 1345 5891 1353 5925
rect 1301 5830 1353 5891
rect 1301 5796 1311 5830
rect 1345 5796 1353 5830
rect 1301 5763 1353 5796
rect 1407 5925 1459 5937
rect 1407 5891 1415 5925
rect 1449 5891 1459 5925
rect 1407 5823 1459 5891
rect 1407 5789 1415 5823
rect 1449 5789 1459 5823
rect 1407 5763 1459 5789
rect 2037 5925 2089 5937
rect 2037 5891 2047 5925
rect 2081 5891 2089 5925
rect 2037 5823 2089 5891
rect 2037 5789 2047 5823
rect 2081 5789 2089 5823
rect 2037 5763 2089 5789
rect 2235 5917 2287 5937
rect 2235 5883 2243 5917
rect 2277 5883 2287 5917
rect 2235 5849 2287 5883
rect 2235 5815 2243 5849
rect 2277 5815 2287 5849
rect 2235 5779 2287 5815
rect 2317 5917 2375 5937
rect 2317 5883 2329 5917
rect 2363 5883 2375 5917
rect 2317 5849 2375 5883
rect 2317 5815 2329 5849
rect 2363 5815 2375 5849
rect 2317 5779 2375 5815
rect 2405 5917 2457 5937
rect 2405 5883 2415 5917
rect 2449 5883 2457 5917
rect 2405 5836 2457 5883
rect 2405 5802 2415 5836
rect 2449 5802 2457 5836
rect 2405 5779 2457 5802
rect 2511 5925 2563 5937
rect 2511 5891 2519 5925
rect 2553 5891 2563 5925
rect 2511 5823 2563 5891
rect 2511 5789 2519 5823
rect 2553 5789 2563 5823
rect 2511 5763 2563 5789
rect 2957 5925 3009 5937
rect 2957 5891 2967 5925
rect 3001 5891 3009 5925
rect 2957 5823 3009 5891
rect 2957 5789 2967 5823
rect 3001 5789 3009 5823
rect 2957 5763 3009 5789
rect 3063 5917 3115 5937
rect 3063 5883 3071 5917
rect 3105 5883 3115 5917
rect 3063 5836 3115 5883
rect 3063 5802 3071 5836
rect 3105 5802 3115 5836
rect 3063 5779 3115 5802
rect 3145 5917 3203 5937
rect 3145 5883 3157 5917
rect 3191 5883 3203 5917
rect 3145 5849 3203 5883
rect 3145 5815 3157 5849
rect 3191 5815 3203 5849
rect 3145 5779 3203 5815
rect 3233 5917 3285 5937
rect 3233 5883 3243 5917
rect 3277 5883 3285 5917
rect 3233 5849 3285 5883
rect 3233 5815 3243 5849
rect 3277 5815 3285 5849
rect 3233 5779 3285 5815
rect 3339 5925 3391 5937
rect 3339 5891 3347 5925
rect 3381 5891 3391 5925
rect 3339 5823 3391 5891
rect 3339 5789 3347 5823
rect 3381 5789 3391 5823
rect 3339 5763 3391 5789
rect 3601 5925 3653 5937
rect 3601 5891 3611 5925
rect 3645 5891 3653 5925
rect 3799 5925 3851 5937
rect 3601 5823 3653 5891
rect 3601 5789 3611 5823
rect 3645 5789 3653 5823
rect 3601 5763 3653 5789
rect 3799 5891 3807 5925
rect 3841 5891 3851 5925
rect 3799 5763 3851 5891
rect 4797 5925 4849 5937
rect 4797 5891 4807 5925
rect 4841 5891 4849 5925
rect 4797 5763 4849 5891
rect 4903 5925 4955 5937
rect 4903 5891 4911 5925
rect 4945 5891 4955 5925
rect 4903 5763 4955 5891
rect 5901 5925 5953 5937
rect 5901 5891 5911 5925
rect 5945 5891 5953 5925
rect 5901 5763 5953 5891
rect 6007 5925 6059 5937
rect 6007 5891 6015 5925
rect 6049 5891 6059 5925
rect 6007 5823 6059 5891
rect 6007 5789 6015 5823
rect 6049 5789 6059 5823
rect 6007 5763 6059 5789
rect 6637 5925 6689 5937
rect 6637 5891 6647 5925
rect 6681 5891 6689 5925
rect 6637 5823 6689 5891
rect 6637 5789 6647 5823
rect 6681 5789 6689 5823
rect 6637 5763 6689 5789
rect 6743 5925 6795 5937
rect 6743 5891 6751 5925
rect 6785 5891 6795 5925
rect 6743 5857 6795 5891
rect 6743 5823 6751 5857
rect 6785 5823 6795 5857
rect 6743 5789 6795 5823
rect 6743 5755 6751 5789
rect 6785 5755 6795 5789
rect 6743 5737 6795 5755
rect 6825 5925 6877 5937
rect 6825 5891 6835 5925
rect 6869 5898 6877 5925
rect 7571 5925 7623 5937
rect 6869 5891 6904 5898
rect 6825 5857 6904 5891
rect 6825 5823 6835 5857
rect 6869 5823 6904 5857
rect 6825 5814 6904 5823
rect 6934 5814 7007 5898
rect 7037 5865 7221 5898
rect 7037 5831 7071 5865
rect 7105 5831 7146 5865
rect 7180 5831 7221 5865
rect 7037 5814 7221 5831
rect 7251 5814 7293 5898
rect 7323 5865 7389 5898
rect 7323 5831 7343 5865
rect 7377 5831 7389 5865
rect 7323 5814 7389 5831
rect 7419 5865 7475 5898
rect 7419 5831 7429 5865
rect 7463 5831 7475 5865
rect 7419 5814 7475 5831
rect 7571 5891 7579 5925
rect 7613 5891 7623 5925
rect 6825 5789 6877 5814
rect 6825 5755 6835 5789
rect 6869 5755 6877 5789
rect 6825 5737 6877 5755
rect 7571 5763 7623 5891
rect 8569 5925 8621 5937
rect 8569 5891 8579 5925
rect 8613 5891 8621 5925
rect 8951 5925 9003 5937
rect 8569 5763 8621 5891
rect 8951 5891 8959 5925
rect 8993 5891 9003 5925
rect 8951 5823 9003 5891
rect 8951 5789 8959 5823
rect 8993 5789 9003 5823
rect 8951 5763 9003 5789
rect 9581 5925 9633 5937
rect 9581 5891 9591 5925
rect 9625 5891 9633 5925
rect 9581 5823 9633 5891
rect 9581 5789 9591 5823
rect 9625 5789 9633 5823
rect 9581 5763 9633 5789
rect 9871 5925 9923 5937
rect 9871 5891 9879 5925
rect 9913 5891 9923 5925
rect 9871 5857 9923 5891
rect 9871 5823 9879 5857
rect 9913 5823 9923 5857
rect 9871 5789 9923 5823
rect 9871 5755 9879 5789
rect 9913 5755 9923 5789
rect 9871 5737 9923 5755
rect 9953 5925 10005 5937
rect 9953 5891 9963 5925
rect 9997 5898 10005 5925
rect 10699 5925 10751 5937
rect 9997 5891 10032 5898
rect 9953 5857 10032 5891
rect 9953 5823 9963 5857
rect 9997 5823 10032 5857
rect 9953 5814 10032 5823
rect 10062 5814 10135 5898
rect 10165 5865 10349 5898
rect 10165 5831 10199 5865
rect 10233 5831 10274 5865
rect 10308 5831 10349 5865
rect 10165 5814 10349 5831
rect 10379 5814 10421 5898
rect 10451 5865 10517 5898
rect 10451 5831 10471 5865
rect 10505 5831 10517 5865
rect 10451 5814 10517 5831
rect 10547 5865 10603 5898
rect 10547 5831 10557 5865
rect 10591 5831 10603 5865
rect 10547 5814 10603 5831
rect 10699 5891 10707 5925
rect 10741 5891 10751 5925
rect 10699 5823 10751 5891
rect 9953 5789 10005 5814
rect 9953 5755 9963 5789
rect 9997 5755 10005 5789
rect 9953 5737 10005 5755
rect 10699 5789 10707 5823
rect 10741 5789 10751 5823
rect 10699 5763 10751 5789
rect 10961 5925 11013 5937
rect 10961 5891 10971 5925
rect 11005 5891 11013 5925
rect 10961 5823 11013 5891
rect 10961 5789 10971 5823
rect 11005 5789 11013 5823
rect 10961 5763 11013 5789
rect 11068 5925 11163 5937
rect 11068 5891 11099 5925
rect 11133 5891 11163 5925
rect 11068 5857 11163 5891
rect 11068 5823 11099 5857
rect 11133 5823 11163 5857
rect 11068 5737 11163 5823
rect 11193 5925 11245 5937
rect 11193 5891 11203 5925
rect 11237 5895 11245 5925
rect 11527 5925 11579 5937
rect 11237 5891 11271 5895
rect 11193 5857 11271 5891
rect 11193 5823 11203 5857
rect 11237 5823 11271 5857
rect 11193 5811 11271 5823
rect 11301 5883 11355 5895
rect 11301 5849 11311 5883
rect 11345 5849 11355 5883
rect 11301 5811 11355 5849
rect 11385 5883 11441 5895
rect 11385 5849 11395 5883
rect 11429 5849 11441 5883
rect 11385 5811 11441 5849
rect 11527 5891 11535 5925
rect 11569 5891 11579 5925
rect 11527 5823 11579 5891
rect 11193 5737 11255 5811
rect 11527 5789 11535 5823
rect 11569 5789 11579 5823
rect 11527 5763 11579 5789
rect 12157 5925 12209 5937
rect 12157 5891 12167 5925
rect 12201 5891 12209 5925
rect 12157 5823 12209 5891
rect 12157 5789 12167 5823
rect 12201 5789 12209 5823
rect 12157 5763 12209 5789
rect 12263 5925 12315 5937
rect 12263 5891 12271 5925
rect 12305 5891 12315 5925
rect 12263 5857 12315 5891
rect 12263 5823 12271 5857
rect 12305 5823 12315 5857
rect 12263 5789 12315 5823
rect 12263 5755 12271 5789
rect 12305 5755 12315 5789
rect 12263 5737 12315 5755
rect 12345 5925 12397 5937
rect 12345 5891 12355 5925
rect 12389 5898 12397 5925
rect 13091 5925 13143 5937
rect 12389 5891 12424 5898
rect 12345 5857 12424 5891
rect 12345 5823 12355 5857
rect 12389 5823 12424 5857
rect 12345 5814 12424 5823
rect 12454 5814 12527 5898
rect 12557 5865 12741 5898
rect 12557 5831 12591 5865
rect 12625 5831 12666 5865
rect 12700 5831 12741 5865
rect 12557 5814 12741 5831
rect 12771 5814 12813 5898
rect 12843 5865 12909 5898
rect 12843 5831 12863 5865
rect 12897 5831 12909 5865
rect 12843 5814 12909 5831
rect 12939 5865 12995 5898
rect 12939 5831 12949 5865
rect 12983 5831 12995 5865
rect 12939 5814 12995 5831
rect 13091 5891 13099 5925
rect 13133 5891 13143 5925
rect 13091 5823 13143 5891
rect 12345 5789 12397 5814
rect 12345 5755 12355 5789
rect 12389 5755 12397 5789
rect 12345 5737 12397 5755
rect 13091 5789 13099 5823
rect 13133 5789 13143 5823
rect 13091 5763 13143 5789
rect 13721 5925 13773 5937
rect 13721 5891 13731 5925
rect 13765 5891 13773 5925
rect 14287 5925 14339 5937
rect 13721 5823 13773 5891
rect 13721 5789 13731 5823
rect 13765 5789 13773 5823
rect 13721 5763 13773 5789
rect 14287 5891 14295 5925
rect 14329 5891 14339 5925
rect 14287 5857 14339 5891
rect 14287 5823 14295 5857
rect 14329 5823 14339 5857
rect 14287 5789 14339 5823
rect 14287 5755 14295 5789
rect 14329 5755 14339 5789
rect 14287 5737 14339 5755
rect 14369 5925 14421 5937
rect 14369 5891 14379 5925
rect 14413 5898 14421 5925
rect 15115 5925 15167 5937
rect 14413 5891 14448 5898
rect 14369 5857 14448 5891
rect 14369 5823 14379 5857
rect 14413 5823 14448 5857
rect 14369 5814 14448 5823
rect 14478 5814 14551 5898
rect 14581 5865 14765 5898
rect 14581 5831 14615 5865
rect 14649 5831 14690 5865
rect 14724 5831 14765 5865
rect 14581 5814 14765 5831
rect 14795 5814 14837 5898
rect 14867 5865 14933 5898
rect 14867 5831 14887 5865
rect 14921 5831 14933 5865
rect 14867 5814 14933 5831
rect 14963 5865 15019 5898
rect 14963 5831 14973 5865
rect 15007 5831 15019 5865
rect 14963 5814 15019 5831
rect 15115 5891 15123 5925
rect 15157 5891 15167 5925
rect 14369 5789 14421 5814
rect 14369 5755 14379 5789
rect 14413 5755 14421 5789
rect 14369 5737 14421 5755
rect 15115 5763 15167 5891
rect 16113 5925 16165 5937
rect 16113 5891 16123 5925
rect 16157 5891 16165 5925
rect 16113 5763 16165 5891
rect 16219 5925 16271 5937
rect 16219 5891 16227 5925
rect 16261 5891 16271 5925
rect 16219 5763 16271 5891
rect 17217 5925 17269 5937
rect 17217 5891 17227 5925
rect 17261 5891 17269 5925
rect 17217 5763 17269 5891
rect 17323 5925 17375 5937
rect 17323 5891 17331 5925
rect 17365 5891 17375 5925
rect 17323 5763 17375 5891
rect 18321 5925 18373 5937
rect 18321 5891 18331 5925
rect 18365 5891 18373 5925
rect 18321 5763 18373 5891
rect 18611 5925 18663 5937
rect 18611 5891 18619 5925
rect 18653 5891 18663 5925
rect 18611 5830 18663 5891
rect 18611 5796 18619 5830
rect 18653 5796 18663 5830
rect 18611 5763 18663 5796
rect 18781 5925 18833 5937
rect 18781 5891 18791 5925
rect 18825 5891 18833 5925
rect 18781 5830 18833 5891
rect 18781 5796 18791 5830
rect 18825 5796 18833 5830
rect 18781 5763 18833 5796
rect 1131 5084 1183 5117
rect 1131 5050 1139 5084
rect 1173 5050 1183 5084
rect 1131 4989 1183 5050
rect 1131 4955 1139 4989
rect 1173 4955 1183 4989
rect 1131 4943 1183 4955
rect 1301 5084 1353 5117
rect 1301 5050 1311 5084
rect 1345 5050 1353 5084
rect 1301 4989 1353 5050
rect 1301 4955 1311 4989
rect 1345 4955 1353 4989
rect 1301 4943 1353 4955
rect 1407 5091 1459 5117
rect 1407 5057 1415 5091
rect 1449 5057 1459 5091
rect 1407 4989 1459 5057
rect 1407 4955 1415 4989
rect 1449 4955 1459 4989
rect 1407 4943 1459 4955
rect 1853 5091 1905 5117
rect 1853 5057 1863 5091
rect 1897 5057 1905 5091
rect 1853 4989 1905 5057
rect 1853 4955 1863 4989
rect 1897 4955 1905 4989
rect 1853 4943 1905 4955
rect 1960 5057 2055 5143
rect 1960 5023 1991 5057
rect 2025 5023 2055 5057
rect 1960 4989 2055 5023
rect 1960 4955 1991 4989
rect 2025 4955 2055 4989
rect 1960 4943 2055 4955
rect 2085 5069 2147 5143
rect 2419 5091 2471 5117
rect 2085 5057 2163 5069
rect 2085 5023 2095 5057
rect 2129 5023 2163 5057
rect 2085 4989 2163 5023
rect 2085 4955 2095 4989
rect 2129 4985 2163 4989
rect 2193 5031 2247 5069
rect 2193 4997 2203 5031
rect 2237 4997 2247 5031
rect 2193 4985 2247 4997
rect 2277 5031 2333 5069
rect 2277 4997 2287 5031
rect 2321 4997 2333 5031
rect 2277 4985 2333 4997
rect 2419 5057 2427 5091
rect 2461 5057 2471 5091
rect 2419 4989 2471 5057
rect 2129 4955 2137 4985
rect 2085 4943 2137 4955
rect 2419 4955 2427 4989
rect 2461 4955 2471 4989
rect 2419 4943 2471 4955
rect 2681 5091 2733 5117
rect 2681 5057 2691 5091
rect 2725 5057 2733 5091
rect 2681 4989 2733 5057
rect 2681 4955 2691 4989
rect 2725 4955 2733 4989
rect 2681 4943 2733 4955
rect 2880 5057 2975 5143
rect 2880 5023 2911 5057
rect 2945 5023 2975 5057
rect 2880 4989 2975 5023
rect 2880 4955 2911 4989
rect 2945 4955 2975 4989
rect 2880 4943 2975 4955
rect 3005 5069 3067 5143
rect 3339 5091 3391 5117
rect 3005 5057 3083 5069
rect 3005 5023 3015 5057
rect 3049 5023 3083 5057
rect 3005 4989 3083 5023
rect 3005 4955 3015 4989
rect 3049 4985 3083 4989
rect 3113 5031 3167 5069
rect 3113 4997 3123 5031
rect 3157 4997 3167 5031
rect 3113 4985 3167 4997
rect 3197 5031 3253 5069
rect 3197 4997 3207 5031
rect 3241 4997 3253 5031
rect 3197 4985 3253 4997
rect 3339 5057 3347 5091
rect 3381 5057 3391 5091
rect 3339 4989 3391 5057
rect 3049 4955 3057 4985
rect 3005 4943 3057 4955
rect 3339 4955 3347 4989
rect 3381 4955 3391 4989
rect 3339 4943 3391 4955
rect 3601 5091 3653 5117
rect 3601 5057 3611 5091
rect 3645 5057 3653 5091
rect 3804 5079 3854 5143
rect 3601 4989 3653 5057
rect 3601 4955 3611 4989
rect 3645 4955 3653 4989
rect 3601 4943 3653 4955
rect 3707 5065 3759 5079
rect 3707 5031 3715 5065
rect 3749 5031 3759 5065
rect 3707 4997 3759 5031
rect 3707 4963 3715 4997
rect 3749 4963 3759 4997
rect 3707 4951 3759 4963
rect 3789 5065 3854 5079
rect 3789 5031 3808 5065
rect 3842 5031 3854 5065
rect 3789 4997 3854 5031
rect 3789 4963 3808 4997
rect 3842 4963 3854 4997
rect 3789 4951 3854 4963
rect 3804 4943 3854 4951
rect 3884 5094 3938 5143
rect 3884 5060 3894 5094
rect 3928 5060 3938 5094
rect 3884 5013 3938 5060
rect 3884 4979 3894 5013
rect 3928 4979 3938 5013
rect 3884 4943 3938 4979
rect 3968 5125 4021 5143
rect 3968 5091 3978 5125
rect 4012 5091 4021 5125
rect 4445 5125 4497 5143
rect 3968 5057 4021 5091
rect 3968 5023 3978 5057
rect 4012 5023 4021 5057
rect 3968 4989 4021 5023
rect 3968 4955 3978 4989
rect 4012 4955 4021 4989
rect 3968 4943 4021 4955
rect 4075 5091 4127 5117
rect 4075 5057 4083 5091
rect 4117 5057 4127 5091
rect 4075 4989 4127 5057
rect 4075 4955 4083 4989
rect 4117 4955 4127 4989
rect 4075 4943 4127 4955
rect 4337 5091 4389 5117
rect 4337 5057 4347 5091
rect 4381 5057 4389 5091
rect 4337 4989 4389 5057
rect 4337 4955 4347 4989
rect 4381 4955 4389 4989
rect 4337 4943 4389 4955
rect 4445 5091 4453 5125
rect 4487 5091 4497 5125
rect 4445 5057 4497 5091
rect 4445 5023 4453 5057
rect 4487 5023 4497 5057
rect 4445 4989 4497 5023
rect 4445 4955 4453 4989
rect 4487 4955 4497 4989
rect 4445 4943 4497 4955
rect 4527 5125 4581 5143
rect 4527 5091 4537 5125
rect 4571 5091 4581 5125
rect 4527 5057 4581 5091
rect 4527 5023 4537 5057
rect 4571 5023 4581 5057
rect 4527 4989 4581 5023
rect 4527 4955 4537 4989
rect 4571 4955 4581 4989
rect 4527 4943 4581 4955
rect 4611 5125 4663 5143
rect 4611 5091 4621 5125
rect 4655 5091 4663 5125
rect 4611 5057 4663 5091
rect 4611 5023 4621 5057
rect 4655 5023 4663 5057
rect 4611 4989 4663 5023
rect 4611 4955 4621 4989
rect 4655 4955 4663 4989
rect 4611 4943 4663 4955
rect 4719 4989 4771 5117
rect 4719 4955 4727 4989
rect 4761 4955 4771 4989
rect 4719 4943 4771 4955
rect 5717 4989 5769 5117
rect 6651 5125 6703 5143
rect 5717 4955 5727 4989
rect 5761 4955 5769 4989
rect 5717 4943 5769 4955
rect 5823 5078 5875 5101
rect 5823 5044 5831 5078
rect 5865 5044 5875 5078
rect 5823 4997 5875 5044
rect 5823 4963 5831 4997
rect 5865 4963 5875 4997
rect 5823 4943 5875 4963
rect 5905 5065 5963 5101
rect 5905 5031 5917 5065
rect 5951 5031 5963 5065
rect 5905 4997 5963 5031
rect 5905 4963 5917 4997
rect 5951 4963 5963 4997
rect 5905 4943 5963 4963
rect 5993 5065 6045 5101
rect 5993 5031 6003 5065
rect 6037 5031 6045 5065
rect 5993 4997 6045 5031
rect 5993 4963 6003 4997
rect 6037 4963 6045 4997
rect 5993 4943 6045 4963
rect 6375 5084 6427 5117
rect 6375 5050 6383 5084
rect 6417 5050 6427 5084
rect 6375 4989 6427 5050
rect 6375 4955 6383 4989
rect 6417 4955 6427 4989
rect 6375 4943 6427 4955
rect 6545 5084 6597 5117
rect 6545 5050 6555 5084
rect 6589 5050 6597 5084
rect 6545 4989 6597 5050
rect 6545 4955 6555 4989
rect 6589 4955 6597 4989
rect 6545 4943 6597 4955
rect 6651 5091 6659 5125
rect 6693 5091 6703 5125
rect 6651 5057 6703 5091
rect 6651 5023 6659 5057
rect 6693 5023 6703 5057
rect 6651 4989 6703 5023
rect 6651 4955 6659 4989
rect 6693 4955 6703 4989
rect 6651 4943 6703 4955
rect 6733 5125 6785 5143
rect 6733 5091 6743 5125
rect 6777 5091 6785 5125
rect 6733 5066 6785 5091
rect 7847 5125 7899 5143
rect 7479 5091 7531 5117
rect 6733 5057 6812 5066
rect 6733 5023 6743 5057
rect 6777 5023 6812 5057
rect 6733 4989 6812 5023
rect 6733 4955 6743 4989
rect 6777 4982 6812 4989
rect 6842 4982 6915 5066
rect 6945 5049 7129 5066
rect 6945 5015 6979 5049
rect 7013 5015 7054 5049
rect 7088 5015 7129 5049
rect 6945 4982 7129 5015
rect 7159 4982 7201 5066
rect 7231 5049 7297 5066
rect 7231 5015 7251 5049
rect 7285 5015 7297 5049
rect 7231 4982 7297 5015
rect 7327 5049 7383 5066
rect 7327 5015 7337 5049
rect 7371 5015 7383 5049
rect 7327 4982 7383 5015
rect 7479 5057 7487 5091
rect 7521 5057 7531 5091
rect 7479 4989 7531 5057
rect 6777 4955 6785 4982
rect 6733 4943 6785 4955
rect 7479 4955 7487 4989
rect 7521 4955 7531 4989
rect 7479 4943 7531 4955
rect 7741 5091 7793 5117
rect 7741 5057 7751 5091
rect 7785 5057 7793 5091
rect 7741 4989 7793 5057
rect 7741 4955 7751 4989
rect 7785 4955 7793 4989
rect 7741 4943 7793 4955
rect 7847 5091 7855 5125
rect 7889 5091 7899 5125
rect 7847 5057 7899 5091
rect 7847 5023 7855 5057
rect 7889 5023 7899 5057
rect 7847 4989 7899 5023
rect 7847 4955 7855 4989
rect 7889 4955 7899 4989
rect 7847 4943 7899 4955
rect 7929 5125 7981 5143
rect 7929 5091 7939 5125
rect 7973 5091 7981 5125
rect 7929 5066 7981 5091
rect 9135 5133 9191 5143
rect 8675 5091 8727 5117
rect 7929 5057 8008 5066
rect 7929 5023 7939 5057
rect 7973 5023 8008 5057
rect 7929 4989 8008 5023
rect 7929 4955 7939 4989
rect 7973 4982 8008 4989
rect 8038 4982 8111 5066
rect 8141 5049 8325 5066
rect 8141 5015 8175 5049
rect 8209 5015 8250 5049
rect 8284 5015 8325 5049
rect 8141 4982 8325 5015
rect 8355 4982 8397 5066
rect 8427 5049 8493 5066
rect 8427 5015 8447 5049
rect 8481 5015 8493 5049
rect 8427 4982 8493 5015
rect 8523 5049 8579 5066
rect 8523 5015 8533 5049
rect 8567 5015 8579 5049
rect 8523 4982 8579 5015
rect 8675 5057 8683 5091
rect 8717 5057 8727 5091
rect 8675 4989 8727 5057
rect 7973 4955 7981 4982
rect 7929 4943 7981 4955
rect 8675 4955 8683 4989
rect 8717 4955 8727 4989
rect 8675 4943 8727 4955
rect 8937 5091 8989 5117
rect 8937 5057 8947 5091
rect 8981 5057 8989 5091
rect 8937 4989 8989 5057
rect 8937 4955 8947 4989
rect 8981 4955 8989 4989
rect 8937 4943 8989 4955
rect 9135 5099 9147 5133
rect 9181 5099 9191 5133
rect 9135 5065 9191 5099
rect 9135 5031 9147 5065
rect 9181 5031 9191 5065
rect 9135 4997 9191 5031
rect 9135 4963 9147 4997
rect 9181 4963 9191 4997
rect 9135 4943 9191 4963
rect 9221 5057 9352 5143
rect 9221 5023 9233 5057
rect 9267 5023 9307 5057
rect 9341 5023 9352 5057
rect 9221 4989 9352 5023
rect 9221 4955 9233 4989
rect 9267 4955 9307 4989
rect 9341 4955 9352 4989
rect 9221 4943 9352 4955
rect 9382 5125 9460 5143
rect 9382 5091 9407 5125
rect 9441 5091 9460 5125
rect 9382 5057 9460 5091
rect 9382 5023 9407 5057
rect 9441 5023 9460 5057
rect 9382 4989 9460 5023
rect 9382 4955 9407 4989
rect 9441 4955 9460 4989
rect 9382 4943 9460 4955
rect 9490 4943 9551 5143
rect 9581 5057 9633 5143
rect 10423 5125 10475 5143
rect 9581 5023 9591 5057
rect 9625 5023 9633 5057
rect 9581 4989 9633 5023
rect 9581 4955 9591 4989
rect 9625 4955 9633 4989
rect 9581 4943 9633 4955
rect 9687 5091 9739 5117
rect 9687 5057 9695 5091
rect 9729 5057 9739 5091
rect 9687 4989 9739 5057
rect 9687 4955 9695 4989
rect 9729 4955 9739 4989
rect 9687 4943 9739 4955
rect 10317 5091 10369 5117
rect 10317 5057 10327 5091
rect 10361 5057 10369 5091
rect 10317 4989 10369 5057
rect 10317 4955 10327 4989
rect 10361 4955 10369 4989
rect 10317 4943 10369 4955
rect 10423 5091 10431 5125
rect 10465 5091 10475 5125
rect 10423 5057 10475 5091
rect 10423 5023 10431 5057
rect 10465 5023 10475 5057
rect 10423 4989 10475 5023
rect 10423 4955 10431 4989
rect 10465 4955 10475 4989
rect 10423 4943 10475 4955
rect 10505 5125 10557 5143
rect 10505 5091 10515 5125
rect 10549 5091 10557 5125
rect 10505 5066 10557 5091
rect 13091 5125 13143 5143
rect 10505 5057 10584 5066
rect 10505 5023 10515 5057
rect 10549 5023 10584 5057
rect 10505 4989 10584 5023
rect 10505 4955 10515 4989
rect 10549 4982 10584 4989
rect 10614 4982 10687 5066
rect 10717 5049 10901 5066
rect 10717 5015 10751 5049
rect 10785 5015 10826 5049
rect 10860 5015 10901 5049
rect 10717 4982 10901 5015
rect 10931 4982 10973 5066
rect 11003 5049 11069 5066
rect 11003 5015 11023 5049
rect 11057 5015 11069 5049
rect 11003 4982 11069 5015
rect 11099 5049 11155 5066
rect 11099 5015 11109 5049
rect 11143 5015 11155 5049
rect 11099 4982 11155 5015
rect 10549 4955 10557 4982
rect 11527 4989 11579 5117
rect 10505 4943 10557 4955
rect 11527 4955 11535 4989
rect 11569 4955 11579 4989
rect 11527 4943 11579 4955
rect 12525 4989 12577 5117
rect 12525 4955 12535 4989
rect 12569 4955 12577 4989
rect 12525 4943 12577 4955
rect 12631 5091 12683 5117
rect 12631 5057 12639 5091
rect 12673 5057 12683 5091
rect 12631 4989 12683 5057
rect 12631 4955 12639 4989
rect 12673 4955 12683 4989
rect 12631 4943 12683 4955
rect 12893 5091 12945 5117
rect 12893 5057 12903 5091
rect 12937 5057 12945 5091
rect 12893 4989 12945 5057
rect 12893 4955 12903 4989
rect 12937 4955 12945 4989
rect 12893 4943 12945 4955
rect 13091 5091 13099 5125
rect 13133 5091 13143 5125
rect 13091 5057 13143 5091
rect 13091 5023 13099 5057
rect 13133 5023 13143 5057
rect 13091 4989 13143 5023
rect 13091 4955 13099 4989
rect 13133 4955 13143 4989
rect 13091 4943 13143 4955
rect 13173 5125 13225 5143
rect 13173 5091 13183 5125
rect 13217 5091 13225 5125
rect 13173 5066 13225 5091
rect 13173 5057 13252 5066
rect 13173 5023 13183 5057
rect 13217 5023 13252 5057
rect 13173 4989 13252 5023
rect 13173 4955 13183 4989
rect 13217 4982 13252 4989
rect 13282 4982 13355 5066
rect 13385 5049 13569 5066
rect 13385 5015 13419 5049
rect 13453 5015 13494 5049
rect 13528 5015 13569 5049
rect 13385 4982 13569 5015
rect 13599 4982 13641 5066
rect 13671 5049 13737 5066
rect 13671 5015 13691 5049
rect 13725 5015 13737 5049
rect 13671 4982 13737 5015
rect 13767 5049 13823 5066
rect 13767 5015 13777 5049
rect 13811 5015 13823 5049
rect 13767 4982 13823 5015
rect 13919 4989 13971 5117
rect 13217 4955 13225 4982
rect 13173 4943 13225 4955
rect 13919 4955 13927 4989
rect 13961 4955 13971 4989
rect 13919 4943 13971 4955
rect 14917 4989 14969 5117
rect 14917 4955 14927 4989
rect 14961 4955 14969 4989
rect 14917 4943 14969 4955
rect 15023 4989 15075 5117
rect 15023 4955 15031 4989
rect 15065 4955 15075 4989
rect 15023 4943 15075 4955
rect 16021 4989 16073 5117
rect 16021 4955 16031 4989
rect 16065 4955 16073 4989
rect 16021 4943 16073 4955
rect 16127 5091 16179 5117
rect 16127 5057 16135 5091
rect 16169 5057 16179 5091
rect 16127 4989 16179 5057
rect 16127 4955 16135 4989
rect 16169 4955 16179 4989
rect 16127 4943 16179 4955
rect 16389 5091 16441 5117
rect 16389 5057 16399 5091
rect 16433 5057 16441 5091
rect 16389 4989 16441 5057
rect 16389 4955 16399 4989
rect 16433 4955 16441 4989
rect 16679 4989 16731 5117
rect 16389 4943 16441 4955
rect 16679 4955 16687 4989
rect 16721 4955 16731 4989
rect 16679 4943 16731 4955
rect 17677 4989 17729 5117
rect 17677 4955 17687 4989
rect 17721 4955 17729 4989
rect 17677 4943 17729 4955
rect 17783 5091 17835 5117
rect 17783 5057 17791 5091
rect 17825 5057 17835 5091
rect 17783 4989 17835 5057
rect 17783 4955 17791 4989
rect 17825 4955 17835 4989
rect 17783 4943 17835 4955
rect 18413 5091 18465 5117
rect 18413 5057 18423 5091
rect 18457 5057 18465 5091
rect 18413 4989 18465 5057
rect 18413 4955 18423 4989
rect 18457 4955 18465 4989
rect 18413 4943 18465 4955
rect 18611 5084 18663 5117
rect 18611 5050 18619 5084
rect 18653 5050 18663 5084
rect 18611 4989 18663 5050
rect 18611 4955 18619 4989
rect 18653 4955 18663 4989
rect 18611 4943 18663 4955
rect 18781 5084 18833 5117
rect 18781 5050 18791 5084
rect 18825 5050 18833 5084
rect 18781 4989 18833 5050
rect 18781 4955 18791 4989
rect 18825 4955 18833 4989
rect 18781 4943 18833 4955
rect 1131 4837 1183 4849
rect 1131 4803 1139 4837
rect 1173 4803 1183 4837
rect 1131 4742 1183 4803
rect 1131 4708 1139 4742
rect 1173 4708 1183 4742
rect 1131 4675 1183 4708
rect 1301 4837 1353 4849
rect 1301 4803 1311 4837
rect 1345 4803 1353 4837
rect 1301 4742 1353 4803
rect 1301 4708 1311 4742
rect 1345 4708 1353 4742
rect 1301 4675 1353 4708
rect 1407 4837 1459 4849
rect 1407 4803 1415 4837
rect 1449 4803 1459 4837
rect 1407 4735 1459 4803
rect 1407 4701 1415 4735
rect 1449 4701 1459 4735
rect 1407 4675 1459 4701
rect 1853 4837 1905 4849
rect 1853 4803 1863 4837
rect 1897 4803 1905 4837
rect 1853 4735 1905 4803
rect 1853 4701 1863 4735
rect 1897 4701 1905 4735
rect 2051 4829 2103 4843
rect 2051 4795 2059 4829
rect 2093 4795 2103 4829
rect 2051 4761 2103 4795
rect 2051 4727 2059 4761
rect 2093 4727 2103 4761
rect 2051 4715 2103 4727
rect 2133 4813 2187 4843
rect 2133 4779 2143 4813
rect 2177 4779 2187 4813
rect 2133 4715 2187 4779
rect 2217 4829 2269 4843
rect 2217 4795 2227 4829
rect 2261 4795 2269 4829
rect 2217 4761 2269 4795
rect 2323 4837 2375 4849
rect 2323 4803 2331 4837
rect 2365 4803 2375 4837
rect 2323 4765 2375 4803
rect 2405 4829 2460 4849
rect 2405 4795 2415 4829
rect 2449 4795 2460 4829
rect 2405 4765 2460 4795
rect 2490 4824 2555 4849
rect 2490 4790 2507 4824
rect 2541 4790 2555 4824
rect 2490 4765 2555 4790
rect 2585 4765 2658 4849
rect 2688 4837 2790 4849
rect 2688 4803 2746 4837
rect 2780 4803 2790 4837
rect 2688 4769 2790 4803
rect 2688 4765 2746 4769
rect 2217 4727 2227 4761
rect 2261 4727 2269 4761
rect 2217 4715 2269 4727
rect 1853 4675 1905 4701
rect 2703 4735 2746 4765
rect 2780 4735 2790 4769
rect 2703 4699 2790 4735
rect 2820 4829 2885 4849
rect 2820 4795 2830 4829
rect 2864 4795 2885 4829
rect 2820 4765 2885 4795
rect 2915 4819 2969 4849
rect 2915 4785 2925 4819
rect 2959 4785 2969 4819
rect 2915 4765 2969 4785
rect 2999 4765 3083 4849
rect 3113 4829 3166 4849
rect 3113 4795 3124 4829
rect 3158 4795 3166 4829
rect 3113 4765 3166 4795
rect 3239 4837 3293 4849
rect 3239 4803 3247 4837
rect 3281 4803 3293 4837
rect 3239 4766 3293 4803
rect 2820 4699 2870 4765
rect 3239 4732 3247 4766
rect 3281 4732 3293 4766
rect 3239 4695 3293 4732
rect 3239 4661 3247 4695
rect 3281 4661 3293 4695
rect 3239 4649 3293 4661
rect 3323 4807 3377 4849
rect 3323 4773 3333 4807
rect 3367 4773 3377 4807
rect 3323 4727 3377 4773
rect 3323 4693 3333 4727
rect 3367 4693 3377 4727
rect 3323 4649 3377 4693
rect 3407 4831 3459 4849
rect 3984 4837 4079 4849
rect 3407 4797 3417 4831
rect 3451 4797 3459 4831
rect 3407 4763 3459 4797
rect 3407 4729 3417 4763
rect 3451 4729 3459 4763
rect 3407 4695 3459 4729
rect 3407 4661 3417 4695
rect 3451 4661 3459 4695
rect 3407 4649 3459 4661
rect 3984 4803 4015 4837
rect 4049 4803 4079 4837
rect 3984 4769 4079 4803
rect 3984 4735 4015 4769
rect 4049 4735 4079 4769
rect 3984 4649 4079 4735
rect 4109 4837 4161 4849
rect 4109 4803 4119 4837
rect 4153 4807 4161 4837
rect 4443 4837 4495 4849
rect 4153 4803 4187 4807
rect 4109 4769 4187 4803
rect 4109 4735 4119 4769
rect 4153 4735 4187 4769
rect 4109 4723 4187 4735
rect 4217 4795 4271 4807
rect 4217 4761 4227 4795
rect 4261 4761 4271 4795
rect 4217 4723 4271 4761
rect 4301 4795 4357 4807
rect 4301 4761 4311 4795
rect 4345 4761 4357 4795
rect 4301 4723 4357 4761
rect 4443 4803 4451 4837
rect 4485 4803 4495 4837
rect 4443 4735 4495 4803
rect 4109 4649 4171 4723
rect 4443 4701 4451 4735
rect 4485 4701 4495 4735
rect 4443 4675 4495 4701
rect 4705 4837 4757 4849
rect 4705 4803 4715 4837
rect 4749 4803 4757 4837
rect 4705 4735 4757 4803
rect 4705 4701 4715 4735
rect 4749 4701 4757 4735
rect 4705 4675 4757 4701
rect 4903 4829 4959 4849
rect 4903 4795 4915 4829
rect 4949 4795 4959 4829
rect 4903 4761 4959 4795
rect 4903 4727 4915 4761
rect 4949 4727 4959 4761
rect 4903 4693 4959 4727
rect 4903 4659 4915 4693
rect 4949 4659 4959 4693
rect 4903 4649 4959 4659
rect 4989 4837 5120 4849
rect 4989 4803 5001 4837
rect 5035 4803 5075 4837
rect 5109 4803 5120 4837
rect 4989 4769 5120 4803
rect 4989 4735 5001 4769
rect 5035 4735 5075 4769
rect 5109 4735 5120 4769
rect 4989 4649 5120 4735
rect 5150 4837 5228 4849
rect 5150 4803 5175 4837
rect 5209 4803 5228 4837
rect 5150 4769 5228 4803
rect 5150 4735 5175 4769
rect 5209 4735 5228 4769
rect 5150 4701 5228 4735
rect 5150 4667 5175 4701
rect 5209 4667 5228 4701
rect 5150 4649 5228 4667
rect 5258 4649 5319 4849
rect 5349 4837 5401 4849
rect 5349 4803 5359 4837
rect 5393 4803 5401 4837
rect 5349 4769 5401 4803
rect 5349 4735 5359 4769
rect 5393 4735 5401 4769
rect 5349 4649 5401 4735
rect 5455 4837 5507 4849
rect 5455 4803 5463 4837
rect 5497 4803 5507 4837
rect 5455 4735 5507 4803
rect 5455 4701 5463 4735
rect 5497 4701 5507 4735
rect 5455 4675 5507 4701
rect 5717 4837 5769 4849
rect 5717 4803 5727 4837
rect 5761 4803 5769 4837
rect 5717 4735 5769 4803
rect 5717 4701 5727 4735
rect 5761 4701 5769 4735
rect 5717 4675 5769 4701
rect 5823 4829 5879 4849
rect 5823 4795 5835 4829
rect 5869 4795 5879 4829
rect 5823 4761 5879 4795
rect 5823 4727 5835 4761
rect 5869 4727 5879 4761
rect 5823 4693 5879 4727
rect 5823 4659 5835 4693
rect 5869 4659 5879 4693
rect 5823 4649 5879 4659
rect 5909 4837 6040 4849
rect 5909 4803 5921 4837
rect 5955 4803 5995 4837
rect 6029 4803 6040 4837
rect 5909 4769 6040 4803
rect 5909 4735 5921 4769
rect 5955 4735 5995 4769
rect 6029 4735 6040 4769
rect 5909 4649 6040 4735
rect 6070 4837 6148 4849
rect 6070 4803 6095 4837
rect 6129 4803 6148 4837
rect 6070 4769 6148 4803
rect 6070 4735 6095 4769
rect 6129 4735 6148 4769
rect 6070 4701 6148 4735
rect 6070 4667 6095 4701
rect 6129 4667 6148 4701
rect 6070 4649 6148 4667
rect 6178 4649 6239 4849
rect 6269 4837 6321 4849
rect 6269 4803 6279 4837
rect 6313 4803 6321 4837
rect 6269 4769 6321 4803
rect 6269 4735 6279 4769
rect 6313 4735 6321 4769
rect 6269 4649 6321 4735
rect 6375 4837 6427 4849
rect 6375 4803 6383 4837
rect 6417 4803 6427 4837
rect 6375 4735 6427 4803
rect 6375 4701 6383 4735
rect 6417 4701 6427 4735
rect 6375 4675 6427 4701
rect 6637 4837 6689 4849
rect 6637 4803 6647 4837
rect 6681 4803 6689 4837
rect 6637 4735 6689 4803
rect 6637 4701 6647 4735
rect 6681 4701 6689 4735
rect 6743 4829 6795 4843
rect 6743 4795 6751 4829
rect 6785 4795 6795 4829
rect 6743 4761 6795 4795
rect 6743 4727 6751 4761
rect 6785 4727 6795 4761
rect 6743 4715 6795 4727
rect 6825 4813 6879 4843
rect 6825 4779 6835 4813
rect 6869 4779 6879 4813
rect 6825 4715 6879 4779
rect 6909 4829 6961 4843
rect 6909 4795 6919 4829
rect 6953 4795 6961 4829
rect 6909 4761 6961 4795
rect 7015 4837 7067 4849
rect 7015 4803 7023 4837
rect 7057 4803 7067 4837
rect 7015 4765 7067 4803
rect 7097 4829 7152 4849
rect 7097 4795 7107 4829
rect 7141 4795 7152 4829
rect 7097 4765 7152 4795
rect 7182 4824 7247 4849
rect 7182 4790 7199 4824
rect 7233 4790 7247 4824
rect 7182 4765 7247 4790
rect 7277 4765 7350 4849
rect 7380 4837 7482 4849
rect 7380 4803 7438 4837
rect 7472 4803 7482 4837
rect 7380 4769 7482 4803
rect 7380 4765 7438 4769
rect 6909 4727 6919 4761
rect 6953 4727 6961 4761
rect 6909 4715 6961 4727
rect 6637 4675 6689 4701
rect 7395 4735 7438 4765
rect 7472 4735 7482 4769
rect 7395 4699 7482 4735
rect 7512 4829 7577 4849
rect 7512 4795 7522 4829
rect 7556 4795 7577 4829
rect 7512 4765 7577 4795
rect 7607 4819 7661 4849
rect 7607 4785 7617 4819
rect 7651 4785 7661 4819
rect 7607 4765 7661 4785
rect 7691 4765 7775 4849
rect 7805 4829 7858 4849
rect 7805 4795 7816 4829
rect 7850 4795 7858 4829
rect 7805 4765 7858 4795
rect 7931 4837 7985 4849
rect 7931 4803 7939 4837
rect 7973 4803 7985 4837
rect 7931 4766 7985 4803
rect 7512 4699 7562 4765
rect 7931 4732 7939 4766
rect 7973 4732 7985 4766
rect 7931 4695 7985 4732
rect 7931 4661 7939 4695
rect 7973 4661 7985 4695
rect 7931 4649 7985 4661
rect 8015 4807 8069 4849
rect 8015 4773 8025 4807
rect 8059 4773 8069 4807
rect 8015 4727 8069 4773
rect 8015 4693 8025 4727
rect 8059 4693 8069 4727
rect 8015 4649 8069 4693
rect 8099 4831 8151 4849
rect 8099 4797 8109 4831
rect 8143 4797 8151 4831
rect 8099 4763 8151 4797
rect 8099 4729 8109 4763
rect 8143 4729 8151 4763
rect 8099 4695 8151 4729
rect 8099 4661 8109 4695
rect 8143 4661 8151 4695
rect 8215 4837 8267 4849
rect 8215 4803 8223 4837
rect 8257 4803 8267 4837
rect 8215 4735 8267 4803
rect 8215 4701 8223 4735
rect 8257 4701 8267 4735
rect 8215 4675 8267 4701
rect 8661 4837 8713 4849
rect 8661 4803 8671 4837
rect 8705 4803 8713 4837
rect 8951 4837 9003 4849
rect 8661 4735 8713 4803
rect 8661 4701 8671 4735
rect 8705 4701 8713 4735
rect 8661 4675 8713 4701
rect 8099 4649 8151 4661
rect 8951 4803 8959 4837
rect 8993 4803 9003 4837
rect 8951 4735 9003 4803
rect 8951 4701 8959 4735
rect 8993 4701 9003 4735
rect 8951 4675 9003 4701
rect 9581 4837 9633 4849
rect 9581 4803 9591 4837
rect 9625 4803 9633 4837
rect 9581 4735 9633 4803
rect 9581 4701 9591 4735
rect 9625 4701 9633 4735
rect 9581 4675 9633 4701
rect 9687 4837 9739 4849
rect 9687 4803 9695 4837
rect 9729 4803 9739 4837
rect 9687 4742 9739 4803
rect 9687 4708 9695 4742
rect 9729 4708 9739 4742
rect 9687 4675 9739 4708
rect 9857 4837 9909 4849
rect 9857 4803 9867 4837
rect 9901 4803 9909 4837
rect 9857 4742 9909 4803
rect 9857 4708 9867 4742
rect 9901 4708 9909 4742
rect 9857 4675 9909 4708
rect 9973 4831 10025 4849
rect 9973 4797 9981 4831
rect 10015 4797 10025 4831
rect 9973 4763 10025 4797
rect 9973 4729 9981 4763
rect 10015 4729 10025 4763
rect 9973 4695 10025 4729
rect 9973 4661 9981 4695
rect 10015 4661 10025 4695
rect 9973 4649 10025 4661
rect 10055 4807 10109 4849
rect 10055 4773 10065 4807
rect 10099 4773 10109 4807
rect 10055 4727 10109 4773
rect 10055 4693 10065 4727
rect 10099 4693 10109 4727
rect 10055 4649 10109 4693
rect 10139 4837 10193 4849
rect 10139 4803 10151 4837
rect 10185 4803 10193 4837
rect 10139 4766 10193 4803
rect 10139 4732 10151 4766
rect 10185 4732 10193 4766
rect 10266 4829 10319 4849
rect 10266 4795 10274 4829
rect 10308 4795 10319 4829
rect 10266 4765 10319 4795
rect 10349 4765 10433 4849
rect 10463 4819 10517 4849
rect 10463 4785 10473 4819
rect 10507 4785 10517 4819
rect 10463 4765 10517 4785
rect 10547 4829 10612 4849
rect 10547 4795 10568 4829
rect 10602 4795 10612 4829
rect 10547 4765 10612 4795
rect 10139 4695 10193 4732
rect 10139 4661 10151 4695
rect 10185 4661 10193 4695
rect 10562 4699 10612 4765
rect 10642 4837 10744 4849
rect 10642 4803 10652 4837
rect 10686 4803 10744 4837
rect 10642 4769 10744 4803
rect 10642 4735 10652 4769
rect 10686 4765 10744 4769
rect 10774 4765 10847 4849
rect 10877 4824 10942 4849
rect 10877 4790 10891 4824
rect 10925 4790 10942 4824
rect 10877 4765 10942 4790
rect 10972 4829 11027 4849
rect 10972 4795 10983 4829
rect 11017 4795 11027 4829
rect 10972 4765 11027 4795
rect 11057 4837 11109 4849
rect 11057 4803 11067 4837
rect 11101 4803 11109 4837
rect 11057 4765 11109 4803
rect 11163 4829 11215 4843
rect 11163 4795 11171 4829
rect 11205 4795 11215 4829
rect 10686 4735 10729 4765
rect 10642 4699 10729 4735
rect 10139 4649 10193 4661
rect 11163 4761 11215 4795
rect 11163 4727 11171 4761
rect 11205 4727 11215 4761
rect 11163 4715 11215 4727
rect 11245 4813 11299 4843
rect 11245 4779 11255 4813
rect 11289 4779 11299 4813
rect 11245 4715 11299 4779
rect 11329 4829 11381 4843
rect 11329 4795 11339 4829
rect 11373 4795 11381 4829
rect 11329 4761 11381 4795
rect 11329 4727 11339 4761
rect 11373 4727 11381 4761
rect 11329 4715 11381 4727
rect 11435 4837 11487 4849
rect 11435 4803 11443 4837
rect 11477 4803 11487 4837
rect 11435 4735 11487 4803
rect 11435 4701 11443 4735
rect 11477 4701 11487 4735
rect 11435 4675 11487 4701
rect 11697 4837 11749 4849
rect 11697 4803 11707 4837
rect 11741 4803 11749 4837
rect 11697 4735 11749 4803
rect 11697 4701 11707 4735
rect 11741 4701 11749 4735
rect 11697 4675 11749 4701
rect 11803 4829 11859 4849
rect 11803 4795 11815 4829
rect 11849 4795 11859 4829
rect 11803 4761 11859 4795
rect 11803 4727 11815 4761
rect 11849 4727 11859 4761
rect 11803 4693 11859 4727
rect 11803 4659 11815 4693
rect 11849 4659 11859 4693
rect 11803 4649 11859 4659
rect 11889 4837 12020 4849
rect 11889 4803 11901 4837
rect 11935 4803 11975 4837
rect 12009 4803 12020 4837
rect 11889 4769 12020 4803
rect 11889 4735 11901 4769
rect 11935 4735 11975 4769
rect 12009 4735 12020 4769
rect 11889 4649 12020 4735
rect 12050 4837 12128 4849
rect 12050 4803 12075 4837
rect 12109 4803 12128 4837
rect 12050 4769 12128 4803
rect 12050 4735 12075 4769
rect 12109 4735 12128 4769
rect 12050 4701 12128 4735
rect 12050 4667 12075 4701
rect 12109 4667 12128 4701
rect 12050 4649 12128 4667
rect 12158 4649 12219 4849
rect 12249 4837 12301 4849
rect 12249 4803 12259 4837
rect 12293 4803 12301 4837
rect 12249 4769 12301 4803
rect 12249 4735 12259 4769
rect 12293 4735 12301 4769
rect 12249 4649 12301 4735
rect 12355 4837 12407 4849
rect 12355 4803 12363 4837
rect 12397 4803 12407 4837
rect 12355 4735 12407 4803
rect 12355 4701 12363 4735
rect 12397 4701 12407 4735
rect 12355 4675 12407 4701
rect 12617 4837 12669 4849
rect 12617 4803 12627 4837
rect 12661 4803 12669 4837
rect 12617 4735 12669 4803
rect 12617 4701 12627 4735
rect 12661 4701 12669 4735
rect 12617 4675 12669 4701
rect 12723 4829 12779 4849
rect 12723 4795 12735 4829
rect 12769 4795 12779 4829
rect 12723 4761 12779 4795
rect 12723 4727 12735 4761
rect 12769 4727 12779 4761
rect 12723 4693 12779 4727
rect 12723 4659 12735 4693
rect 12769 4659 12779 4693
rect 12723 4649 12779 4659
rect 12809 4837 12940 4849
rect 12809 4803 12821 4837
rect 12855 4803 12895 4837
rect 12929 4803 12940 4837
rect 12809 4769 12940 4803
rect 12809 4735 12821 4769
rect 12855 4735 12895 4769
rect 12929 4735 12940 4769
rect 12809 4649 12940 4735
rect 12970 4837 13048 4849
rect 12970 4803 12995 4837
rect 13029 4803 13048 4837
rect 12970 4769 13048 4803
rect 12970 4735 12995 4769
rect 13029 4735 13048 4769
rect 12970 4701 13048 4735
rect 12970 4667 12995 4701
rect 13029 4667 13048 4701
rect 12970 4649 13048 4667
rect 13078 4649 13139 4849
rect 13169 4837 13221 4849
rect 13169 4803 13179 4837
rect 13213 4803 13221 4837
rect 13169 4769 13221 4803
rect 13169 4735 13179 4769
rect 13213 4735 13221 4769
rect 13169 4649 13221 4735
rect 13275 4837 13327 4849
rect 13275 4803 13283 4837
rect 13317 4803 13327 4837
rect 13275 4735 13327 4803
rect 13275 4701 13283 4735
rect 13317 4701 13327 4735
rect 13275 4675 13327 4701
rect 13905 4837 13957 4849
rect 13905 4803 13915 4837
rect 13949 4803 13957 4837
rect 14103 4837 14155 4849
rect 13905 4735 13957 4803
rect 13905 4701 13915 4735
rect 13949 4701 13957 4735
rect 13905 4675 13957 4701
rect 14103 4803 14111 4837
rect 14145 4803 14155 4837
rect 14103 4742 14155 4803
rect 14103 4708 14111 4742
rect 14145 4708 14155 4742
rect 14103 4675 14155 4708
rect 14273 4837 14325 4849
rect 14273 4803 14283 4837
rect 14317 4803 14325 4837
rect 14607 4837 14659 4849
rect 14607 4807 14615 4837
rect 14273 4742 14325 4803
rect 14273 4708 14283 4742
rect 14317 4708 14325 4742
rect 14411 4795 14467 4807
rect 14411 4761 14423 4795
rect 14457 4761 14467 4795
rect 14411 4723 14467 4761
rect 14497 4795 14551 4807
rect 14497 4761 14507 4795
rect 14541 4761 14551 4795
rect 14497 4723 14551 4761
rect 14581 4803 14615 4807
rect 14649 4803 14659 4837
rect 14581 4769 14659 4803
rect 14581 4735 14615 4769
rect 14649 4735 14659 4769
rect 14581 4723 14659 4735
rect 14273 4675 14325 4708
rect 14597 4649 14659 4723
rect 14689 4837 14784 4849
rect 14689 4803 14719 4837
rect 14753 4803 14784 4837
rect 14689 4769 14784 4803
rect 14689 4735 14719 4769
rect 14753 4735 14784 4769
rect 14689 4649 14784 4735
rect 14839 4837 14891 4849
rect 14839 4803 14847 4837
rect 14881 4803 14891 4837
rect 14839 4675 14891 4803
rect 15837 4837 15889 4849
rect 15837 4803 15847 4837
rect 15881 4803 15889 4837
rect 15837 4675 15889 4803
rect 15943 4837 15995 4849
rect 15943 4803 15951 4837
rect 15985 4803 15995 4837
rect 15943 4675 15995 4803
rect 16941 4837 16993 4849
rect 16941 4803 16951 4837
rect 16985 4803 16993 4837
rect 16941 4675 16993 4803
rect 17047 4837 17099 4849
rect 17047 4803 17055 4837
rect 17089 4803 17099 4837
rect 17047 4675 17099 4803
rect 18045 4837 18097 4849
rect 18045 4803 18055 4837
rect 18089 4803 18097 4837
rect 18045 4675 18097 4803
rect 18151 4837 18203 4849
rect 18151 4803 18159 4837
rect 18193 4803 18203 4837
rect 18151 4735 18203 4803
rect 18151 4701 18159 4735
rect 18193 4701 18203 4735
rect 18151 4675 18203 4701
rect 18413 4837 18465 4849
rect 18413 4803 18423 4837
rect 18457 4803 18465 4837
rect 18413 4735 18465 4803
rect 18413 4701 18423 4735
rect 18457 4701 18465 4735
rect 18413 4675 18465 4701
rect 18611 4837 18663 4849
rect 18611 4803 18619 4837
rect 18653 4803 18663 4837
rect 18611 4742 18663 4803
rect 18611 4708 18619 4742
rect 18653 4708 18663 4742
rect 18611 4675 18663 4708
rect 18781 4837 18833 4849
rect 18781 4803 18791 4837
rect 18825 4803 18833 4837
rect 18781 4742 18833 4803
rect 18781 4708 18791 4742
rect 18825 4708 18833 4742
rect 18781 4675 18833 4708
rect 1131 3996 1183 4029
rect 1131 3962 1139 3996
rect 1173 3962 1183 3996
rect 1131 3901 1183 3962
rect 1131 3867 1139 3901
rect 1173 3867 1183 3901
rect 1131 3855 1183 3867
rect 1301 3996 1353 4029
rect 1301 3962 1311 3996
rect 1345 3962 1353 3996
rect 1301 3901 1353 3962
rect 1301 3867 1311 3901
rect 1345 3867 1353 3901
rect 1301 3855 1353 3867
rect 1407 4003 1459 4029
rect 1407 3969 1415 4003
rect 1449 3969 1459 4003
rect 1407 3901 1459 3969
rect 1407 3867 1415 3901
rect 1449 3867 1459 3901
rect 1407 3855 1459 3867
rect 1853 4003 1905 4029
rect 2613 4043 2665 4055
rect 1853 3969 1863 4003
rect 1897 3969 1905 4003
rect 1853 3901 1905 3969
rect 1853 3867 1863 3901
rect 1897 3867 1905 3901
rect 1853 3855 1905 3867
rect 1959 3977 2011 4013
rect 1959 3943 1967 3977
rect 2001 3943 2011 3977
rect 1959 3909 2011 3943
rect 1959 3875 1967 3909
rect 2001 3875 2011 3909
rect 1959 3855 2011 3875
rect 2041 3977 2099 4013
rect 2041 3943 2053 3977
rect 2087 3943 2099 3977
rect 2041 3909 2099 3943
rect 2041 3875 2053 3909
rect 2087 3875 2099 3909
rect 2041 3855 2099 3875
rect 2129 3990 2181 4013
rect 2129 3956 2139 3990
rect 2173 3956 2181 3990
rect 2129 3909 2181 3956
rect 2129 3875 2139 3909
rect 2173 3875 2181 3909
rect 2129 3855 2181 3875
rect 2235 4003 2287 4029
rect 2235 3969 2243 4003
rect 2277 3969 2287 4003
rect 2235 3901 2287 3969
rect 2235 3867 2243 3901
rect 2277 3867 2287 3901
rect 2235 3855 2287 3867
rect 2497 4003 2549 4029
rect 2497 3969 2507 4003
rect 2541 3969 2549 4003
rect 2497 3901 2549 3969
rect 2497 3867 2507 3901
rect 2541 3867 2549 3901
rect 2497 3855 2549 3867
rect 2613 4009 2621 4043
rect 2655 4009 2665 4043
rect 2613 3975 2665 4009
rect 2613 3941 2621 3975
rect 2655 3941 2665 3975
rect 2613 3907 2665 3941
rect 2613 3873 2621 3907
rect 2655 3873 2665 3907
rect 2613 3855 2665 3873
rect 2695 4011 2749 4055
rect 2695 3977 2705 4011
rect 2739 3977 2749 4011
rect 2695 3931 2749 3977
rect 2695 3897 2705 3931
rect 2739 3897 2749 3931
rect 2695 3855 2749 3897
rect 2779 4043 2833 4055
rect 2779 4009 2791 4043
rect 2825 4009 2833 4043
rect 2779 3972 2833 4009
rect 2779 3938 2791 3972
rect 2825 3938 2833 3972
rect 3202 3939 3252 4005
rect 2779 3901 2833 3938
rect 2779 3867 2791 3901
rect 2825 3867 2833 3901
rect 2779 3855 2833 3867
rect 2906 3909 2959 3939
rect 2906 3875 2914 3909
rect 2948 3875 2959 3909
rect 2906 3855 2959 3875
rect 2989 3855 3073 3939
rect 3103 3919 3157 3939
rect 3103 3885 3113 3919
rect 3147 3885 3157 3919
rect 3103 3855 3157 3885
rect 3187 3909 3252 3939
rect 3187 3875 3208 3909
rect 3242 3875 3252 3909
rect 3187 3855 3252 3875
rect 3282 3969 3369 4005
rect 3282 3935 3292 3969
rect 3326 3939 3369 3969
rect 4637 4043 4689 4055
rect 4075 4003 4127 4029
rect 3803 3977 3855 3989
rect 3803 3943 3811 3977
rect 3845 3943 3855 3977
rect 3326 3935 3384 3939
rect 3282 3901 3384 3935
rect 3282 3867 3292 3901
rect 3326 3867 3384 3901
rect 3282 3855 3384 3867
rect 3414 3855 3487 3939
rect 3517 3914 3582 3939
rect 3517 3880 3531 3914
rect 3565 3880 3582 3914
rect 3517 3855 3582 3880
rect 3612 3909 3667 3939
rect 3612 3875 3623 3909
rect 3657 3875 3667 3909
rect 3612 3855 3667 3875
rect 3697 3901 3749 3939
rect 3697 3867 3707 3901
rect 3741 3867 3749 3901
rect 3697 3855 3749 3867
rect 3803 3909 3855 3943
rect 3803 3875 3811 3909
rect 3845 3875 3855 3909
rect 3803 3861 3855 3875
rect 3885 3925 3939 3989
rect 3885 3891 3895 3925
rect 3929 3891 3939 3925
rect 3885 3861 3939 3891
rect 3969 3977 4021 3989
rect 3969 3943 3979 3977
rect 4013 3943 4021 3977
rect 3969 3909 4021 3943
rect 3969 3875 3979 3909
rect 4013 3875 4021 3909
rect 3969 3861 4021 3875
rect 4075 3969 4083 4003
rect 4117 3969 4127 4003
rect 4075 3901 4127 3969
rect 4075 3867 4083 3901
rect 4117 3867 4127 3901
rect 4075 3855 4127 3867
rect 4521 4003 4573 4029
rect 4521 3969 4531 4003
rect 4565 3969 4573 4003
rect 4521 3901 4573 3969
rect 4521 3867 4531 3901
rect 4565 3867 4573 3901
rect 4521 3855 4573 3867
rect 4637 4009 4645 4043
rect 4679 4009 4689 4043
rect 4637 3975 4689 4009
rect 4637 3941 4645 3975
rect 4679 3941 4689 3975
rect 4637 3907 4689 3941
rect 4637 3873 4645 3907
rect 4679 3873 4689 3907
rect 4637 3855 4689 3873
rect 4719 4011 4773 4055
rect 4719 3977 4729 4011
rect 4763 3977 4773 4011
rect 4719 3931 4773 3977
rect 4719 3897 4729 3931
rect 4763 3897 4773 3931
rect 4719 3855 4773 3897
rect 4803 4043 4857 4055
rect 4803 4009 4815 4043
rect 4849 4009 4857 4043
rect 4803 3972 4857 4009
rect 4803 3938 4815 3972
rect 4849 3938 4857 3972
rect 5226 3939 5276 4005
rect 4803 3901 4857 3938
rect 4803 3867 4815 3901
rect 4849 3867 4857 3901
rect 4803 3855 4857 3867
rect 4930 3909 4983 3939
rect 4930 3875 4938 3909
rect 4972 3875 4983 3909
rect 4930 3855 4983 3875
rect 5013 3855 5097 3939
rect 5127 3919 5181 3939
rect 5127 3885 5137 3919
rect 5171 3885 5181 3919
rect 5127 3855 5181 3885
rect 5211 3909 5276 3939
rect 5211 3875 5232 3909
rect 5266 3875 5276 3909
rect 5211 3855 5276 3875
rect 5306 3969 5393 4005
rect 5306 3935 5316 3969
rect 5350 3939 5393 3969
rect 6927 4045 6983 4055
rect 5827 3977 5879 3989
rect 5827 3943 5835 3977
rect 5869 3943 5879 3977
rect 5350 3935 5408 3939
rect 5306 3901 5408 3935
rect 5306 3867 5316 3901
rect 5350 3867 5408 3901
rect 5306 3855 5408 3867
rect 5438 3855 5511 3939
rect 5541 3914 5606 3939
rect 5541 3880 5555 3914
rect 5589 3880 5606 3914
rect 5541 3855 5606 3880
rect 5636 3909 5691 3939
rect 5636 3875 5647 3909
rect 5681 3875 5691 3909
rect 5636 3855 5691 3875
rect 5721 3901 5773 3939
rect 5721 3867 5731 3901
rect 5765 3867 5773 3901
rect 5721 3855 5773 3867
rect 5827 3909 5879 3943
rect 5827 3875 5835 3909
rect 5869 3875 5879 3909
rect 5827 3861 5879 3875
rect 5909 3925 5963 3989
rect 5909 3891 5919 3925
rect 5953 3891 5963 3925
rect 5909 3861 5963 3891
rect 5993 3977 6045 3989
rect 5993 3943 6003 3977
rect 6037 3943 6045 3977
rect 5993 3909 6045 3943
rect 5993 3875 6003 3909
rect 6037 3875 6045 3909
rect 5993 3861 6045 3875
rect 6375 4003 6427 4029
rect 6375 3969 6383 4003
rect 6417 3969 6427 4003
rect 6375 3901 6427 3969
rect 6375 3867 6383 3901
rect 6417 3867 6427 3901
rect 6375 3855 6427 3867
rect 6821 4003 6873 4029
rect 6821 3969 6831 4003
rect 6865 3969 6873 4003
rect 6821 3901 6873 3969
rect 6821 3867 6831 3901
rect 6865 3867 6873 3901
rect 6821 3855 6873 3867
rect 6927 4011 6939 4045
rect 6973 4011 6983 4045
rect 6927 3977 6983 4011
rect 6927 3943 6939 3977
rect 6973 3943 6983 3977
rect 6927 3909 6983 3943
rect 6927 3875 6939 3909
rect 6973 3875 6983 3909
rect 6927 3855 6983 3875
rect 7013 3969 7144 4055
rect 7013 3935 7025 3969
rect 7059 3935 7099 3969
rect 7133 3935 7144 3969
rect 7013 3901 7144 3935
rect 7013 3867 7025 3901
rect 7059 3867 7099 3901
rect 7133 3867 7144 3901
rect 7013 3855 7144 3867
rect 7174 4037 7252 4055
rect 7174 4003 7199 4037
rect 7233 4003 7252 4037
rect 7174 3969 7252 4003
rect 7174 3935 7199 3969
rect 7233 3935 7252 3969
rect 7174 3901 7252 3935
rect 7174 3867 7199 3901
rect 7233 3867 7252 3901
rect 7174 3855 7252 3867
rect 7282 3855 7343 4055
rect 7373 3969 7425 4055
rect 7373 3935 7383 3969
rect 7417 3935 7425 3969
rect 7373 3901 7425 3935
rect 7373 3867 7383 3901
rect 7417 3867 7425 3901
rect 7373 3855 7425 3867
rect 7479 4003 7531 4029
rect 7479 3969 7487 4003
rect 7521 3969 7531 4003
rect 7479 3901 7531 3969
rect 7479 3867 7487 3901
rect 7521 3867 7531 3901
rect 7479 3855 7531 3867
rect 7741 4003 7793 4029
rect 7741 3969 7751 4003
rect 7785 3969 7793 4003
rect 7741 3901 7793 3969
rect 7741 3867 7751 3901
rect 7785 3867 7793 3901
rect 7741 3855 7793 3867
rect 7847 3969 7900 4055
rect 7847 3935 7855 3969
rect 7889 3935 7900 3969
rect 7847 3901 7900 3935
rect 7847 3867 7855 3901
rect 7889 3867 7900 3901
rect 7847 3855 7900 3867
rect 7930 3977 7986 4055
rect 7930 3943 7941 3977
rect 7975 3943 7986 3977
rect 7930 3909 7986 3943
rect 7930 3875 7941 3909
rect 7975 3875 7986 3909
rect 7930 3855 7986 3875
rect 8016 3969 8072 4055
rect 8016 3935 8027 3969
rect 8061 3935 8072 3969
rect 8016 3901 8072 3935
rect 8016 3867 8027 3901
rect 8061 3867 8072 3901
rect 8016 3855 8072 3867
rect 8102 3985 8158 4055
rect 8102 3951 8113 3985
rect 8147 3951 8158 3985
rect 8102 3917 8158 3951
rect 8102 3883 8113 3917
rect 8147 3883 8158 3917
rect 8102 3855 8158 3883
rect 8188 3969 8244 4055
rect 8188 3935 8199 3969
rect 8233 3935 8244 3969
rect 8188 3901 8244 3935
rect 8188 3867 8199 3901
rect 8233 3867 8244 3901
rect 8188 3855 8244 3867
rect 8274 4031 8330 4055
rect 8274 3997 8285 4031
rect 8319 3997 8330 4031
rect 8274 3945 8330 3997
rect 8274 3911 8285 3945
rect 8319 3911 8330 3945
rect 8274 3855 8330 3911
rect 8360 3925 8416 4055
rect 8360 3891 8371 3925
rect 8405 3891 8416 3925
rect 8360 3855 8416 3891
rect 8446 4031 8502 4055
rect 8446 3997 8457 4031
rect 8491 3997 8502 4031
rect 8446 3945 8502 3997
rect 8446 3911 8457 3945
rect 8491 3911 8502 3945
rect 8446 3855 8502 3911
rect 8532 3925 8588 4055
rect 8532 3891 8543 3925
rect 8577 3891 8588 3925
rect 8532 3855 8588 3891
rect 8618 4031 8674 4055
rect 8618 3997 8629 4031
rect 8663 3997 8674 4031
rect 8618 3945 8674 3997
rect 8618 3911 8629 3945
rect 8663 3911 8674 3945
rect 8618 3855 8674 3911
rect 8704 3925 8760 4055
rect 8704 3891 8715 3925
rect 8749 3891 8760 3925
rect 8704 3855 8760 3891
rect 8790 4031 8846 4055
rect 8790 3997 8801 4031
rect 8835 3997 8846 4031
rect 8790 3945 8846 3997
rect 8790 3911 8801 3945
rect 8835 3911 8846 3945
rect 8790 3855 8846 3911
rect 8876 3925 8931 4055
rect 8876 3891 8887 3925
rect 8921 3891 8931 3925
rect 8876 3855 8931 3891
rect 8961 4031 9017 4055
rect 8961 3997 8972 4031
rect 9006 3997 9017 4031
rect 8961 3945 9017 3997
rect 8961 3911 8972 3945
rect 9006 3911 9017 3945
rect 8961 3855 9017 3911
rect 9047 3925 9103 4055
rect 9047 3891 9058 3925
rect 9092 3891 9103 3925
rect 9047 3855 9103 3891
rect 9133 4031 9189 4055
rect 9133 3997 9144 4031
rect 9178 3997 9189 4031
rect 9133 3945 9189 3997
rect 9133 3911 9144 3945
rect 9178 3911 9189 3945
rect 9133 3855 9189 3911
rect 9219 3925 9275 4055
rect 9219 3891 9230 3925
rect 9264 3891 9275 3925
rect 9219 3855 9275 3891
rect 9305 4031 9361 4055
rect 9305 3997 9316 4031
rect 9350 3997 9361 4031
rect 9305 3945 9361 3997
rect 9305 3911 9316 3945
rect 9350 3911 9361 3945
rect 9305 3855 9361 3911
rect 9391 3925 9447 4055
rect 9391 3891 9402 3925
rect 9436 3891 9447 3925
rect 9391 3855 9447 3891
rect 9477 4031 9533 4055
rect 9477 3997 9488 4031
rect 9522 3997 9533 4031
rect 9477 3945 9533 3997
rect 9477 3911 9488 3945
rect 9522 3911 9533 3945
rect 9477 3855 9533 3911
rect 9563 3925 9616 4055
rect 10515 4045 10571 4055
rect 9563 3891 9574 3925
rect 9608 3891 9616 3925
rect 9563 3855 9616 3891
rect 9687 4003 9739 4029
rect 9687 3969 9695 4003
rect 9729 3969 9739 4003
rect 9687 3901 9739 3969
rect 9687 3867 9695 3901
rect 9729 3867 9739 3901
rect 9687 3855 9739 3867
rect 10317 4003 10369 4029
rect 10317 3969 10327 4003
rect 10361 3969 10369 4003
rect 10317 3901 10369 3969
rect 10317 3867 10327 3901
rect 10361 3867 10369 3901
rect 10317 3855 10369 3867
rect 10515 4011 10527 4045
rect 10561 4011 10571 4045
rect 10515 3977 10571 4011
rect 10515 3943 10527 3977
rect 10561 3943 10571 3977
rect 10515 3909 10571 3943
rect 10515 3875 10527 3909
rect 10561 3875 10571 3909
rect 10515 3855 10571 3875
rect 10601 3969 10732 4055
rect 10601 3935 10613 3969
rect 10647 3935 10687 3969
rect 10721 3935 10732 3969
rect 10601 3901 10732 3935
rect 10601 3867 10613 3901
rect 10647 3867 10687 3901
rect 10721 3867 10732 3901
rect 10601 3855 10732 3867
rect 10762 4037 10840 4055
rect 10762 4003 10787 4037
rect 10821 4003 10840 4037
rect 10762 3969 10840 4003
rect 10762 3935 10787 3969
rect 10821 3935 10840 3969
rect 10762 3901 10840 3935
rect 10762 3867 10787 3901
rect 10821 3867 10840 3901
rect 10762 3855 10840 3867
rect 10870 3855 10931 4055
rect 10961 3969 11013 4055
rect 10961 3935 10971 3969
rect 11005 3935 11013 3969
rect 10961 3901 11013 3935
rect 10961 3867 10971 3901
rect 11005 3867 11013 3901
rect 10961 3855 11013 3867
rect 11067 4003 11119 4029
rect 11067 3969 11075 4003
rect 11109 3969 11119 4003
rect 11067 3901 11119 3969
rect 11067 3867 11075 3901
rect 11109 3867 11119 3901
rect 11067 3855 11119 3867
rect 11329 4003 11381 4029
rect 11329 3969 11339 4003
rect 11373 3969 11381 4003
rect 11329 3901 11381 3969
rect 11329 3867 11339 3901
rect 11373 3867 11381 3901
rect 11711 3977 11763 3989
rect 11711 3943 11719 3977
rect 11753 3943 11763 3977
rect 11711 3909 11763 3943
rect 11711 3875 11719 3909
rect 11753 3875 11763 3909
rect 11329 3855 11381 3867
rect 11711 3861 11763 3875
rect 11793 3925 11847 3989
rect 11793 3891 11803 3925
rect 11837 3891 11847 3925
rect 11793 3861 11847 3891
rect 11877 3977 11929 3989
rect 11877 3943 11887 3977
rect 11921 3943 11929 3977
rect 11877 3909 11929 3943
rect 12899 4043 12953 4055
rect 12363 3969 12450 4005
rect 12363 3939 12406 3969
rect 11877 3875 11887 3909
rect 11921 3875 11929 3909
rect 11877 3861 11929 3875
rect 11983 3901 12035 3939
rect 11983 3867 11991 3901
rect 12025 3867 12035 3901
rect 11983 3855 12035 3867
rect 12065 3909 12120 3939
rect 12065 3875 12075 3909
rect 12109 3875 12120 3909
rect 12065 3855 12120 3875
rect 12150 3914 12215 3939
rect 12150 3880 12167 3914
rect 12201 3880 12215 3914
rect 12150 3855 12215 3880
rect 12245 3855 12318 3939
rect 12348 3935 12406 3939
rect 12440 3935 12450 3969
rect 12348 3901 12450 3935
rect 12348 3867 12406 3901
rect 12440 3867 12450 3901
rect 12348 3855 12450 3867
rect 12480 3939 12530 4005
rect 12899 4009 12907 4043
rect 12941 4009 12953 4043
rect 12899 3972 12953 4009
rect 12480 3909 12545 3939
rect 12480 3875 12490 3909
rect 12524 3875 12545 3909
rect 12480 3855 12545 3875
rect 12575 3919 12629 3939
rect 12575 3885 12585 3919
rect 12619 3885 12629 3919
rect 12575 3855 12629 3885
rect 12659 3855 12743 3939
rect 12773 3909 12826 3939
rect 12773 3875 12784 3909
rect 12818 3875 12826 3909
rect 12773 3855 12826 3875
rect 12899 3938 12907 3972
rect 12941 3938 12953 3972
rect 12899 3901 12953 3938
rect 12899 3867 12907 3901
rect 12941 3867 12953 3901
rect 12899 3855 12953 3867
rect 12983 4011 13037 4055
rect 12983 3977 12993 4011
rect 13027 3977 13037 4011
rect 12983 3931 13037 3977
rect 12983 3897 12993 3931
rect 13027 3897 13037 3931
rect 12983 3855 13037 3897
rect 13067 4043 13119 4055
rect 13067 4009 13077 4043
rect 13111 4009 13119 4043
rect 13067 3975 13119 4009
rect 13067 3941 13077 3975
rect 13111 3941 13119 3975
rect 13067 3907 13119 3941
rect 13067 3873 13077 3907
rect 13111 3873 13119 3907
rect 13067 3855 13119 3873
rect 13183 3901 13235 4029
rect 13183 3867 13191 3901
rect 13225 3867 13235 3901
rect 13183 3855 13235 3867
rect 14181 3901 14233 4029
rect 14181 3867 14191 3901
rect 14225 3867 14233 3901
rect 14181 3855 14233 3867
rect 14287 3901 14339 4029
rect 14287 3867 14295 3901
rect 14329 3867 14339 3901
rect 14287 3855 14339 3867
rect 15285 3901 15337 4029
rect 15285 3867 15295 3901
rect 15329 3867 15337 3901
rect 15285 3855 15337 3867
rect 15483 3990 15535 4013
rect 15483 3956 15491 3990
rect 15525 3956 15535 3990
rect 15483 3909 15535 3956
rect 15483 3875 15491 3909
rect 15525 3875 15535 3909
rect 15483 3855 15535 3875
rect 15565 3977 15623 4013
rect 15565 3943 15577 3977
rect 15611 3943 15623 3977
rect 15565 3909 15623 3943
rect 15565 3875 15577 3909
rect 15611 3875 15623 3909
rect 15565 3855 15623 3875
rect 15653 3977 15705 4013
rect 15653 3943 15663 3977
rect 15697 3943 15705 3977
rect 15653 3909 15705 3943
rect 15653 3875 15663 3909
rect 15697 3875 15705 3909
rect 15653 3855 15705 3875
rect 15759 4003 15811 4029
rect 15759 3969 15767 4003
rect 15801 3969 15811 4003
rect 15759 3901 15811 3969
rect 15759 3867 15767 3901
rect 15801 3867 15811 3901
rect 15759 3855 15811 3867
rect 16389 4003 16441 4029
rect 16389 3969 16399 4003
rect 16433 3969 16441 4003
rect 16389 3901 16441 3969
rect 16389 3867 16399 3901
rect 16433 3867 16441 3901
rect 17081 3981 17143 4055
rect 16895 3943 16951 3981
rect 16895 3909 16907 3943
rect 16941 3909 16951 3943
rect 16895 3897 16951 3909
rect 16981 3943 17035 3981
rect 16981 3909 16991 3943
rect 17025 3909 17035 3943
rect 16981 3897 17035 3909
rect 17065 3969 17143 3981
rect 17065 3935 17099 3969
rect 17133 3935 17143 3969
rect 17065 3901 17143 3935
rect 17065 3897 17099 3901
rect 16389 3855 16441 3867
rect 17091 3867 17099 3897
rect 17133 3867 17143 3901
rect 17091 3855 17143 3867
rect 17173 3969 17268 4055
rect 17173 3935 17203 3969
rect 17237 3935 17268 3969
rect 17173 3901 17268 3935
rect 17173 3867 17203 3901
rect 17237 3867 17268 3901
rect 17173 3855 17268 3867
rect 17323 3901 17375 4029
rect 17323 3867 17331 3901
rect 17365 3867 17375 3901
rect 17323 3855 17375 3867
rect 18321 3901 18373 4029
rect 18321 3867 18331 3901
rect 18365 3867 18373 3901
rect 18321 3855 18373 3867
rect 18611 3996 18663 4029
rect 18611 3962 18619 3996
rect 18653 3962 18663 3996
rect 18611 3901 18663 3962
rect 18611 3867 18619 3901
rect 18653 3867 18663 3901
rect 18611 3855 18663 3867
rect 18781 3996 18833 4029
rect 18781 3962 18791 3996
rect 18825 3962 18833 3996
rect 18781 3901 18833 3962
rect 18781 3867 18791 3901
rect 18825 3867 18833 3901
rect 18781 3855 18833 3867
rect 1131 3749 1183 3761
rect 1131 3715 1139 3749
rect 1173 3715 1183 3749
rect 1131 3654 1183 3715
rect 1131 3620 1139 3654
rect 1173 3620 1183 3654
rect 1131 3587 1183 3620
rect 1301 3749 1353 3761
rect 1301 3715 1311 3749
rect 1345 3715 1353 3749
rect 1301 3654 1353 3715
rect 1301 3620 1311 3654
rect 1345 3620 1353 3654
rect 1301 3587 1353 3620
rect 1407 3749 1459 3761
rect 1407 3715 1415 3749
rect 1449 3715 1459 3749
rect 1407 3647 1459 3715
rect 1407 3613 1415 3647
rect 1449 3613 1459 3647
rect 1407 3587 1459 3613
rect 1853 3749 1905 3761
rect 1853 3715 1863 3749
rect 1897 3715 1905 3749
rect 1853 3647 1905 3715
rect 1853 3613 1863 3647
rect 1897 3613 1905 3647
rect 2051 3741 2103 3755
rect 2051 3707 2059 3741
rect 2093 3707 2103 3741
rect 2051 3673 2103 3707
rect 2051 3639 2059 3673
rect 2093 3639 2103 3673
rect 2051 3627 2103 3639
rect 2133 3725 2187 3755
rect 2133 3691 2143 3725
rect 2177 3691 2187 3725
rect 2133 3627 2187 3691
rect 2217 3741 2269 3755
rect 2217 3707 2227 3741
rect 2261 3707 2269 3741
rect 2217 3673 2269 3707
rect 2323 3749 2375 3761
rect 2323 3715 2331 3749
rect 2365 3715 2375 3749
rect 2323 3677 2375 3715
rect 2405 3741 2460 3761
rect 2405 3707 2415 3741
rect 2449 3707 2460 3741
rect 2405 3677 2460 3707
rect 2490 3736 2555 3761
rect 2490 3702 2507 3736
rect 2541 3702 2555 3736
rect 2490 3677 2555 3702
rect 2585 3677 2658 3761
rect 2688 3749 2790 3761
rect 2688 3715 2746 3749
rect 2780 3715 2790 3749
rect 2688 3681 2790 3715
rect 2688 3677 2746 3681
rect 2217 3639 2227 3673
rect 2261 3639 2269 3673
rect 2217 3627 2269 3639
rect 1853 3587 1905 3613
rect 2703 3647 2746 3677
rect 2780 3647 2790 3681
rect 2703 3611 2790 3647
rect 2820 3741 2885 3761
rect 2820 3707 2830 3741
rect 2864 3707 2885 3741
rect 2820 3677 2885 3707
rect 2915 3731 2969 3761
rect 2915 3697 2925 3731
rect 2959 3697 2969 3731
rect 2915 3677 2969 3697
rect 2999 3677 3083 3761
rect 3113 3741 3166 3761
rect 3113 3707 3124 3741
rect 3158 3707 3166 3741
rect 3113 3677 3166 3707
rect 3239 3749 3293 3761
rect 3239 3715 3247 3749
rect 3281 3715 3293 3749
rect 3239 3678 3293 3715
rect 2820 3611 2870 3677
rect 3239 3644 3247 3678
rect 3281 3644 3293 3678
rect 3239 3607 3293 3644
rect 3239 3573 3247 3607
rect 3281 3573 3293 3607
rect 3239 3561 3293 3573
rect 3323 3719 3377 3761
rect 3323 3685 3333 3719
rect 3367 3685 3377 3719
rect 3323 3639 3377 3685
rect 3323 3605 3333 3639
rect 3367 3605 3377 3639
rect 3323 3561 3377 3605
rect 3407 3743 3459 3761
rect 3407 3709 3417 3743
rect 3451 3709 3459 3743
rect 3407 3675 3459 3709
rect 3407 3641 3417 3675
rect 3451 3641 3459 3675
rect 3407 3607 3459 3641
rect 3407 3573 3417 3607
rect 3451 3573 3459 3607
rect 3407 3561 3459 3573
rect 3983 3741 4035 3755
rect 3983 3707 3991 3741
rect 4025 3707 4035 3741
rect 3983 3673 4035 3707
rect 3983 3639 3991 3673
rect 4025 3639 4035 3673
rect 3983 3627 4035 3639
rect 4065 3725 4119 3755
rect 4065 3691 4075 3725
rect 4109 3691 4119 3725
rect 4065 3627 4119 3691
rect 4149 3741 4201 3755
rect 4149 3707 4159 3741
rect 4193 3707 4201 3741
rect 4149 3673 4201 3707
rect 4255 3749 4307 3761
rect 4255 3715 4263 3749
rect 4297 3715 4307 3749
rect 4255 3677 4307 3715
rect 4337 3741 4392 3761
rect 4337 3707 4347 3741
rect 4381 3707 4392 3741
rect 4337 3677 4392 3707
rect 4422 3736 4487 3761
rect 4422 3702 4439 3736
rect 4473 3702 4487 3736
rect 4422 3677 4487 3702
rect 4517 3677 4590 3761
rect 4620 3749 4722 3761
rect 4620 3715 4678 3749
rect 4712 3715 4722 3749
rect 4620 3681 4722 3715
rect 4620 3677 4678 3681
rect 4149 3639 4159 3673
rect 4193 3639 4201 3673
rect 4149 3627 4201 3639
rect 4635 3647 4678 3677
rect 4712 3647 4722 3681
rect 4635 3611 4722 3647
rect 4752 3741 4817 3761
rect 4752 3707 4762 3741
rect 4796 3707 4817 3741
rect 4752 3677 4817 3707
rect 4847 3731 4901 3761
rect 4847 3697 4857 3731
rect 4891 3697 4901 3731
rect 4847 3677 4901 3697
rect 4931 3677 5015 3761
rect 5045 3741 5098 3761
rect 5045 3707 5056 3741
rect 5090 3707 5098 3741
rect 5045 3677 5098 3707
rect 5171 3749 5225 3761
rect 5171 3715 5179 3749
rect 5213 3715 5225 3749
rect 5171 3678 5225 3715
rect 4752 3611 4802 3677
rect 5171 3644 5179 3678
rect 5213 3644 5225 3678
rect 5171 3607 5225 3644
rect 5171 3573 5179 3607
rect 5213 3573 5225 3607
rect 5171 3561 5225 3573
rect 5255 3719 5309 3761
rect 5255 3685 5265 3719
rect 5299 3685 5309 3719
rect 5255 3639 5309 3685
rect 5255 3605 5265 3639
rect 5299 3605 5309 3639
rect 5255 3561 5309 3605
rect 5339 3743 5391 3761
rect 5339 3709 5349 3743
rect 5383 3709 5391 3743
rect 5339 3675 5391 3709
rect 5339 3641 5349 3675
rect 5383 3641 5391 3675
rect 5339 3607 5391 3641
rect 5339 3573 5349 3607
rect 5383 3573 5391 3607
rect 5455 3749 5507 3761
rect 5455 3715 5463 3749
rect 5497 3715 5507 3749
rect 5455 3647 5507 3715
rect 5455 3613 5463 3647
rect 5497 3613 5507 3647
rect 5455 3587 5507 3613
rect 6085 3749 6137 3761
rect 6085 3715 6095 3749
rect 6129 3715 6137 3749
rect 6085 3647 6137 3715
rect 6085 3613 6095 3647
rect 6129 3613 6137 3647
rect 6085 3587 6137 3613
rect 6283 3741 6339 3761
rect 6283 3707 6295 3741
rect 6329 3707 6339 3741
rect 6283 3673 6339 3707
rect 6283 3639 6295 3673
rect 6329 3639 6339 3673
rect 6283 3605 6339 3639
rect 5339 3561 5391 3573
rect 6283 3571 6295 3605
rect 6329 3571 6339 3605
rect 6283 3561 6339 3571
rect 6369 3749 6500 3761
rect 6369 3715 6381 3749
rect 6415 3715 6455 3749
rect 6489 3715 6500 3749
rect 6369 3681 6500 3715
rect 6369 3647 6381 3681
rect 6415 3647 6455 3681
rect 6489 3647 6500 3681
rect 6369 3561 6500 3647
rect 6530 3749 6608 3761
rect 6530 3715 6555 3749
rect 6589 3715 6608 3749
rect 6530 3681 6608 3715
rect 6530 3647 6555 3681
rect 6589 3647 6608 3681
rect 6530 3613 6608 3647
rect 6530 3579 6555 3613
rect 6589 3579 6608 3613
rect 6530 3561 6608 3579
rect 6638 3561 6699 3761
rect 6729 3749 6781 3761
rect 6729 3715 6739 3749
rect 6773 3715 6781 3749
rect 6729 3681 6781 3715
rect 6729 3647 6739 3681
rect 6773 3647 6781 3681
rect 6729 3561 6781 3647
rect 6835 3749 6887 3761
rect 6835 3715 6843 3749
rect 6877 3715 6887 3749
rect 6835 3647 6887 3715
rect 6835 3613 6843 3647
rect 6877 3613 6887 3647
rect 6835 3587 6887 3613
rect 7097 3749 7149 3761
rect 7097 3715 7107 3749
rect 7141 3715 7149 3749
rect 7097 3647 7149 3715
rect 7097 3613 7107 3647
rect 7141 3613 7149 3647
rect 7203 3741 7255 3755
rect 7203 3707 7211 3741
rect 7245 3707 7255 3741
rect 7203 3673 7255 3707
rect 7203 3639 7211 3673
rect 7245 3639 7255 3673
rect 7203 3627 7255 3639
rect 7285 3725 7339 3755
rect 7285 3691 7295 3725
rect 7329 3691 7339 3725
rect 7285 3627 7339 3691
rect 7369 3741 7421 3755
rect 7369 3707 7379 3741
rect 7413 3707 7421 3741
rect 7369 3673 7421 3707
rect 7475 3749 7527 3761
rect 7475 3715 7483 3749
rect 7517 3715 7527 3749
rect 7475 3677 7527 3715
rect 7557 3741 7612 3761
rect 7557 3707 7567 3741
rect 7601 3707 7612 3741
rect 7557 3677 7612 3707
rect 7642 3736 7707 3761
rect 7642 3702 7659 3736
rect 7693 3702 7707 3736
rect 7642 3677 7707 3702
rect 7737 3677 7810 3761
rect 7840 3749 7942 3761
rect 7840 3715 7898 3749
rect 7932 3715 7942 3749
rect 7840 3681 7942 3715
rect 7840 3677 7898 3681
rect 7369 3639 7379 3673
rect 7413 3639 7421 3673
rect 7369 3627 7421 3639
rect 7097 3587 7149 3613
rect 7855 3647 7898 3677
rect 7932 3647 7942 3681
rect 7855 3611 7942 3647
rect 7972 3741 8037 3761
rect 7972 3707 7982 3741
rect 8016 3707 8037 3741
rect 7972 3677 8037 3707
rect 8067 3731 8121 3761
rect 8067 3697 8077 3731
rect 8111 3697 8121 3731
rect 8067 3677 8121 3697
rect 8151 3677 8235 3761
rect 8265 3741 8318 3761
rect 8265 3707 8276 3741
rect 8310 3707 8318 3741
rect 8265 3677 8318 3707
rect 8391 3749 8445 3761
rect 8391 3715 8399 3749
rect 8433 3715 8445 3749
rect 8391 3678 8445 3715
rect 7972 3611 8022 3677
rect 8391 3644 8399 3678
rect 8433 3644 8445 3678
rect 8391 3607 8445 3644
rect 8391 3573 8399 3607
rect 8433 3573 8445 3607
rect 8391 3561 8445 3573
rect 8475 3719 8529 3761
rect 8475 3685 8485 3719
rect 8519 3685 8529 3719
rect 8475 3639 8529 3685
rect 8475 3605 8485 3639
rect 8519 3605 8529 3639
rect 8475 3561 8529 3605
rect 8559 3743 8611 3761
rect 8951 3749 9003 3761
rect 8559 3709 8569 3743
rect 8603 3709 8611 3743
rect 8559 3675 8611 3709
rect 8559 3641 8569 3675
rect 8603 3641 8611 3675
rect 8559 3607 8611 3641
rect 8559 3573 8569 3607
rect 8603 3573 8611 3607
rect 8559 3561 8611 3573
rect 8951 3715 8959 3749
rect 8993 3715 9003 3749
rect 8951 3647 9003 3715
rect 8951 3613 8959 3647
rect 8993 3613 9003 3647
rect 8951 3587 9003 3613
rect 9581 3749 9633 3761
rect 9581 3715 9591 3749
rect 9625 3715 9633 3749
rect 9581 3647 9633 3715
rect 9581 3613 9591 3647
rect 9625 3613 9633 3647
rect 9779 3741 9831 3755
rect 9779 3707 9787 3741
rect 9821 3707 9831 3741
rect 9779 3673 9831 3707
rect 9779 3639 9787 3673
rect 9821 3639 9831 3673
rect 9779 3627 9831 3639
rect 9861 3725 9915 3755
rect 9861 3691 9871 3725
rect 9905 3691 9915 3725
rect 9861 3627 9915 3691
rect 9945 3741 9997 3755
rect 9945 3707 9955 3741
rect 9989 3707 9997 3741
rect 9945 3673 9997 3707
rect 10051 3749 10103 3761
rect 10051 3715 10059 3749
rect 10093 3715 10103 3749
rect 10051 3677 10103 3715
rect 10133 3741 10188 3761
rect 10133 3707 10143 3741
rect 10177 3707 10188 3741
rect 10133 3677 10188 3707
rect 10218 3736 10283 3761
rect 10218 3702 10235 3736
rect 10269 3702 10283 3736
rect 10218 3677 10283 3702
rect 10313 3677 10386 3761
rect 10416 3749 10518 3761
rect 10416 3715 10474 3749
rect 10508 3715 10518 3749
rect 10416 3681 10518 3715
rect 10416 3677 10474 3681
rect 9945 3639 9955 3673
rect 9989 3639 9997 3673
rect 9945 3627 9997 3639
rect 9581 3587 9633 3613
rect 10431 3647 10474 3677
rect 10508 3647 10518 3681
rect 10431 3611 10518 3647
rect 10548 3741 10613 3761
rect 10548 3707 10558 3741
rect 10592 3707 10613 3741
rect 10548 3677 10613 3707
rect 10643 3731 10697 3761
rect 10643 3697 10653 3731
rect 10687 3697 10697 3731
rect 10643 3677 10697 3697
rect 10727 3677 10811 3761
rect 10841 3741 10894 3761
rect 10841 3707 10852 3741
rect 10886 3707 10894 3741
rect 10841 3677 10894 3707
rect 10967 3749 11021 3761
rect 10967 3715 10975 3749
rect 11009 3715 11021 3749
rect 10967 3678 11021 3715
rect 10548 3611 10598 3677
rect 10967 3644 10975 3678
rect 11009 3644 11021 3678
rect 10967 3607 11021 3644
rect 10967 3573 10975 3607
rect 11009 3573 11021 3607
rect 10967 3561 11021 3573
rect 11051 3719 11105 3761
rect 11051 3685 11061 3719
rect 11095 3685 11105 3719
rect 11051 3639 11105 3685
rect 11051 3605 11061 3639
rect 11095 3605 11105 3639
rect 11051 3561 11105 3605
rect 11135 3743 11187 3761
rect 11135 3709 11145 3743
rect 11179 3709 11187 3743
rect 11135 3675 11187 3709
rect 11135 3641 11145 3675
rect 11179 3641 11187 3675
rect 11135 3607 11187 3641
rect 11135 3573 11145 3607
rect 11179 3573 11187 3607
rect 11251 3749 11303 3761
rect 11251 3715 11259 3749
rect 11293 3715 11303 3749
rect 11251 3647 11303 3715
rect 11251 3613 11259 3647
rect 11293 3613 11303 3647
rect 11251 3587 11303 3613
rect 11697 3749 11749 3761
rect 11697 3715 11707 3749
rect 11741 3715 11749 3749
rect 11697 3647 11749 3715
rect 11697 3613 11707 3647
rect 11741 3613 11749 3647
rect 11803 3741 11855 3755
rect 11803 3707 11811 3741
rect 11845 3707 11855 3741
rect 11803 3673 11855 3707
rect 11803 3639 11811 3673
rect 11845 3639 11855 3673
rect 11803 3627 11855 3639
rect 11885 3725 11939 3755
rect 11885 3691 11895 3725
rect 11929 3691 11939 3725
rect 11885 3627 11939 3691
rect 11969 3741 12021 3755
rect 11969 3707 11979 3741
rect 12013 3707 12021 3741
rect 11969 3673 12021 3707
rect 12075 3749 12127 3761
rect 12075 3715 12083 3749
rect 12117 3715 12127 3749
rect 12075 3677 12127 3715
rect 12157 3741 12212 3761
rect 12157 3707 12167 3741
rect 12201 3707 12212 3741
rect 12157 3677 12212 3707
rect 12242 3736 12307 3761
rect 12242 3702 12259 3736
rect 12293 3702 12307 3736
rect 12242 3677 12307 3702
rect 12337 3677 12410 3761
rect 12440 3749 12542 3761
rect 12440 3715 12498 3749
rect 12532 3715 12542 3749
rect 12440 3681 12542 3715
rect 12440 3677 12498 3681
rect 11969 3639 11979 3673
rect 12013 3639 12021 3673
rect 11969 3627 12021 3639
rect 11697 3587 11749 3613
rect 11135 3561 11187 3573
rect 12455 3647 12498 3677
rect 12532 3647 12542 3681
rect 12455 3611 12542 3647
rect 12572 3741 12637 3761
rect 12572 3707 12582 3741
rect 12616 3707 12637 3741
rect 12572 3677 12637 3707
rect 12667 3731 12721 3761
rect 12667 3697 12677 3731
rect 12711 3697 12721 3731
rect 12667 3677 12721 3697
rect 12751 3677 12835 3761
rect 12865 3741 12918 3761
rect 12865 3707 12876 3741
rect 12910 3707 12918 3741
rect 12865 3677 12918 3707
rect 12991 3749 13045 3761
rect 12991 3715 12999 3749
rect 13033 3715 13045 3749
rect 12991 3678 13045 3715
rect 12572 3611 12622 3677
rect 12991 3644 12999 3678
rect 13033 3644 13045 3678
rect 12991 3607 13045 3644
rect 12991 3573 12999 3607
rect 13033 3573 13045 3607
rect 12991 3561 13045 3573
rect 13075 3719 13129 3761
rect 13075 3685 13085 3719
rect 13119 3685 13129 3719
rect 13075 3639 13129 3685
rect 13075 3605 13085 3639
rect 13119 3605 13129 3639
rect 13075 3561 13129 3605
rect 13159 3743 13211 3761
rect 13159 3709 13169 3743
rect 13203 3709 13211 3743
rect 13159 3675 13211 3709
rect 13159 3641 13169 3675
rect 13203 3641 13211 3675
rect 13159 3607 13211 3641
rect 13159 3573 13169 3607
rect 13203 3573 13211 3607
rect 13275 3749 13327 3761
rect 13275 3715 13283 3749
rect 13317 3715 13327 3749
rect 13275 3647 13327 3715
rect 13275 3613 13283 3647
rect 13317 3613 13327 3647
rect 13275 3587 13327 3613
rect 13905 3749 13957 3761
rect 13905 3715 13915 3749
rect 13949 3715 13957 3749
rect 14103 3749 14155 3761
rect 13905 3647 13957 3715
rect 13905 3613 13915 3647
rect 13949 3613 13957 3647
rect 13905 3587 13957 3613
rect 13159 3561 13211 3573
rect 14103 3715 14111 3749
rect 14145 3715 14155 3749
rect 14103 3587 14155 3715
rect 15101 3749 15153 3761
rect 15101 3715 15111 3749
rect 15145 3715 15153 3749
rect 15101 3587 15153 3715
rect 15207 3749 15259 3761
rect 15207 3715 15215 3749
rect 15249 3715 15259 3749
rect 15207 3647 15259 3715
rect 15207 3613 15215 3647
rect 15249 3613 15259 3647
rect 15207 3587 15259 3613
rect 15653 3749 15705 3761
rect 15653 3715 15663 3749
rect 15697 3715 15705 3749
rect 15653 3647 15705 3715
rect 15653 3613 15663 3647
rect 15697 3613 15705 3647
rect 15653 3587 15705 3613
rect 15759 3741 15811 3761
rect 15759 3707 15767 3741
rect 15801 3707 15811 3741
rect 15759 3660 15811 3707
rect 15759 3626 15767 3660
rect 15801 3626 15811 3660
rect 15759 3603 15811 3626
rect 15841 3741 15899 3761
rect 15841 3707 15853 3741
rect 15887 3707 15899 3741
rect 15841 3673 15899 3707
rect 15841 3639 15853 3673
rect 15887 3639 15899 3673
rect 15841 3603 15899 3639
rect 15929 3741 15981 3761
rect 15929 3707 15939 3741
rect 15973 3707 15981 3741
rect 15929 3673 15981 3707
rect 15929 3639 15939 3673
rect 15973 3639 15981 3673
rect 15929 3603 15981 3639
rect 16035 3749 16087 3761
rect 16035 3715 16043 3749
rect 16077 3715 16087 3749
rect 16035 3647 16087 3715
rect 16035 3613 16043 3647
rect 16077 3613 16087 3647
rect 16035 3587 16087 3613
rect 16297 3749 16349 3761
rect 16297 3715 16307 3749
rect 16341 3715 16349 3749
rect 16297 3647 16349 3715
rect 16297 3613 16307 3647
rect 16341 3613 16349 3647
rect 16297 3587 16349 3613
rect 16404 3749 16499 3761
rect 16404 3715 16435 3749
rect 16469 3715 16499 3749
rect 16404 3681 16499 3715
rect 16404 3647 16435 3681
rect 16469 3647 16499 3681
rect 16404 3561 16499 3647
rect 16529 3749 16581 3761
rect 16529 3715 16539 3749
rect 16573 3719 16581 3749
rect 16863 3749 16915 3761
rect 16573 3715 16607 3719
rect 16529 3681 16607 3715
rect 16529 3647 16539 3681
rect 16573 3647 16607 3681
rect 16529 3635 16607 3647
rect 16637 3707 16691 3719
rect 16637 3673 16647 3707
rect 16681 3673 16691 3707
rect 16637 3635 16691 3673
rect 16721 3707 16777 3719
rect 16721 3673 16731 3707
rect 16765 3673 16777 3707
rect 16721 3635 16777 3673
rect 16863 3715 16871 3749
rect 16905 3715 16915 3749
rect 16863 3647 16915 3715
rect 16529 3561 16591 3635
rect 16863 3613 16871 3647
rect 16905 3613 16915 3647
rect 16863 3587 16915 3613
rect 17125 3749 17177 3761
rect 17125 3715 17135 3749
rect 17169 3715 17177 3749
rect 17125 3647 17177 3715
rect 17125 3613 17135 3647
rect 17169 3613 17177 3647
rect 17125 3587 17177 3613
rect 17232 3749 17327 3761
rect 17232 3715 17263 3749
rect 17297 3715 17327 3749
rect 17232 3681 17327 3715
rect 17232 3647 17263 3681
rect 17297 3647 17327 3681
rect 17232 3561 17327 3647
rect 17357 3749 17409 3761
rect 17357 3715 17367 3749
rect 17401 3719 17409 3749
rect 17691 3749 17743 3761
rect 17401 3715 17435 3719
rect 17357 3681 17435 3715
rect 17357 3647 17367 3681
rect 17401 3647 17435 3681
rect 17357 3635 17435 3647
rect 17465 3707 17519 3719
rect 17465 3673 17475 3707
rect 17509 3673 17519 3707
rect 17465 3635 17519 3673
rect 17549 3707 17605 3719
rect 17549 3673 17559 3707
rect 17593 3673 17605 3707
rect 17549 3635 17605 3673
rect 17691 3715 17699 3749
rect 17733 3715 17743 3749
rect 17691 3647 17743 3715
rect 17357 3561 17419 3635
rect 17691 3613 17699 3647
rect 17733 3613 17743 3647
rect 17691 3587 17743 3613
rect 18321 3749 18373 3761
rect 18321 3715 18331 3749
rect 18365 3715 18373 3749
rect 18321 3647 18373 3715
rect 18321 3613 18331 3647
rect 18365 3613 18373 3647
rect 18321 3587 18373 3613
rect 18611 3749 18663 3761
rect 18611 3715 18619 3749
rect 18653 3715 18663 3749
rect 18611 3654 18663 3715
rect 18611 3620 18619 3654
rect 18653 3620 18663 3654
rect 18611 3587 18663 3620
rect 18781 3749 18833 3761
rect 18781 3715 18791 3749
rect 18825 3715 18833 3749
rect 18781 3654 18833 3715
rect 18781 3620 18791 3654
rect 18825 3620 18833 3654
rect 18781 3587 18833 3620
rect 1131 2908 1183 2941
rect 1131 2874 1139 2908
rect 1173 2874 1183 2908
rect 1131 2813 1183 2874
rect 1131 2779 1139 2813
rect 1173 2779 1183 2813
rect 1131 2767 1183 2779
rect 1301 2908 1353 2941
rect 1301 2874 1311 2908
rect 1345 2874 1353 2908
rect 1301 2813 1353 2874
rect 1301 2779 1311 2813
rect 1345 2779 1353 2813
rect 1301 2767 1353 2779
rect 1407 2915 1459 2941
rect 1407 2881 1415 2915
rect 1449 2881 1459 2915
rect 1407 2813 1459 2881
rect 1407 2779 1415 2813
rect 1449 2779 1459 2813
rect 1407 2767 1459 2779
rect 1669 2915 1721 2941
rect 1669 2881 1679 2915
rect 1713 2881 1721 2915
rect 1669 2813 1721 2881
rect 1669 2779 1679 2813
rect 1713 2779 1721 2813
rect 1669 2767 1721 2779
rect 1867 2932 1920 2967
rect 1867 2898 1875 2932
rect 1909 2898 1920 2932
rect 1867 2827 1920 2898
rect 1867 2793 1875 2827
rect 1909 2793 1920 2827
rect 1867 2767 1920 2793
rect 1950 2893 2015 2967
rect 1950 2859 1961 2893
rect 1995 2859 2015 2893
rect 1950 2825 2015 2859
rect 1950 2791 1961 2825
rect 1995 2791 2015 2825
rect 1950 2767 2015 2791
rect 2045 2827 2099 2967
rect 2045 2793 2055 2827
rect 2089 2793 2099 2827
rect 2045 2767 2099 2793
rect 2129 2822 2181 2967
rect 2129 2788 2139 2822
rect 2173 2788 2181 2822
rect 2129 2767 2181 2788
rect 2235 2915 2287 2941
rect 2235 2881 2243 2915
rect 2277 2881 2287 2915
rect 2235 2813 2287 2881
rect 2235 2779 2243 2813
rect 2277 2779 2287 2813
rect 2235 2767 2287 2779
rect 2497 2915 2549 2941
rect 2497 2881 2507 2915
rect 2541 2881 2549 2915
rect 2497 2813 2549 2881
rect 2497 2779 2507 2813
rect 2541 2779 2549 2813
rect 2497 2767 2549 2779
rect 2620 2837 2673 2967
rect 2620 2803 2628 2837
rect 2662 2803 2673 2837
rect 2620 2767 2673 2803
rect 2703 2943 2759 2967
rect 2703 2909 2714 2943
rect 2748 2909 2759 2943
rect 2703 2857 2759 2909
rect 2703 2823 2714 2857
rect 2748 2823 2759 2857
rect 2703 2767 2759 2823
rect 2789 2837 2845 2967
rect 2789 2803 2800 2837
rect 2834 2803 2845 2837
rect 2789 2767 2845 2803
rect 2875 2943 2931 2967
rect 2875 2909 2886 2943
rect 2920 2909 2931 2943
rect 2875 2857 2931 2909
rect 2875 2823 2886 2857
rect 2920 2823 2931 2857
rect 2875 2767 2931 2823
rect 2961 2837 3017 2967
rect 2961 2803 2972 2837
rect 3006 2803 3017 2837
rect 2961 2767 3017 2803
rect 3047 2943 3103 2967
rect 3047 2909 3058 2943
rect 3092 2909 3103 2943
rect 3047 2857 3103 2909
rect 3047 2823 3058 2857
rect 3092 2823 3103 2857
rect 3047 2767 3103 2823
rect 3133 2837 3189 2967
rect 3133 2803 3144 2837
rect 3178 2803 3189 2837
rect 3133 2767 3189 2803
rect 3219 2943 3275 2967
rect 3219 2909 3230 2943
rect 3264 2909 3275 2943
rect 3219 2857 3275 2909
rect 3219 2823 3230 2857
rect 3264 2823 3275 2857
rect 3219 2767 3275 2823
rect 3305 2837 3360 2967
rect 3305 2803 3315 2837
rect 3349 2803 3360 2837
rect 3305 2767 3360 2803
rect 3390 2943 3446 2967
rect 3390 2909 3401 2943
rect 3435 2909 3446 2943
rect 3390 2857 3446 2909
rect 3390 2823 3401 2857
rect 3435 2823 3446 2857
rect 3390 2767 3446 2823
rect 3476 2837 3532 2967
rect 3476 2803 3487 2837
rect 3521 2803 3532 2837
rect 3476 2767 3532 2803
rect 3562 2943 3618 2967
rect 3562 2909 3573 2943
rect 3607 2909 3618 2943
rect 3562 2857 3618 2909
rect 3562 2823 3573 2857
rect 3607 2823 3618 2857
rect 3562 2767 3618 2823
rect 3648 2837 3704 2967
rect 3648 2803 3659 2837
rect 3693 2803 3704 2837
rect 3648 2767 3704 2803
rect 3734 2943 3790 2967
rect 3734 2909 3745 2943
rect 3779 2909 3790 2943
rect 3734 2857 3790 2909
rect 3734 2823 3745 2857
rect 3779 2823 3790 2857
rect 3734 2767 3790 2823
rect 3820 2837 3876 2967
rect 3820 2803 3831 2837
rect 3865 2803 3876 2837
rect 3820 2767 3876 2803
rect 3906 2943 3962 2967
rect 3906 2909 3917 2943
rect 3951 2909 3962 2943
rect 3906 2857 3962 2909
rect 3906 2823 3917 2857
rect 3951 2823 3962 2857
rect 3906 2767 3962 2823
rect 3992 2881 4048 2967
rect 3992 2847 4003 2881
rect 4037 2847 4048 2881
rect 3992 2813 4048 2847
rect 3992 2779 4003 2813
rect 4037 2779 4048 2813
rect 3992 2767 4048 2779
rect 4078 2897 4134 2967
rect 4078 2863 4089 2897
rect 4123 2863 4134 2897
rect 4078 2829 4134 2863
rect 4078 2795 4089 2829
rect 4123 2795 4134 2829
rect 4078 2767 4134 2795
rect 4164 2881 4220 2967
rect 4164 2847 4175 2881
rect 4209 2847 4220 2881
rect 4164 2813 4220 2847
rect 4164 2779 4175 2813
rect 4209 2779 4220 2813
rect 4164 2767 4220 2779
rect 4250 2889 4306 2967
rect 4250 2855 4261 2889
rect 4295 2855 4306 2889
rect 4250 2821 4306 2855
rect 4250 2787 4261 2821
rect 4295 2787 4306 2821
rect 4250 2767 4306 2787
rect 4336 2881 4389 2967
rect 4336 2847 4347 2881
rect 4381 2847 4389 2881
rect 4336 2813 4389 2847
rect 4336 2779 4347 2813
rect 4381 2779 4389 2813
rect 4336 2767 4389 2779
rect 4443 2813 4495 2941
rect 4443 2779 4451 2813
rect 4485 2779 4495 2813
rect 4443 2767 4495 2779
rect 5441 2813 5493 2941
rect 5441 2779 5451 2813
rect 5485 2779 5493 2813
rect 5441 2767 5493 2779
rect 5547 2915 5599 2941
rect 5547 2881 5555 2915
rect 5589 2881 5599 2915
rect 5547 2813 5599 2881
rect 5547 2779 5555 2813
rect 5589 2779 5599 2813
rect 5547 2767 5599 2779
rect 6177 2915 6229 2941
rect 6177 2881 6187 2915
rect 6221 2881 6229 2915
rect 6177 2813 6229 2881
rect 6177 2779 6187 2813
rect 6221 2779 6229 2813
rect 6375 2915 6427 2941
rect 6375 2881 6383 2915
rect 6417 2881 6427 2915
rect 6375 2813 6427 2881
rect 6177 2767 6229 2779
rect 6375 2779 6383 2813
rect 6417 2779 6427 2813
rect 6375 2767 6427 2779
rect 7005 2915 7057 2941
rect 7005 2881 7015 2915
rect 7049 2881 7057 2915
rect 7005 2813 7057 2881
rect 7005 2779 7015 2813
rect 7049 2779 7057 2813
rect 7005 2767 7057 2779
rect 7387 2915 7439 2941
rect 7387 2881 7395 2915
rect 7429 2881 7439 2915
rect 7387 2813 7439 2881
rect 7387 2779 7395 2813
rect 7429 2779 7439 2813
rect 7387 2767 7439 2779
rect 7649 2915 7701 2941
rect 7649 2881 7659 2915
rect 7693 2881 7701 2915
rect 7649 2813 7701 2881
rect 7649 2779 7659 2813
rect 7693 2779 7701 2813
rect 7649 2767 7701 2779
rect 7755 2881 7808 2967
rect 7755 2847 7763 2881
rect 7797 2847 7808 2881
rect 7755 2813 7808 2847
rect 7755 2779 7763 2813
rect 7797 2779 7808 2813
rect 7755 2767 7808 2779
rect 7838 2889 7894 2967
rect 7838 2855 7849 2889
rect 7883 2855 7894 2889
rect 7838 2821 7894 2855
rect 7838 2787 7849 2821
rect 7883 2787 7894 2821
rect 7838 2767 7894 2787
rect 7924 2881 7980 2967
rect 7924 2847 7935 2881
rect 7969 2847 7980 2881
rect 7924 2813 7980 2847
rect 7924 2779 7935 2813
rect 7969 2779 7980 2813
rect 7924 2767 7980 2779
rect 8010 2897 8066 2967
rect 8010 2863 8021 2897
rect 8055 2863 8066 2897
rect 8010 2829 8066 2863
rect 8010 2795 8021 2829
rect 8055 2795 8066 2829
rect 8010 2767 8066 2795
rect 8096 2881 8152 2967
rect 8096 2847 8107 2881
rect 8141 2847 8152 2881
rect 8096 2813 8152 2847
rect 8096 2779 8107 2813
rect 8141 2779 8152 2813
rect 8096 2767 8152 2779
rect 8182 2943 8238 2967
rect 8182 2909 8193 2943
rect 8227 2909 8238 2943
rect 8182 2857 8238 2909
rect 8182 2823 8193 2857
rect 8227 2823 8238 2857
rect 8182 2767 8238 2823
rect 8268 2837 8324 2967
rect 8268 2803 8279 2837
rect 8313 2803 8324 2837
rect 8268 2767 8324 2803
rect 8354 2943 8410 2967
rect 8354 2909 8365 2943
rect 8399 2909 8410 2943
rect 8354 2857 8410 2909
rect 8354 2823 8365 2857
rect 8399 2823 8410 2857
rect 8354 2767 8410 2823
rect 8440 2837 8496 2967
rect 8440 2803 8451 2837
rect 8485 2803 8496 2837
rect 8440 2767 8496 2803
rect 8526 2943 8582 2967
rect 8526 2909 8537 2943
rect 8571 2909 8582 2943
rect 8526 2857 8582 2909
rect 8526 2823 8537 2857
rect 8571 2823 8582 2857
rect 8526 2767 8582 2823
rect 8612 2837 8668 2967
rect 8612 2803 8623 2837
rect 8657 2803 8668 2837
rect 8612 2767 8668 2803
rect 8698 2943 8754 2967
rect 8698 2909 8709 2943
rect 8743 2909 8754 2943
rect 8698 2857 8754 2909
rect 8698 2823 8709 2857
rect 8743 2823 8754 2857
rect 8698 2767 8754 2823
rect 8784 2837 8839 2967
rect 8784 2803 8795 2837
rect 8829 2803 8839 2837
rect 8784 2767 8839 2803
rect 8869 2943 8925 2967
rect 8869 2909 8880 2943
rect 8914 2909 8925 2943
rect 8869 2857 8925 2909
rect 8869 2823 8880 2857
rect 8914 2823 8925 2857
rect 8869 2767 8925 2823
rect 8955 2837 9011 2967
rect 8955 2803 8966 2837
rect 9000 2803 9011 2837
rect 8955 2767 9011 2803
rect 9041 2943 9097 2967
rect 9041 2909 9052 2943
rect 9086 2909 9097 2943
rect 9041 2857 9097 2909
rect 9041 2823 9052 2857
rect 9086 2823 9097 2857
rect 9041 2767 9097 2823
rect 9127 2837 9183 2967
rect 9127 2803 9138 2837
rect 9172 2803 9183 2837
rect 9127 2767 9183 2803
rect 9213 2943 9269 2967
rect 9213 2909 9224 2943
rect 9258 2909 9269 2943
rect 9213 2857 9269 2909
rect 9213 2823 9224 2857
rect 9258 2823 9269 2857
rect 9213 2767 9269 2823
rect 9299 2837 9355 2967
rect 9299 2803 9310 2837
rect 9344 2803 9355 2837
rect 9299 2767 9355 2803
rect 9385 2943 9441 2967
rect 9385 2909 9396 2943
rect 9430 2909 9441 2943
rect 9385 2857 9441 2909
rect 9385 2823 9396 2857
rect 9430 2823 9441 2857
rect 9385 2767 9441 2823
rect 9471 2837 9524 2967
rect 9471 2803 9482 2837
rect 9516 2803 9524 2837
rect 9471 2767 9524 2803
rect 9595 2813 9647 2941
rect 9595 2779 9603 2813
rect 9637 2779 9647 2813
rect 9595 2767 9647 2779
rect 10593 2813 10645 2941
rect 10593 2779 10603 2813
rect 10637 2779 10645 2813
rect 10593 2767 10645 2779
rect 10699 2915 10751 2941
rect 10699 2881 10707 2915
rect 10741 2881 10751 2915
rect 10699 2813 10751 2881
rect 10699 2779 10707 2813
rect 10741 2779 10751 2813
rect 10699 2767 10751 2779
rect 11329 2915 11381 2941
rect 11329 2881 11339 2915
rect 11373 2881 11381 2915
rect 11329 2813 11381 2881
rect 11329 2779 11339 2813
rect 11373 2779 11381 2813
rect 11711 2889 11763 2901
rect 11711 2855 11719 2889
rect 11753 2855 11763 2889
rect 11711 2821 11763 2855
rect 11711 2787 11719 2821
rect 11753 2787 11763 2821
rect 11329 2767 11381 2779
rect 11711 2773 11763 2787
rect 11793 2837 11847 2901
rect 11793 2803 11803 2837
rect 11837 2803 11847 2837
rect 11793 2773 11847 2803
rect 11877 2889 11929 2901
rect 11877 2855 11887 2889
rect 11921 2855 11929 2889
rect 11877 2821 11929 2855
rect 12899 2955 12953 2967
rect 12363 2881 12450 2917
rect 12363 2851 12406 2881
rect 11877 2787 11887 2821
rect 11921 2787 11929 2821
rect 11877 2773 11929 2787
rect 11983 2813 12035 2851
rect 11983 2779 11991 2813
rect 12025 2779 12035 2813
rect 11983 2767 12035 2779
rect 12065 2821 12120 2851
rect 12065 2787 12075 2821
rect 12109 2787 12120 2821
rect 12065 2767 12120 2787
rect 12150 2826 12215 2851
rect 12150 2792 12167 2826
rect 12201 2792 12215 2826
rect 12150 2767 12215 2792
rect 12245 2767 12318 2851
rect 12348 2847 12406 2851
rect 12440 2847 12450 2881
rect 12348 2813 12450 2847
rect 12348 2779 12406 2813
rect 12440 2779 12450 2813
rect 12348 2767 12450 2779
rect 12480 2851 12530 2917
rect 12899 2921 12907 2955
rect 12941 2921 12953 2955
rect 12899 2884 12953 2921
rect 12480 2821 12545 2851
rect 12480 2787 12490 2821
rect 12524 2787 12545 2821
rect 12480 2767 12545 2787
rect 12575 2831 12629 2851
rect 12575 2797 12585 2831
rect 12619 2797 12629 2831
rect 12575 2767 12629 2797
rect 12659 2767 12743 2851
rect 12773 2821 12826 2851
rect 12773 2787 12784 2821
rect 12818 2787 12826 2821
rect 12773 2767 12826 2787
rect 12899 2850 12907 2884
rect 12941 2850 12953 2884
rect 12899 2813 12953 2850
rect 12899 2779 12907 2813
rect 12941 2779 12953 2813
rect 12899 2767 12953 2779
rect 12983 2923 13037 2967
rect 12983 2889 12993 2923
rect 13027 2889 13037 2923
rect 12983 2843 13037 2889
rect 12983 2809 12993 2843
rect 13027 2809 13037 2843
rect 12983 2767 13037 2809
rect 13067 2955 13119 2967
rect 13067 2921 13077 2955
rect 13111 2921 13119 2955
rect 13067 2887 13119 2921
rect 13067 2853 13077 2887
rect 13111 2853 13119 2887
rect 13067 2819 13119 2853
rect 13067 2785 13077 2819
rect 13111 2785 13119 2819
rect 13067 2767 13119 2785
rect 13183 2813 13235 2941
rect 13183 2779 13191 2813
rect 13225 2779 13235 2813
rect 13183 2767 13235 2779
rect 14181 2813 14233 2941
rect 14181 2779 14191 2813
rect 14225 2779 14233 2813
rect 14181 2767 14233 2779
rect 14287 2813 14339 2941
rect 14287 2779 14295 2813
rect 14329 2779 14339 2813
rect 14287 2767 14339 2779
rect 15285 2813 15337 2941
rect 15285 2779 15295 2813
rect 15329 2779 15337 2813
rect 15285 2767 15337 2779
rect 15391 2813 15443 2941
rect 15391 2779 15399 2813
rect 15433 2779 15443 2813
rect 15391 2767 15443 2779
rect 16389 2813 16441 2941
rect 16389 2779 16399 2813
rect 16433 2779 16441 2813
rect 16863 2902 16915 2925
rect 16863 2868 16871 2902
rect 16905 2868 16915 2902
rect 16863 2821 16915 2868
rect 16863 2787 16871 2821
rect 16905 2787 16915 2821
rect 16389 2767 16441 2779
rect 16863 2767 16915 2787
rect 16945 2889 17003 2925
rect 16945 2855 16957 2889
rect 16991 2855 17003 2889
rect 16945 2821 17003 2855
rect 16945 2787 16957 2821
rect 16991 2787 17003 2821
rect 16945 2767 17003 2787
rect 17033 2889 17085 2925
rect 17033 2855 17043 2889
rect 17077 2855 17085 2889
rect 17033 2821 17085 2855
rect 17033 2787 17043 2821
rect 17077 2787 17085 2821
rect 17033 2767 17085 2787
rect 17139 2813 17191 2941
rect 17139 2779 17147 2813
rect 17181 2779 17191 2813
rect 17139 2767 17191 2779
rect 18137 2813 18189 2941
rect 18137 2779 18147 2813
rect 18181 2779 18189 2813
rect 18137 2767 18189 2779
rect 18243 2915 18295 2941
rect 18243 2881 18251 2915
rect 18285 2881 18295 2915
rect 18243 2813 18295 2881
rect 18243 2779 18251 2813
rect 18285 2779 18295 2813
rect 18243 2767 18295 2779
rect 18505 2915 18557 2941
rect 18505 2881 18515 2915
rect 18549 2881 18557 2915
rect 18505 2813 18557 2881
rect 18505 2779 18515 2813
rect 18549 2779 18557 2813
rect 18505 2767 18557 2779
rect 18611 2908 18663 2941
rect 18611 2874 18619 2908
rect 18653 2874 18663 2908
rect 18611 2813 18663 2874
rect 18611 2779 18619 2813
rect 18653 2779 18663 2813
rect 18611 2767 18663 2779
rect 18781 2908 18833 2941
rect 18781 2874 18791 2908
rect 18825 2874 18833 2908
rect 18781 2813 18833 2874
rect 18781 2779 18791 2813
rect 18825 2779 18833 2813
rect 18781 2767 18833 2779
rect 1131 2661 1183 2673
rect 1131 2627 1139 2661
rect 1173 2627 1183 2661
rect 1131 2566 1183 2627
rect 1131 2532 1139 2566
rect 1173 2532 1183 2566
rect 1131 2499 1183 2532
rect 1301 2661 1353 2673
rect 1301 2627 1311 2661
rect 1345 2627 1353 2661
rect 1301 2566 1353 2627
rect 1301 2532 1311 2566
rect 1345 2532 1353 2566
rect 1301 2499 1353 2532
rect 1407 2661 1459 2673
rect 1407 2627 1415 2661
rect 1449 2627 1459 2661
rect 1407 2559 1459 2627
rect 1407 2525 1415 2559
rect 1449 2525 1459 2559
rect 1407 2499 1459 2525
rect 1853 2661 1905 2673
rect 1853 2627 1863 2661
rect 1897 2627 1905 2661
rect 1853 2559 1905 2627
rect 1853 2525 1863 2559
rect 1897 2525 1905 2559
rect 1853 2499 1905 2525
rect 2061 2655 2113 2673
rect 2061 2621 2069 2655
rect 2103 2621 2113 2655
rect 2061 2587 2113 2621
rect 2061 2553 2069 2587
rect 2103 2553 2113 2587
rect 2061 2519 2113 2553
rect 2061 2485 2069 2519
rect 2103 2485 2113 2519
rect 2061 2473 2113 2485
rect 2143 2631 2197 2673
rect 2143 2597 2153 2631
rect 2187 2597 2197 2631
rect 2143 2551 2197 2597
rect 2143 2517 2153 2551
rect 2187 2517 2197 2551
rect 2143 2473 2197 2517
rect 2227 2661 2281 2673
rect 2227 2627 2239 2661
rect 2273 2627 2281 2661
rect 2227 2590 2281 2627
rect 2227 2556 2239 2590
rect 2273 2556 2281 2590
rect 2354 2653 2407 2673
rect 2354 2619 2362 2653
rect 2396 2619 2407 2653
rect 2354 2589 2407 2619
rect 2437 2589 2521 2673
rect 2551 2643 2605 2673
rect 2551 2609 2561 2643
rect 2595 2609 2605 2643
rect 2551 2589 2605 2609
rect 2635 2653 2700 2673
rect 2635 2619 2656 2653
rect 2690 2619 2700 2653
rect 2635 2589 2700 2619
rect 2227 2519 2281 2556
rect 2227 2485 2239 2519
rect 2273 2485 2281 2519
rect 2650 2523 2700 2589
rect 2730 2661 2832 2673
rect 2730 2627 2740 2661
rect 2774 2627 2832 2661
rect 2730 2593 2832 2627
rect 2730 2559 2740 2593
rect 2774 2589 2832 2593
rect 2862 2589 2935 2673
rect 2965 2648 3030 2673
rect 2965 2614 2979 2648
rect 3013 2614 3030 2648
rect 2965 2589 3030 2614
rect 3060 2653 3115 2673
rect 3060 2619 3071 2653
rect 3105 2619 3115 2653
rect 3060 2589 3115 2619
rect 3145 2661 3197 2673
rect 3145 2627 3155 2661
rect 3189 2627 3197 2661
rect 3145 2589 3197 2627
rect 3251 2653 3303 2667
rect 3251 2619 3259 2653
rect 3293 2619 3303 2653
rect 2774 2559 2817 2589
rect 2730 2523 2817 2559
rect 2227 2473 2281 2485
rect 3251 2585 3303 2619
rect 3251 2551 3259 2585
rect 3293 2551 3303 2585
rect 3251 2539 3303 2551
rect 3333 2637 3387 2667
rect 3333 2603 3343 2637
rect 3377 2603 3387 2637
rect 3333 2539 3387 2603
rect 3417 2653 3469 2667
rect 4167 2661 4219 2673
rect 3417 2619 3427 2653
rect 3461 2619 3469 2653
rect 3417 2585 3469 2619
rect 3417 2551 3427 2585
rect 3461 2551 3469 2585
rect 3417 2539 3469 2551
rect 4167 2627 4175 2661
rect 4209 2627 4219 2661
rect 4167 2559 4219 2627
rect 4167 2525 4175 2559
rect 4209 2525 4219 2559
rect 4167 2499 4219 2525
rect 4429 2661 4481 2673
rect 4429 2627 4439 2661
rect 4473 2627 4481 2661
rect 4429 2559 4481 2627
rect 4429 2525 4439 2559
rect 4473 2525 4481 2559
rect 4627 2653 4679 2667
rect 4627 2619 4635 2653
rect 4669 2619 4679 2653
rect 4627 2585 4679 2619
rect 4627 2551 4635 2585
rect 4669 2551 4679 2585
rect 4627 2539 4679 2551
rect 4709 2637 4763 2667
rect 4709 2603 4719 2637
rect 4753 2603 4763 2637
rect 4709 2539 4763 2603
rect 4793 2653 4845 2667
rect 4793 2619 4803 2653
rect 4837 2619 4845 2653
rect 4793 2585 4845 2619
rect 4899 2661 4951 2673
rect 4899 2627 4907 2661
rect 4941 2627 4951 2661
rect 4899 2589 4951 2627
rect 4981 2653 5036 2673
rect 4981 2619 4991 2653
rect 5025 2619 5036 2653
rect 4981 2589 5036 2619
rect 5066 2648 5131 2673
rect 5066 2614 5083 2648
rect 5117 2614 5131 2648
rect 5066 2589 5131 2614
rect 5161 2589 5234 2673
rect 5264 2661 5366 2673
rect 5264 2627 5322 2661
rect 5356 2627 5366 2661
rect 5264 2593 5366 2627
rect 5264 2589 5322 2593
rect 4793 2551 4803 2585
rect 4837 2551 4845 2585
rect 4793 2539 4845 2551
rect 4429 2499 4481 2525
rect 5279 2559 5322 2589
rect 5356 2559 5366 2593
rect 5279 2523 5366 2559
rect 5396 2653 5461 2673
rect 5396 2619 5406 2653
rect 5440 2619 5461 2653
rect 5396 2589 5461 2619
rect 5491 2643 5545 2673
rect 5491 2609 5501 2643
rect 5535 2609 5545 2643
rect 5491 2589 5545 2609
rect 5575 2589 5659 2673
rect 5689 2653 5742 2673
rect 5689 2619 5700 2653
rect 5734 2619 5742 2653
rect 5689 2589 5742 2619
rect 5815 2661 5869 2673
rect 5815 2627 5823 2661
rect 5857 2627 5869 2661
rect 5815 2590 5869 2627
rect 5396 2523 5446 2589
rect 5815 2556 5823 2590
rect 5857 2556 5869 2590
rect 5815 2519 5869 2556
rect 5815 2485 5823 2519
rect 5857 2485 5869 2519
rect 5815 2473 5869 2485
rect 5899 2631 5953 2673
rect 5899 2597 5909 2631
rect 5943 2597 5953 2631
rect 5899 2551 5953 2597
rect 5899 2517 5909 2551
rect 5943 2517 5953 2551
rect 5899 2473 5953 2517
rect 5983 2655 6035 2673
rect 6375 2661 6427 2673
rect 5983 2621 5993 2655
rect 6027 2621 6035 2655
rect 5983 2587 6035 2621
rect 5983 2553 5993 2587
rect 6027 2553 6035 2587
rect 5983 2519 6035 2553
rect 5983 2485 5993 2519
rect 6027 2485 6035 2519
rect 5983 2473 6035 2485
rect 6375 2627 6383 2661
rect 6417 2627 6427 2661
rect 6375 2559 6427 2627
rect 6375 2525 6383 2559
rect 6417 2525 6427 2559
rect 6375 2499 6427 2525
rect 7005 2661 7057 2673
rect 7005 2627 7015 2661
rect 7049 2627 7057 2661
rect 7005 2559 7057 2627
rect 7005 2525 7015 2559
rect 7049 2525 7057 2559
rect 7005 2499 7057 2525
rect 7213 2655 7265 2673
rect 7213 2621 7221 2655
rect 7255 2621 7265 2655
rect 7213 2587 7265 2621
rect 7213 2553 7221 2587
rect 7255 2553 7265 2587
rect 7213 2519 7265 2553
rect 7213 2485 7221 2519
rect 7255 2485 7265 2519
rect 7213 2473 7265 2485
rect 7295 2631 7349 2673
rect 7295 2597 7305 2631
rect 7339 2597 7349 2631
rect 7295 2551 7349 2597
rect 7295 2517 7305 2551
rect 7339 2517 7349 2551
rect 7295 2473 7349 2517
rect 7379 2661 7433 2673
rect 7379 2627 7391 2661
rect 7425 2627 7433 2661
rect 7379 2590 7433 2627
rect 7379 2556 7391 2590
rect 7425 2556 7433 2590
rect 7506 2653 7559 2673
rect 7506 2619 7514 2653
rect 7548 2619 7559 2653
rect 7506 2589 7559 2619
rect 7589 2589 7673 2673
rect 7703 2643 7757 2673
rect 7703 2609 7713 2643
rect 7747 2609 7757 2643
rect 7703 2589 7757 2609
rect 7787 2653 7852 2673
rect 7787 2619 7808 2653
rect 7842 2619 7852 2653
rect 7787 2589 7852 2619
rect 7379 2519 7433 2556
rect 7379 2485 7391 2519
rect 7425 2485 7433 2519
rect 7802 2523 7852 2589
rect 7882 2661 7984 2673
rect 7882 2627 7892 2661
rect 7926 2627 7984 2661
rect 7882 2593 7984 2627
rect 7882 2559 7892 2593
rect 7926 2589 7984 2593
rect 8014 2589 8087 2673
rect 8117 2648 8182 2673
rect 8117 2614 8131 2648
rect 8165 2614 8182 2648
rect 8117 2589 8182 2614
rect 8212 2653 8267 2673
rect 8212 2619 8223 2653
rect 8257 2619 8267 2653
rect 8212 2589 8267 2619
rect 8297 2661 8349 2673
rect 8297 2627 8307 2661
rect 8341 2627 8349 2661
rect 8297 2589 8349 2627
rect 8403 2653 8455 2667
rect 8403 2619 8411 2653
rect 8445 2619 8455 2653
rect 7926 2559 7969 2589
rect 7882 2523 7969 2559
rect 7379 2473 7433 2485
rect 8403 2585 8455 2619
rect 8403 2551 8411 2585
rect 8445 2551 8455 2585
rect 8403 2539 8455 2551
rect 8485 2637 8539 2667
rect 8485 2603 8495 2637
rect 8529 2603 8539 2637
rect 8485 2539 8539 2603
rect 8569 2653 8621 2667
rect 8951 2661 9003 2673
rect 8569 2619 8579 2653
rect 8613 2619 8621 2653
rect 8569 2585 8621 2619
rect 8569 2551 8579 2585
rect 8613 2551 8621 2585
rect 8569 2539 8621 2551
rect 8951 2627 8959 2661
rect 8993 2627 9003 2661
rect 8951 2559 9003 2627
rect 8951 2525 8959 2559
rect 8993 2525 9003 2559
rect 8951 2499 9003 2525
rect 9581 2661 9633 2673
rect 9581 2627 9591 2661
rect 9625 2627 9633 2661
rect 9581 2559 9633 2627
rect 9581 2525 9591 2559
rect 9625 2525 9633 2559
rect 9779 2653 9831 2667
rect 9779 2619 9787 2653
rect 9821 2619 9831 2653
rect 9779 2585 9831 2619
rect 9779 2551 9787 2585
rect 9821 2551 9831 2585
rect 9779 2539 9831 2551
rect 9861 2637 9915 2667
rect 9861 2603 9871 2637
rect 9905 2603 9915 2637
rect 9861 2539 9915 2603
rect 9945 2653 9997 2667
rect 9945 2619 9955 2653
rect 9989 2619 9997 2653
rect 9945 2585 9997 2619
rect 10051 2661 10103 2673
rect 10051 2627 10059 2661
rect 10093 2627 10103 2661
rect 10051 2589 10103 2627
rect 10133 2653 10188 2673
rect 10133 2619 10143 2653
rect 10177 2619 10188 2653
rect 10133 2589 10188 2619
rect 10218 2648 10283 2673
rect 10218 2614 10235 2648
rect 10269 2614 10283 2648
rect 10218 2589 10283 2614
rect 10313 2589 10386 2673
rect 10416 2661 10518 2673
rect 10416 2627 10474 2661
rect 10508 2627 10518 2661
rect 10416 2593 10518 2627
rect 10416 2589 10474 2593
rect 9945 2551 9955 2585
rect 9989 2551 9997 2585
rect 9945 2539 9997 2551
rect 9581 2499 9633 2525
rect 10431 2559 10474 2589
rect 10508 2559 10518 2593
rect 10431 2523 10518 2559
rect 10548 2653 10613 2673
rect 10548 2619 10558 2653
rect 10592 2619 10613 2653
rect 10548 2589 10613 2619
rect 10643 2643 10697 2673
rect 10643 2609 10653 2643
rect 10687 2609 10697 2643
rect 10643 2589 10697 2609
rect 10727 2589 10811 2673
rect 10841 2653 10894 2673
rect 10841 2619 10852 2653
rect 10886 2619 10894 2653
rect 10841 2589 10894 2619
rect 10967 2661 11021 2673
rect 10967 2627 10975 2661
rect 11009 2627 11021 2661
rect 10967 2590 11021 2627
rect 10548 2523 10598 2589
rect 10967 2556 10975 2590
rect 11009 2556 11021 2590
rect 10967 2519 11021 2556
rect 10967 2485 10975 2519
rect 11009 2485 11021 2519
rect 10967 2473 11021 2485
rect 11051 2631 11105 2673
rect 11051 2597 11061 2631
rect 11095 2597 11105 2631
rect 11051 2551 11105 2597
rect 11051 2517 11061 2551
rect 11095 2517 11105 2551
rect 11051 2473 11105 2517
rect 11135 2655 11187 2673
rect 11527 2661 11579 2673
rect 11135 2621 11145 2655
rect 11179 2621 11187 2655
rect 11135 2587 11187 2621
rect 11135 2553 11145 2587
rect 11179 2553 11187 2587
rect 11135 2519 11187 2553
rect 11135 2485 11145 2519
rect 11179 2485 11187 2519
rect 11135 2473 11187 2485
rect 11527 2627 11535 2661
rect 11569 2627 11579 2661
rect 11527 2559 11579 2627
rect 11527 2525 11535 2559
rect 11569 2525 11579 2559
rect 11527 2499 11579 2525
rect 11789 2661 11841 2673
rect 11789 2627 11799 2661
rect 11833 2627 11841 2661
rect 11789 2559 11841 2627
rect 11789 2525 11799 2559
rect 11833 2525 11841 2559
rect 11789 2499 11841 2525
rect 11905 2655 11957 2673
rect 11905 2621 11913 2655
rect 11947 2621 11957 2655
rect 11905 2587 11957 2621
rect 11905 2553 11913 2587
rect 11947 2553 11957 2587
rect 11905 2519 11957 2553
rect 11905 2485 11913 2519
rect 11947 2485 11957 2519
rect 11905 2473 11957 2485
rect 11987 2631 12041 2673
rect 11987 2597 11997 2631
rect 12031 2597 12041 2631
rect 11987 2551 12041 2597
rect 11987 2517 11997 2551
rect 12031 2517 12041 2551
rect 11987 2473 12041 2517
rect 12071 2661 12125 2673
rect 12071 2627 12083 2661
rect 12117 2627 12125 2661
rect 12071 2590 12125 2627
rect 12071 2556 12083 2590
rect 12117 2556 12125 2590
rect 12198 2653 12251 2673
rect 12198 2619 12206 2653
rect 12240 2619 12251 2653
rect 12198 2589 12251 2619
rect 12281 2589 12365 2673
rect 12395 2643 12449 2673
rect 12395 2609 12405 2643
rect 12439 2609 12449 2643
rect 12395 2589 12449 2609
rect 12479 2653 12544 2673
rect 12479 2619 12500 2653
rect 12534 2619 12544 2653
rect 12479 2589 12544 2619
rect 12071 2519 12125 2556
rect 12071 2485 12083 2519
rect 12117 2485 12125 2519
rect 12494 2523 12544 2589
rect 12574 2661 12676 2673
rect 12574 2627 12584 2661
rect 12618 2627 12676 2661
rect 12574 2593 12676 2627
rect 12574 2559 12584 2593
rect 12618 2589 12676 2593
rect 12706 2589 12779 2673
rect 12809 2648 12874 2673
rect 12809 2614 12823 2648
rect 12857 2614 12874 2648
rect 12809 2589 12874 2614
rect 12904 2653 12959 2673
rect 12904 2619 12915 2653
rect 12949 2619 12959 2653
rect 12904 2589 12959 2619
rect 12989 2661 13041 2673
rect 12989 2627 12999 2661
rect 13033 2627 13041 2661
rect 12989 2589 13041 2627
rect 13095 2653 13147 2667
rect 13095 2619 13103 2653
rect 13137 2619 13147 2653
rect 12618 2559 12661 2589
rect 12574 2523 12661 2559
rect 12071 2473 12125 2485
rect 13095 2585 13147 2619
rect 13095 2551 13103 2585
rect 13137 2551 13147 2585
rect 13095 2539 13147 2551
rect 13177 2637 13231 2667
rect 13177 2603 13187 2637
rect 13221 2603 13231 2637
rect 13177 2539 13231 2603
rect 13261 2653 13313 2667
rect 13261 2619 13271 2653
rect 13305 2619 13313 2653
rect 13261 2585 13313 2619
rect 13261 2551 13271 2585
rect 13305 2551 13313 2585
rect 13261 2539 13313 2551
rect 13367 2661 13419 2673
rect 13367 2627 13375 2661
rect 13409 2627 13419 2661
rect 13367 2559 13419 2627
rect 13367 2525 13375 2559
rect 13409 2525 13419 2559
rect 13367 2499 13419 2525
rect 13813 2661 13865 2673
rect 13813 2627 13823 2661
rect 13857 2627 13865 2661
rect 13813 2559 13865 2627
rect 13813 2525 13823 2559
rect 13857 2525 13865 2559
rect 13813 2499 13865 2525
rect 14563 2661 14615 2673
rect 14563 2627 14571 2661
rect 14605 2627 14615 2661
rect 14563 2499 14615 2627
rect 15561 2661 15613 2673
rect 15561 2627 15571 2661
rect 15605 2627 15613 2661
rect 15561 2499 15613 2627
rect 15667 2661 15719 2673
rect 15667 2627 15675 2661
rect 15709 2627 15719 2661
rect 15667 2559 15719 2627
rect 15667 2525 15675 2559
rect 15709 2525 15719 2559
rect 15667 2499 15719 2525
rect 16297 2661 16349 2673
rect 16297 2627 16307 2661
rect 16341 2627 16349 2661
rect 16297 2559 16349 2627
rect 16297 2525 16307 2559
rect 16341 2525 16349 2559
rect 16297 2499 16349 2525
rect 16863 2653 16915 2673
rect 16863 2619 16871 2653
rect 16905 2619 16915 2653
rect 16863 2572 16915 2619
rect 16863 2538 16871 2572
rect 16905 2538 16915 2572
rect 16863 2515 16915 2538
rect 16945 2653 17003 2673
rect 16945 2619 16957 2653
rect 16991 2619 17003 2653
rect 16945 2585 17003 2619
rect 16945 2551 16957 2585
rect 16991 2551 17003 2585
rect 16945 2515 17003 2551
rect 17033 2653 17085 2673
rect 17033 2619 17043 2653
rect 17077 2619 17085 2653
rect 17033 2585 17085 2619
rect 17033 2551 17043 2585
rect 17077 2551 17085 2585
rect 17033 2515 17085 2551
rect 17139 2661 17191 2673
rect 17139 2627 17147 2661
rect 17181 2627 17191 2661
rect 17139 2559 17191 2627
rect 17139 2525 17147 2559
rect 17181 2525 17191 2559
rect 17139 2499 17191 2525
rect 17401 2661 17453 2673
rect 17604 2665 17654 2673
rect 17401 2627 17411 2661
rect 17445 2627 17453 2661
rect 17401 2559 17453 2627
rect 17401 2525 17411 2559
rect 17445 2525 17453 2559
rect 17507 2653 17559 2665
rect 17507 2619 17515 2653
rect 17549 2619 17559 2653
rect 17507 2585 17559 2619
rect 17507 2551 17515 2585
rect 17549 2551 17559 2585
rect 17507 2537 17559 2551
rect 17589 2653 17654 2665
rect 17589 2619 17608 2653
rect 17642 2619 17654 2653
rect 17589 2585 17654 2619
rect 17589 2551 17608 2585
rect 17642 2551 17654 2585
rect 17589 2537 17654 2551
rect 17401 2499 17453 2525
rect 17604 2473 17654 2537
rect 17684 2637 17738 2673
rect 17684 2603 17694 2637
rect 17728 2603 17738 2637
rect 17684 2556 17738 2603
rect 17684 2522 17694 2556
rect 17728 2522 17738 2556
rect 17684 2473 17738 2522
rect 17768 2661 17821 2673
rect 17768 2627 17778 2661
rect 17812 2627 17821 2661
rect 17768 2593 17821 2627
rect 17768 2559 17778 2593
rect 17812 2559 17821 2593
rect 17768 2525 17821 2559
rect 17768 2491 17778 2525
rect 17812 2491 17821 2525
rect 17875 2661 17927 2673
rect 17875 2627 17883 2661
rect 17917 2627 17927 2661
rect 17875 2559 17927 2627
rect 17875 2525 17883 2559
rect 17917 2525 17927 2559
rect 17875 2499 17927 2525
rect 18505 2661 18557 2673
rect 18505 2627 18515 2661
rect 18549 2627 18557 2661
rect 18505 2559 18557 2627
rect 18505 2525 18515 2559
rect 18549 2525 18557 2559
rect 18505 2499 18557 2525
rect 18611 2661 18663 2673
rect 18611 2627 18619 2661
rect 18653 2627 18663 2661
rect 18611 2566 18663 2627
rect 18611 2532 18619 2566
rect 18653 2532 18663 2566
rect 18611 2499 18663 2532
rect 18781 2661 18833 2673
rect 18781 2627 18791 2661
rect 18825 2627 18833 2661
rect 18781 2566 18833 2627
rect 18781 2532 18791 2566
rect 18825 2532 18833 2566
rect 18781 2499 18833 2532
rect 17768 2473 17821 2491
<< ndiffc >>
rect 1139 7502 1173 7536
rect 1311 7502 1345 7536
rect 1600 7519 1634 7553
rect 1600 7451 1634 7485
rect 1684 7493 1718 7527
rect 1770 7523 1804 7557
rect 1863 7510 1897 7544
rect 1967 7504 2001 7538
rect 2967 7504 3001 7538
rect 3071 7504 3105 7538
rect 3519 7504 3553 7538
rect 3992 7519 4026 7553
rect 3992 7451 4026 7485
rect 4076 7493 4110 7527
rect 4162 7523 4196 7557
rect 4255 7510 4289 7544
rect 4359 7504 4393 7538
rect 5359 7504 5393 7538
rect 5648 7519 5682 7553
rect 5648 7451 5682 7485
rect 5732 7493 5766 7527
rect 5818 7523 5852 7557
rect 5911 7510 5945 7544
rect 6015 7502 6049 7536
rect 6187 7502 6221 7536
rect 6383 7504 6417 7538
rect 7383 7504 7417 7538
rect 7487 7497 7521 7531
rect 7751 7497 7785 7531
rect 7855 7510 7889 7544
rect 7948 7523 7982 7557
rect 8034 7493 8068 7527
rect 8118 7519 8152 7553
rect 8118 7451 8152 7485
rect 8223 7504 8257 7538
rect 8671 7504 8705 7538
rect 8959 7504 8993 7538
rect 9407 7504 9441 7538
rect 9695 7497 9729 7531
rect 9959 7497 9993 7531
rect 10063 7515 10097 7549
rect 10149 7519 10183 7553
rect 10243 7515 10277 7549
rect 10327 7519 10361 7553
rect 10431 7504 10465 7538
rect 11063 7504 11097 7538
rect 11167 7502 11201 7536
rect 11339 7502 11373 7536
rect 11535 7504 11569 7538
rect 12167 7504 12201 7538
rect 12271 7510 12305 7544
rect 12364 7523 12398 7557
rect 12450 7493 12484 7527
rect 12534 7519 12568 7553
rect 12534 7451 12568 7485
rect 12639 7504 12673 7538
rect 13639 7504 13673 7538
rect 13743 7502 13777 7536
rect 13915 7502 13949 7536
rect 14111 7497 14145 7531
rect 14375 7497 14409 7531
rect 14479 7510 14513 7544
rect 14572 7523 14606 7557
rect 14658 7493 14692 7527
rect 14742 7519 14776 7553
rect 14742 7451 14776 7485
rect 14847 7504 14881 7538
rect 15847 7504 15881 7538
rect 15951 7504 15985 7538
rect 16399 7504 16433 7538
rect 16871 7510 16905 7544
rect 16964 7523 16998 7557
rect 17050 7493 17084 7527
rect 17134 7519 17168 7553
rect 17134 7451 17168 7485
rect 17239 7504 17273 7538
rect 17871 7504 17905 7538
rect 18067 7510 18101 7544
rect 18160 7523 18194 7557
rect 18246 7493 18280 7527
rect 18330 7519 18364 7553
rect 18330 7451 18364 7485
rect 18619 7502 18653 7536
rect 18791 7502 18825 7536
rect 1139 6608 1173 6642
rect 1311 6608 1345 6642
rect 1415 6606 1449 6640
rect 2415 6606 2449 6640
rect 2519 6606 2553 6640
rect 3519 6606 3553 6640
rect 3807 6606 3841 6640
rect 4807 6606 4841 6640
rect 4911 6606 4945 6640
rect 5911 6606 5945 6640
rect 6015 6606 6049 6640
rect 7015 6606 7049 6640
rect 7119 6606 7153 6640
rect 8119 6606 8153 6640
rect 8223 6606 8257 6640
rect 8671 6606 8705 6640
rect 8959 6606 8993 6640
rect 9959 6606 9993 6640
rect 10063 6606 10097 6640
rect 11063 6606 11097 6640
rect 11167 6606 11201 6640
rect 12167 6606 12201 6640
rect 12271 6606 12305 6640
rect 13271 6606 13305 6640
rect 13375 6606 13409 6640
rect 13823 6606 13857 6640
rect 14111 6606 14145 6640
rect 15111 6606 15145 6640
rect 15215 6606 15249 6640
rect 16215 6606 16249 6640
rect 16319 6606 16353 6640
rect 17319 6606 17353 6640
rect 17423 6606 17457 6640
rect 18423 6606 18457 6640
rect 18619 6608 18653 6642
rect 18791 6608 18825 6642
rect 1139 6414 1173 6448
rect 1311 6414 1345 6448
rect 1415 6416 1449 6450
rect 2415 6416 2449 6450
rect 2519 6416 2553 6450
rect 3519 6416 3553 6450
rect 3623 6416 3657 6450
rect 4623 6416 4657 6450
rect 4727 6416 4761 6450
rect 5727 6416 5761 6450
rect 5831 6409 5865 6443
rect 6095 6409 6129 6443
rect 6383 6416 6417 6450
rect 7383 6416 7417 6450
rect 7487 6416 7521 6450
rect 8487 6416 8521 6450
rect 8591 6416 8625 6450
rect 9591 6416 9625 6450
rect 9695 6416 9729 6450
rect 10695 6416 10729 6450
rect 10799 6416 10833 6450
rect 11247 6416 11281 6450
rect 11535 6416 11569 6450
rect 12535 6416 12569 6450
rect 12639 6416 12673 6450
rect 13639 6416 13673 6450
rect 13743 6416 13777 6450
rect 14743 6416 14777 6450
rect 14847 6416 14881 6450
rect 15847 6416 15881 6450
rect 15951 6416 15985 6450
rect 16399 6416 16433 6450
rect 16687 6416 16721 6450
rect 17687 6416 17721 6450
rect 17791 6416 17825 6450
rect 18423 6416 18457 6450
rect 18619 6414 18653 6448
rect 18791 6414 18825 6448
rect 1139 5520 1173 5554
rect 1311 5520 1345 5554
rect 1415 5518 1449 5552
rect 2047 5518 2081 5552
rect 2243 5512 2277 5546
rect 2329 5499 2363 5533
rect 2415 5529 2449 5563
rect 2519 5518 2553 5552
rect 2967 5518 3001 5552
rect 3071 5529 3105 5563
rect 3157 5499 3191 5533
rect 3243 5512 3277 5546
rect 3347 5525 3381 5559
rect 3611 5525 3645 5559
rect 3807 5518 3841 5552
rect 4807 5518 4841 5552
rect 4911 5518 4945 5552
rect 5911 5518 5945 5552
rect 6015 5518 6049 5552
rect 6647 5518 6681 5552
rect 6751 5518 6785 5552
rect 6835 5499 6869 5533
rect 7042 5514 7076 5548
rect 7277 5514 7311 5548
rect 7345 5514 7379 5548
rect 7429 5514 7463 5548
rect 7579 5518 7613 5552
rect 8579 5518 8613 5552
rect 8959 5518 8993 5552
rect 9591 5518 9625 5552
rect 9879 5518 9913 5552
rect 9963 5499 9997 5533
rect 10170 5514 10204 5548
rect 10405 5514 10439 5548
rect 10473 5514 10507 5548
rect 10557 5514 10591 5548
rect 10707 5525 10741 5559
rect 10971 5525 11005 5559
rect 11119 5499 11153 5533
rect 11203 5499 11237 5533
rect 11395 5527 11429 5561
rect 11535 5518 11569 5552
rect 12167 5518 12201 5552
rect 12271 5518 12305 5552
rect 12355 5499 12389 5533
rect 12562 5514 12596 5548
rect 12797 5514 12831 5548
rect 12865 5514 12899 5548
rect 12949 5514 12983 5548
rect 13099 5518 13133 5552
rect 13731 5518 13765 5552
rect 14295 5518 14329 5552
rect 14379 5499 14413 5533
rect 14586 5514 14620 5548
rect 14821 5514 14855 5548
rect 14889 5514 14923 5548
rect 14973 5514 15007 5548
rect 15123 5518 15157 5552
rect 16123 5518 16157 5552
rect 16227 5518 16261 5552
rect 17227 5518 17261 5552
rect 17331 5518 17365 5552
rect 18331 5518 18365 5552
rect 18619 5520 18653 5554
rect 18791 5520 18825 5554
rect 1139 5326 1173 5360
rect 1311 5326 1345 5360
rect 1415 5328 1449 5362
rect 1863 5328 1897 5362
rect 2011 5347 2045 5381
rect 2095 5347 2129 5381
rect 2287 5319 2321 5353
rect 2427 5321 2461 5355
rect 2691 5321 2725 5355
rect 2931 5347 2965 5381
rect 3015 5347 3049 5381
rect 3207 5319 3241 5353
rect 3347 5321 3381 5355
rect 3611 5321 3645 5355
rect 3715 5334 3749 5368
rect 3808 5347 3842 5381
rect 3894 5317 3928 5351
rect 3978 5343 4012 5377
rect 3978 5275 4012 5309
rect 4083 5321 4117 5355
rect 4347 5321 4381 5355
rect 4453 5347 4487 5381
rect 4453 5275 4487 5309
rect 4537 5347 4571 5381
rect 4537 5275 4571 5309
rect 4621 5347 4655 5381
rect 4621 5275 4655 5309
rect 4727 5328 4761 5362
rect 5727 5328 5761 5362
rect 5831 5317 5865 5351
rect 5917 5347 5951 5381
rect 6003 5334 6037 5368
rect 6383 5326 6417 5360
rect 6555 5326 6589 5360
rect 6659 5328 6693 5362
rect 6743 5347 6777 5381
rect 6950 5332 6984 5366
rect 7185 5332 7219 5366
rect 7253 5332 7287 5366
rect 7337 5332 7371 5366
rect 7487 5321 7521 5355
rect 7751 5321 7785 5355
rect 7855 5328 7889 5362
rect 7939 5347 7973 5381
rect 8146 5332 8180 5366
rect 8381 5332 8415 5366
rect 8449 5332 8483 5366
rect 8533 5332 8567 5366
rect 8683 5321 8717 5355
rect 8947 5321 8981 5355
rect 9143 5344 9177 5378
rect 9143 5276 9177 5310
rect 9227 5347 9261 5381
rect 9331 5343 9365 5377
rect 9331 5275 9365 5309
rect 9423 5279 9457 5313
rect 9507 5347 9541 5381
rect 9591 5343 9625 5377
rect 9591 5275 9625 5309
rect 9695 5328 9729 5362
rect 10327 5328 10361 5362
rect 10431 5328 10465 5362
rect 10515 5347 10549 5381
rect 10722 5332 10756 5366
rect 10957 5332 10991 5366
rect 11025 5332 11059 5366
rect 11109 5332 11143 5366
rect 11535 5328 11569 5362
rect 12535 5328 12569 5362
rect 12639 5321 12673 5355
rect 12903 5321 12937 5355
rect 13099 5328 13133 5362
rect 13183 5347 13217 5381
rect 13390 5332 13424 5366
rect 13625 5332 13659 5366
rect 13693 5332 13727 5366
rect 13777 5332 13811 5366
rect 13927 5328 13961 5362
rect 14927 5328 14961 5362
rect 15031 5328 15065 5362
rect 16031 5328 16065 5362
rect 16135 5321 16169 5355
rect 16399 5321 16433 5355
rect 16687 5328 16721 5362
rect 17687 5328 17721 5362
rect 17791 5328 17825 5362
rect 18423 5328 18457 5362
rect 18619 5326 18653 5360
rect 18791 5326 18825 5360
rect 1139 4432 1173 4466
rect 1311 4432 1345 4466
rect 1415 4430 1449 4464
rect 1863 4430 1897 4464
rect 2059 4437 2093 4471
rect 2143 4411 2177 4445
rect 2227 4437 2261 4471
rect 2331 4411 2365 4445
rect 2416 4425 2450 4459
rect 2527 4425 2561 4459
rect 2726 4419 2760 4453
rect 2845 4425 2879 4459
rect 2948 4425 2982 4459
rect 3146 4425 3180 4459
rect 3251 4480 3285 4514
rect 3251 4412 3285 4446
rect 3335 4441 3369 4475
rect 3419 4482 3453 4516
rect 3419 4414 3453 4448
rect 4035 4411 4069 4445
rect 4119 4411 4153 4445
rect 4311 4439 4345 4473
rect 4451 4437 4485 4471
rect 4715 4437 4749 4471
rect 4911 4482 4945 4516
rect 4911 4414 4945 4448
rect 4995 4411 5029 4445
rect 5099 4483 5133 4517
rect 5099 4415 5133 4449
rect 5191 4479 5225 4513
rect 5275 4411 5309 4445
rect 5359 4483 5393 4517
rect 5359 4415 5393 4449
rect 5463 4437 5497 4471
rect 5727 4437 5761 4471
rect 5831 4482 5865 4516
rect 5831 4414 5865 4448
rect 5915 4411 5949 4445
rect 6019 4483 6053 4517
rect 6019 4415 6053 4449
rect 6111 4479 6145 4513
rect 6195 4411 6229 4445
rect 6279 4483 6313 4517
rect 6279 4415 6313 4449
rect 6383 4437 6417 4471
rect 6647 4437 6681 4471
rect 6751 4437 6785 4471
rect 6835 4411 6869 4445
rect 6919 4437 6953 4471
rect 7023 4411 7057 4445
rect 7108 4425 7142 4459
rect 7219 4425 7253 4459
rect 7418 4419 7452 4453
rect 7537 4425 7571 4459
rect 7640 4425 7674 4459
rect 7838 4425 7872 4459
rect 7943 4480 7977 4514
rect 7943 4412 7977 4446
rect 8027 4441 8061 4475
rect 8111 4482 8145 4516
rect 8111 4414 8145 4448
rect 8223 4430 8257 4464
rect 8671 4430 8705 4464
rect 8959 4430 8993 4464
rect 9591 4430 9625 4464
rect 9695 4432 9729 4466
rect 9867 4432 9901 4466
rect 9979 4482 10013 4516
rect 9979 4414 10013 4448
rect 10063 4441 10097 4475
rect 10147 4480 10181 4514
rect 10147 4412 10181 4446
rect 10252 4425 10286 4459
rect 10450 4425 10484 4459
rect 10553 4425 10587 4459
rect 10672 4419 10706 4453
rect 10871 4425 10905 4459
rect 10982 4425 11016 4459
rect 11067 4411 11101 4445
rect 11171 4437 11205 4471
rect 11255 4411 11289 4445
rect 11339 4437 11373 4471
rect 11443 4437 11477 4471
rect 11707 4437 11741 4471
rect 11811 4482 11845 4516
rect 11811 4414 11845 4448
rect 11895 4411 11929 4445
rect 11999 4483 12033 4517
rect 11999 4415 12033 4449
rect 12091 4479 12125 4513
rect 12175 4411 12209 4445
rect 12259 4483 12293 4517
rect 12259 4415 12293 4449
rect 12363 4437 12397 4471
rect 12627 4437 12661 4471
rect 12731 4482 12765 4516
rect 12731 4414 12765 4448
rect 12815 4411 12849 4445
rect 12919 4483 12953 4517
rect 12919 4415 12953 4449
rect 13011 4479 13045 4513
rect 13095 4411 13129 4445
rect 13179 4483 13213 4517
rect 13179 4415 13213 4449
rect 13283 4430 13317 4464
rect 13915 4430 13949 4464
rect 14111 4432 14145 4466
rect 14283 4432 14317 4466
rect 14423 4439 14457 4473
rect 14615 4411 14649 4445
rect 14699 4411 14733 4445
rect 14847 4430 14881 4464
rect 15847 4430 15881 4464
rect 15951 4430 15985 4464
rect 16951 4430 16985 4464
rect 17055 4430 17089 4464
rect 18055 4430 18089 4464
rect 18159 4437 18193 4471
rect 18423 4437 18457 4471
rect 18619 4432 18653 4466
rect 18791 4432 18825 4466
rect 1139 4238 1173 4272
rect 1311 4238 1345 4272
rect 1415 4240 1449 4274
rect 1863 4240 1897 4274
rect 1967 4246 2001 4280
rect 2053 4259 2087 4293
rect 2139 4229 2173 4263
rect 2243 4233 2277 4267
rect 2507 4233 2541 4267
rect 2619 4256 2653 4290
rect 2619 4188 2653 4222
rect 2703 4229 2737 4263
rect 2787 4258 2821 4292
rect 2787 4190 2821 4224
rect 2892 4245 2926 4279
rect 3090 4245 3124 4279
rect 3193 4245 3227 4279
rect 3312 4251 3346 4285
rect 3511 4245 3545 4279
rect 3622 4245 3656 4279
rect 3707 4259 3741 4293
rect 3811 4233 3845 4267
rect 3895 4259 3929 4293
rect 3979 4233 4013 4267
rect 4083 4240 4117 4274
rect 4531 4240 4565 4274
rect 4643 4256 4677 4290
rect 4643 4188 4677 4222
rect 4727 4229 4761 4263
rect 4811 4258 4845 4292
rect 4811 4190 4845 4224
rect 4916 4245 4950 4279
rect 5114 4245 5148 4279
rect 5217 4245 5251 4279
rect 5336 4251 5370 4285
rect 5535 4245 5569 4279
rect 5646 4245 5680 4279
rect 5731 4259 5765 4293
rect 5835 4233 5869 4267
rect 5919 4259 5953 4293
rect 6003 4233 6037 4267
rect 6383 4240 6417 4274
rect 6831 4240 6865 4274
rect 6935 4256 6969 4290
rect 6935 4188 6969 4222
rect 7019 4259 7053 4293
rect 7123 4255 7157 4289
rect 7123 4187 7157 4221
rect 7215 4191 7249 4225
rect 7299 4259 7333 4293
rect 7383 4255 7417 4289
rect 7383 4187 7417 4221
rect 7487 4233 7521 4267
rect 7751 4233 7785 4267
rect 7855 4259 7889 4293
rect 7941 4246 7975 4280
rect 8027 4246 8061 4280
rect 8113 4246 8147 4280
rect 8199 4246 8233 4280
rect 8285 4246 8319 4280
rect 8371 4255 8405 4289
rect 8457 4246 8491 4280
rect 8543 4255 8577 4289
rect 8629 4246 8663 4280
rect 8715 4255 8749 4289
rect 8801 4246 8835 4280
rect 8887 4255 8921 4289
rect 8972 4246 9006 4280
rect 9058 4255 9092 4289
rect 9144 4246 9178 4280
rect 9230 4255 9264 4289
rect 9316 4246 9350 4280
rect 9402 4255 9436 4289
rect 9488 4246 9522 4280
rect 9574 4255 9608 4289
rect 9695 4240 9729 4274
rect 10327 4240 10361 4274
rect 10523 4256 10557 4290
rect 10523 4188 10557 4222
rect 10607 4259 10641 4293
rect 10711 4255 10745 4289
rect 10711 4187 10745 4221
rect 10803 4191 10837 4225
rect 10887 4259 10921 4293
rect 10971 4255 11005 4289
rect 10971 4187 11005 4221
rect 11075 4233 11109 4267
rect 11339 4233 11373 4267
rect 11719 4233 11753 4267
rect 11803 4259 11837 4293
rect 11887 4233 11921 4267
rect 11991 4259 12025 4293
rect 12076 4245 12110 4279
rect 12187 4245 12221 4279
rect 12386 4251 12420 4285
rect 12505 4245 12539 4279
rect 12608 4245 12642 4279
rect 12806 4245 12840 4279
rect 12911 4258 12945 4292
rect 12911 4190 12945 4224
rect 12995 4229 13029 4263
rect 13079 4256 13113 4290
rect 13079 4188 13113 4222
rect 13191 4240 13225 4274
rect 14191 4240 14225 4274
rect 14295 4240 14329 4274
rect 15295 4240 15329 4274
rect 15491 4229 15525 4263
rect 15577 4259 15611 4293
rect 15663 4246 15697 4280
rect 15767 4240 15801 4274
rect 16399 4240 16433 4274
rect 16907 4231 16941 4265
rect 17099 4259 17133 4293
rect 17183 4259 17217 4293
rect 17331 4240 17365 4274
rect 18331 4240 18365 4274
rect 18619 4238 18653 4272
rect 18791 4238 18825 4272
rect 1139 3344 1173 3378
rect 1311 3344 1345 3378
rect 1415 3342 1449 3376
rect 1863 3342 1897 3376
rect 2059 3349 2093 3383
rect 2143 3323 2177 3357
rect 2227 3349 2261 3383
rect 2331 3323 2365 3357
rect 2416 3337 2450 3371
rect 2527 3337 2561 3371
rect 2726 3331 2760 3365
rect 2845 3337 2879 3371
rect 2948 3337 2982 3371
rect 3146 3337 3180 3371
rect 3251 3392 3285 3426
rect 3251 3324 3285 3358
rect 3335 3353 3369 3387
rect 3419 3394 3453 3428
rect 3419 3326 3453 3360
rect 3991 3349 4025 3383
rect 4075 3323 4109 3357
rect 4159 3349 4193 3383
rect 4263 3323 4297 3357
rect 4348 3337 4382 3371
rect 4459 3337 4493 3371
rect 4658 3331 4692 3365
rect 4777 3337 4811 3371
rect 4880 3337 4914 3371
rect 5078 3337 5112 3371
rect 5183 3392 5217 3426
rect 5183 3324 5217 3358
rect 5267 3353 5301 3387
rect 5351 3394 5385 3428
rect 5351 3326 5385 3360
rect 5463 3342 5497 3376
rect 6095 3342 6129 3376
rect 6291 3394 6325 3428
rect 6291 3326 6325 3360
rect 6375 3323 6409 3357
rect 6479 3395 6513 3429
rect 6479 3327 6513 3361
rect 6571 3391 6605 3425
rect 6655 3323 6689 3357
rect 6739 3395 6773 3429
rect 6739 3327 6773 3361
rect 6843 3349 6877 3383
rect 7107 3349 7141 3383
rect 7211 3349 7245 3383
rect 7295 3323 7329 3357
rect 7379 3349 7413 3383
rect 7483 3323 7517 3357
rect 7568 3337 7602 3371
rect 7679 3337 7713 3371
rect 7878 3331 7912 3365
rect 7997 3337 8031 3371
rect 8100 3337 8134 3371
rect 8298 3337 8332 3371
rect 8403 3392 8437 3426
rect 8403 3324 8437 3358
rect 8487 3353 8521 3387
rect 8571 3394 8605 3428
rect 8571 3326 8605 3360
rect 8959 3342 8993 3376
rect 9591 3342 9625 3376
rect 9787 3349 9821 3383
rect 9871 3323 9905 3357
rect 9955 3349 9989 3383
rect 10059 3323 10093 3357
rect 10144 3337 10178 3371
rect 10255 3337 10289 3371
rect 10454 3331 10488 3365
rect 10573 3337 10607 3371
rect 10676 3337 10710 3371
rect 10874 3337 10908 3371
rect 10979 3392 11013 3426
rect 10979 3324 11013 3358
rect 11063 3353 11097 3387
rect 11147 3394 11181 3428
rect 11147 3326 11181 3360
rect 11259 3342 11293 3376
rect 11707 3342 11741 3376
rect 11811 3349 11845 3383
rect 11895 3323 11929 3357
rect 11979 3349 12013 3383
rect 12083 3323 12117 3357
rect 12168 3337 12202 3371
rect 12279 3337 12313 3371
rect 12478 3331 12512 3365
rect 12597 3337 12631 3371
rect 12700 3337 12734 3371
rect 12898 3337 12932 3371
rect 13003 3392 13037 3426
rect 13003 3324 13037 3358
rect 13087 3353 13121 3387
rect 13171 3394 13205 3428
rect 13171 3326 13205 3360
rect 13283 3342 13317 3376
rect 13915 3342 13949 3376
rect 14111 3342 14145 3376
rect 15111 3342 15145 3376
rect 15215 3342 15249 3376
rect 15663 3342 15697 3376
rect 15767 3353 15801 3387
rect 15853 3323 15887 3357
rect 15939 3336 15973 3370
rect 16043 3349 16077 3383
rect 16307 3349 16341 3383
rect 16455 3323 16489 3357
rect 16539 3323 16573 3357
rect 16731 3351 16765 3385
rect 16871 3349 16905 3383
rect 17135 3349 17169 3383
rect 17283 3323 17317 3357
rect 17367 3323 17401 3357
rect 17559 3351 17593 3385
rect 17699 3342 17733 3376
rect 18331 3342 18365 3376
rect 18619 3344 18653 3378
rect 18791 3344 18825 3378
rect 1139 3150 1173 3184
rect 1311 3150 1345 3184
rect 1415 3145 1449 3179
rect 1679 3145 1713 3179
rect 1875 3163 1909 3197
rect 1961 3167 1995 3201
rect 2055 3163 2089 3197
rect 2139 3167 2173 3201
rect 2243 3145 2277 3179
rect 2507 3145 2541 3179
rect 2628 3167 2662 3201
rect 2714 3158 2748 3192
rect 2800 3167 2834 3201
rect 2886 3158 2920 3192
rect 2972 3167 3006 3201
rect 3058 3158 3092 3192
rect 3144 3167 3178 3201
rect 3230 3158 3264 3192
rect 3315 3167 3349 3201
rect 3401 3158 3435 3192
rect 3487 3167 3521 3201
rect 3573 3158 3607 3192
rect 3659 3167 3693 3201
rect 3745 3158 3779 3192
rect 3831 3167 3865 3201
rect 3917 3158 3951 3192
rect 4003 3158 4037 3192
rect 4089 3158 4123 3192
rect 4175 3158 4209 3192
rect 4261 3158 4295 3192
rect 4347 3171 4381 3205
rect 4451 3152 4485 3186
rect 5451 3152 5485 3186
rect 5555 3152 5589 3186
rect 6187 3152 6221 3186
rect 6383 3152 6417 3186
rect 7015 3152 7049 3186
rect 7395 3145 7429 3179
rect 7659 3145 7693 3179
rect 7763 3171 7797 3205
rect 7849 3158 7883 3192
rect 7935 3158 7969 3192
rect 8021 3158 8055 3192
rect 8107 3158 8141 3192
rect 8193 3158 8227 3192
rect 8279 3167 8313 3201
rect 8365 3158 8399 3192
rect 8451 3167 8485 3201
rect 8537 3158 8571 3192
rect 8623 3167 8657 3201
rect 8709 3158 8743 3192
rect 8795 3167 8829 3201
rect 8880 3158 8914 3192
rect 8966 3167 9000 3201
rect 9052 3158 9086 3192
rect 9138 3167 9172 3201
rect 9224 3158 9258 3192
rect 9310 3167 9344 3201
rect 9396 3158 9430 3192
rect 9482 3167 9516 3201
rect 9603 3152 9637 3186
rect 10603 3152 10637 3186
rect 10707 3152 10741 3186
rect 11339 3152 11373 3186
rect 11719 3145 11753 3179
rect 11803 3171 11837 3205
rect 11887 3145 11921 3179
rect 11991 3171 12025 3205
rect 12076 3157 12110 3191
rect 12187 3157 12221 3191
rect 12386 3163 12420 3197
rect 12505 3157 12539 3191
rect 12608 3157 12642 3191
rect 12806 3157 12840 3191
rect 12911 3170 12945 3204
rect 12911 3102 12945 3136
rect 12995 3141 13029 3175
rect 13079 3168 13113 3202
rect 13079 3100 13113 3134
rect 13191 3152 13225 3186
rect 14191 3152 14225 3186
rect 14295 3152 14329 3186
rect 15295 3152 15329 3186
rect 15399 3152 15433 3186
rect 16399 3152 16433 3186
rect 16871 3141 16905 3175
rect 16957 3171 16991 3205
rect 17043 3158 17077 3192
rect 17147 3152 17181 3186
rect 18147 3152 18181 3186
rect 18251 3145 18285 3179
rect 18515 3145 18549 3179
rect 18619 3150 18653 3184
rect 18791 3150 18825 3184
rect 1139 2256 1173 2290
rect 1311 2256 1345 2290
rect 1415 2254 1449 2288
rect 1863 2254 1897 2288
rect 2067 2306 2101 2340
rect 2067 2238 2101 2272
rect 2151 2265 2185 2299
rect 2235 2304 2269 2338
rect 2235 2236 2269 2270
rect 2340 2249 2374 2283
rect 2538 2249 2572 2283
rect 2641 2249 2675 2283
rect 2760 2243 2794 2277
rect 2959 2249 2993 2283
rect 3070 2249 3104 2283
rect 3155 2235 3189 2269
rect 3259 2261 3293 2295
rect 3343 2235 3377 2269
rect 3427 2261 3461 2295
rect 4175 2261 4209 2295
rect 4439 2261 4473 2295
rect 4635 2261 4669 2295
rect 4719 2235 4753 2269
rect 4803 2261 4837 2295
rect 4907 2235 4941 2269
rect 4992 2249 5026 2283
rect 5103 2249 5137 2283
rect 5302 2243 5336 2277
rect 5421 2249 5455 2283
rect 5524 2249 5558 2283
rect 5722 2249 5756 2283
rect 5827 2304 5861 2338
rect 5827 2236 5861 2270
rect 5911 2265 5945 2299
rect 5995 2306 6029 2340
rect 5995 2238 6029 2272
rect 6383 2254 6417 2288
rect 7015 2254 7049 2288
rect 7219 2306 7253 2340
rect 7219 2238 7253 2272
rect 7303 2265 7337 2299
rect 7387 2304 7421 2338
rect 7387 2236 7421 2270
rect 7492 2249 7526 2283
rect 7690 2249 7724 2283
rect 7793 2249 7827 2283
rect 7912 2243 7946 2277
rect 8111 2249 8145 2283
rect 8222 2249 8256 2283
rect 8307 2235 8341 2269
rect 8411 2261 8445 2295
rect 8495 2235 8529 2269
rect 8579 2261 8613 2295
rect 8959 2254 8993 2288
rect 9591 2254 9625 2288
rect 9787 2261 9821 2295
rect 9871 2235 9905 2269
rect 9955 2261 9989 2295
rect 10059 2235 10093 2269
rect 10144 2249 10178 2283
rect 10255 2249 10289 2283
rect 10454 2243 10488 2277
rect 10573 2249 10607 2283
rect 10676 2249 10710 2283
rect 10874 2249 10908 2283
rect 10979 2304 11013 2338
rect 10979 2236 11013 2270
rect 11063 2265 11097 2299
rect 11147 2306 11181 2340
rect 11147 2238 11181 2272
rect 11535 2261 11569 2295
rect 11799 2261 11833 2295
rect 11911 2306 11945 2340
rect 11911 2238 11945 2272
rect 11995 2265 12029 2299
rect 12079 2304 12113 2338
rect 12079 2236 12113 2270
rect 12184 2249 12218 2283
rect 12382 2249 12416 2283
rect 12485 2249 12519 2283
rect 12604 2243 12638 2277
rect 12803 2249 12837 2283
rect 12914 2249 12948 2283
rect 12999 2235 13033 2269
rect 13103 2261 13137 2295
rect 13187 2235 13221 2269
rect 13271 2261 13305 2295
rect 13375 2254 13409 2288
rect 13823 2254 13857 2288
rect 14571 2254 14605 2288
rect 15571 2254 15605 2288
rect 15675 2254 15709 2288
rect 16307 2254 16341 2288
rect 16871 2265 16905 2299
rect 16957 2235 16991 2269
rect 17043 2248 17077 2282
rect 17147 2261 17181 2295
rect 17411 2261 17445 2295
rect 17515 2248 17549 2282
rect 17608 2235 17642 2269
rect 17694 2265 17728 2299
rect 17778 2307 17812 2341
rect 17778 2239 17812 2273
rect 17883 2254 17917 2288
rect 18515 2254 18549 2288
rect 18619 2256 18653 2290
rect 18791 2256 18825 2290
<< pdiffc >>
rect 1139 7226 1173 7260
rect 1139 7131 1173 7165
rect 1311 7226 1345 7260
rect 1311 7131 1345 7165
rect 1600 7267 1634 7301
rect 1600 7199 1634 7233
rect 1600 7131 1634 7165
rect 1684 7236 1718 7270
rect 1684 7155 1718 7189
rect 1770 7207 1804 7241
rect 1770 7139 1804 7173
rect 1863 7207 1897 7241
rect 1863 7139 1897 7173
rect 1967 7131 2001 7165
rect 2967 7131 3001 7165
rect 3071 7233 3105 7267
rect 3071 7131 3105 7165
rect 3519 7233 3553 7267
rect 3519 7131 3553 7165
rect 3992 7267 4026 7301
rect 3992 7199 4026 7233
rect 3992 7131 4026 7165
rect 4076 7236 4110 7270
rect 4076 7155 4110 7189
rect 4162 7207 4196 7241
rect 4162 7139 4196 7173
rect 4255 7207 4289 7241
rect 4255 7139 4289 7173
rect 4359 7131 4393 7165
rect 5359 7131 5393 7165
rect 5648 7267 5682 7301
rect 5648 7199 5682 7233
rect 5648 7131 5682 7165
rect 5732 7236 5766 7270
rect 5732 7155 5766 7189
rect 5818 7207 5852 7241
rect 5818 7139 5852 7173
rect 5911 7207 5945 7241
rect 5911 7139 5945 7173
rect 6015 7226 6049 7260
rect 6015 7131 6049 7165
rect 6187 7226 6221 7260
rect 6187 7131 6221 7165
rect 6383 7131 6417 7165
rect 7383 7131 7417 7165
rect 7487 7233 7521 7267
rect 7487 7131 7521 7165
rect 7751 7233 7785 7267
rect 7751 7131 7785 7165
rect 7855 7207 7889 7241
rect 7855 7139 7889 7173
rect 7948 7207 7982 7241
rect 7948 7139 7982 7173
rect 8034 7236 8068 7270
rect 8034 7155 8068 7189
rect 8118 7267 8152 7301
rect 8118 7199 8152 7233
rect 8118 7131 8152 7165
rect 8223 7233 8257 7267
rect 8223 7131 8257 7165
rect 8671 7233 8705 7267
rect 8671 7131 8705 7165
rect 8959 7233 8993 7267
rect 8959 7131 8993 7165
rect 9407 7233 9441 7267
rect 9407 7131 9441 7165
rect 9695 7233 9729 7267
rect 9695 7131 9729 7165
rect 9959 7233 9993 7267
rect 9959 7131 9993 7165
rect 10063 7250 10097 7284
rect 10063 7145 10097 7179
rect 10149 7211 10183 7245
rect 10149 7143 10183 7177
rect 10243 7145 10277 7179
rect 10327 7140 10361 7174
rect 10431 7233 10465 7267
rect 10431 7131 10465 7165
rect 11063 7233 11097 7267
rect 11063 7131 11097 7165
rect 11167 7226 11201 7260
rect 11167 7131 11201 7165
rect 11339 7226 11373 7260
rect 11339 7131 11373 7165
rect 11535 7233 11569 7267
rect 11535 7131 11569 7165
rect 12167 7233 12201 7267
rect 12167 7131 12201 7165
rect 12271 7207 12305 7241
rect 12271 7139 12305 7173
rect 12364 7207 12398 7241
rect 12364 7139 12398 7173
rect 12450 7236 12484 7270
rect 12450 7155 12484 7189
rect 12534 7267 12568 7301
rect 12534 7199 12568 7233
rect 12534 7131 12568 7165
rect 12639 7131 12673 7165
rect 13639 7131 13673 7165
rect 13743 7226 13777 7260
rect 13743 7131 13777 7165
rect 13915 7226 13949 7260
rect 13915 7131 13949 7165
rect 14111 7233 14145 7267
rect 14111 7131 14145 7165
rect 14375 7233 14409 7267
rect 14375 7131 14409 7165
rect 14479 7207 14513 7241
rect 14479 7139 14513 7173
rect 14572 7207 14606 7241
rect 14572 7139 14606 7173
rect 14658 7236 14692 7270
rect 14658 7155 14692 7189
rect 14742 7267 14776 7301
rect 14742 7199 14776 7233
rect 14742 7131 14776 7165
rect 14847 7131 14881 7165
rect 15847 7131 15881 7165
rect 15951 7233 15985 7267
rect 15951 7131 15985 7165
rect 16399 7233 16433 7267
rect 16399 7131 16433 7165
rect 16871 7207 16905 7241
rect 16871 7139 16905 7173
rect 16964 7207 16998 7241
rect 16964 7139 16998 7173
rect 17050 7236 17084 7270
rect 17050 7155 17084 7189
rect 17134 7267 17168 7301
rect 17134 7199 17168 7233
rect 17134 7131 17168 7165
rect 17239 7233 17273 7267
rect 17239 7131 17273 7165
rect 17871 7233 17905 7267
rect 17871 7131 17905 7165
rect 18067 7207 18101 7241
rect 18067 7139 18101 7173
rect 18160 7207 18194 7241
rect 18160 7139 18194 7173
rect 18246 7236 18280 7270
rect 18246 7155 18280 7189
rect 18330 7267 18364 7301
rect 18330 7199 18364 7233
rect 18330 7131 18364 7165
rect 18619 7226 18653 7260
rect 18619 7131 18653 7165
rect 18791 7226 18825 7260
rect 18791 7131 18825 7165
rect 1139 6979 1173 7013
rect 1139 6884 1173 6918
rect 1311 6979 1345 7013
rect 1311 6884 1345 6918
rect 1415 6979 1449 7013
rect 2415 6979 2449 7013
rect 2519 6979 2553 7013
rect 3519 6979 3553 7013
rect 3807 6979 3841 7013
rect 4807 6979 4841 7013
rect 4911 6979 4945 7013
rect 5911 6979 5945 7013
rect 6015 6979 6049 7013
rect 7015 6979 7049 7013
rect 7119 6979 7153 7013
rect 8119 6979 8153 7013
rect 8223 6979 8257 7013
rect 8223 6877 8257 6911
rect 8671 6979 8705 7013
rect 8671 6877 8705 6911
rect 8959 6979 8993 7013
rect 9959 6979 9993 7013
rect 10063 6979 10097 7013
rect 11063 6979 11097 7013
rect 11167 6979 11201 7013
rect 12167 6979 12201 7013
rect 12271 6979 12305 7013
rect 13271 6979 13305 7013
rect 13375 6979 13409 7013
rect 13375 6877 13409 6911
rect 13823 6979 13857 7013
rect 13823 6877 13857 6911
rect 14111 6979 14145 7013
rect 15111 6979 15145 7013
rect 15215 6979 15249 7013
rect 16215 6979 16249 7013
rect 16319 6979 16353 7013
rect 17319 6979 17353 7013
rect 17423 6979 17457 7013
rect 18423 6979 18457 7013
rect 18619 6979 18653 7013
rect 18619 6884 18653 6918
rect 18791 6979 18825 7013
rect 18791 6884 18825 6918
rect 1139 6138 1173 6172
rect 1139 6043 1173 6077
rect 1311 6138 1345 6172
rect 1311 6043 1345 6077
rect 1415 6043 1449 6077
rect 2415 6043 2449 6077
rect 2519 6043 2553 6077
rect 3519 6043 3553 6077
rect 3623 6043 3657 6077
rect 4623 6043 4657 6077
rect 4727 6043 4761 6077
rect 5727 6043 5761 6077
rect 5831 6145 5865 6179
rect 5831 6043 5865 6077
rect 6095 6145 6129 6179
rect 6095 6043 6129 6077
rect 6383 6043 6417 6077
rect 7383 6043 7417 6077
rect 7487 6043 7521 6077
rect 8487 6043 8521 6077
rect 8591 6043 8625 6077
rect 9591 6043 9625 6077
rect 9695 6043 9729 6077
rect 10695 6043 10729 6077
rect 10799 6145 10833 6179
rect 10799 6043 10833 6077
rect 11247 6145 11281 6179
rect 11247 6043 11281 6077
rect 11535 6043 11569 6077
rect 12535 6043 12569 6077
rect 12639 6043 12673 6077
rect 13639 6043 13673 6077
rect 13743 6043 13777 6077
rect 14743 6043 14777 6077
rect 14847 6043 14881 6077
rect 15847 6043 15881 6077
rect 15951 6145 15985 6179
rect 15951 6043 15985 6077
rect 16399 6145 16433 6179
rect 16399 6043 16433 6077
rect 16687 6043 16721 6077
rect 17687 6043 17721 6077
rect 17791 6145 17825 6179
rect 17791 6043 17825 6077
rect 18423 6145 18457 6179
rect 18423 6043 18457 6077
rect 18619 6138 18653 6172
rect 18619 6043 18653 6077
rect 18791 6138 18825 6172
rect 18791 6043 18825 6077
rect 1139 5891 1173 5925
rect 1139 5796 1173 5830
rect 1311 5891 1345 5925
rect 1311 5796 1345 5830
rect 1415 5891 1449 5925
rect 1415 5789 1449 5823
rect 2047 5891 2081 5925
rect 2047 5789 2081 5823
rect 2243 5883 2277 5917
rect 2243 5815 2277 5849
rect 2329 5883 2363 5917
rect 2329 5815 2363 5849
rect 2415 5883 2449 5917
rect 2415 5802 2449 5836
rect 2519 5891 2553 5925
rect 2519 5789 2553 5823
rect 2967 5891 3001 5925
rect 2967 5789 3001 5823
rect 3071 5883 3105 5917
rect 3071 5802 3105 5836
rect 3157 5883 3191 5917
rect 3157 5815 3191 5849
rect 3243 5883 3277 5917
rect 3243 5815 3277 5849
rect 3347 5891 3381 5925
rect 3347 5789 3381 5823
rect 3611 5891 3645 5925
rect 3611 5789 3645 5823
rect 3807 5891 3841 5925
rect 4807 5891 4841 5925
rect 4911 5891 4945 5925
rect 5911 5891 5945 5925
rect 6015 5891 6049 5925
rect 6015 5789 6049 5823
rect 6647 5891 6681 5925
rect 6647 5789 6681 5823
rect 6751 5891 6785 5925
rect 6751 5823 6785 5857
rect 6751 5755 6785 5789
rect 6835 5891 6869 5925
rect 6835 5823 6869 5857
rect 7071 5831 7105 5865
rect 7146 5831 7180 5865
rect 7343 5831 7377 5865
rect 7429 5831 7463 5865
rect 7579 5891 7613 5925
rect 6835 5755 6869 5789
rect 8579 5891 8613 5925
rect 8959 5891 8993 5925
rect 8959 5789 8993 5823
rect 9591 5891 9625 5925
rect 9591 5789 9625 5823
rect 9879 5891 9913 5925
rect 9879 5823 9913 5857
rect 9879 5755 9913 5789
rect 9963 5891 9997 5925
rect 9963 5823 9997 5857
rect 10199 5831 10233 5865
rect 10274 5831 10308 5865
rect 10471 5831 10505 5865
rect 10557 5831 10591 5865
rect 10707 5891 10741 5925
rect 9963 5755 9997 5789
rect 10707 5789 10741 5823
rect 10971 5891 11005 5925
rect 10971 5789 11005 5823
rect 11099 5891 11133 5925
rect 11099 5823 11133 5857
rect 11203 5891 11237 5925
rect 11203 5823 11237 5857
rect 11311 5849 11345 5883
rect 11395 5849 11429 5883
rect 11535 5891 11569 5925
rect 11535 5789 11569 5823
rect 12167 5891 12201 5925
rect 12167 5789 12201 5823
rect 12271 5891 12305 5925
rect 12271 5823 12305 5857
rect 12271 5755 12305 5789
rect 12355 5891 12389 5925
rect 12355 5823 12389 5857
rect 12591 5831 12625 5865
rect 12666 5831 12700 5865
rect 12863 5831 12897 5865
rect 12949 5831 12983 5865
rect 13099 5891 13133 5925
rect 12355 5755 12389 5789
rect 13099 5789 13133 5823
rect 13731 5891 13765 5925
rect 13731 5789 13765 5823
rect 14295 5891 14329 5925
rect 14295 5823 14329 5857
rect 14295 5755 14329 5789
rect 14379 5891 14413 5925
rect 14379 5823 14413 5857
rect 14615 5831 14649 5865
rect 14690 5831 14724 5865
rect 14887 5831 14921 5865
rect 14973 5831 15007 5865
rect 15123 5891 15157 5925
rect 14379 5755 14413 5789
rect 16123 5891 16157 5925
rect 16227 5891 16261 5925
rect 17227 5891 17261 5925
rect 17331 5891 17365 5925
rect 18331 5891 18365 5925
rect 18619 5891 18653 5925
rect 18619 5796 18653 5830
rect 18791 5891 18825 5925
rect 18791 5796 18825 5830
rect 1139 5050 1173 5084
rect 1139 4955 1173 4989
rect 1311 5050 1345 5084
rect 1311 4955 1345 4989
rect 1415 5057 1449 5091
rect 1415 4955 1449 4989
rect 1863 5057 1897 5091
rect 1863 4955 1897 4989
rect 1991 5023 2025 5057
rect 1991 4955 2025 4989
rect 2095 5023 2129 5057
rect 2095 4955 2129 4989
rect 2203 4997 2237 5031
rect 2287 4997 2321 5031
rect 2427 5057 2461 5091
rect 2427 4955 2461 4989
rect 2691 5057 2725 5091
rect 2691 4955 2725 4989
rect 2911 5023 2945 5057
rect 2911 4955 2945 4989
rect 3015 5023 3049 5057
rect 3015 4955 3049 4989
rect 3123 4997 3157 5031
rect 3207 4997 3241 5031
rect 3347 5057 3381 5091
rect 3347 4955 3381 4989
rect 3611 5057 3645 5091
rect 3611 4955 3645 4989
rect 3715 5031 3749 5065
rect 3715 4963 3749 4997
rect 3808 5031 3842 5065
rect 3808 4963 3842 4997
rect 3894 5060 3928 5094
rect 3894 4979 3928 5013
rect 3978 5091 4012 5125
rect 3978 5023 4012 5057
rect 3978 4955 4012 4989
rect 4083 5057 4117 5091
rect 4083 4955 4117 4989
rect 4347 5057 4381 5091
rect 4347 4955 4381 4989
rect 4453 5091 4487 5125
rect 4453 5023 4487 5057
rect 4453 4955 4487 4989
rect 4537 5091 4571 5125
rect 4537 5023 4571 5057
rect 4537 4955 4571 4989
rect 4621 5091 4655 5125
rect 4621 5023 4655 5057
rect 4621 4955 4655 4989
rect 4727 4955 4761 4989
rect 5727 4955 5761 4989
rect 5831 5044 5865 5078
rect 5831 4963 5865 4997
rect 5917 5031 5951 5065
rect 5917 4963 5951 4997
rect 6003 5031 6037 5065
rect 6003 4963 6037 4997
rect 6383 5050 6417 5084
rect 6383 4955 6417 4989
rect 6555 5050 6589 5084
rect 6555 4955 6589 4989
rect 6659 5091 6693 5125
rect 6659 5023 6693 5057
rect 6659 4955 6693 4989
rect 6743 5091 6777 5125
rect 6743 5023 6777 5057
rect 6743 4955 6777 4989
rect 6979 5015 7013 5049
rect 7054 5015 7088 5049
rect 7251 5015 7285 5049
rect 7337 5015 7371 5049
rect 7487 5057 7521 5091
rect 7487 4955 7521 4989
rect 7751 5057 7785 5091
rect 7751 4955 7785 4989
rect 7855 5091 7889 5125
rect 7855 5023 7889 5057
rect 7855 4955 7889 4989
rect 7939 5091 7973 5125
rect 7939 5023 7973 5057
rect 7939 4955 7973 4989
rect 8175 5015 8209 5049
rect 8250 5015 8284 5049
rect 8447 5015 8481 5049
rect 8533 5015 8567 5049
rect 8683 5057 8717 5091
rect 8683 4955 8717 4989
rect 8947 5057 8981 5091
rect 8947 4955 8981 4989
rect 9147 5099 9181 5133
rect 9147 5031 9181 5065
rect 9147 4963 9181 4997
rect 9233 5023 9267 5057
rect 9307 5023 9341 5057
rect 9233 4955 9267 4989
rect 9307 4955 9341 4989
rect 9407 5091 9441 5125
rect 9407 5023 9441 5057
rect 9407 4955 9441 4989
rect 9591 5023 9625 5057
rect 9591 4955 9625 4989
rect 9695 5057 9729 5091
rect 9695 4955 9729 4989
rect 10327 5057 10361 5091
rect 10327 4955 10361 4989
rect 10431 5091 10465 5125
rect 10431 5023 10465 5057
rect 10431 4955 10465 4989
rect 10515 5091 10549 5125
rect 10515 5023 10549 5057
rect 10515 4955 10549 4989
rect 10751 5015 10785 5049
rect 10826 5015 10860 5049
rect 11023 5015 11057 5049
rect 11109 5015 11143 5049
rect 11535 4955 11569 4989
rect 12535 4955 12569 4989
rect 12639 5057 12673 5091
rect 12639 4955 12673 4989
rect 12903 5057 12937 5091
rect 12903 4955 12937 4989
rect 13099 5091 13133 5125
rect 13099 5023 13133 5057
rect 13099 4955 13133 4989
rect 13183 5091 13217 5125
rect 13183 5023 13217 5057
rect 13183 4955 13217 4989
rect 13419 5015 13453 5049
rect 13494 5015 13528 5049
rect 13691 5015 13725 5049
rect 13777 5015 13811 5049
rect 13927 4955 13961 4989
rect 14927 4955 14961 4989
rect 15031 4955 15065 4989
rect 16031 4955 16065 4989
rect 16135 5057 16169 5091
rect 16135 4955 16169 4989
rect 16399 5057 16433 5091
rect 16399 4955 16433 4989
rect 16687 4955 16721 4989
rect 17687 4955 17721 4989
rect 17791 5057 17825 5091
rect 17791 4955 17825 4989
rect 18423 5057 18457 5091
rect 18423 4955 18457 4989
rect 18619 5050 18653 5084
rect 18619 4955 18653 4989
rect 18791 5050 18825 5084
rect 18791 4955 18825 4989
rect 1139 4803 1173 4837
rect 1139 4708 1173 4742
rect 1311 4803 1345 4837
rect 1311 4708 1345 4742
rect 1415 4803 1449 4837
rect 1415 4701 1449 4735
rect 1863 4803 1897 4837
rect 1863 4701 1897 4735
rect 2059 4795 2093 4829
rect 2059 4727 2093 4761
rect 2143 4779 2177 4813
rect 2227 4795 2261 4829
rect 2331 4803 2365 4837
rect 2415 4795 2449 4829
rect 2507 4790 2541 4824
rect 2746 4803 2780 4837
rect 2227 4727 2261 4761
rect 2746 4735 2780 4769
rect 2830 4795 2864 4829
rect 2925 4785 2959 4819
rect 3124 4795 3158 4829
rect 3247 4803 3281 4837
rect 3247 4732 3281 4766
rect 3247 4661 3281 4695
rect 3333 4773 3367 4807
rect 3333 4693 3367 4727
rect 3417 4797 3451 4831
rect 3417 4729 3451 4763
rect 3417 4661 3451 4695
rect 4015 4803 4049 4837
rect 4015 4735 4049 4769
rect 4119 4803 4153 4837
rect 4119 4735 4153 4769
rect 4227 4761 4261 4795
rect 4311 4761 4345 4795
rect 4451 4803 4485 4837
rect 4451 4701 4485 4735
rect 4715 4803 4749 4837
rect 4715 4701 4749 4735
rect 4915 4795 4949 4829
rect 4915 4727 4949 4761
rect 4915 4659 4949 4693
rect 5001 4803 5035 4837
rect 5075 4803 5109 4837
rect 5001 4735 5035 4769
rect 5075 4735 5109 4769
rect 5175 4803 5209 4837
rect 5175 4735 5209 4769
rect 5175 4667 5209 4701
rect 5359 4803 5393 4837
rect 5359 4735 5393 4769
rect 5463 4803 5497 4837
rect 5463 4701 5497 4735
rect 5727 4803 5761 4837
rect 5727 4701 5761 4735
rect 5835 4795 5869 4829
rect 5835 4727 5869 4761
rect 5835 4659 5869 4693
rect 5921 4803 5955 4837
rect 5995 4803 6029 4837
rect 5921 4735 5955 4769
rect 5995 4735 6029 4769
rect 6095 4803 6129 4837
rect 6095 4735 6129 4769
rect 6095 4667 6129 4701
rect 6279 4803 6313 4837
rect 6279 4735 6313 4769
rect 6383 4803 6417 4837
rect 6383 4701 6417 4735
rect 6647 4803 6681 4837
rect 6647 4701 6681 4735
rect 6751 4795 6785 4829
rect 6751 4727 6785 4761
rect 6835 4779 6869 4813
rect 6919 4795 6953 4829
rect 7023 4803 7057 4837
rect 7107 4795 7141 4829
rect 7199 4790 7233 4824
rect 7438 4803 7472 4837
rect 6919 4727 6953 4761
rect 7438 4735 7472 4769
rect 7522 4795 7556 4829
rect 7617 4785 7651 4819
rect 7816 4795 7850 4829
rect 7939 4803 7973 4837
rect 7939 4732 7973 4766
rect 7939 4661 7973 4695
rect 8025 4773 8059 4807
rect 8025 4693 8059 4727
rect 8109 4797 8143 4831
rect 8109 4729 8143 4763
rect 8109 4661 8143 4695
rect 8223 4803 8257 4837
rect 8223 4701 8257 4735
rect 8671 4803 8705 4837
rect 8671 4701 8705 4735
rect 8959 4803 8993 4837
rect 8959 4701 8993 4735
rect 9591 4803 9625 4837
rect 9591 4701 9625 4735
rect 9695 4803 9729 4837
rect 9695 4708 9729 4742
rect 9867 4803 9901 4837
rect 9867 4708 9901 4742
rect 9981 4797 10015 4831
rect 9981 4729 10015 4763
rect 9981 4661 10015 4695
rect 10065 4773 10099 4807
rect 10065 4693 10099 4727
rect 10151 4803 10185 4837
rect 10151 4732 10185 4766
rect 10274 4795 10308 4829
rect 10473 4785 10507 4819
rect 10568 4795 10602 4829
rect 10151 4661 10185 4695
rect 10652 4803 10686 4837
rect 10652 4735 10686 4769
rect 10891 4790 10925 4824
rect 10983 4795 11017 4829
rect 11067 4803 11101 4837
rect 11171 4795 11205 4829
rect 11171 4727 11205 4761
rect 11255 4779 11289 4813
rect 11339 4795 11373 4829
rect 11339 4727 11373 4761
rect 11443 4803 11477 4837
rect 11443 4701 11477 4735
rect 11707 4803 11741 4837
rect 11707 4701 11741 4735
rect 11815 4795 11849 4829
rect 11815 4727 11849 4761
rect 11815 4659 11849 4693
rect 11901 4803 11935 4837
rect 11975 4803 12009 4837
rect 11901 4735 11935 4769
rect 11975 4735 12009 4769
rect 12075 4803 12109 4837
rect 12075 4735 12109 4769
rect 12075 4667 12109 4701
rect 12259 4803 12293 4837
rect 12259 4735 12293 4769
rect 12363 4803 12397 4837
rect 12363 4701 12397 4735
rect 12627 4803 12661 4837
rect 12627 4701 12661 4735
rect 12735 4795 12769 4829
rect 12735 4727 12769 4761
rect 12735 4659 12769 4693
rect 12821 4803 12855 4837
rect 12895 4803 12929 4837
rect 12821 4735 12855 4769
rect 12895 4735 12929 4769
rect 12995 4803 13029 4837
rect 12995 4735 13029 4769
rect 12995 4667 13029 4701
rect 13179 4803 13213 4837
rect 13179 4735 13213 4769
rect 13283 4803 13317 4837
rect 13283 4701 13317 4735
rect 13915 4803 13949 4837
rect 13915 4701 13949 4735
rect 14111 4803 14145 4837
rect 14111 4708 14145 4742
rect 14283 4803 14317 4837
rect 14283 4708 14317 4742
rect 14423 4761 14457 4795
rect 14507 4761 14541 4795
rect 14615 4803 14649 4837
rect 14615 4735 14649 4769
rect 14719 4803 14753 4837
rect 14719 4735 14753 4769
rect 14847 4803 14881 4837
rect 15847 4803 15881 4837
rect 15951 4803 15985 4837
rect 16951 4803 16985 4837
rect 17055 4803 17089 4837
rect 18055 4803 18089 4837
rect 18159 4803 18193 4837
rect 18159 4701 18193 4735
rect 18423 4803 18457 4837
rect 18423 4701 18457 4735
rect 18619 4803 18653 4837
rect 18619 4708 18653 4742
rect 18791 4803 18825 4837
rect 18791 4708 18825 4742
rect 1139 3962 1173 3996
rect 1139 3867 1173 3901
rect 1311 3962 1345 3996
rect 1311 3867 1345 3901
rect 1415 3969 1449 4003
rect 1415 3867 1449 3901
rect 1863 3969 1897 4003
rect 1863 3867 1897 3901
rect 1967 3943 2001 3977
rect 1967 3875 2001 3909
rect 2053 3943 2087 3977
rect 2053 3875 2087 3909
rect 2139 3956 2173 3990
rect 2139 3875 2173 3909
rect 2243 3969 2277 4003
rect 2243 3867 2277 3901
rect 2507 3969 2541 4003
rect 2507 3867 2541 3901
rect 2621 4009 2655 4043
rect 2621 3941 2655 3975
rect 2621 3873 2655 3907
rect 2705 3977 2739 4011
rect 2705 3897 2739 3931
rect 2791 4009 2825 4043
rect 2791 3938 2825 3972
rect 2791 3867 2825 3901
rect 2914 3875 2948 3909
rect 3113 3885 3147 3919
rect 3208 3875 3242 3909
rect 3292 3935 3326 3969
rect 3811 3943 3845 3977
rect 3292 3867 3326 3901
rect 3531 3880 3565 3914
rect 3623 3875 3657 3909
rect 3707 3867 3741 3901
rect 3811 3875 3845 3909
rect 3895 3891 3929 3925
rect 3979 3943 4013 3977
rect 3979 3875 4013 3909
rect 4083 3969 4117 4003
rect 4083 3867 4117 3901
rect 4531 3969 4565 4003
rect 4531 3867 4565 3901
rect 4645 4009 4679 4043
rect 4645 3941 4679 3975
rect 4645 3873 4679 3907
rect 4729 3977 4763 4011
rect 4729 3897 4763 3931
rect 4815 4009 4849 4043
rect 4815 3938 4849 3972
rect 4815 3867 4849 3901
rect 4938 3875 4972 3909
rect 5137 3885 5171 3919
rect 5232 3875 5266 3909
rect 5316 3935 5350 3969
rect 5835 3943 5869 3977
rect 5316 3867 5350 3901
rect 5555 3880 5589 3914
rect 5647 3875 5681 3909
rect 5731 3867 5765 3901
rect 5835 3875 5869 3909
rect 5919 3891 5953 3925
rect 6003 3943 6037 3977
rect 6003 3875 6037 3909
rect 6383 3969 6417 4003
rect 6383 3867 6417 3901
rect 6831 3969 6865 4003
rect 6831 3867 6865 3901
rect 6939 4011 6973 4045
rect 6939 3943 6973 3977
rect 6939 3875 6973 3909
rect 7025 3935 7059 3969
rect 7099 3935 7133 3969
rect 7025 3867 7059 3901
rect 7099 3867 7133 3901
rect 7199 4003 7233 4037
rect 7199 3935 7233 3969
rect 7199 3867 7233 3901
rect 7383 3935 7417 3969
rect 7383 3867 7417 3901
rect 7487 3969 7521 4003
rect 7487 3867 7521 3901
rect 7751 3969 7785 4003
rect 7751 3867 7785 3901
rect 7855 3935 7889 3969
rect 7855 3867 7889 3901
rect 7941 3943 7975 3977
rect 7941 3875 7975 3909
rect 8027 3935 8061 3969
rect 8027 3867 8061 3901
rect 8113 3951 8147 3985
rect 8113 3883 8147 3917
rect 8199 3935 8233 3969
rect 8199 3867 8233 3901
rect 8285 3997 8319 4031
rect 8285 3911 8319 3945
rect 8371 3891 8405 3925
rect 8457 3997 8491 4031
rect 8457 3911 8491 3945
rect 8543 3891 8577 3925
rect 8629 3997 8663 4031
rect 8629 3911 8663 3945
rect 8715 3891 8749 3925
rect 8801 3997 8835 4031
rect 8801 3911 8835 3945
rect 8887 3891 8921 3925
rect 8972 3997 9006 4031
rect 8972 3911 9006 3945
rect 9058 3891 9092 3925
rect 9144 3997 9178 4031
rect 9144 3911 9178 3945
rect 9230 3891 9264 3925
rect 9316 3997 9350 4031
rect 9316 3911 9350 3945
rect 9402 3891 9436 3925
rect 9488 3997 9522 4031
rect 9488 3911 9522 3945
rect 9574 3891 9608 3925
rect 9695 3969 9729 4003
rect 9695 3867 9729 3901
rect 10327 3969 10361 4003
rect 10327 3867 10361 3901
rect 10527 4011 10561 4045
rect 10527 3943 10561 3977
rect 10527 3875 10561 3909
rect 10613 3935 10647 3969
rect 10687 3935 10721 3969
rect 10613 3867 10647 3901
rect 10687 3867 10721 3901
rect 10787 4003 10821 4037
rect 10787 3935 10821 3969
rect 10787 3867 10821 3901
rect 10971 3935 11005 3969
rect 10971 3867 11005 3901
rect 11075 3969 11109 4003
rect 11075 3867 11109 3901
rect 11339 3969 11373 4003
rect 11339 3867 11373 3901
rect 11719 3943 11753 3977
rect 11719 3875 11753 3909
rect 11803 3891 11837 3925
rect 11887 3943 11921 3977
rect 11887 3875 11921 3909
rect 11991 3867 12025 3901
rect 12075 3875 12109 3909
rect 12167 3880 12201 3914
rect 12406 3935 12440 3969
rect 12406 3867 12440 3901
rect 12907 4009 12941 4043
rect 12490 3875 12524 3909
rect 12585 3885 12619 3919
rect 12784 3875 12818 3909
rect 12907 3938 12941 3972
rect 12907 3867 12941 3901
rect 12993 3977 13027 4011
rect 12993 3897 13027 3931
rect 13077 4009 13111 4043
rect 13077 3941 13111 3975
rect 13077 3873 13111 3907
rect 13191 3867 13225 3901
rect 14191 3867 14225 3901
rect 14295 3867 14329 3901
rect 15295 3867 15329 3901
rect 15491 3956 15525 3990
rect 15491 3875 15525 3909
rect 15577 3943 15611 3977
rect 15577 3875 15611 3909
rect 15663 3943 15697 3977
rect 15663 3875 15697 3909
rect 15767 3969 15801 4003
rect 15767 3867 15801 3901
rect 16399 3969 16433 4003
rect 16399 3867 16433 3901
rect 16907 3909 16941 3943
rect 16991 3909 17025 3943
rect 17099 3935 17133 3969
rect 17099 3867 17133 3901
rect 17203 3935 17237 3969
rect 17203 3867 17237 3901
rect 17331 3867 17365 3901
rect 18331 3867 18365 3901
rect 18619 3962 18653 3996
rect 18619 3867 18653 3901
rect 18791 3962 18825 3996
rect 18791 3867 18825 3901
rect 1139 3715 1173 3749
rect 1139 3620 1173 3654
rect 1311 3715 1345 3749
rect 1311 3620 1345 3654
rect 1415 3715 1449 3749
rect 1415 3613 1449 3647
rect 1863 3715 1897 3749
rect 1863 3613 1897 3647
rect 2059 3707 2093 3741
rect 2059 3639 2093 3673
rect 2143 3691 2177 3725
rect 2227 3707 2261 3741
rect 2331 3715 2365 3749
rect 2415 3707 2449 3741
rect 2507 3702 2541 3736
rect 2746 3715 2780 3749
rect 2227 3639 2261 3673
rect 2746 3647 2780 3681
rect 2830 3707 2864 3741
rect 2925 3697 2959 3731
rect 3124 3707 3158 3741
rect 3247 3715 3281 3749
rect 3247 3644 3281 3678
rect 3247 3573 3281 3607
rect 3333 3685 3367 3719
rect 3333 3605 3367 3639
rect 3417 3709 3451 3743
rect 3417 3641 3451 3675
rect 3417 3573 3451 3607
rect 3991 3707 4025 3741
rect 3991 3639 4025 3673
rect 4075 3691 4109 3725
rect 4159 3707 4193 3741
rect 4263 3715 4297 3749
rect 4347 3707 4381 3741
rect 4439 3702 4473 3736
rect 4678 3715 4712 3749
rect 4159 3639 4193 3673
rect 4678 3647 4712 3681
rect 4762 3707 4796 3741
rect 4857 3697 4891 3731
rect 5056 3707 5090 3741
rect 5179 3715 5213 3749
rect 5179 3644 5213 3678
rect 5179 3573 5213 3607
rect 5265 3685 5299 3719
rect 5265 3605 5299 3639
rect 5349 3709 5383 3743
rect 5349 3641 5383 3675
rect 5349 3573 5383 3607
rect 5463 3715 5497 3749
rect 5463 3613 5497 3647
rect 6095 3715 6129 3749
rect 6095 3613 6129 3647
rect 6295 3707 6329 3741
rect 6295 3639 6329 3673
rect 6295 3571 6329 3605
rect 6381 3715 6415 3749
rect 6455 3715 6489 3749
rect 6381 3647 6415 3681
rect 6455 3647 6489 3681
rect 6555 3715 6589 3749
rect 6555 3647 6589 3681
rect 6555 3579 6589 3613
rect 6739 3715 6773 3749
rect 6739 3647 6773 3681
rect 6843 3715 6877 3749
rect 6843 3613 6877 3647
rect 7107 3715 7141 3749
rect 7107 3613 7141 3647
rect 7211 3707 7245 3741
rect 7211 3639 7245 3673
rect 7295 3691 7329 3725
rect 7379 3707 7413 3741
rect 7483 3715 7517 3749
rect 7567 3707 7601 3741
rect 7659 3702 7693 3736
rect 7898 3715 7932 3749
rect 7379 3639 7413 3673
rect 7898 3647 7932 3681
rect 7982 3707 8016 3741
rect 8077 3697 8111 3731
rect 8276 3707 8310 3741
rect 8399 3715 8433 3749
rect 8399 3644 8433 3678
rect 8399 3573 8433 3607
rect 8485 3685 8519 3719
rect 8485 3605 8519 3639
rect 8569 3709 8603 3743
rect 8569 3641 8603 3675
rect 8569 3573 8603 3607
rect 8959 3715 8993 3749
rect 8959 3613 8993 3647
rect 9591 3715 9625 3749
rect 9591 3613 9625 3647
rect 9787 3707 9821 3741
rect 9787 3639 9821 3673
rect 9871 3691 9905 3725
rect 9955 3707 9989 3741
rect 10059 3715 10093 3749
rect 10143 3707 10177 3741
rect 10235 3702 10269 3736
rect 10474 3715 10508 3749
rect 9955 3639 9989 3673
rect 10474 3647 10508 3681
rect 10558 3707 10592 3741
rect 10653 3697 10687 3731
rect 10852 3707 10886 3741
rect 10975 3715 11009 3749
rect 10975 3644 11009 3678
rect 10975 3573 11009 3607
rect 11061 3685 11095 3719
rect 11061 3605 11095 3639
rect 11145 3709 11179 3743
rect 11145 3641 11179 3675
rect 11145 3573 11179 3607
rect 11259 3715 11293 3749
rect 11259 3613 11293 3647
rect 11707 3715 11741 3749
rect 11707 3613 11741 3647
rect 11811 3707 11845 3741
rect 11811 3639 11845 3673
rect 11895 3691 11929 3725
rect 11979 3707 12013 3741
rect 12083 3715 12117 3749
rect 12167 3707 12201 3741
rect 12259 3702 12293 3736
rect 12498 3715 12532 3749
rect 11979 3639 12013 3673
rect 12498 3647 12532 3681
rect 12582 3707 12616 3741
rect 12677 3697 12711 3731
rect 12876 3707 12910 3741
rect 12999 3715 13033 3749
rect 12999 3644 13033 3678
rect 12999 3573 13033 3607
rect 13085 3685 13119 3719
rect 13085 3605 13119 3639
rect 13169 3709 13203 3743
rect 13169 3641 13203 3675
rect 13169 3573 13203 3607
rect 13283 3715 13317 3749
rect 13283 3613 13317 3647
rect 13915 3715 13949 3749
rect 13915 3613 13949 3647
rect 14111 3715 14145 3749
rect 15111 3715 15145 3749
rect 15215 3715 15249 3749
rect 15215 3613 15249 3647
rect 15663 3715 15697 3749
rect 15663 3613 15697 3647
rect 15767 3707 15801 3741
rect 15767 3626 15801 3660
rect 15853 3707 15887 3741
rect 15853 3639 15887 3673
rect 15939 3707 15973 3741
rect 15939 3639 15973 3673
rect 16043 3715 16077 3749
rect 16043 3613 16077 3647
rect 16307 3715 16341 3749
rect 16307 3613 16341 3647
rect 16435 3715 16469 3749
rect 16435 3647 16469 3681
rect 16539 3715 16573 3749
rect 16539 3647 16573 3681
rect 16647 3673 16681 3707
rect 16731 3673 16765 3707
rect 16871 3715 16905 3749
rect 16871 3613 16905 3647
rect 17135 3715 17169 3749
rect 17135 3613 17169 3647
rect 17263 3715 17297 3749
rect 17263 3647 17297 3681
rect 17367 3715 17401 3749
rect 17367 3647 17401 3681
rect 17475 3673 17509 3707
rect 17559 3673 17593 3707
rect 17699 3715 17733 3749
rect 17699 3613 17733 3647
rect 18331 3715 18365 3749
rect 18331 3613 18365 3647
rect 18619 3715 18653 3749
rect 18619 3620 18653 3654
rect 18791 3715 18825 3749
rect 18791 3620 18825 3654
rect 1139 2874 1173 2908
rect 1139 2779 1173 2813
rect 1311 2874 1345 2908
rect 1311 2779 1345 2813
rect 1415 2881 1449 2915
rect 1415 2779 1449 2813
rect 1679 2881 1713 2915
rect 1679 2779 1713 2813
rect 1875 2898 1909 2932
rect 1875 2793 1909 2827
rect 1961 2859 1995 2893
rect 1961 2791 1995 2825
rect 2055 2793 2089 2827
rect 2139 2788 2173 2822
rect 2243 2881 2277 2915
rect 2243 2779 2277 2813
rect 2507 2881 2541 2915
rect 2507 2779 2541 2813
rect 2628 2803 2662 2837
rect 2714 2909 2748 2943
rect 2714 2823 2748 2857
rect 2800 2803 2834 2837
rect 2886 2909 2920 2943
rect 2886 2823 2920 2857
rect 2972 2803 3006 2837
rect 3058 2909 3092 2943
rect 3058 2823 3092 2857
rect 3144 2803 3178 2837
rect 3230 2909 3264 2943
rect 3230 2823 3264 2857
rect 3315 2803 3349 2837
rect 3401 2909 3435 2943
rect 3401 2823 3435 2857
rect 3487 2803 3521 2837
rect 3573 2909 3607 2943
rect 3573 2823 3607 2857
rect 3659 2803 3693 2837
rect 3745 2909 3779 2943
rect 3745 2823 3779 2857
rect 3831 2803 3865 2837
rect 3917 2909 3951 2943
rect 3917 2823 3951 2857
rect 4003 2847 4037 2881
rect 4003 2779 4037 2813
rect 4089 2863 4123 2897
rect 4089 2795 4123 2829
rect 4175 2847 4209 2881
rect 4175 2779 4209 2813
rect 4261 2855 4295 2889
rect 4261 2787 4295 2821
rect 4347 2847 4381 2881
rect 4347 2779 4381 2813
rect 4451 2779 4485 2813
rect 5451 2779 5485 2813
rect 5555 2881 5589 2915
rect 5555 2779 5589 2813
rect 6187 2881 6221 2915
rect 6187 2779 6221 2813
rect 6383 2881 6417 2915
rect 6383 2779 6417 2813
rect 7015 2881 7049 2915
rect 7015 2779 7049 2813
rect 7395 2881 7429 2915
rect 7395 2779 7429 2813
rect 7659 2881 7693 2915
rect 7659 2779 7693 2813
rect 7763 2847 7797 2881
rect 7763 2779 7797 2813
rect 7849 2855 7883 2889
rect 7849 2787 7883 2821
rect 7935 2847 7969 2881
rect 7935 2779 7969 2813
rect 8021 2863 8055 2897
rect 8021 2795 8055 2829
rect 8107 2847 8141 2881
rect 8107 2779 8141 2813
rect 8193 2909 8227 2943
rect 8193 2823 8227 2857
rect 8279 2803 8313 2837
rect 8365 2909 8399 2943
rect 8365 2823 8399 2857
rect 8451 2803 8485 2837
rect 8537 2909 8571 2943
rect 8537 2823 8571 2857
rect 8623 2803 8657 2837
rect 8709 2909 8743 2943
rect 8709 2823 8743 2857
rect 8795 2803 8829 2837
rect 8880 2909 8914 2943
rect 8880 2823 8914 2857
rect 8966 2803 9000 2837
rect 9052 2909 9086 2943
rect 9052 2823 9086 2857
rect 9138 2803 9172 2837
rect 9224 2909 9258 2943
rect 9224 2823 9258 2857
rect 9310 2803 9344 2837
rect 9396 2909 9430 2943
rect 9396 2823 9430 2857
rect 9482 2803 9516 2837
rect 9603 2779 9637 2813
rect 10603 2779 10637 2813
rect 10707 2881 10741 2915
rect 10707 2779 10741 2813
rect 11339 2881 11373 2915
rect 11339 2779 11373 2813
rect 11719 2855 11753 2889
rect 11719 2787 11753 2821
rect 11803 2803 11837 2837
rect 11887 2855 11921 2889
rect 11887 2787 11921 2821
rect 11991 2779 12025 2813
rect 12075 2787 12109 2821
rect 12167 2792 12201 2826
rect 12406 2847 12440 2881
rect 12406 2779 12440 2813
rect 12907 2921 12941 2955
rect 12490 2787 12524 2821
rect 12585 2797 12619 2831
rect 12784 2787 12818 2821
rect 12907 2850 12941 2884
rect 12907 2779 12941 2813
rect 12993 2889 13027 2923
rect 12993 2809 13027 2843
rect 13077 2921 13111 2955
rect 13077 2853 13111 2887
rect 13077 2785 13111 2819
rect 13191 2779 13225 2813
rect 14191 2779 14225 2813
rect 14295 2779 14329 2813
rect 15295 2779 15329 2813
rect 15399 2779 15433 2813
rect 16399 2779 16433 2813
rect 16871 2868 16905 2902
rect 16871 2787 16905 2821
rect 16957 2855 16991 2889
rect 16957 2787 16991 2821
rect 17043 2855 17077 2889
rect 17043 2787 17077 2821
rect 17147 2779 17181 2813
rect 18147 2779 18181 2813
rect 18251 2881 18285 2915
rect 18251 2779 18285 2813
rect 18515 2881 18549 2915
rect 18515 2779 18549 2813
rect 18619 2874 18653 2908
rect 18619 2779 18653 2813
rect 18791 2874 18825 2908
rect 18791 2779 18825 2813
rect 1139 2627 1173 2661
rect 1139 2532 1173 2566
rect 1311 2627 1345 2661
rect 1311 2532 1345 2566
rect 1415 2627 1449 2661
rect 1415 2525 1449 2559
rect 1863 2627 1897 2661
rect 1863 2525 1897 2559
rect 2069 2621 2103 2655
rect 2069 2553 2103 2587
rect 2069 2485 2103 2519
rect 2153 2597 2187 2631
rect 2153 2517 2187 2551
rect 2239 2627 2273 2661
rect 2239 2556 2273 2590
rect 2362 2619 2396 2653
rect 2561 2609 2595 2643
rect 2656 2619 2690 2653
rect 2239 2485 2273 2519
rect 2740 2627 2774 2661
rect 2740 2559 2774 2593
rect 2979 2614 3013 2648
rect 3071 2619 3105 2653
rect 3155 2627 3189 2661
rect 3259 2619 3293 2653
rect 3259 2551 3293 2585
rect 3343 2603 3377 2637
rect 3427 2619 3461 2653
rect 3427 2551 3461 2585
rect 4175 2627 4209 2661
rect 4175 2525 4209 2559
rect 4439 2627 4473 2661
rect 4439 2525 4473 2559
rect 4635 2619 4669 2653
rect 4635 2551 4669 2585
rect 4719 2603 4753 2637
rect 4803 2619 4837 2653
rect 4907 2627 4941 2661
rect 4991 2619 5025 2653
rect 5083 2614 5117 2648
rect 5322 2627 5356 2661
rect 4803 2551 4837 2585
rect 5322 2559 5356 2593
rect 5406 2619 5440 2653
rect 5501 2609 5535 2643
rect 5700 2619 5734 2653
rect 5823 2627 5857 2661
rect 5823 2556 5857 2590
rect 5823 2485 5857 2519
rect 5909 2597 5943 2631
rect 5909 2517 5943 2551
rect 5993 2621 6027 2655
rect 5993 2553 6027 2587
rect 5993 2485 6027 2519
rect 6383 2627 6417 2661
rect 6383 2525 6417 2559
rect 7015 2627 7049 2661
rect 7015 2525 7049 2559
rect 7221 2621 7255 2655
rect 7221 2553 7255 2587
rect 7221 2485 7255 2519
rect 7305 2597 7339 2631
rect 7305 2517 7339 2551
rect 7391 2627 7425 2661
rect 7391 2556 7425 2590
rect 7514 2619 7548 2653
rect 7713 2609 7747 2643
rect 7808 2619 7842 2653
rect 7391 2485 7425 2519
rect 7892 2627 7926 2661
rect 7892 2559 7926 2593
rect 8131 2614 8165 2648
rect 8223 2619 8257 2653
rect 8307 2627 8341 2661
rect 8411 2619 8445 2653
rect 8411 2551 8445 2585
rect 8495 2603 8529 2637
rect 8579 2619 8613 2653
rect 8579 2551 8613 2585
rect 8959 2627 8993 2661
rect 8959 2525 8993 2559
rect 9591 2627 9625 2661
rect 9591 2525 9625 2559
rect 9787 2619 9821 2653
rect 9787 2551 9821 2585
rect 9871 2603 9905 2637
rect 9955 2619 9989 2653
rect 10059 2627 10093 2661
rect 10143 2619 10177 2653
rect 10235 2614 10269 2648
rect 10474 2627 10508 2661
rect 9955 2551 9989 2585
rect 10474 2559 10508 2593
rect 10558 2619 10592 2653
rect 10653 2609 10687 2643
rect 10852 2619 10886 2653
rect 10975 2627 11009 2661
rect 10975 2556 11009 2590
rect 10975 2485 11009 2519
rect 11061 2597 11095 2631
rect 11061 2517 11095 2551
rect 11145 2621 11179 2655
rect 11145 2553 11179 2587
rect 11145 2485 11179 2519
rect 11535 2627 11569 2661
rect 11535 2525 11569 2559
rect 11799 2627 11833 2661
rect 11799 2525 11833 2559
rect 11913 2621 11947 2655
rect 11913 2553 11947 2587
rect 11913 2485 11947 2519
rect 11997 2597 12031 2631
rect 11997 2517 12031 2551
rect 12083 2627 12117 2661
rect 12083 2556 12117 2590
rect 12206 2619 12240 2653
rect 12405 2609 12439 2643
rect 12500 2619 12534 2653
rect 12083 2485 12117 2519
rect 12584 2627 12618 2661
rect 12584 2559 12618 2593
rect 12823 2614 12857 2648
rect 12915 2619 12949 2653
rect 12999 2627 13033 2661
rect 13103 2619 13137 2653
rect 13103 2551 13137 2585
rect 13187 2603 13221 2637
rect 13271 2619 13305 2653
rect 13271 2551 13305 2585
rect 13375 2627 13409 2661
rect 13375 2525 13409 2559
rect 13823 2627 13857 2661
rect 13823 2525 13857 2559
rect 14571 2627 14605 2661
rect 15571 2627 15605 2661
rect 15675 2627 15709 2661
rect 15675 2525 15709 2559
rect 16307 2627 16341 2661
rect 16307 2525 16341 2559
rect 16871 2619 16905 2653
rect 16871 2538 16905 2572
rect 16957 2619 16991 2653
rect 16957 2551 16991 2585
rect 17043 2619 17077 2653
rect 17043 2551 17077 2585
rect 17147 2627 17181 2661
rect 17147 2525 17181 2559
rect 17411 2627 17445 2661
rect 17411 2525 17445 2559
rect 17515 2619 17549 2653
rect 17515 2551 17549 2585
rect 17608 2619 17642 2653
rect 17608 2551 17642 2585
rect 17694 2603 17728 2637
rect 17694 2522 17728 2556
rect 17778 2627 17812 2661
rect 17778 2559 17812 2593
rect 17778 2491 17812 2525
rect 17883 2627 17917 2661
rect 17883 2525 17917 2559
rect 18515 2627 18549 2661
rect 18515 2525 18549 2559
rect 18619 2627 18653 2661
rect 18619 2532 18653 2566
rect 18791 2627 18825 2661
rect 18791 2532 18825 2566
<< psubdiff >>
rect 3709 7505 3743 7552
rect 3709 7447 3743 7471
rect 6285 7505 6319 7552
rect 6285 7447 6319 7471
rect 8861 7505 8895 7552
rect 8861 7447 8895 7471
rect 11437 7505 11471 7552
rect 11437 7447 11471 7471
rect 14013 7505 14047 7552
rect 14013 7447 14047 7471
rect 16589 7505 16623 7552
rect 16589 7447 16623 7471
rect 3709 6673 3743 6697
rect 3709 6592 3743 6639
rect 8861 6673 8895 6697
rect 8861 6592 8895 6639
rect 14013 6673 14047 6697
rect 14013 6592 14047 6639
rect 6285 6417 6319 6464
rect 6285 6359 6319 6383
rect 11437 6417 11471 6464
rect 11437 6359 11471 6383
rect 16589 6417 16623 6464
rect 16589 6359 16623 6383
rect 3709 5585 3743 5609
rect 3709 5504 3743 5551
rect 8861 5585 8895 5609
rect 8861 5504 8895 5551
rect 14013 5585 14047 5609
rect 14013 5504 14047 5551
rect 6285 5329 6319 5376
rect 6285 5271 6319 5295
rect 11437 5329 11471 5376
rect 11437 5271 11471 5295
rect 16589 5329 16623 5376
rect 16589 5271 16623 5295
rect 3709 4497 3743 4521
rect 3709 4416 3743 4463
rect 8861 4497 8895 4521
rect 8861 4416 8895 4463
rect 14013 4497 14047 4521
rect 14013 4416 14047 4463
rect 6285 4241 6319 4288
rect 6285 4183 6319 4207
rect 11437 4241 11471 4288
rect 11437 4183 11471 4207
rect 16589 4241 16623 4288
rect 16589 4183 16623 4207
rect 3709 3409 3743 3433
rect 3709 3328 3743 3375
rect 8861 3409 8895 3433
rect 8861 3328 8895 3375
rect 14013 3409 14047 3433
rect 14013 3328 14047 3375
rect 6285 3153 6319 3200
rect 6285 3095 6319 3119
rect 11437 3153 11471 3200
rect 11437 3095 11471 3119
rect 16589 3153 16623 3200
rect 16589 3095 16623 3119
rect 3709 2321 3743 2345
rect 3709 2240 3743 2287
rect 6285 2321 6319 2345
rect 6285 2240 6319 2287
rect 8861 2321 8895 2345
rect 8861 2240 8895 2287
rect 11437 2321 11471 2345
rect 11437 2240 11471 2287
rect 14013 2321 14047 2345
rect 14013 2240 14047 2287
rect 16589 2321 16623 2345
rect 16589 2240 16623 2287
<< nsubdiff >>
rect 3709 7287 3743 7311
rect 3709 7194 3743 7253
rect 3709 7136 3743 7160
rect 6285 7287 6319 7311
rect 6285 7194 6319 7253
rect 6285 7136 6319 7160
rect 8861 7287 8895 7311
rect 8861 7194 8895 7253
rect 8861 7136 8895 7160
rect 11437 7287 11471 7311
rect 11437 7194 11471 7253
rect 11437 7136 11471 7160
rect 14013 7287 14047 7311
rect 14013 7194 14047 7253
rect 14013 7136 14047 7160
rect 16589 7287 16623 7311
rect 16589 7194 16623 7253
rect 16589 7136 16623 7160
rect 3709 6984 3743 7008
rect 3709 6891 3743 6950
rect 3709 6833 3743 6857
rect 8861 6984 8895 7008
rect 8861 6891 8895 6950
rect 8861 6833 8895 6857
rect 14013 6984 14047 7008
rect 14013 6891 14047 6950
rect 14013 6833 14047 6857
rect 6285 6199 6319 6223
rect 6285 6106 6319 6165
rect 6285 6048 6319 6072
rect 11437 6199 11471 6223
rect 11437 6106 11471 6165
rect 11437 6048 11471 6072
rect 16589 6199 16623 6223
rect 16589 6106 16623 6165
rect 16589 6048 16623 6072
rect 3709 5896 3743 5920
rect 3709 5803 3743 5862
rect 3709 5745 3743 5769
rect 8861 5896 8895 5920
rect 8861 5803 8895 5862
rect 8861 5745 8895 5769
rect 14013 5896 14047 5920
rect 14013 5803 14047 5862
rect 14013 5745 14047 5769
rect 6285 5111 6319 5135
rect 6285 5018 6319 5077
rect 6285 4960 6319 4984
rect 11437 5111 11471 5135
rect 11437 5018 11471 5077
rect 11437 4960 11471 4984
rect 16589 5111 16623 5135
rect 16589 5018 16623 5077
rect 16589 4960 16623 4984
rect 3709 4808 3743 4832
rect 3709 4715 3743 4774
rect 3709 4657 3743 4681
rect 8861 4808 8895 4832
rect 8861 4715 8895 4774
rect 8861 4657 8895 4681
rect 14013 4808 14047 4832
rect 14013 4715 14047 4774
rect 14013 4657 14047 4681
rect 6285 4023 6319 4047
rect 6285 3930 6319 3989
rect 6285 3872 6319 3896
rect 11437 4023 11471 4047
rect 11437 3930 11471 3989
rect 11437 3872 11471 3896
rect 16589 4023 16623 4047
rect 16589 3930 16623 3989
rect 16589 3872 16623 3896
rect 3709 3720 3743 3744
rect 3709 3627 3743 3686
rect 3709 3569 3743 3593
rect 8861 3720 8895 3744
rect 8861 3627 8895 3686
rect 8861 3569 8895 3593
rect 14013 3720 14047 3744
rect 14013 3627 14047 3686
rect 14013 3569 14047 3593
rect 6285 2935 6319 2959
rect 6285 2842 6319 2901
rect 6285 2784 6319 2808
rect 11437 2935 11471 2959
rect 11437 2842 11471 2901
rect 11437 2784 11471 2808
rect 16589 2935 16623 2959
rect 16589 2842 16623 2901
rect 16589 2784 16623 2808
rect 3709 2632 3743 2656
rect 3709 2539 3743 2598
rect 3709 2481 3743 2505
rect 6285 2632 6319 2656
rect 6285 2539 6319 2598
rect 6285 2481 6319 2505
rect 8861 2632 8895 2656
rect 8861 2539 8895 2598
rect 8861 2481 8895 2505
rect 11437 2632 11471 2656
rect 11437 2539 11471 2598
rect 11437 2481 11471 2505
rect 14013 2632 14047 2656
rect 14013 2539 14047 2598
rect 14013 2481 14047 2505
rect 16589 2632 16623 2656
rect 16589 2539 16623 2598
rect 16589 2481 16623 2505
<< psubdiffcont >>
rect 3709 7471 3743 7505
rect 6285 7471 6319 7505
rect 8861 7471 8895 7505
rect 11437 7471 11471 7505
rect 14013 7471 14047 7505
rect 16589 7471 16623 7505
rect 3709 6639 3743 6673
rect 8861 6639 8895 6673
rect 14013 6639 14047 6673
rect 6285 6383 6319 6417
rect 11437 6383 11471 6417
rect 16589 6383 16623 6417
rect 3709 5551 3743 5585
rect 8861 5551 8895 5585
rect 14013 5551 14047 5585
rect 6285 5295 6319 5329
rect 11437 5295 11471 5329
rect 16589 5295 16623 5329
rect 3709 4463 3743 4497
rect 8861 4463 8895 4497
rect 14013 4463 14047 4497
rect 6285 4207 6319 4241
rect 11437 4207 11471 4241
rect 16589 4207 16623 4241
rect 3709 3375 3743 3409
rect 8861 3375 8895 3409
rect 14013 3375 14047 3409
rect 6285 3119 6319 3153
rect 11437 3119 11471 3153
rect 16589 3119 16623 3153
rect 3709 2287 3743 2321
rect 6285 2287 6319 2321
rect 8861 2287 8895 2321
rect 11437 2287 11471 2321
rect 14013 2287 14047 2321
rect 16589 2287 16623 2321
<< nsubdiffcont >>
rect 3709 7253 3743 7287
rect 3709 7160 3743 7194
rect 6285 7253 6319 7287
rect 6285 7160 6319 7194
rect 8861 7253 8895 7287
rect 8861 7160 8895 7194
rect 11437 7253 11471 7287
rect 11437 7160 11471 7194
rect 14013 7253 14047 7287
rect 14013 7160 14047 7194
rect 16589 7253 16623 7287
rect 16589 7160 16623 7194
rect 3709 6950 3743 6984
rect 3709 6857 3743 6891
rect 8861 6950 8895 6984
rect 8861 6857 8895 6891
rect 14013 6950 14047 6984
rect 14013 6857 14047 6891
rect 6285 6165 6319 6199
rect 6285 6072 6319 6106
rect 11437 6165 11471 6199
rect 11437 6072 11471 6106
rect 16589 6165 16623 6199
rect 16589 6072 16623 6106
rect 3709 5862 3743 5896
rect 3709 5769 3743 5803
rect 8861 5862 8895 5896
rect 8861 5769 8895 5803
rect 14013 5862 14047 5896
rect 14013 5769 14047 5803
rect 6285 5077 6319 5111
rect 6285 4984 6319 5018
rect 11437 5077 11471 5111
rect 11437 4984 11471 5018
rect 16589 5077 16623 5111
rect 16589 4984 16623 5018
rect 3709 4774 3743 4808
rect 3709 4681 3743 4715
rect 8861 4774 8895 4808
rect 8861 4681 8895 4715
rect 14013 4774 14047 4808
rect 14013 4681 14047 4715
rect 6285 3989 6319 4023
rect 6285 3896 6319 3930
rect 11437 3989 11471 4023
rect 11437 3896 11471 3930
rect 16589 3989 16623 4023
rect 16589 3896 16623 3930
rect 3709 3686 3743 3720
rect 3709 3593 3743 3627
rect 8861 3686 8895 3720
rect 8861 3593 8895 3627
rect 14013 3686 14047 3720
rect 14013 3593 14047 3627
rect 6285 2901 6319 2935
rect 6285 2808 6319 2842
rect 11437 2901 11471 2935
rect 11437 2808 11471 2842
rect 16589 2901 16623 2935
rect 16589 2808 16623 2842
rect 3709 2598 3743 2632
rect 3709 2505 3743 2539
rect 6285 2598 6319 2632
rect 6285 2505 6319 2539
rect 8861 2598 8895 2632
rect 8861 2505 8895 2539
rect 11437 2598 11471 2632
rect 11437 2505 11471 2539
rect 14013 2598 14047 2632
rect 14013 2505 14047 2539
rect 16589 2598 16623 2632
rect 16589 2505 16623 2539
<< poly >>
rect 1183 7569 1301 7595
rect 1644 7569 1674 7595
rect 1728 7569 1758 7595
rect 1823 7569 1853 7595
rect 2011 7569 2957 7595
rect 3115 7569 3509 7595
rect 4036 7569 4066 7595
rect 4120 7569 4150 7595
rect 4215 7569 4245 7595
rect 4403 7569 5349 7595
rect 5692 7569 5722 7595
rect 5776 7569 5806 7595
rect 5871 7569 5901 7595
rect 6059 7569 6177 7595
rect 6427 7569 7373 7595
rect 7531 7569 7741 7595
rect 7899 7569 7929 7595
rect 7994 7569 8024 7595
rect 8078 7569 8108 7595
rect 8267 7569 8661 7595
rect 9003 7569 9397 7595
rect 1183 7433 1301 7459
rect 1263 7431 1301 7433
rect 1263 7415 1329 7431
rect 1155 7375 1221 7391
rect 1155 7341 1171 7375
rect 1205 7341 1221 7375
rect 1263 7381 1279 7415
rect 1313 7381 1329 7415
rect 1263 7365 1329 7381
rect 1644 7417 1674 7439
rect 1728 7417 1758 7439
rect 1823 7417 1853 7485
rect 2011 7433 2957 7459
rect 3115 7433 3509 7459
rect 1644 7401 1781 7417
rect 1644 7367 1737 7401
rect 1771 7367 1781 7401
rect 1155 7325 1221 7341
rect 1183 7323 1221 7325
rect 1644 7351 1781 7367
rect 1823 7401 1905 7417
rect 1823 7367 1861 7401
rect 1895 7367 1905 7401
rect 2503 7411 2957 7433
rect 1823 7351 1905 7367
rect 2011 7375 2461 7391
rect 1183 7293 1301 7323
rect 1644 7319 1674 7351
rect 1728 7319 1758 7351
rect 1823 7255 1853 7351
rect 2011 7341 2283 7375
rect 2317 7341 2461 7375
rect 2503 7377 2647 7411
rect 2681 7377 2957 7411
rect 3333 7411 3509 7433
rect 2503 7361 2957 7377
rect 3115 7375 3291 7391
rect 2011 7319 2461 7341
rect 3115 7341 3131 7375
rect 3165 7341 3241 7375
rect 3275 7341 3291 7375
rect 3333 7377 3349 7411
rect 3383 7377 3459 7411
rect 3493 7377 3509 7411
rect 3333 7361 3509 7377
rect 4036 7417 4066 7439
rect 4120 7417 4150 7439
rect 4215 7417 4245 7485
rect 4403 7433 5349 7459
rect 4036 7401 4173 7417
rect 4036 7367 4129 7401
rect 4163 7367 4173 7401
rect 3115 7319 3291 7341
rect 4036 7351 4173 7367
rect 4215 7401 4297 7417
rect 4215 7367 4253 7401
rect 4287 7367 4297 7401
rect 4895 7411 5349 7433
rect 4215 7351 4297 7367
rect 4403 7375 4853 7391
rect 4036 7319 4066 7351
rect 4120 7319 4150 7351
rect 2011 7293 2957 7319
rect 3115 7293 3509 7319
rect 1183 7093 1301 7119
rect 1644 7093 1674 7119
rect 1728 7093 1758 7119
rect 1823 7101 1853 7127
rect 4215 7255 4245 7351
rect 4403 7341 4675 7375
rect 4709 7341 4853 7375
rect 4895 7377 5039 7411
rect 5073 7377 5349 7411
rect 4895 7361 5349 7377
rect 5692 7417 5722 7439
rect 5776 7417 5806 7439
rect 5871 7417 5901 7485
rect 6059 7433 6177 7459
rect 6427 7433 7373 7459
rect 7531 7433 7741 7459
rect 6139 7431 6177 7433
rect 5692 7401 5829 7417
rect 5692 7367 5785 7401
rect 5819 7367 5829 7401
rect 4403 7319 4853 7341
rect 5692 7351 5829 7367
rect 5871 7401 5953 7417
rect 5871 7367 5909 7401
rect 5943 7367 5953 7401
rect 6139 7415 6205 7431
rect 5871 7351 5953 7367
rect 6031 7375 6097 7391
rect 5692 7319 5722 7351
rect 5776 7319 5806 7351
rect 4403 7293 5349 7319
rect 2011 7093 2957 7119
rect 3115 7093 3509 7119
rect 4036 7093 4066 7119
rect 4120 7093 4150 7119
rect 4215 7101 4245 7127
rect 5871 7255 5901 7351
rect 6031 7341 6047 7375
rect 6081 7341 6097 7375
rect 6139 7381 6155 7415
rect 6189 7381 6205 7415
rect 6919 7411 7373 7433
rect 6139 7365 6205 7381
rect 6427 7375 6877 7391
rect 6031 7325 6097 7341
rect 6059 7323 6097 7325
rect 6427 7341 6699 7375
rect 6733 7341 6877 7375
rect 6919 7377 7063 7411
rect 7097 7377 7373 7411
rect 7657 7427 7741 7433
rect 7657 7411 7799 7427
rect 7899 7417 7929 7485
rect 7994 7417 8024 7439
rect 8078 7417 8108 7439
rect 8267 7433 8661 7459
rect 9739 7569 9949 7595
rect 10108 7569 10138 7595
rect 10203 7569 10233 7595
rect 10287 7569 10317 7595
rect 10475 7569 11053 7595
rect 11211 7569 11329 7595
rect 11579 7569 12157 7595
rect 12315 7569 12345 7595
rect 12410 7569 12440 7595
rect 12494 7569 12524 7595
rect 12683 7569 13629 7595
rect 13787 7569 13905 7595
rect 14155 7569 14365 7595
rect 14523 7569 14553 7595
rect 14618 7569 14648 7595
rect 14702 7569 14732 7595
rect 14891 7569 15837 7595
rect 15995 7569 16389 7595
rect 16915 7569 16945 7595
rect 17010 7569 17040 7595
rect 17094 7569 17124 7595
rect 17283 7569 17861 7595
rect 18111 7569 18141 7595
rect 18206 7569 18236 7595
rect 18290 7569 18320 7595
rect 18663 7569 18781 7595
rect 9003 7433 9397 7459
rect 9739 7433 9949 7459
rect 6919 7361 7373 7377
rect 7473 7375 7615 7391
rect 6059 7293 6177 7323
rect 6427 7319 6877 7341
rect 7473 7341 7489 7375
rect 7523 7341 7615 7375
rect 7657 7377 7749 7411
rect 7783 7377 7799 7411
rect 7657 7361 7799 7377
rect 7847 7401 7929 7417
rect 7847 7367 7857 7401
rect 7891 7367 7929 7401
rect 7847 7351 7929 7367
rect 7971 7401 8108 7417
rect 7971 7367 7981 7401
rect 8015 7367 8108 7401
rect 8485 7411 8661 7433
rect 7971 7351 8108 7367
rect 7473 7325 7615 7341
rect 7531 7319 7615 7325
rect 4403 7093 5349 7119
rect 5692 7093 5722 7119
rect 5776 7093 5806 7119
rect 5871 7101 5901 7127
rect 6427 7293 7373 7319
rect 7531 7293 7741 7319
rect 7899 7255 7929 7351
rect 7994 7319 8024 7351
rect 8078 7319 8108 7351
rect 8267 7375 8443 7391
rect 8267 7341 8283 7375
rect 8317 7341 8393 7375
rect 8427 7341 8443 7375
rect 8485 7377 8501 7411
rect 8535 7377 8611 7411
rect 8645 7377 8661 7411
rect 9221 7411 9397 7433
rect 8485 7361 8661 7377
rect 9003 7375 9179 7391
rect 8267 7319 8443 7341
rect 9003 7341 9019 7375
rect 9053 7341 9129 7375
rect 9163 7341 9179 7375
rect 9221 7377 9237 7411
rect 9271 7377 9347 7411
rect 9381 7377 9397 7411
rect 9865 7427 9949 7433
rect 10108 7436 10138 7485
rect 10203 7467 10233 7485
rect 10287 7467 10317 7485
rect 9865 7411 10007 7427
rect 10108 7421 10161 7436
rect 9221 7361 9397 7377
rect 9681 7375 9823 7391
rect 9003 7319 9179 7341
rect 9681 7341 9697 7375
rect 9731 7341 9823 7375
rect 9865 7377 9957 7411
rect 9991 7377 10007 7411
rect 9865 7361 10007 7377
rect 10097 7401 10161 7421
rect 10097 7367 10117 7401
rect 10151 7367 10161 7401
rect 9681 7325 9823 7341
rect 10097 7337 10161 7367
rect 10203 7401 10317 7467
rect 10475 7433 11053 7459
rect 11211 7433 11329 7459
rect 11579 7433 12157 7459
rect 10203 7367 10221 7401
rect 10255 7367 10317 7401
rect 10781 7411 11053 7433
rect 10203 7337 10317 7367
rect 9739 7319 9823 7325
rect 10108 7319 10138 7337
rect 10203 7319 10233 7337
rect 10287 7319 10317 7337
rect 10475 7375 10739 7391
rect 10475 7341 10491 7375
rect 10525 7341 10590 7375
rect 10624 7341 10689 7375
rect 10723 7341 10739 7375
rect 10781 7377 10797 7411
rect 10831 7377 10900 7411
rect 10934 7377 11003 7411
rect 11037 7377 11053 7411
rect 11291 7431 11329 7433
rect 11291 7415 11357 7431
rect 10781 7361 11053 7377
rect 11183 7375 11249 7391
rect 10475 7319 10739 7341
rect 11183 7341 11199 7375
rect 11233 7341 11249 7375
rect 11291 7381 11307 7415
rect 11341 7381 11357 7415
rect 11885 7411 12157 7433
rect 12315 7417 12345 7485
rect 12410 7417 12440 7439
rect 12494 7417 12524 7439
rect 12683 7433 13629 7459
rect 13787 7433 13905 7459
rect 14155 7433 14365 7459
rect 11291 7365 11357 7381
rect 11579 7375 11843 7391
rect 11183 7325 11249 7341
rect 11211 7323 11249 7325
rect 11579 7341 11595 7375
rect 11629 7341 11694 7375
rect 11728 7341 11793 7375
rect 11827 7341 11843 7375
rect 11885 7377 11901 7411
rect 11935 7377 12004 7411
rect 12038 7377 12107 7411
rect 12141 7377 12157 7411
rect 11885 7361 12157 7377
rect 12263 7401 12345 7417
rect 12263 7367 12273 7401
rect 12307 7367 12345 7401
rect 12263 7351 12345 7367
rect 12387 7401 12524 7417
rect 12387 7367 12397 7401
rect 12431 7367 12524 7401
rect 13175 7411 13629 7433
rect 12387 7351 12524 7367
rect 6059 7093 6177 7119
rect 6427 7093 7373 7119
rect 7531 7093 7741 7119
rect 7899 7101 7929 7127
rect 8267 7293 8661 7319
rect 9003 7293 9397 7319
rect 9739 7293 9949 7319
rect 10475 7293 11053 7319
rect 11211 7293 11329 7323
rect 11579 7319 11843 7341
rect 11579 7293 12157 7319
rect 12315 7255 12345 7351
rect 12410 7319 12440 7351
rect 12494 7319 12524 7351
rect 12683 7375 13133 7391
rect 12683 7341 12955 7375
rect 12989 7341 13133 7375
rect 13175 7377 13319 7411
rect 13353 7377 13629 7411
rect 13867 7431 13905 7433
rect 13867 7415 13933 7431
rect 13175 7361 13629 7377
rect 13759 7375 13825 7391
rect 12683 7319 13133 7341
rect 13759 7341 13775 7375
rect 13809 7341 13825 7375
rect 13867 7381 13883 7415
rect 13917 7381 13933 7415
rect 14281 7427 14365 7433
rect 14281 7411 14423 7427
rect 14523 7417 14553 7485
rect 14618 7417 14648 7439
rect 14702 7417 14732 7439
rect 14891 7433 15837 7459
rect 15995 7433 16389 7459
rect 13867 7365 13933 7381
rect 14097 7375 14239 7391
rect 13759 7325 13825 7341
rect 14097 7341 14113 7375
rect 14147 7341 14239 7375
rect 14281 7377 14373 7411
rect 14407 7377 14423 7411
rect 14281 7361 14423 7377
rect 14471 7401 14553 7417
rect 14471 7367 14481 7401
rect 14515 7367 14553 7401
rect 14471 7351 14553 7367
rect 14595 7401 14732 7417
rect 14595 7367 14605 7401
rect 14639 7367 14732 7401
rect 15383 7411 15837 7433
rect 14595 7351 14732 7367
rect 14097 7325 14239 7341
rect 13787 7323 13825 7325
rect 7994 7093 8024 7119
rect 8078 7093 8108 7119
rect 8267 7093 8661 7119
rect 9003 7093 9397 7119
rect 9739 7093 9949 7119
rect 10108 7093 10138 7119
rect 10203 7093 10233 7119
rect 10287 7093 10317 7119
rect 10475 7093 11053 7119
rect 11211 7093 11329 7119
rect 11579 7093 12157 7119
rect 12315 7101 12345 7127
rect 12683 7293 13629 7319
rect 13787 7293 13905 7323
rect 14155 7319 14239 7325
rect 14155 7293 14365 7319
rect 14523 7255 14553 7351
rect 14618 7319 14648 7351
rect 14702 7319 14732 7351
rect 14891 7375 15341 7391
rect 14891 7341 15163 7375
rect 15197 7341 15341 7375
rect 15383 7377 15527 7411
rect 15561 7377 15837 7411
rect 16213 7411 16389 7433
rect 16915 7417 16945 7485
rect 17010 7417 17040 7439
rect 17094 7417 17124 7439
rect 17283 7433 17861 7459
rect 15383 7361 15837 7377
rect 15995 7375 16171 7391
rect 14891 7319 15341 7341
rect 15995 7341 16011 7375
rect 16045 7341 16121 7375
rect 16155 7341 16171 7375
rect 16213 7377 16229 7411
rect 16263 7377 16339 7411
rect 16373 7377 16389 7411
rect 16213 7361 16389 7377
rect 16863 7401 16945 7417
rect 16863 7367 16873 7401
rect 16907 7367 16945 7401
rect 16863 7351 16945 7367
rect 16987 7401 17124 7417
rect 16987 7367 16997 7401
rect 17031 7367 17124 7401
rect 17589 7411 17861 7433
rect 18111 7417 18141 7485
rect 18206 7417 18236 7439
rect 18290 7417 18320 7439
rect 18663 7433 18781 7459
rect 18663 7431 18701 7433
rect 16987 7351 17124 7367
rect 15995 7319 16171 7341
rect 12410 7093 12440 7119
rect 12494 7093 12524 7119
rect 12683 7093 13629 7119
rect 13787 7093 13905 7119
rect 14155 7093 14365 7119
rect 14523 7101 14553 7127
rect 14891 7293 15837 7319
rect 15995 7293 16389 7319
rect 16915 7255 16945 7351
rect 17010 7319 17040 7351
rect 17094 7319 17124 7351
rect 17283 7375 17547 7391
rect 17283 7341 17299 7375
rect 17333 7341 17398 7375
rect 17432 7341 17497 7375
rect 17531 7341 17547 7375
rect 17589 7377 17605 7411
rect 17639 7377 17708 7411
rect 17742 7377 17811 7411
rect 17845 7377 17861 7411
rect 17589 7361 17861 7377
rect 18059 7401 18141 7417
rect 18059 7367 18069 7401
rect 18103 7367 18141 7401
rect 18059 7351 18141 7367
rect 18183 7401 18320 7417
rect 18183 7367 18193 7401
rect 18227 7367 18320 7401
rect 18183 7351 18320 7367
rect 18635 7415 18701 7431
rect 18635 7381 18651 7415
rect 18685 7381 18701 7415
rect 18635 7365 18701 7381
rect 18743 7375 18809 7391
rect 17283 7319 17547 7341
rect 14618 7093 14648 7119
rect 14702 7093 14732 7119
rect 14891 7093 15837 7119
rect 15995 7093 16389 7119
rect 16915 7101 16945 7127
rect 17283 7293 17861 7319
rect 18111 7255 18141 7351
rect 18206 7319 18236 7351
rect 18290 7319 18320 7351
rect 18743 7341 18759 7375
rect 18793 7341 18809 7375
rect 18743 7325 18809 7341
rect 18743 7323 18781 7325
rect 17010 7093 17040 7119
rect 17094 7093 17124 7119
rect 17283 7093 17861 7119
rect 18111 7101 18141 7127
rect 18663 7293 18781 7323
rect 18206 7093 18236 7119
rect 18290 7093 18320 7119
rect 18663 7093 18781 7119
rect 1183 7025 1301 7051
rect 1459 7025 2405 7051
rect 2563 7025 3509 7051
rect 3851 7025 4797 7051
rect 4955 7025 5901 7051
rect 6059 7025 7005 7051
rect 7163 7025 8109 7051
rect 8267 7025 8661 7051
rect 9003 7025 9949 7051
rect 10107 7025 11053 7051
rect 11211 7025 12157 7051
rect 12315 7025 13261 7051
rect 13419 7025 13813 7051
rect 14155 7025 15101 7051
rect 15259 7025 16205 7051
rect 16363 7025 17309 7051
rect 17467 7025 18413 7051
rect 18663 7025 18781 7051
rect 1183 6821 1301 6851
rect 1459 6825 2405 6851
rect 2563 6825 3509 6851
rect 3851 6825 4797 6851
rect 4955 6825 5901 6851
rect 6059 6825 7005 6851
rect 7163 6825 8109 6851
rect 8267 6825 8661 6851
rect 9003 6825 9949 6851
rect 10107 6825 11053 6851
rect 11211 6825 12157 6851
rect 12315 6825 13261 6851
rect 13419 6825 13813 6851
rect 14155 6825 15101 6851
rect 15259 6825 16205 6851
rect 16363 6825 17309 6851
rect 17467 6825 18413 6851
rect 1183 6819 1221 6821
rect 1155 6803 1221 6819
rect 1155 6769 1171 6803
rect 1205 6769 1221 6803
rect 1459 6803 1909 6825
rect 1155 6753 1221 6769
rect 1263 6763 1329 6779
rect 1263 6729 1279 6763
rect 1313 6729 1329 6763
rect 1459 6769 1731 6803
rect 1765 6769 1909 6803
rect 2563 6803 3013 6825
rect 1459 6753 1909 6769
rect 1951 6767 2405 6783
rect 1263 6713 1329 6729
rect 1951 6733 2095 6767
rect 2129 6733 2405 6767
rect 2563 6769 2835 6803
rect 2869 6769 3013 6803
rect 3851 6803 4301 6825
rect 2563 6753 3013 6769
rect 3055 6767 3509 6783
rect 1263 6711 1301 6713
rect 1951 6711 2405 6733
rect 3055 6733 3199 6767
rect 3233 6733 3509 6767
rect 3851 6769 4123 6803
rect 4157 6769 4301 6803
rect 4955 6803 5405 6825
rect 3851 6753 4301 6769
rect 4343 6767 4797 6783
rect 3055 6711 3509 6733
rect 4343 6733 4487 6767
rect 4521 6733 4797 6767
rect 4955 6769 5227 6803
rect 5261 6769 5405 6803
rect 6059 6803 6509 6825
rect 4955 6753 5405 6769
rect 5447 6767 5901 6783
rect 4343 6711 4797 6733
rect 5447 6733 5591 6767
rect 5625 6733 5901 6767
rect 6059 6769 6331 6803
rect 6365 6769 6509 6803
rect 7163 6803 7613 6825
rect 6059 6753 6509 6769
rect 6551 6767 7005 6783
rect 5447 6711 5901 6733
rect 6551 6733 6695 6767
rect 6729 6733 7005 6767
rect 7163 6769 7435 6803
rect 7469 6769 7613 6803
rect 8267 6803 8443 6825
rect 7163 6753 7613 6769
rect 7655 6767 8109 6783
rect 6551 6711 7005 6733
rect 7655 6733 7799 6767
rect 7833 6733 8109 6767
rect 8267 6769 8283 6803
rect 8317 6769 8393 6803
rect 8427 6769 8443 6803
rect 9003 6803 9453 6825
rect 8267 6753 8443 6769
rect 8485 6767 8661 6783
rect 7655 6711 8109 6733
rect 8485 6733 8501 6767
rect 8535 6733 8611 6767
rect 8645 6733 8661 6767
rect 9003 6769 9275 6803
rect 9309 6769 9453 6803
rect 10107 6803 10557 6825
rect 9003 6753 9453 6769
rect 9495 6767 9949 6783
rect 8485 6711 8661 6733
rect 9495 6733 9639 6767
rect 9673 6733 9949 6767
rect 10107 6769 10379 6803
rect 10413 6769 10557 6803
rect 11211 6803 11661 6825
rect 10107 6753 10557 6769
rect 10599 6767 11053 6783
rect 9495 6711 9949 6733
rect 10599 6733 10743 6767
rect 10777 6733 11053 6767
rect 11211 6769 11483 6803
rect 11517 6769 11661 6803
rect 12315 6803 12765 6825
rect 11211 6753 11661 6769
rect 11703 6767 12157 6783
rect 10599 6711 11053 6733
rect 11703 6733 11847 6767
rect 11881 6733 12157 6767
rect 12315 6769 12587 6803
rect 12621 6769 12765 6803
rect 13419 6803 13595 6825
rect 12315 6753 12765 6769
rect 12807 6767 13261 6783
rect 11703 6711 12157 6733
rect 12807 6733 12951 6767
rect 12985 6733 13261 6767
rect 13419 6769 13435 6803
rect 13469 6769 13545 6803
rect 13579 6769 13595 6803
rect 14155 6803 14605 6825
rect 13419 6753 13595 6769
rect 13637 6767 13813 6783
rect 12807 6711 13261 6733
rect 13637 6733 13653 6767
rect 13687 6733 13763 6767
rect 13797 6733 13813 6767
rect 14155 6769 14427 6803
rect 14461 6769 14605 6803
rect 15259 6803 15709 6825
rect 14155 6753 14605 6769
rect 14647 6767 15101 6783
rect 13637 6711 13813 6733
rect 14647 6733 14791 6767
rect 14825 6733 15101 6767
rect 15259 6769 15531 6803
rect 15565 6769 15709 6803
rect 16363 6803 16813 6825
rect 15259 6753 15709 6769
rect 15751 6767 16205 6783
rect 14647 6711 15101 6733
rect 15751 6733 15895 6767
rect 15929 6733 16205 6767
rect 16363 6769 16635 6803
rect 16669 6769 16813 6803
rect 17467 6803 17917 6825
rect 18663 6821 18781 6851
rect 16363 6753 16813 6769
rect 16855 6767 17309 6783
rect 15751 6711 16205 6733
rect 16855 6733 16999 6767
rect 17033 6733 17309 6767
rect 17467 6769 17739 6803
rect 17773 6769 17917 6803
rect 18743 6819 18781 6821
rect 18743 6803 18809 6819
rect 17467 6753 17917 6769
rect 17959 6767 18413 6783
rect 16855 6711 17309 6733
rect 17959 6733 18103 6767
rect 18137 6733 18413 6767
rect 17959 6711 18413 6733
rect 18635 6763 18701 6779
rect 18635 6729 18651 6763
rect 18685 6729 18701 6763
rect 18743 6769 18759 6803
rect 18793 6769 18809 6803
rect 18743 6753 18809 6769
rect 18635 6713 18701 6729
rect 1183 6685 1301 6711
rect 1459 6685 2405 6711
rect 2563 6685 3509 6711
rect 3851 6685 4797 6711
rect 4955 6685 5901 6711
rect 6059 6685 7005 6711
rect 7163 6685 8109 6711
rect 8267 6685 8661 6711
rect 9003 6685 9949 6711
rect 10107 6685 11053 6711
rect 11211 6685 12157 6711
rect 12315 6685 13261 6711
rect 13419 6685 13813 6711
rect 14155 6685 15101 6711
rect 15259 6685 16205 6711
rect 16363 6685 17309 6711
rect 17467 6685 18413 6711
rect 18663 6711 18701 6713
rect 18663 6685 18781 6711
rect 1183 6549 1301 6575
rect 1459 6549 2405 6575
rect 2563 6549 3509 6575
rect 3851 6549 4797 6575
rect 4955 6549 5901 6575
rect 6059 6549 7005 6575
rect 7163 6549 8109 6575
rect 8267 6549 8661 6575
rect 9003 6549 9949 6575
rect 10107 6549 11053 6575
rect 11211 6549 12157 6575
rect 12315 6549 13261 6575
rect 13419 6549 13813 6575
rect 14155 6549 15101 6575
rect 15259 6549 16205 6575
rect 16363 6549 17309 6575
rect 17467 6549 18413 6575
rect 18663 6549 18781 6575
rect 1183 6481 1301 6507
rect 1459 6481 2405 6507
rect 2563 6481 3509 6507
rect 3667 6481 4613 6507
rect 4771 6481 5717 6507
rect 5875 6481 6085 6507
rect 6427 6481 7373 6507
rect 7531 6481 8477 6507
rect 8635 6481 9581 6507
rect 9739 6481 10685 6507
rect 10843 6481 11237 6507
rect 11579 6481 12525 6507
rect 12683 6481 13629 6507
rect 13787 6481 14733 6507
rect 14891 6481 15837 6507
rect 15995 6481 16389 6507
rect 16731 6481 17677 6507
rect 17835 6481 18413 6507
rect 18663 6481 18781 6507
rect 1183 6345 1301 6371
rect 1459 6345 2405 6371
rect 2563 6345 3509 6371
rect 3667 6345 4613 6371
rect 4771 6345 5717 6371
rect 5875 6345 6085 6371
rect 6427 6345 7373 6371
rect 7531 6345 8477 6371
rect 8635 6345 9581 6371
rect 9739 6345 10685 6371
rect 10843 6345 11237 6371
rect 11579 6345 12525 6371
rect 12683 6345 13629 6371
rect 13787 6345 14733 6371
rect 14891 6345 15837 6371
rect 15995 6345 16389 6371
rect 16731 6345 17677 6371
rect 17835 6345 18413 6371
rect 1263 6343 1301 6345
rect 1263 6327 1329 6343
rect 1155 6287 1221 6303
rect 1155 6253 1171 6287
rect 1205 6253 1221 6287
rect 1263 6293 1279 6327
rect 1313 6293 1329 6327
rect 1951 6323 2405 6345
rect 1263 6277 1329 6293
rect 1459 6287 1909 6303
rect 1155 6237 1221 6253
rect 1183 6235 1221 6237
rect 1459 6253 1731 6287
rect 1765 6253 1909 6287
rect 1951 6289 2095 6323
rect 2129 6289 2405 6323
rect 3055 6323 3509 6345
rect 1951 6273 2405 6289
rect 2563 6287 3013 6303
rect 1183 6205 1301 6235
rect 1459 6231 1909 6253
rect 2563 6253 2835 6287
rect 2869 6253 3013 6287
rect 3055 6289 3199 6323
rect 3233 6289 3509 6323
rect 4159 6323 4613 6345
rect 3055 6273 3509 6289
rect 3667 6287 4117 6303
rect 2563 6231 3013 6253
rect 3667 6253 3939 6287
rect 3973 6253 4117 6287
rect 4159 6289 4303 6323
rect 4337 6289 4613 6323
rect 5263 6323 5717 6345
rect 4159 6273 4613 6289
rect 4771 6287 5221 6303
rect 3667 6231 4117 6253
rect 4771 6253 5043 6287
rect 5077 6253 5221 6287
rect 5263 6289 5407 6323
rect 5441 6289 5717 6323
rect 6001 6339 6085 6345
rect 6001 6323 6143 6339
rect 5263 6273 5717 6289
rect 5817 6287 5959 6303
rect 4771 6231 5221 6253
rect 5817 6253 5833 6287
rect 5867 6253 5959 6287
rect 6001 6289 6093 6323
rect 6127 6289 6143 6323
rect 6919 6323 7373 6345
rect 6001 6273 6143 6289
rect 6427 6287 6877 6303
rect 5817 6237 5959 6253
rect 5875 6231 5959 6237
rect 6427 6253 6699 6287
rect 6733 6253 6877 6287
rect 6919 6289 7063 6323
rect 7097 6289 7373 6323
rect 8023 6323 8477 6345
rect 6919 6273 7373 6289
rect 7531 6287 7981 6303
rect 6427 6231 6877 6253
rect 7531 6253 7803 6287
rect 7837 6253 7981 6287
rect 8023 6289 8167 6323
rect 8201 6289 8477 6323
rect 9127 6323 9581 6345
rect 8023 6273 8477 6289
rect 8635 6287 9085 6303
rect 7531 6231 7981 6253
rect 8635 6253 8907 6287
rect 8941 6253 9085 6287
rect 9127 6289 9271 6323
rect 9305 6289 9581 6323
rect 10231 6323 10685 6345
rect 9127 6273 9581 6289
rect 9739 6287 10189 6303
rect 8635 6231 9085 6253
rect 9739 6253 10011 6287
rect 10045 6253 10189 6287
rect 10231 6289 10375 6323
rect 10409 6289 10685 6323
rect 11061 6323 11237 6345
rect 10231 6273 10685 6289
rect 10843 6287 11019 6303
rect 9739 6231 10189 6253
rect 10843 6253 10859 6287
rect 10893 6253 10969 6287
rect 11003 6253 11019 6287
rect 11061 6289 11077 6323
rect 11111 6289 11187 6323
rect 11221 6289 11237 6323
rect 12071 6323 12525 6345
rect 11061 6273 11237 6289
rect 11579 6287 12029 6303
rect 10843 6231 11019 6253
rect 11579 6253 11851 6287
rect 11885 6253 12029 6287
rect 12071 6289 12215 6323
rect 12249 6289 12525 6323
rect 13175 6323 13629 6345
rect 12071 6273 12525 6289
rect 12683 6287 13133 6303
rect 11579 6231 12029 6253
rect 12683 6253 12955 6287
rect 12989 6253 13133 6287
rect 13175 6289 13319 6323
rect 13353 6289 13629 6323
rect 14279 6323 14733 6345
rect 13175 6273 13629 6289
rect 13787 6287 14237 6303
rect 12683 6231 13133 6253
rect 13787 6253 14059 6287
rect 14093 6253 14237 6287
rect 14279 6289 14423 6323
rect 14457 6289 14733 6323
rect 15383 6323 15837 6345
rect 14279 6273 14733 6289
rect 14891 6287 15341 6303
rect 13787 6231 14237 6253
rect 14891 6253 15163 6287
rect 15197 6253 15341 6287
rect 15383 6289 15527 6323
rect 15561 6289 15837 6323
rect 16213 6323 16389 6345
rect 15383 6273 15837 6289
rect 15995 6287 16171 6303
rect 14891 6231 15341 6253
rect 15995 6253 16011 6287
rect 16045 6253 16121 6287
rect 16155 6253 16171 6287
rect 16213 6289 16229 6323
rect 16263 6289 16339 6323
rect 16373 6289 16389 6323
rect 17223 6323 17677 6345
rect 16213 6273 16389 6289
rect 16731 6287 17181 6303
rect 15995 6231 16171 6253
rect 16731 6253 17003 6287
rect 17037 6253 17181 6287
rect 17223 6289 17367 6323
rect 17401 6289 17677 6323
rect 18141 6323 18413 6345
rect 18663 6345 18781 6371
rect 18663 6343 18701 6345
rect 17223 6273 17677 6289
rect 17835 6287 18099 6303
rect 16731 6231 17181 6253
rect 17835 6253 17851 6287
rect 17885 6253 17950 6287
rect 17984 6253 18049 6287
rect 18083 6253 18099 6287
rect 18141 6289 18157 6323
rect 18191 6289 18260 6323
rect 18294 6289 18363 6323
rect 18397 6289 18413 6323
rect 18141 6273 18413 6289
rect 18635 6327 18701 6343
rect 18635 6293 18651 6327
rect 18685 6293 18701 6327
rect 18635 6277 18701 6293
rect 18743 6287 18809 6303
rect 17835 6231 18099 6253
rect 18743 6253 18759 6287
rect 18793 6253 18809 6287
rect 18743 6237 18809 6253
rect 18743 6235 18781 6237
rect 1459 6205 2405 6231
rect 2563 6205 3509 6231
rect 3667 6205 4613 6231
rect 4771 6205 5717 6231
rect 5875 6205 6085 6231
rect 6427 6205 7373 6231
rect 7531 6205 8477 6231
rect 8635 6205 9581 6231
rect 9739 6205 10685 6231
rect 10843 6205 11237 6231
rect 11579 6205 12525 6231
rect 12683 6205 13629 6231
rect 13787 6205 14733 6231
rect 14891 6205 15837 6231
rect 15995 6205 16389 6231
rect 16731 6205 17677 6231
rect 17835 6205 18413 6231
rect 18663 6205 18781 6235
rect 1183 6005 1301 6031
rect 1459 6005 2405 6031
rect 2563 6005 3509 6031
rect 3667 6005 4613 6031
rect 4771 6005 5717 6031
rect 5875 6005 6085 6031
rect 6427 6005 7373 6031
rect 7531 6005 8477 6031
rect 8635 6005 9581 6031
rect 9739 6005 10685 6031
rect 10843 6005 11237 6031
rect 11579 6005 12525 6031
rect 12683 6005 13629 6031
rect 13787 6005 14733 6031
rect 14891 6005 15837 6031
rect 15995 6005 16389 6031
rect 16731 6005 17677 6031
rect 17835 6005 18413 6031
rect 18663 6005 18781 6031
rect 1183 5937 1301 5963
rect 1459 5937 2037 5963
rect 2287 5937 2317 5963
rect 2375 5937 2405 5963
rect 2563 5937 2957 5963
rect 3115 5937 3145 5963
rect 3203 5937 3233 5963
rect 3391 5937 3601 5963
rect 3851 5937 4797 5963
rect 4955 5937 5901 5963
rect 6059 5937 6637 5963
rect 6795 5937 6825 5963
rect 7623 5937 8569 5963
rect 9003 5937 9581 5963
rect 9923 5937 9953 5963
rect 10751 5937 10961 5963
rect 11163 5937 11193 5963
rect 11579 5937 12157 5963
rect 12315 5937 12345 5963
rect 13143 5937 13721 5963
rect 14339 5937 14369 5963
rect 15167 5937 16113 5963
rect 16271 5937 17217 5963
rect 17375 5937 18321 5963
rect 18663 5937 18781 5963
rect 2287 5764 2317 5779
rect 1183 5733 1301 5763
rect 1459 5737 2037 5763
rect 2281 5740 2317 5764
rect 1183 5731 1221 5733
rect 1155 5715 1221 5731
rect 1155 5681 1171 5715
rect 1205 5681 1221 5715
rect 1459 5715 1723 5737
rect 1155 5665 1221 5681
rect 1263 5675 1329 5691
rect 1263 5641 1279 5675
rect 1313 5641 1329 5675
rect 1459 5681 1475 5715
rect 1509 5681 1574 5715
rect 1608 5681 1673 5715
rect 1707 5681 1723 5715
rect 2281 5705 2311 5740
rect 2375 5718 2405 5779
rect 2563 5737 2957 5763
rect 1459 5665 1723 5681
rect 1765 5679 2037 5695
rect 1263 5625 1329 5641
rect 1765 5645 1781 5679
rect 1815 5645 1884 5679
rect 1918 5645 1987 5679
rect 2021 5645 2037 5679
rect 1263 5623 1301 5625
rect 1765 5623 2037 5645
rect 2235 5689 2311 5705
rect 2235 5655 2245 5689
rect 2279 5655 2311 5689
rect 2235 5639 2311 5655
rect 2355 5702 2409 5718
rect 2355 5668 2365 5702
rect 2399 5668 2409 5702
rect 2355 5652 2409 5668
rect 2563 5715 2739 5737
rect 3115 5718 3145 5779
rect 3203 5764 3233 5779
rect 3203 5740 3239 5764
rect 2563 5681 2579 5715
rect 2613 5681 2689 5715
rect 2723 5681 2739 5715
rect 3111 5702 3165 5718
rect 2563 5665 2739 5681
rect 2781 5679 2957 5695
rect 1183 5597 1301 5623
rect 1459 5597 2037 5623
rect 2281 5630 2311 5639
rect 2281 5606 2317 5630
rect 2287 5591 2317 5606
rect 2375 5591 2405 5652
rect 2781 5645 2797 5679
rect 2831 5645 2907 5679
rect 2941 5645 2957 5679
rect 3111 5668 3121 5702
rect 3155 5668 3165 5702
rect 3111 5652 3165 5668
rect 3209 5705 3239 5740
rect 3391 5737 3601 5763
rect 3851 5737 4797 5763
rect 4955 5737 5901 5763
rect 6059 5737 6637 5763
rect 6904 5898 6934 5924
rect 7007 5898 7037 5924
rect 7221 5898 7251 5924
rect 7293 5898 7323 5924
rect 7389 5898 7419 5924
rect 3391 5731 3475 5737
rect 3333 5715 3475 5731
rect 3209 5689 3285 5705
rect 3209 5655 3241 5689
rect 3275 5655 3285 5689
rect 3333 5681 3349 5715
rect 3383 5681 3475 5715
rect 3851 5715 4301 5737
rect 3333 5665 3475 5681
rect 3517 5679 3659 5695
rect 2781 5623 2957 5645
rect 2563 5597 2957 5623
rect 3115 5591 3145 5652
rect 3209 5639 3285 5655
rect 3517 5645 3609 5679
rect 3643 5645 3659 5679
rect 3851 5681 4123 5715
rect 4157 5681 4301 5715
rect 4955 5715 5405 5737
rect 3851 5665 4301 5681
rect 4343 5679 4797 5695
rect 3209 5630 3239 5639
rect 3203 5606 3239 5630
rect 3517 5629 3659 5645
rect 4343 5645 4487 5679
rect 4521 5645 4797 5679
rect 4955 5681 5227 5715
rect 5261 5681 5405 5715
rect 6059 5715 6323 5737
rect 4955 5665 5405 5681
rect 5447 5679 5901 5695
rect 3517 5623 3601 5629
rect 4343 5623 4797 5645
rect 5447 5645 5591 5679
rect 5625 5645 5901 5679
rect 6059 5681 6075 5715
rect 6109 5681 6174 5715
rect 6208 5681 6273 5715
rect 6307 5681 6323 5715
rect 6795 5705 6825 5737
rect 6904 5705 6934 5814
rect 7007 5799 7037 5814
rect 7007 5769 7155 5799
rect 7221 5782 7251 5814
rect 6059 5665 6323 5681
rect 6365 5679 6637 5695
rect 5447 5623 5901 5645
rect 6365 5645 6381 5679
rect 6415 5645 6484 5679
rect 6518 5645 6587 5679
rect 6621 5645 6637 5679
rect 6365 5623 6637 5645
rect 6792 5689 6846 5705
rect 6792 5655 6802 5689
rect 6836 5655 6846 5689
rect 6792 5639 6846 5655
rect 6888 5689 6942 5705
rect 6888 5655 6898 5689
rect 6932 5655 6942 5689
rect 7125 5669 7155 5769
rect 7197 5766 7251 5782
rect 7197 5732 7207 5766
rect 7241 5732 7251 5766
rect 7197 5716 7251 5732
rect 6888 5639 6942 5655
rect 7000 5653 7083 5669
rect 3203 5591 3233 5606
rect 3391 5597 3601 5623
rect 3851 5597 4797 5623
rect 4955 5597 5901 5623
rect 6059 5597 6637 5623
rect 6795 5617 6825 5639
rect 6904 5571 6934 5639
rect 7000 5619 7039 5653
rect 7073 5619 7083 5653
rect 7000 5603 7083 5619
rect 7125 5653 7179 5669
rect 7293 5663 7323 5814
rect 7389 5782 7419 5814
rect 7365 5766 7419 5782
rect 7365 5732 7375 5766
rect 7409 5732 7419 5766
rect 7365 5716 7419 5732
rect 7125 5619 7135 5653
rect 7169 5619 7179 5653
rect 7281 5653 7347 5663
rect 7281 5639 7297 5653
rect 7125 5603 7179 5619
rect 7221 5619 7297 5639
rect 7331 5619 7347 5653
rect 7221 5609 7347 5619
rect 7000 5571 7030 5603
rect 7125 5571 7155 5603
rect 7221 5571 7251 5609
rect 7389 5571 7419 5716
rect 7623 5737 8569 5763
rect 9003 5737 9581 5763
rect 10032 5898 10062 5924
rect 10135 5898 10165 5924
rect 10349 5898 10379 5924
rect 10421 5898 10451 5924
rect 10517 5898 10547 5924
rect 7623 5715 8073 5737
rect 7623 5681 7895 5715
rect 7929 5681 8073 5715
rect 9003 5715 9267 5737
rect 7623 5665 8073 5681
rect 8115 5679 8569 5695
rect 8115 5645 8259 5679
rect 8293 5645 8569 5679
rect 9003 5681 9019 5715
rect 9053 5681 9118 5715
rect 9152 5681 9217 5715
rect 9251 5681 9267 5715
rect 9923 5705 9953 5737
rect 10032 5705 10062 5814
rect 10135 5799 10165 5814
rect 10135 5769 10283 5799
rect 10349 5782 10379 5814
rect 9003 5665 9267 5681
rect 9309 5679 9581 5695
rect 8115 5623 8569 5645
rect 9309 5645 9325 5679
rect 9359 5645 9428 5679
rect 9462 5645 9531 5679
rect 9565 5645 9581 5679
rect 9309 5623 9581 5645
rect 9920 5689 9974 5705
rect 9920 5655 9930 5689
rect 9964 5655 9974 5689
rect 9920 5639 9974 5655
rect 10016 5689 10070 5705
rect 10016 5655 10026 5689
rect 10060 5655 10070 5689
rect 10253 5669 10283 5769
rect 10325 5766 10379 5782
rect 10325 5732 10335 5766
rect 10369 5732 10379 5766
rect 10325 5716 10379 5732
rect 10016 5639 10070 5655
rect 10128 5653 10211 5669
rect 7623 5597 8569 5623
rect 9003 5597 9581 5623
rect 9923 5617 9953 5639
rect 10032 5571 10062 5639
rect 10128 5619 10167 5653
rect 10201 5619 10211 5653
rect 10128 5603 10211 5619
rect 10253 5653 10307 5669
rect 10421 5663 10451 5814
rect 10517 5782 10547 5814
rect 10493 5766 10547 5782
rect 10493 5732 10503 5766
rect 10537 5732 10547 5766
rect 10493 5716 10547 5732
rect 10751 5737 10961 5763
rect 11271 5895 11301 5921
rect 11355 5895 11385 5921
rect 10751 5731 10835 5737
rect 10253 5619 10263 5653
rect 10297 5619 10307 5653
rect 10409 5653 10475 5663
rect 10409 5639 10425 5653
rect 10253 5603 10307 5619
rect 10349 5619 10425 5639
rect 10459 5619 10475 5653
rect 10349 5609 10475 5619
rect 10128 5571 10158 5603
rect 10253 5571 10283 5603
rect 10349 5571 10379 5609
rect 10517 5571 10547 5716
rect 10693 5715 10835 5731
rect 10693 5681 10709 5715
rect 10743 5681 10835 5715
rect 11163 5705 11193 5737
rect 11271 5705 11301 5811
rect 10693 5665 10835 5681
rect 10877 5679 11019 5695
rect 10877 5645 10969 5679
rect 11003 5645 11019 5679
rect 10877 5629 11019 5645
rect 11127 5689 11193 5705
rect 11127 5655 11143 5689
rect 11177 5655 11193 5689
rect 11127 5639 11193 5655
rect 11235 5689 11301 5705
rect 11235 5655 11251 5689
rect 11285 5655 11301 5689
rect 11235 5639 11301 5655
rect 10877 5623 10961 5629
rect 10751 5597 10961 5623
rect 11163 5617 11193 5639
rect 11271 5599 11301 5639
rect 11355 5705 11385 5811
rect 11579 5737 12157 5763
rect 12424 5898 12454 5924
rect 12527 5898 12557 5924
rect 12741 5898 12771 5924
rect 12813 5898 12843 5924
rect 12909 5898 12939 5924
rect 11579 5715 11843 5737
rect 11355 5689 11442 5705
rect 11355 5655 11392 5689
rect 11426 5655 11442 5689
rect 11579 5681 11595 5715
rect 11629 5681 11694 5715
rect 11728 5681 11793 5715
rect 11827 5681 11843 5715
rect 12315 5705 12345 5737
rect 12424 5705 12454 5814
rect 12527 5799 12557 5814
rect 12527 5769 12675 5799
rect 12741 5782 12771 5814
rect 11579 5665 11843 5681
rect 11885 5679 12157 5695
rect 11355 5639 11442 5655
rect 11885 5645 11901 5679
rect 11935 5645 12004 5679
rect 12038 5645 12107 5679
rect 12141 5645 12157 5679
rect 11355 5599 11385 5639
rect 11885 5623 12157 5645
rect 12312 5689 12366 5705
rect 12312 5655 12322 5689
rect 12356 5655 12366 5689
rect 12312 5639 12366 5655
rect 12408 5689 12462 5705
rect 12408 5655 12418 5689
rect 12452 5655 12462 5689
rect 12645 5669 12675 5769
rect 12717 5766 12771 5782
rect 12717 5732 12727 5766
rect 12761 5732 12771 5766
rect 12717 5716 12771 5732
rect 12408 5639 12462 5655
rect 12520 5653 12603 5669
rect 11579 5597 12157 5623
rect 12315 5617 12345 5639
rect 11271 5489 11301 5515
rect 11355 5489 11385 5515
rect 12424 5571 12454 5639
rect 12520 5619 12559 5653
rect 12593 5619 12603 5653
rect 12520 5603 12603 5619
rect 12645 5653 12699 5669
rect 12813 5663 12843 5814
rect 12909 5782 12939 5814
rect 12885 5766 12939 5782
rect 12885 5732 12895 5766
rect 12929 5732 12939 5766
rect 12885 5716 12939 5732
rect 12645 5619 12655 5653
rect 12689 5619 12699 5653
rect 12801 5653 12867 5663
rect 12801 5639 12817 5653
rect 12645 5603 12699 5619
rect 12741 5619 12817 5639
rect 12851 5619 12867 5653
rect 12741 5609 12867 5619
rect 12520 5571 12550 5603
rect 12645 5571 12675 5603
rect 12741 5571 12771 5609
rect 12909 5571 12939 5716
rect 13143 5737 13721 5763
rect 14448 5898 14478 5924
rect 14551 5898 14581 5924
rect 14765 5898 14795 5924
rect 14837 5898 14867 5924
rect 14933 5898 14963 5924
rect 13143 5715 13407 5737
rect 13143 5681 13159 5715
rect 13193 5681 13258 5715
rect 13292 5681 13357 5715
rect 13391 5681 13407 5715
rect 14339 5705 14369 5737
rect 14448 5705 14478 5814
rect 14551 5799 14581 5814
rect 14551 5769 14699 5799
rect 14765 5782 14795 5814
rect 13143 5665 13407 5681
rect 13449 5679 13721 5695
rect 13449 5645 13465 5679
rect 13499 5645 13568 5679
rect 13602 5645 13671 5679
rect 13705 5645 13721 5679
rect 13449 5623 13721 5645
rect 14336 5689 14390 5705
rect 14336 5655 14346 5689
rect 14380 5655 14390 5689
rect 14336 5639 14390 5655
rect 14432 5689 14486 5705
rect 14432 5655 14442 5689
rect 14476 5655 14486 5689
rect 14669 5669 14699 5769
rect 14741 5766 14795 5782
rect 14741 5732 14751 5766
rect 14785 5732 14795 5766
rect 14741 5716 14795 5732
rect 14432 5639 14486 5655
rect 14544 5653 14627 5669
rect 13143 5597 13721 5623
rect 14339 5617 14369 5639
rect 14448 5571 14478 5639
rect 14544 5619 14583 5653
rect 14617 5619 14627 5653
rect 14544 5603 14627 5619
rect 14669 5653 14723 5669
rect 14837 5663 14867 5814
rect 14933 5782 14963 5814
rect 14909 5766 14963 5782
rect 14909 5732 14919 5766
rect 14953 5732 14963 5766
rect 14909 5716 14963 5732
rect 14669 5619 14679 5653
rect 14713 5619 14723 5653
rect 14825 5653 14891 5663
rect 14825 5639 14841 5653
rect 14669 5603 14723 5619
rect 14765 5619 14841 5639
rect 14875 5619 14891 5653
rect 14765 5609 14891 5619
rect 14544 5571 14574 5603
rect 14669 5571 14699 5603
rect 14765 5571 14795 5609
rect 14933 5571 14963 5716
rect 15167 5737 16113 5763
rect 16271 5737 17217 5763
rect 17375 5737 18321 5763
rect 15167 5715 15617 5737
rect 15167 5681 15439 5715
rect 15473 5681 15617 5715
rect 16271 5715 16721 5737
rect 15167 5665 15617 5681
rect 15659 5679 16113 5695
rect 15659 5645 15803 5679
rect 15837 5645 16113 5679
rect 16271 5681 16543 5715
rect 16577 5681 16721 5715
rect 17375 5715 17825 5737
rect 18663 5733 18781 5763
rect 16271 5665 16721 5681
rect 16763 5679 17217 5695
rect 15659 5623 16113 5645
rect 16763 5645 16907 5679
rect 16941 5645 17217 5679
rect 17375 5681 17647 5715
rect 17681 5681 17825 5715
rect 18743 5731 18781 5733
rect 18743 5715 18809 5731
rect 17375 5665 17825 5681
rect 17867 5679 18321 5695
rect 16763 5623 17217 5645
rect 17867 5645 18011 5679
rect 18045 5645 18321 5679
rect 17867 5623 18321 5645
rect 18635 5675 18701 5691
rect 18635 5641 18651 5675
rect 18685 5641 18701 5675
rect 18743 5681 18759 5715
rect 18793 5681 18809 5715
rect 18743 5665 18809 5681
rect 18635 5625 18701 5641
rect 15167 5597 16113 5623
rect 16271 5597 17217 5623
rect 17375 5597 18321 5623
rect 18663 5623 18701 5625
rect 18663 5597 18781 5623
rect 1183 5461 1301 5487
rect 1459 5461 2037 5487
rect 2287 5461 2317 5487
rect 2375 5461 2405 5487
rect 2563 5461 2957 5487
rect 3115 5461 3145 5487
rect 3203 5461 3233 5487
rect 3391 5461 3601 5487
rect 3851 5461 4797 5487
rect 4955 5461 5901 5487
rect 6059 5461 6637 5487
rect 6795 5461 6825 5487
rect 6904 5461 6934 5487
rect 7000 5461 7030 5487
rect 7125 5461 7155 5487
rect 7221 5461 7251 5487
rect 7389 5461 7419 5487
rect 7623 5461 8569 5487
rect 9003 5461 9581 5487
rect 9923 5461 9953 5487
rect 10032 5461 10062 5487
rect 10128 5461 10158 5487
rect 10253 5461 10283 5487
rect 10349 5461 10379 5487
rect 10517 5461 10547 5487
rect 10751 5461 10961 5487
rect 11163 5461 11193 5487
rect 11579 5461 12157 5487
rect 12315 5461 12345 5487
rect 12424 5461 12454 5487
rect 12520 5461 12550 5487
rect 12645 5461 12675 5487
rect 12741 5461 12771 5487
rect 12909 5461 12939 5487
rect 13143 5461 13721 5487
rect 14339 5461 14369 5487
rect 14448 5461 14478 5487
rect 14544 5461 14574 5487
rect 14669 5461 14699 5487
rect 14765 5461 14795 5487
rect 14933 5461 14963 5487
rect 15167 5461 16113 5487
rect 16271 5461 17217 5487
rect 17375 5461 18321 5487
rect 18663 5461 18781 5487
rect 1183 5393 1301 5419
rect 1459 5393 1853 5419
rect 2055 5393 2085 5419
rect 2471 5393 2681 5419
rect 2975 5393 3005 5419
rect 3391 5393 3601 5419
rect 3759 5393 3789 5419
rect 3854 5393 3884 5419
rect 3938 5393 3968 5419
rect 4127 5393 4337 5419
rect 4497 5393 4527 5419
rect 4581 5393 4611 5419
rect 4771 5393 5717 5419
rect 5875 5393 5905 5419
rect 5963 5393 5993 5419
rect 6427 5393 6545 5419
rect 6703 5393 6733 5419
rect 6812 5393 6842 5419
rect 6908 5393 6938 5419
rect 7033 5393 7063 5419
rect 7129 5393 7159 5419
rect 7297 5393 7327 5419
rect 7531 5393 7741 5419
rect 7899 5393 7929 5419
rect 8008 5393 8038 5419
rect 8104 5393 8134 5419
rect 8229 5393 8259 5419
rect 8325 5393 8355 5419
rect 8493 5393 8523 5419
rect 8727 5393 8937 5419
rect 9187 5393 9217 5419
rect 9375 5393 9405 5419
rect 9467 5393 9497 5419
rect 9551 5393 9581 5419
rect 9739 5393 10317 5419
rect 10475 5393 10505 5419
rect 10584 5393 10614 5419
rect 10680 5393 10710 5419
rect 10805 5393 10835 5419
rect 10901 5393 10931 5419
rect 11069 5393 11099 5419
rect 11579 5393 12525 5419
rect 12683 5393 12893 5419
rect 13143 5393 13173 5419
rect 13252 5393 13282 5419
rect 13348 5393 13378 5419
rect 13473 5393 13503 5419
rect 13569 5393 13599 5419
rect 13737 5393 13767 5419
rect 13971 5393 14917 5419
rect 15075 5393 16021 5419
rect 16179 5393 16389 5419
rect 16731 5393 17677 5419
rect 17835 5393 18413 5419
rect 18663 5393 18781 5419
rect 1183 5257 1301 5283
rect 1459 5257 1853 5283
rect 2163 5365 2193 5391
rect 2247 5365 2277 5391
rect 1263 5255 1301 5257
rect 1263 5239 1329 5255
rect 1155 5199 1221 5215
rect 1155 5165 1171 5199
rect 1205 5165 1221 5199
rect 1263 5205 1279 5239
rect 1313 5205 1329 5239
rect 1677 5235 1853 5257
rect 2055 5241 2085 5263
rect 2163 5241 2193 5281
rect 1263 5189 1329 5205
rect 1459 5199 1635 5215
rect 1155 5149 1221 5165
rect 1183 5147 1221 5149
rect 1459 5165 1475 5199
rect 1509 5165 1585 5199
rect 1619 5165 1635 5199
rect 1677 5201 1693 5235
rect 1727 5201 1803 5235
rect 1837 5201 1853 5235
rect 1677 5185 1853 5201
rect 2019 5225 2085 5241
rect 2019 5191 2035 5225
rect 2069 5191 2085 5225
rect 2019 5175 2085 5191
rect 2127 5225 2193 5241
rect 2127 5191 2143 5225
rect 2177 5191 2193 5225
rect 2127 5175 2193 5191
rect 1183 5117 1301 5147
rect 1459 5143 1635 5165
rect 2055 5143 2085 5175
rect 1459 5117 1853 5143
rect 2163 5069 2193 5175
rect 2247 5241 2277 5281
rect 2471 5257 2681 5283
rect 3083 5365 3113 5391
rect 3167 5365 3197 5391
rect 2597 5251 2681 5257
rect 2247 5225 2334 5241
rect 2247 5191 2284 5225
rect 2318 5191 2334 5225
rect 2597 5235 2739 5251
rect 2975 5241 3005 5263
rect 3083 5241 3113 5281
rect 2247 5175 2334 5191
rect 2413 5199 2555 5215
rect 2247 5069 2277 5175
rect 2413 5165 2429 5199
rect 2463 5165 2555 5199
rect 2597 5201 2689 5235
rect 2723 5201 2739 5235
rect 2597 5185 2739 5201
rect 2939 5225 3005 5241
rect 2939 5191 2955 5225
rect 2989 5191 3005 5225
rect 2939 5175 3005 5191
rect 3047 5225 3113 5241
rect 3047 5191 3063 5225
rect 3097 5191 3113 5225
rect 3047 5175 3113 5191
rect 2413 5149 2555 5165
rect 2471 5143 2555 5149
rect 2975 5143 3005 5175
rect 2471 5117 2681 5143
rect 2163 4959 2193 4985
rect 2247 4959 2277 4985
rect 3083 5069 3113 5175
rect 3167 5241 3197 5281
rect 3391 5257 3601 5283
rect 3517 5251 3601 5257
rect 3167 5225 3254 5241
rect 3167 5191 3204 5225
rect 3238 5191 3254 5225
rect 3517 5235 3659 5251
rect 3759 5241 3789 5309
rect 3854 5241 3884 5263
rect 3938 5241 3968 5263
rect 4127 5257 4337 5283
rect 3167 5175 3254 5191
rect 3333 5199 3475 5215
rect 3167 5069 3197 5175
rect 3333 5165 3349 5199
rect 3383 5165 3475 5199
rect 3517 5201 3609 5235
rect 3643 5201 3659 5235
rect 3517 5185 3659 5201
rect 3707 5225 3789 5241
rect 3707 5191 3717 5225
rect 3751 5191 3789 5225
rect 3707 5175 3789 5191
rect 3831 5225 3968 5241
rect 3831 5191 3841 5225
rect 3875 5191 3968 5225
rect 4253 5251 4337 5257
rect 4253 5235 4395 5251
rect 4497 5241 4527 5263
rect 4581 5241 4611 5263
rect 4771 5257 5717 5283
rect 3831 5175 3968 5191
rect 3333 5149 3475 5165
rect 3391 5143 3475 5149
rect 3391 5117 3601 5143
rect 3083 4959 3113 4985
rect 3167 4959 3197 4985
rect 3759 5079 3789 5175
rect 3854 5143 3884 5175
rect 3938 5143 3968 5175
rect 4069 5199 4211 5215
rect 4069 5165 4085 5199
rect 4119 5165 4211 5199
rect 4253 5201 4345 5235
rect 4379 5201 4395 5235
rect 4253 5185 4395 5201
rect 4437 5225 4611 5241
rect 4437 5191 4453 5225
rect 4487 5191 4611 5225
rect 5263 5235 5717 5257
rect 4437 5175 4611 5191
rect 4069 5149 4211 5165
rect 4127 5143 4211 5149
rect 4497 5143 4527 5175
rect 4581 5143 4611 5175
rect 4771 5199 5221 5215
rect 4771 5165 5043 5199
rect 5077 5165 5221 5199
rect 5263 5201 5407 5235
rect 5441 5201 5717 5235
rect 5875 5228 5905 5289
rect 5963 5274 5993 5289
rect 5963 5250 5999 5274
rect 6427 5257 6545 5283
rect 5969 5241 5999 5250
rect 6507 5255 6545 5257
rect 5263 5185 5717 5201
rect 5871 5212 5925 5228
rect 4771 5143 5221 5165
rect 5871 5178 5881 5212
rect 5915 5178 5925 5212
rect 5871 5162 5925 5178
rect 5969 5225 6045 5241
rect 5969 5191 6001 5225
rect 6035 5191 6045 5225
rect 6507 5239 6573 5255
rect 6703 5241 6733 5263
rect 6812 5241 6842 5309
rect 6908 5277 6938 5309
rect 7033 5277 7063 5309
rect 6908 5261 6991 5277
rect 5969 5175 6045 5191
rect 6399 5199 6465 5215
rect 1183 4917 1301 4943
rect 1459 4917 1853 4943
rect 2055 4917 2085 4943
rect 2471 4917 2681 4943
rect 2975 4917 3005 4943
rect 3391 4917 3601 4943
rect 3759 4925 3789 4951
rect 4127 5117 4337 5143
rect 4771 5117 5717 5143
rect 5875 5101 5905 5162
rect 5969 5140 5999 5175
rect 6399 5165 6415 5199
rect 6449 5165 6465 5199
rect 6507 5205 6523 5239
rect 6557 5205 6573 5239
rect 6507 5189 6573 5205
rect 6700 5225 6754 5241
rect 6700 5191 6710 5225
rect 6744 5191 6754 5225
rect 6700 5175 6754 5191
rect 6796 5225 6850 5241
rect 6796 5191 6806 5225
rect 6840 5191 6850 5225
rect 6908 5227 6947 5261
rect 6981 5227 6991 5261
rect 6908 5211 6991 5227
rect 7033 5261 7087 5277
rect 7033 5227 7043 5261
rect 7077 5227 7087 5261
rect 7129 5271 7159 5309
rect 7129 5261 7255 5271
rect 7129 5241 7205 5261
rect 7033 5211 7087 5227
rect 7189 5227 7205 5241
rect 7239 5227 7255 5261
rect 7189 5217 7255 5227
rect 6796 5175 6850 5191
rect 6399 5149 6465 5165
rect 5963 5116 5999 5140
rect 6427 5147 6465 5149
rect 5963 5101 5993 5116
rect 6427 5117 6545 5147
rect 6703 5143 6733 5175
rect 6812 5066 6842 5175
rect 7033 5111 7063 5211
rect 6915 5081 7063 5111
rect 7105 5148 7159 5164
rect 7105 5114 7115 5148
rect 7149 5114 7159 5148
rect 7105 5098 7159 5114
rect 6915 5066 6945 5081
rect 7129 5066 7159 5098
rect 7201 5066 7231 5217
rect 7297 5164 7327 5309
rect 7531 5257 7741 5283
rect 7657 5251 7741 5257
rect 7657 5235 7799 5251
rect 7899 5241 7929 5263
rect 8008 5241 8038 5309
rect 8104 5277 8134 5309
rect 8229 5277 8259 5309
rect 8104 5261 8187 5277
rect 7273 5148 7327 5164
rect 7473 5199 7615 5215
rect 7473 5165 7489 5199
rect 7523 5165 7615 5199
rect 7657 5201 7749 5235
rect 7783 5201 7799 5235
rect 7657 5185 7799 5201
rect 7896 5225 7950 5241
rect 7896 5191 7906 5225
rect 7940 5191 7950 5225
rect 7896 5175 7950 5191
rect 7992 5225 8046 5241
rect 7992 5191 8002 5225
rect 8036 5191 8046 5225
rect 8104 5227 8143 5261
rect 8177 5227 8187 5261
rect 8104 5211 8187 5227
rect 8229 5261 8283 5277
rect 8229 5227 8239 5261
rect 8273 5227 8283 5261
rect 8325 5271 8355 5309
rect 8325 5261 8451 5271
rect 8325 5241 8401 5261
rect 8229 5211 8283 5227
rect 8385 5227 8401 5241
rect 8435 5227 8451 5261
rect 8385 5217 8451 5227
rect 7992 5175 8046 5191
rect 7473 5149 7615 5165
rect 7273 5114 7283 5148
rect 7317 5114 7327 5148
rect 7531 5143 7615 5149
rect 7899 5143 7929 5175
rect 7531 5117 7741 5143
rect 7273 5098 7327 5114
rect 7297 5066 7327 5098
rect 6812 4956 6842 4982
rect 6915 4956 6945 4982
rect 7129 4956 7159 4982
rect 7201 4956 7231 4982
rect 7297 4956 7327 4982
rect 8008 5066 8038 5175
rect 8229 5111 8259 5211
rect 8111 5081 8259 5111
rect 8301 5148 8355 5164
rect 8301 5114 8311 5148
rect 8345 5114 8355 5148
rect 8301 5098 8355 5114
rect 8111 5066 8141 5081
rect 8325 5066 8355 5098
rect 8397 5066 8427 5217
rect 8493 5164 8523 5309
rect 8727 5257 8937 5283
rect 8853 5251 8937 5257
rect 8853 5235 8995 5251
rect 8469 5148 8523 5164
rect 8669 5199 8811 5215
rect 8669 5165 8685 5199
rect 8719 5165 8811 5199
rect 8853 5201 8945 5235
rect 8979 5201 8995 5235
rect 8853 5185 8995 5201
rect 9187 5241 9217 5263
rect 9375 5241 9405 5263
rect 9467 5241 9497 5263
rect 9551 5241 9581 5263
rect 9739 5257 10317 5283
rect 9187 5225 9271 5241
rect 9187 5191 9227 5225
rect 9261 5191 9271 5225
rect 9187 5175 9271 5191
rect 9352 5225 9409 5241
rect 9352 5191 9365 5225
rect 9399 5191 9409 5225
rect 9352 5175 9409 5191
rect 9455 5225 9509 5241
rect 9455 5191 9465 5225
rect 9499 5191 9509 5225
rect 9455 5175 9509 5191
rect 9551 5225 9637 5241
rect 9551 5191 9593 5225
rect 9627 5191 9637 5225
rect 10045 5235 10317 5257
rect 10475 5241 10505 5263
rect 10584 5241 10614 5309
rect 10680 5277 10710 5309
rect 10805 5277 10835 5309
rect 10680 5261 10763 5277
rect 8669 5149 8811 5165
rect 8469 5114 8479 5148
rect 8513 5114 8523 5148
rect 8727 5143 8811 5149
rect 9191 5143 9221 5175
rect 9352 5143 9382 5175
rect 9460 5143 9490 5175
rect 9551 5171 9637 5191
rect 9739 5199 10003 5215
rect 9551 5143 9581 5171
rect 9739 5165 9755 5199
rect 9789 5165 9854 5199
rect 9888 5165 9953 5199
rect 9987 5165 10003 5199
rect 10045 5201 10061 5235
rect 10095 5201 10164 5235
rect 10198 5201 10267 5235
rect 10301 5201 10317 5235
rect 10045 5185 10317 5201
rect 10472 5225 10526 5241
rect 10472 5191 10482 5225
rect 10516 5191 10526 5225
rect 10472 5175 10526 5191
rect 10568 5225 10622 5241
rect 10568 5191 10578 5225
rect 10612 5191 10622 5225
rect 10680 5227 10719 5261
rect 10753 5227 10763 5261
rect 10680 5211 10763 5227
rect 10805 5261 10859 5277
rect 10805 5227 10815 5261
rect 10849 5227 10859 5261
rect 10901 5271 10931 5309
rect 10901 5261 11027 5271
rect 10901 5241 10977 5261
rect 10805 5211 10859 5227
rect 10961 5227 10977 5241
rect 11011 5227 11027 5261
rect 10961 5217 11027 5227
rect 10568 5175 10622 5191
rect 9739 5143 10003 5165
rect 10475 5143 10505 5175
rect 8727 5117 8937 5143
rect 8469 5098 8523 5114
rect 8493 5066 8523 5098
rect 8008 4956 8038 4982
rect 8111 4956 8141 4982
rect 8325 4956 8355 4982
rect 8397 4956 8427 4982
rect 8493 4956 8523 4982
rect 9739 5117 10317 5143
rect 10584 5066 10614 5175
rect 10805 5111 10835 5211
rect 10687 5081 10835 5111
rect 10877 5148 10931 5164
rect 10877 5114 10887 5148
rect 10921 5114 10931 5148
rect 10877 5098 10931 5114
rect 10687 5066 10717 5081
rect 10901 5066 10931 5098
rect 10973 5066 11003 5217
rect 11069 5164 11099 5309
rect 11579 5257 12525 5283
rect 12683 5257 12893 5283
rect 12071 5235 12525 5257
rect 11045 5148 11099 5164
rect 11045 5114 11055 5148
rect 11089 5114 11099 5148
rect 11579 5199 12029 5215
rect 11579 5165 11851 5199
rect 11885 5165 12029 5199
rect 12071 5201 12215 5235
rect 12249 5201 12525 5235
rect 12809 5251 12893 5257
rect 12809 5235 12951 5251
rect 13143 5241 13173 5263
rect 13252 5241 13282 5309
rect 13348 5277 13378 5309
rect 13473 5277 13503 5309
rect 13348 5261 13431 5277
rect 12071 5185 12525 5201
rect 12625 5199 12767 5215
rect 11579 5143 12029 5165
rect 12625 5165 12641 5199
rect 12675 5165 12767 5199
rect 12809 5201 12901 5235
rect 12935 5201 12951 5235
rect 12809 5185 12951 5201
rect 13140 5225 13194 5241
rect 13140 5191 13150 5225
rect 13184 5191 13194 5225
rect 13140 5175 13194 5191
rect 13236 5225 13290 5241
rect 13236 5191 13246 5225
rect 13280 5191 13290 5225
rect 13348 5227 13387 5261
rect 13421 5227 13431 5261
rect 13348 5211 13431 5227
rect 13473 5261 13527 5277
rect 13473 5227 13483 5261
rect 13517 5227 13527 5261
rect 13569 5271 13599 5309
rect 13569 5261 13695 5271
rect 13569 5241 13645 5261
rect 13473 5211 13527 5227
rect 13629 5227 13645 5241
rect 13679 5227 13695 5261
rect 13629 5217 13695 5227
rect 13236 5175 13290 5191
rect 12625 5149 12767 5165
rect 12683 5143 12767 5149
rect 13143 5143 13173 5175
rect 11045 5098 11099 5114
rect 11069 5066 11099 5098
rect 11579 5117 12525 5143
rect 12683 5117 12893 5143
rect 10584 4956 10614 4982
rect 10687 4956 10717 4982
rect 10901 4956 10931 4982
rect 10973 4956 11003 4982
rect 11069 4956 11099 4982
rect 13252 5066 13282 5175
rect 13473 5111 13503 5211
rect 13355 5081 13503 5111
rect 13545 5148 13599 5164
rect 13545 5114 13555 5148
rect 13589 5114 13599 5148
rect 13545 5098 13599 5114
rect 13355 5066 13385 5081
rect 13569 5066 13599 5098
rect 13641 5066 13671 5217
rect 13737 5164 13767 5309
rect 13971 5257 14917 5283
rect 15075 5257 16021 5283
rect 16179 5257 16389 5283
rect 16731 5257 17677 5283
rect 17835 5257 18413 5283
rect 14463 5235 14917 5257
rect 13713 5148 13767 5164
rect 13713 5114 13723 5148
rect 13757 5114 13767 5148
rect 13971 5199 14421 5215
rect 13971 5165 14243 5199
rect 14277 5165 14421 5199
rect 14463 5201 14607 5235
rect 14641 5201 14917 5235
rect 15567 5235 16021 5257
rect 14463 5185 14917 5201
rect 15075 5199 15525 5215
rect 13971 5143 14421 5165
rect 15075 5165 15347 5199
rect 15381 5165 15525 5199
rect 15567 5201 15711 5235
rect 15745 5201 16021 5235
rect 16305 5251 16389 5257
rect 16305 5235 16447 5251
rect 15567 5185 16021 5201
rect 16121 5199 16263 5215
rect 15075 5143 15525 5165
rect 16121 5165 16137 5199
rect 16171 5165 16263 5199
rect 16305 5201 16397 5235
rect 16431 5201 16447 5235
rect 17223 5235 17677 5257
rect 16305 5185 16447 5201
rect 16731 5199 17181 5215
rect 16121 5149 16263 5165
rect 16179 5143 16263 5149
rect 16731 5165 17003 5199
rect 17037 5165 17181 5199
rect 17223 5201 17367 5235
rect 17401 5201 17677 5235
rect 18141 5235 18413 5257
rect 18663 5257 18781 5283
rect 18663 5255 18701 5257
rect 17223 5185 17677 5201
rect 17835 5199 18099 5215
rect 16731 5143 17181 5165
rect 17835 5165 17851 5199
rect 17885 5165 17950 5199
rect 17984 5165 18049 5199
rect 18083 5165 18099 5199
rect 18141 5201 18157 5235
rect 18191 5201 18260 5235
rect 18294 5201 18363 5235
rect 18397 5201 18413 5235
rect 18141 5185 18413 5201
rect 18635 5239 18701 5255
rect 18635 5205 18651 5239
rect 18685 5205 18701 5239
rect 18635 5189 18701 5205
rect 18743 5199 18809 5215
rect 17835 5143 18099 5165
rect 18743 5165 18759 5199
rect 18793 5165 18809 5199
rect 18743 5149 18809 5165
rect 18743 5147 18781 5149
rect 13971 5117 14917 5143
rect 15075 5117 16021 5143
rect 16179 5117 16389 5143
rect 13713 5098 13767 5114
rect 13737 5066 13767 5098
rect 13252 4956 13282 4982
rect 13355 4956 13385 4982
rect 13569 4956 13599 4982
rect 13641 4956 13671 4982
rect 13737 4956 13767 4982
rect 16731 5117 17677 5143
rect 17835 5117 18413 5143
rect 18663 5117 18781 5147
rect 3854 4917 3884 4943
rect 3938 4917 3968 4943
rect 4127 4917 4337 4943
rect 4497 4917 4527 4943
rect 4581 4917 4611 4943
rect 4771 4917 5717 4943
rect 5875 4917 5905 4943
rect 5963 4917 5993 4943
rect 6427 4917 6545 4943
rect 6703 4917 6733 4943
rect 7531 4917 7741 4943
rect 7899 4917 7929 4943
rect 8727 4917 8937 4943
rect 9191 4917 9221 4943
rect 9352 4917 9382 4943
rect 9460 4917 9490 4943
rect 9551 4917 9581 4943
rect 9739 4917 10317 4943
rect 10475 4917 10505 4943
rect 11579 4917 12525 4943
rect 12683 4917 12893 4943
rect 13143 4917 13173 4943
rect 13971 4917 14917 4943
rect 15075 4917 16021 4943
rect 16179 4917 16389 4943
rect 16731 4917 17677 4943
rect 17835 4917 18413 4943
rect 18663 4917 18781 4943
rect 1183 4849 1301 4875
rect 1459 4849 1853 4875
rect 2103 4843 2133 4869
rect 2187 4843 2217 4869
rect 2375 4849 2405 4875
rect 2460 4849 2490 4875
rect 2555 4849 2585 4875
rect 2658 4849 2688 4875
rect 2790 4849 2820 4875
rect 2885 4849 2915 4875
rect 2969 4849 2999 4875
rect 3083 4849 3113 4875
rect 3293 4849 3323 4875
rect 3377 4849 3407 4875
rect 4079 4849 4109 4875
rect 4495 4849 4705 4875
rect 4959 4849 4989 4875
rect 5120 4849 5150 4875
rect 5228 4849 5258 4875
rect 5319 4849 5349 4875
rect 5507 4849 5717 4875
rect 5879 4849 5909 4875
rect 6040 4849 6070 4875
rect 6148 4849 6178 4875
rect 6239 4849 6269 4875
rect 6427 4849 6637 4875
rect 2103 4700 2133 4715
rect 1183 4645 1301 4675
rect 1459 4649 1853 4675
rect 2070 4670 2133 4700
rect 1183 4643 1221 4645
rect 1155 4627 1221 4643
rect 1155 4593 1171 4627
rect 1205 4593 1221 4627
rect 1459 4627 1635 4649
rect 1155 4577 1221 4593
rect 1263 4587 1329 4603
rect 1263 4553 1279 4587
rect 1313 4553 1329 4587
rect 1459 4593 1475 4627
rect 1509 4593 1585 4627
rect 1619 4593 1635 4627
rect 2070 4617 2100 4670
rect 2187 4626 2217 4715
rect 2375 4685 2405 4765
rect 1459 4577 1635 4593
rect 1677 4591 1853 4607
rect 1263 4537 1329 4553
rect 1677 4557 1693 4591
rect 1727 4557 1803 4591
rect 1837 4557 1853 4591
rect 1263 4535 1301 4537
rect 1677 4535 1853 4557
rect 2046 4601 2100 4617
rect 2046 4567 2056 4601
rect 2090 4567 2100 4601
rect 2142 4616 2217 4626
rect 2310 4669 2405 4685
rect 2310 4635 2320 4669
rect 2354 4635 2405 4669
rect 2460 4649 2490 4765
rect 2555 4733 2585 4765
rect 2555 4717 2616 4733
rect 2555 4683 2572 4717
rect 2606 4683 2616 4717
rect 2555 4667 2616 4683
rect 2310 4619 2405 4635
rect 2142 4582 2158 4616
rect 2192 4582 2217 4616
rect 2142 4572 2217 4582
rect 2046 4551 2100 4567
rect 1183 4509 1301 4535
rect 1459 4509 1853 4535
rect 2070 4528 2100 4551
rect 2070 4498 2133 4528
rect 2103 4483 2133 4498
rect 2187 4483 2217 4572
rect 2375 4483 2405 4619
rect 2447 4639 2513 4649
rect 2447 4605 2463 4639
rect 2497 4625 2513 4639
rect 2497 4605 2616 4625
rect 2447 4595 2616 4605
rect 2467 4543 2533 4553
rect 2467 4509 2483 4543
rect 2517 4509 2533 4543
rect 2467 4499 2533 4509
rect 2487 4471 2517 4499
rect 2586 4471 2616 4595
rect 2658 4565 2688 4765
rect 2790 4661 2820 4699
rect 2885 4667 2915 4765
rect 2969 4727 2999 4765
rect 3083 4733 3113 4765
rect 2968 4717 3034 4727
rect 2968 4683 2984 4717
rect 3018 4683 3034 4717
rect 2968 4673 3034 4683
rect 3083 4717 3164 4733
rect 3083 4683 3120 4717
rect 3154 4683 3164 4717
rect 3083 4667 3164 4683
rect 2730 4651 2820 4661
rect 2730 4617 2746 4651
rect 2780 4617 2820 4651
rect 2730 4607 2820 4617
rect 2790 4572 2820 4607
rect 2872 4651 2926 4667
rect 2872 4617 2882 4651
rect 2916 4631 2926 4651
rect 2916 4617 3041 4631
rect 2872 4601 3041 4617
rect 2658 4555 2732 4565
rect 2658 4521 2682 4555
rect 2716 4521 2732 4555
rect 2790 4542 2834 4572
rect 2804 4527 2834 4542
rect 2905 4543 2969 4559
rect 2658 4511 2732 4521
rect 2685 4483 2715 4511
rect 2905 4509 2925 4543
rect 2959 4509 2969 4543
rect 2905 4493 2969 4509
rect 2905 4471 2935 4493
rect 3011 4471 3041 4601
rect 3106 4483 3136 4667
rect 4187 4807 4217 4833
rect 4271 4807 4301 4833
rect 3293 4617 3323 4649
rect 3377 4617 3407 4649
rect 4079 4617 4109 4649
rect 4187 4617 4217 4723
rect 3183 4601 3325 4617
rect 3183 4567 3193 4601
rect 3227 4567 3325 4601
rect 3183 4551 3325 4567
rect 3367 4601 3421 4617
rect 3367 4567 3377 4601
rect 3411 4567 3421 4601
rect 3367 4551 3421 4567
rect 4043 4601 4109 4617
rect 4043 4567 4059 4601
rect 4093 4567 4109 4601
rect 4043 4551 4109 4567
rect 4151 4601 4217 4617
rect 4151 4567 4167 4601
rect 4201 4567 4217 4601
rect 4151 4551 4217 4567
rect 3295 4529 3325 4551
rect 3379 4529 3409 4551
rect 4079 4529 4109 4551
rect 4187 4511 4217 4551
rect 4271 4617 4301 4723
rect 4495 4649 4705 4675
rect 5507 4649 5717 4675
rect 6795 4843 6825 4869
rect 6879 4843 6909 4869
rect 7067 4849 7097 4875
rect 7152 4849 7182 4875
rect 7247 4849 7277 4875
rect 7350 4849 7380 4875
rect 7482 4849 7512 4875
rect 7577 4849 7607 4875
rect 7661 4849 7691 4875
rect 7775 4849 7805 4875
rect 7985 4849 8015 4875
rect 8069 4849 8099 4875
rect 8267 4849 8661 4875
rect 9003 4849 9581 4875
rect 9739 4849 9857 4875
rect 10025 4849 10055 4875
rect 10109 4849 10139 4875
rect 10319 4849 10349 4875
rect 10433 4849 10463 4875
rect 10517 4849 10547 4875
rect 10612 4849 10642 4875
rect 10744 4849 10774 4875
rect 10847 4849 10877 4875
rect 10942 4849 10972 4875
rect 11027 4849 11057 4875
rect 6795 4700 6825 4715
rect 6427 4649 6637 4675
rect 6762 4670 6825 4700
rect 4495 4643 4579 4649
rect 4437 4627 4579 4643
rect 4271 4601 4358 4617
rect 4271 4567 4308 4601
rect 4342 4567 4358 4601
rect 4437 4593 4453 4627
rect 4487 4593 4579 4627
rect 4959 4617 4989 4649
rect 5120 4617 5150 4649
rect 5228 4617 5258 4649
rect 5319 4621 5349 4649
rect 5507 4643 5591 4649
rect 5449 4627 5591 4643
rect 4437 4577 4579 4593
rect 4621 4591 4763 4607
rect 4271 4551 4358 4567
rect 4621 4557 4713 4591
rect 4747 4557 4763 4591
rect 4271 4511 4301 4551
rect 4621 4541 4763 4557
rect 4955 4601 5039 4617
rect 4955 4567 4995 4601
rect 5029 4567 5039 4601
rect 4955 4551 5039 4567
rect 5120 4601 5177 4617
rect 5120 4567 5133 4601
rect 5167 4567 5177 4601
rect 5120 4551 5177 4567
rect 5223 4601 5277 4617
rect 5223 4567 5233 4601
rect 5267 4567 5277 4601
rect 5223 4551 5277 4567
rect 5319 4601 5405 4621
rect 5319 4567 5361 4601
rect 5395 4567 5405 4601
rect 5449 4593 5465 4627
rect 5499 4593 5591 4627
rect 5879 4617 5909 4649
rect 6040 4617 6070 4649
rect 6148 4617 6178 4649
rect 6239 4621 6269 4649
rect 6427 4643 6511 4649
rect 6369 4627 6511 4643
rect 5449 4577 5591 4593
rect 5633 4591 5775 4607
rect 5319 4551 5405 4567
rect 5633 4557 5725 4591
rect 5759 4557 5775 4591
rect 4621 4535 4705 4541
rect 4495 4509 4705 4535
rect 4955 4529 4985 4551
rect 5143 4529 5173 4551
rect 5235 4529 5265 4551
rect 5319 4529 5349 4551
rect 5633 4541 5775 4557
rect 5875 4601 5959 4617
rect 5875 4567 5915 4601
rect 5949 4567 5959 4601
rect 5875 4551 5959 4567
rect 6040 4601 6097 4617
rect 6040 4567 6053 4601
rect 6087 4567 6097 4601
rect 6040 4551 6097 4567
rect 6143 4601 6197 4617
rect 6143 4567 6153 4601
rect 6187 4567 6197 4601
rect 6143 4551 6197 4567
rect 6239 4601 6325 4621
rect 6239 4567 6281 4601
rect 6315 4567 6325 4601
rect 6369 4593 6385 4627
rect 6419 4593 6511 4627
rect 6762 4617 6792 4670
rect 6879 4626 6909 4715
rect 7067 4685 7097 4765
rect 6369 4577 6511 4593
rect 6553 4591 6695 4607
rect 6239 4551 6325 4567
rect 6553 4557 6645 4591
rect 6679 4557 6695 4591
rect 5633 4535 5717 4541
rect 4187 4401 4217 4427
rect 4271 4401 4301 4427
rect 5507 4509 5717 4535
rect 5875 4529 5905 4551
rect 6063 4529 6093 4551
rect 6155 4529 6185 4551
rect 6239 4529 6269 4551
rect 6553 4541 6695 4557
rect 6738 4601 6792 4617
rect 6738 4567 6748 4601
rect 6782 4567 6792 4601
rect 6834 4616 6909 4626
rect 7002 4669 7097 4685
rect 7002 4635 7012 4669
rect 7046 4635 7097 4669
rect 7152 4649 7182 4765
rect 7247 4733 7277 4765
rect 7247 4717 7308 4733
rect 7247 4683 7264 4717
rect 7298 4683 7308 4717
rect 7247 4667 7308 4683
rect 7002 4619 7097 4635
rect 6834 4582 6850 4616
rect 6884 4582 6909 4616
rect 6834 4572 6909 4582
rect 6738 4551 6792 4567
rect 6553 4535 6637 4541
rect 6427 4509 6637 4535
rect 6762 4528 6792 4551
rect 6762 4498 6825 4528
rect 6795 4483 6825 4498
rect 6879 4483 6909 4572
rect 7067 4483 7097 4619
rect 7139 4639 7205 4649
rect 7139 4605 7155 4639
rect 7189 4625 7205 4639
rect 7189 4605 7308 4625
rect 7139 4595 7308 4605
rect 7159 4543 7225 4553
rect 7159 4509 7175 4543
rect 7209 4509 7225 4543
rect 7159 4499 7225 4509
rect 7179 4471 7209 4499
rect 7278 4471 7308 4595
rect 7350 4565 7380 4765
rect 7482 4661 7512 4699
rect 7577 4667 7607 4765
rect 7661 4727 7691 4765
rect 7775 4733 7805 4765
rect 7660 4717 7726 4727
rect 7660 4683 7676 4717
rect 7710 4683 7726 4717
rect 7660 4673 7726 4683
rect 7775 4717 7856 4733
rect 7775 4683 7812 4717
rect 7846 4683 7856 4717
rect 7775 4667 7856 4683
rect 7422 4651 7512 4661
rect 7422 4617 7438 4651
rect 7472 4617 7512 4651
rect 7422 4607 7512 4617
rect 7482 4572 7512 4607
rect 7564 4651 7618 4667
rect 7564 4617 7574 4651
rect 7608 4631 7618 4651
rect 7608 4617 7733 4631
rect 7564 4601 7733 4617
rect 7350 4555 7424 4565
rect 7350 4521 7374 4555
rect 7408 4521 7424 4555
rect 7482 4542 7526 4572
rect 7496 4527 7526 4542
rect 7597 4543 7661 4559
rect 7350 4511 7424 4521
rect 7377 4483 7407 4511
rect 7597 4509 7617 4543
rect 7651 4509 7661 4543
rect 7597 4493 7661 4509
rect 7597 4471 7627 4493
rect 7703 4471 7733 4601
rect 7798 4483 7828 4667
rect 8267 4649 8661 4675
rect 9003 4649 9581 4675
rect 7985 4617 8015 4649
rect 8069 4617 8099 4649
rect 8267 4627 8443 4649
rect 7875 4601 8017 4617
rect 7875 4567 7885 4601
rect 7919 4567 8017 4601
rect 7875 4551 8017 4567
rect 8059 4601 8113 4617
rect 8059 4567 8069 4601
rect 8103 4567 8113 4601
rect 8267 4593 8283 4627
rect 8317 4593 8393 4627
rect 8427 4593 8443 4627
rect 9003 4627 9267 4649
rect 9739 4645 9857 4675
rect 10319 4733 10349 4765
rect 10268 4717 10349 4733
rect 10433 4727 10463 4765
rect 10268 4683 10278 4717
rect 10312 4683 10349 4717
rect 10268 4667 10349 4683
rect 10398 4717 10464 4727
rect 10398 4683 10414 4717
rect 10448 4683 10464 4717
rect 10398 4673 10464 4683
rect 10517 4667 10547 4765
rect 11215 4843 11245 4869
rect 11299 4843 11329 4869
rect 11487 4849 11697 4875
rect 11859 4849 11889 4875
rect 12020 4849 12050 4875
rect 12128 4849 12158 4875
rect 12219 4849 12249 4875
rect 12407 4849 12617 4875
rect 12779 4849 12809 4875
rect 12940 4849 12970 4875
rect 13048 4849 13078 4875
rect 13139 4849 13169 4875
rect 13327 4849 13905 4875
rect 14155 4849 14273 4875
rect 14659 4849 14689 4875
rect 14891 4849 15837 4875
rect 15995 4849 16941 4875
rect 17099 4849 18045 4875
rect 18203 4849 18413 4875
rect 18663 4849 18781 4875
rect 9739 4643 9777 4645
rect 8267 4577 8443 4593
rect 8485 4591 8661 4607
rect 8059 4551 8113 4567
rect 8485 4557 8501 4591
rect 8535 4557 8611 4591
rect 8645 4557 8661 4591
rect 9003 4593 9019 4627
rect 9053 4593 9118 4627
rect 9152 4593 9217 4627
rect 9251 4593 9267 4627
rect 9711 4627 9777 4643
rect 9003 4577 9267 4593
rect 9309 4591 9581 4607
rect 7987 4529 8017 4551
rect 8071 4529 8101 4551
rect 8485 4535 8661 4557
rect 9309 4557 9325 4591
rect 9359 4557 9428 4591
rect 9462 4557 9531 4591
rect 9565 4557 9581 4591
rect 9711 4593 9727 4627
rect 9761 4593 9777 4627
rect 10025 4617 10055 4649
rect 10109 4617 10139 4649
rect 9711 4577 9777 4593
rect 9819 4587 9885 4603
rect 9309 4535 9581 4557
rect 9819 4553 9835 4587
rect 9869 4553 9885 4587
rect 9819 4537 9885 4553
rect 10011 4601 10065 4617
rect 10011 4567 10021 4601
rect 10055 4567 10065 4601
rect 10011 4551 10065 4567
rect 10107 4601 10249 4617
rect 10107 4567 10205 4601
rect 10239 4567 10249 4601
rect 10107 4551 10249 4567
rect 9819 4535 9857 4537
rect 8267 4509 8661 4535
rect 9003 4509 9581 4535
rect 9739 4509 9857 4535
rect 10023 4529 10053 4551
rect 10107 4529 10137 4551
rect 10296 4483 10326 4667
rect 10506 4651 10560 4667
rect 10506 4631 10516 4651
rect 10391 4617 10516 4631
rect 10550 4617 10560 4651
rect 10391 4601 10560 4617
rect 10612 4661 10642 4699
rect 10612 4651 10702 4661
rect 10612 4617 10652 4651
rect 10686 4617 10702 4651
rect 10612 4607 10702 4617
rect 10391 4471 10421 4601
rect 10612 4572 10642 4607
rect 10463 4543 10527 4559
rect 10463 4509 10473 4543
rect 10507 4509 10527 4543
rect 10598 4542 10642 4572
rect 10744 4565 10774 4765
rect 10847 4733 10877 4765
rect 10816 4717 10877 4733
rect 10816 4683 10826 4717
rect 10860 4683 10877 4717
rect 10816 4667 10877 4683
rect 10942 4649 10972 4765
rect 11027 4685 11057 4765
rect 11027 4669 11122 4685
rect 10919 4639 10985 4649
rect 10919 4625 10935 4639
rect 10700 4555 10774 4565
rect 10598 4527 10628 4542
rect 10463 4493 10527 4509
rect 10497 4471 10527 4493
rect 10700 4521 10716 4555
rect 10750 4521 10774 4555
rect 10700 4511 10774 4521
rect 10816 4605 10935 4625
rect 10969 4605 10985 4639
rect 10816 4595 10985 4605
rect 11027 4635 11078 4669
rect 11112 4635 11122 4669
rect 11027 4619 11122 4635
rect 11215 4626 11245 4715
rect 11299 4700 11329 4715
rect 11299 4670 11362 4700
rect 10717 4483 10747 4511
rect 10816 4471 10846 4595
rect 10899 4543 10965 4553
rect 10899 4509 10915 4543
rect 10949 4509 10965 4543
rect 10899 4499 10965 4509
rect 10915 4471 10945 4499
rect 11027 4483 11057 4619
rect 11215 4616 11290 4626
rect 11215 4582 11240 4616
rect 11274 4582 11290 4616
rect 11215 4572 11290 4582
rect 11332 4617 11362 4670
rect 11487 4649 11697 4675
rect 12407 4649 12617 4675
rect 13327 4649 13905 4675
rect 14467 4807 14497 4833
rect 14551 4807 14581 4833
rect 11487 4643 11571 4649
rect 11429 4627 11571 4643
rect 11332 4601 11386 4617
rect 11215 4483 11245 4572
rect 11332 4567 11342 4601
rect 11376 4567 11386 4601
rect 11429 4593 11445 4627
rect 11479 4593 11571 4627
rect 11859 4617 11889 4649
rect 12020 4617 12050 4649
rect 12128 4617 12158 4649
rect 12219 4621 12249 4649
rect 12407 4643 12491 4649
rect 12349 4627 12491 4643
rect 11429 4577 11571 4593
rect 11613 4591 11755 4607
rect 11332 4551 11386 4567
rect 11613 4557 11705 4591
rect 11739 4557 11755 4591
rect 11332 4528 11362 4551
rect 11613 4541 11755 4557
rect 11855 4601 11939 4617
rect 11855 4567 11895 4601
rect 11929 4567 11939 4601
rect 11855 4551 11939 4567
rect 12020 4601 12077 4617
rect 12020 4567 12033 4601
rect 12067 4567 12077 4601
rect 12020 4551 12077 4567
rect 12123 4601 12177 4617
rect 12123 4567 12133 4601
rect 12167 4567 12177 4601
rect 12123 4551 12177 4567
rect 12219 4601 12305 4621
rect 12219 4567 12261 4601
rect 12295 4567 12305 4601
rect 12349 4593 12365 4627
rect 12399 4593 12491 4627
rect 12779 4617 12809 4649
rect 12940 4617 12970 4649
rect 13048 4617 13078 4649
rect 13139 4621 13169 4649
rect 13327 4627 13591 4649
rect 14155 4645 14273 4675
rect 14155 4643 14193 4645
rect 12349 4577 12491 4593
rect 12533 4591 12675 4607
rect 12219 4551 12305 4567
rect 12533 4557 12625 4591
rect 12659 4557 12675 4591
rect 11613 4535 11697 4541
rect 11299 4498 11362 4528
rect 11487 4509 11697 4535
rect 11855 4529 11885 4551
rect 12043 4529 12073 4551
rect 12135 4529 12165 4551
rect 12219 4529 12249 4551
rect 12533 4541 12675 4557
rect 12775 4601 12859 4617
rect 12775 4567 12815 4601
rect 12849 4567 12859 4601
rect 12775 4551 12859 4567
rect 12940 4601 12997 4617
rect 12940 4567 12953 4601
rect 12987 4567 12997 4601
rect 12940 4551 12997 4567
rect 13043 4601 13097 4617
rect 13043 4567 13053 4601
rect 13087 4567 13097 4601
rect 13043 4551 13097 4567
rect 13139 4601 13225 4621
rect 13139 4567 13181 4601
rect 13215 4567 13225 4601
rect 13327 4593 13343 4627
rect 13377 4593 13442 4627
rect 13476 4593 13541 4627
rect 13575 4593 13591 4627
rect 14127 4627 14193 4643
rect 13327 4577 13591 4593
rect 13633 4591 13905 4607
rect 13139 4551 13225 4567
rect 13633 4557 13649 4591
rect 13683 4557 13752 4591
rect 13786 4557 13855 4591
rect 13889 4557 13905 4591
rect 14127 4593 14143 4627
rect 14177 4593 14193 4627
rect 14467 4617 14497 4723
rect 14127 4577 14193 4593
rect 14235 4587 14301 4603
rect 12533 4535 12617 4541
rect 11299 4483 11329 4498
rect 12407 4509 12617 4535
rect 12775 4529 12805 4551
rect 12963 4529 12993 4551
rect 13055 4529 13085 4551
rect 13139 4529 13169 4551
rect 13633 4535 13905 4557
rect 14235 4553 14251 4587
rect 14285 4553 14301 4587
rect 14235 4537 14301 4553
rect 14410 4601 14497 4617
rect 14410 4567 14426 4601
rect 14460 4567 14497 4601
rect 14410 4551 14497 4567
rect 14235 4535 14273 4537
rect 13327 4509 13905 4535
rect 14155 4509 14273 4535
rect 14467 4511 14497 4551
rect 14551 4617 14581 4723
rect 14891 4649 15837 4675
rect 15995 4649 16941 4675
rect 17099 4649 18045 4675
rect 18203 4649 18413 4675
rect 14659 4617 14689 4649
rect 14891 4627 15341 4649
rect 14551 4601 14617 4617
rect 14551 4567 14567 4601
rect 14601 4567 14617 4601
rect 14551 4551 14617 4567
rect 14659 4601 14725 4617
rect 14659 4567 14675 4601
rect 14709 4567 14725 4601
rect 14891 4593 15163 4627
rect 15197 4593 15341 4627
rect 15995 4627 16445 4649
rect 14891 4577 15341 4593
rect 15383 4591 15837 4607
rect 14659 4551 14725 4567
rect 15383 4557 15527 4591
rect 15561 4557 15837 4591
rect 15995 4593 16267 4627
rect 16301 4593 16445 4627
rect 17099 4627 17549 4649
rect 18203 4643 18287 4649
rect 18663 4645 18781 4675
rect 15995 4577 16445 4593
rect 16487 4591 16941 4607
rect 14551 4511 14581 4551
rect 14659 4529 14689 4551
rect 15383 4535 15837 4557
rect 16487 4557 16631 4591
rect 16665 4557 16941 4591
rect 17099 4593 17371 4627
rect 17405 4593 17549 4627
rect 18145 4627 18287 4643
rect 17099 4577 17549 4593
rect 17591 4591 18045 4607
rect 16487 4535 16941 4557
rect 17591 4557 17735 4591
rect 17769 4557 18045 4591
rect 18145 4593 18161 4627
rect 18195 4593 18287 4627
rect 18743 4643 18781 4645
rect 18743 4627 18809 4643
rect 18145 4577 18287 4593
rect 18329 4591 18471 4607
rect 17591 4535 18045 4557
rect 18329 4557 18421 4591
rect 18455 4557 18471 4591
rect 18329 4541 18471 4557
rect 18635 4587 18701 4603
rect 18635 4553 18651 4587
rect 18685 4553 18701 4587
rect 18743 4593 18759 4627
rect 18793 4593 18809 4627
rect 18743 4577 18809 4593
rect 18329 4535 18413 4541
rect 18635 4537 18701 4553
rect 14467 4401 14497 4427
rect 14551 4401 14581 4427
rect 14891 4509 15837 4535
rect 15995 4509 16941 4535
rect 17099 4509 18045 4535
rect 18203 4509 18413 4535
rect 18663 4535 18701 4537
rect 18663 4509 18781 4535
rect 1183 4373 1301 4399
rect 1459 4373 1853 4399
rect 2103 4373 2133 4399
rect 2187 4373 2217 4399
rect 2375 4373 2405 4399
rect 2487 4373 2517 4399
rect 2586 4373 2616 4399
rect 2685 4373 2715 4399
rect 2804 4373 2834 4399
rect 2905 4373 2935 4399
rect 3011 4373 3041 4399
rect 3106 4373 3136 4399
rect 3295 4373 3325 4399
rect 3379 4373 3409 4399
rect 4079 4373 4109 4399
rect 4495 4373 4705 4399
rect 4955 4373 4985 4399
rect 5143 4373 5173 4399
rect 5235 4373 5265 4399
rect 5319 4373 5349 4399
rect 5507 4373 5717 4399
rect 5875 4373 5905 4399
rect 6063 4373 6093 4399
rect 6155 4373 6185 4399
rect 6239 4373 6269 4399
rect 6427 4373 6637 4399
rect 6795 4373 6825 4399
rect 6879 4373 6909 4399
rect 7067 4373 7097 4399
rect 7179 4373 7209 4399
rect 7278 4373 7308 4399
rect 7377 4373 7407 4399
rect 7496 4373 7526 4399
rect 7597 4373 7627 4399
rect 7703 4373 7733 4399
rect 7798 4373 7828 4399
rect 7987 4373 8017 4399
rect 8071 4373 8101 4399
rect 8267 4373 8661 4399
rect 9003 4373 9581 4399
rect 9739 4373 9857 4399
rect 10023 4373 10053 4399
rect 10107 4373 10137 4399
rect 10296 4373 10326 4399
rect 10391 4373 10421 4399
rect 10497 4373 10527 4399
rect 10598 4373 10628 4399
rect 10717 4373 10747 4399
rect 10816 4373 10846 4399
rect 10915 4373 10945 4399
rect 11027 4373 11057 4399
rect 11215 4373 11245 4399
rect 11299 4373 11329 4399
rect 11487 4373 11697 4399
rect 11855 4373 11885 4399
rect 12043 4373 12073 4399
rect 12135 4373 12165 4399
rect 12219 4373 12249 4399
rect 12407 4373 12617 4399
rect 12775 4373 12805 4399
rect 12963 4373 12993 4399
rect 13055 4373 13085 4399
rect 13139 4373 13169 4399
rect 13327 4373 13905 4399
rect 14155 4373 14273 4399
rect 14659 4373 14689 4399
rect 14891 4373 15837 4399
rect 15995 4373 16941 4399
rect 17099 4373 18045 4399
rect 18203 4373 18413 4399
rect 18663 4373 18781 4399
rect 1183 4305 1301 4331
rect 1459 4305 1853 4331
rect 2011 4305 2041 4331
rect 2099 4305 2129 4331
rect 2287 4305 2497 4331
rect 2663 4305 2693 4331
rect 2747 4305 2777 4331
rect 2936 4305 2966 4331
rect 3031 4305 3061 4331
rect 3137 4305 3167 4331
rect 3238 4305 3268 4331
rect 3357 4305 3387 4331
rect 3456 4305 3486 4331
rect 3555 4305 3585 4331
rect 3667 4305 3697 4331
rect 3855 4305 3885 4331
rect 3939 4305 3969 4331
rect 4127 4305 4521 4331
rect 4687 4305 4717 4331
rect 4771 4305 4801 4331
rect 4960 4305 4990 4331
rect 5055 4305 5085 4331
rect 5161 4305 5191 4331
rect 5262 4305 5292 4331
rect 5381 4305 5411 4331
rect 5480 4305 5510 4331
rect 5579 4305 5609 4331
rect 5691 4305 5721 4331
rect 5879 4305 5909 4331
rect 5963 4305 5993 4331
rect 6427 4305 6821 4331
rect 6979 4305 7009 4331
rect 7167 4305 7197 4331
rect 7259 4305 7289 4331
rect 7343 4305 7373 4331
rect 7531 4305 7741 4331
rect 7900 4305 7930 4331
rect 7986 4305 8016 4331
rect 8072 4305 8102 4331
rect 8158 4305 8188 4331
rect 8244 4305 8274 4331
rect 8330 4305 8360 4331
rect 8416 4305 8446 4331
rect 8502 4305 8532 4331
rect 8588 4305 8618 4331
rect 8674 4305 8704 4331
rect 8760 4305 8790 4331
rect 8846 4305 8876 4331
rect 8931 4305 8961 4331
rect 9017 4305 9047 4331
rect 9103 4305 9133 4331
rect 9189 4305 9219 4331
rect 9275 4305 9305 4331
rect 9361 4305 9391 4331
rect 9447 4305 9477 4331
rect 9533 4305 9563 4331
rect 9739 4305 10317 4331
rect 10567 4305 10597 4331
rect 10755 4305 10785 4331
rect 10847 4305 10877 4331
rect 10931 4305 10961 4331
rect 11119 4305 11329 4331
rect 11763 4305 11793 4331
rect 11847 4305 11877 4331
rect 12035 4305 12065 4331
rect 12147 4305 12177 4331
rect 12246 4305 12276 4331
rect 12345 4305 12375 4331
rect 12464 4305 12494 4331
rect 12565 4305 12595 4331
rect 12671 4305 12701 4331
rect 12766 4305 12796 4331
rect 12955 4305 12985 4331
rect 13039 4305 13069 4331
rect 13235 4305 14181 4331
rect 14339 4305 15285 4331
rect 15535 4305 15565 4331
rect 15623 4305 15653 4331
rect 15811 4305 16389 4331
rect 17143 4305 17173 4331
rect 17375 4305 18321 4331
rect 18663 4305 18781 4331
rect 1183 4169 1301 4195
rect 1459 4169 1853 4195
rect 2011 4186 2041 4201
rect 1263 4167 1301 4169
rect 1263 4151 1329 4167
rect 1155 4111 1221 4127
rect 1155 4077 1171 4111
rect 1205 4077 1221 4111
rect 1263 4117 1279 4151
rect 1313 4117 1329 4151
rect 1677 4147 1853 4169
rect 2005 4162 2041 4186
rect 2005 4153 2035 4162
rect 1263 4101 1329 4117
rect 1459 4111 1635 4127
rect 1155 4061 1221 4077
rect 1183 4059 1221 4061
rect 1459 4077 1475 4111
rect 1509 4077 1585 4111
rect 1619 4077 1635 4111
rect 1677 4113 1693 4147
rect 1727 4113 1803 4147
rect 1837 4113 1853 4147
rect 1677 4097 1853 4113
rect 1959 4137 2035 4153
rect 2099 4140 2129 4201
rect 2287 4169 2497 4195
rect 2413 4163 2497 4169
rect 2413 4147 2555 4163
rect 2663 4153 2693 4175
rect 2747 4153 2777 4175
rect 1959 4103 1969 4137
rect 2003 4103 2035 4137
rect 1959 4087 2035 4103
rect 1183 4029 1301 4059
rect 1459 4055 1635 4077
rect 1459 4029 1853 4055
rect 2005 4052 2035 4087
rect 2079 4124 2133 4140
rect 2079 4090 2089 4124
rect 2123 4090 2133 4124
rect 2079 4074 2133 4090
rect 2229 4111 2371 4127
rect 2229 4077 2245 4111
rect 2279 4077 2371 4111
rect 2413 4113 2505 4147
rect 2539 4113 2555 4147
rect 2413 4097 2555 4113
rect 2651 4137 2705 4153
rect 2651 4103 2661 4137
rect 2695 4103 2705 4137
rect 2651 4087 2705 4103
rect 2747 4137 2889 4153
rect 2747 4103 2845 4137
rect 2879 4103 2889 4137
rect 2747 4087 2889 4103
rect 2005 4028 2041 4052
rect 2011 4013 2041 4028
rect 2099 4013 2129 4074
rect 2229 4061 2371 4077
rect 2287 4055 2371 4061
rect 2665 4055 2695 4087
rect 2749 4055 2779 4087
rect 2287 4029 2497 4055
rect 2936 4037 2966 4221
rect 3031 4103 3061 4233
rect 3137 4211 3167 4233
rect 3103 4195 3167 4211
rect 3103 4161 3113 4195
rect 3147 4161 3167 4195
rect 3357 4193 3387 4221
rect 3340 4183 3414 4193
rect 3103 4145 3167 4161
rect 3238 4162 3268 4177
rect 3238 4132 3282 4162
rect 3340 4149 3356 4183
rect 3390 4149 3414 4183
rect 3340 4139 3414 4149
rect 3031 4087 3200 4103
rect 3031 4073 3156 4087
rect 3146 4053 3156 4073
rect 3190 4053 3200 4087
rect 3146 4037 3200 4053
rect 3252 4097 3282 4132
rect 3252 4087 3342 4097
rect 3252 4053 3292 4087
rect 3326 4053 3342 4087
rect 3252 4043 3342 4053
rect 2908 4021 2989 4037
rect 2908 3987 2918 4021
rect 2952 3987 2989 4021
rect 2908 3971 2989 3987
rect 3038 4021 3104 4031
rect 3038 3987 3054 4021
rect 3088 3987 3104 4021
rect 3038 3977 3104 3987
rect 2959 3939 2989 3971
rect 3073 3939 3103 3977
rect 3157 3939 3187 4037
rect 3252 4005 3282 4043
rect 3384 3939 3414 4139
rect 3456 4109 3486 4233
rect 3555 4205 3585 4233
rect 3539 4195 3605 4205
rect 3539 4161 3555 4195
rect 3589 4161 3605 4195
rect 3539 4151 3605 4161
rect 3456 4099 3625 4109
rect 3456 4079 3575 4099
rect 3559 4065 3575 4079
rect 3609 4065 3625 4099
rect 3559 4055 3625 4065
rect 3667 4085 3697 4221
rect 3855 4132 3885 4221
rect 3939 4206 3969 4221
rect 3939 4176 4002 4206
rect 3972 4153 4002 4176
rect 4127 4169 4521 4195
rect 3972 4137 4026 4153
rect 3855 4122 3930 4132
rect 3855 4088 3880 4122
rect 3914 4088 3930 4122
rect 3667 4069 3762 4085
rect 3456 4021 3517 4037
rect 3456 3987 3466 4021
rect 3500 3987 3517 4021
rect 3456 3971 3517 3987
rect 3487 3939 3517 3971
rect 3582 3939 3612 4055
rect 3667 4035 3718 4069
rect 3752 4035 3762 4069
rect 3667 4019 3762 4035
rect 3855 4078 3930 4088
rect 3972 4103 3982 4137
rect 4016 4103 4026 4137
rect 4345 4147 4521 4169
rect 4687 4153 4717 4175
rect 4771 4153 4801 4175
rect 3972 4087 4026 4103
rect 4127 4111 4303 4127
rect 3667 3939 3697 4019
rect 3855 3989 3885 4078
rect 3972 4034 4002 4087
rect 3939 4004 4002 4034
rect 4127 4077 4143 4111
rect 4177 4077 4253 4111
rect 4287 4077 4303 4111
rect 4345 4113 4361 4147
rect 4395 4113 4471 4147
rect 4505 4113 4521 4147
rect 4345 4097 4521 4113
rect 4675 4137 4729 4153
rect 4675 4103 4685 4137
rect 4719 4103 4729 4137
rect 4675 4087 4729 4103
rect 4771 4137 4913 4153
rect 4771 4103 4869 4137
rect 4903 4103 4913 4137
rect 4771 4087 4913 4103
rect 4127 4055 4303 4077
rect 4689 4055 4719 4087
rect 4773 4055 4803 4087
rect 4127 4029 4521 4055
rect 3939 3989 3969 4004
rect 1183 3829 1301 3855
rect 1459 3829 1853 3855
rect 2011 3829 2041 3855
rect 2099 3829 2129 3855
rect 2287 3829 2497 3855
rect 2665 3829 2695 3855
rect 2749 3829 2779 3855
rect 2959 3829 2989 3855
rect 3073 3829 3103 3855
rect 3157 3829 3187 3855
rect 3252 3829 3282 3855
rect 3384 3829 3414 3855
rect 3487 3829 3517 3855
rect 3582 3829 3612 3855
rect 3667 3829 3697 3855
rect 3855 3835 3885 3861
rect 3939 3835 3969 3861
rect 4960 4037 4990 4221
rect 5055 4103 5085 4233
rect 5161 4211 5191 4233
rect 5127 4195 5191 4211
rect 5127 4161 5137 4195
rect 5171 4161 5191 4195
rect 5381 4193 5411 4221
rect 5364 4183 5438 4193
rect 5127 4145 5191 4161
rect 5262 4162 5292 4177
rect 5262 4132 5306 4162
rect 5364 4149 5380 4183
rect 5414 4149 5438 4183
rect 5364 4139 5438 4149
rect 5055 4087 5224 4103
rect 5055 4073 5180 4087
rect 5170 4053 5180 4073
rect 5214 4053 5224 4087
rect 5170 4037 5224 4053
rect 5276 4097 5306 4132
rect 5276 4087 5366 4097
rect 5276 4053 5316 4087
rect 5350 4053 5366 4087
rect 5276 4043 5366 4053
rect 4932 4021 5013 4037
rect 4932 3987 4942 4021
rect 4976 3987 5013 4021
rect 4932 3971 5013 3987
rect 5062 4021 5128 4031
rect 5062 3987 5078 4021
rect 5112 3987 5128 4021
rect 5062 3977 5128 3987
rect 4983 3939 5013 3971
rect 5097 3939 5127 3977
rect 5181 3939 5211 4037
rect 5276 4005 5306 4043
rect 5408 3939 5438 4139
rect 5480 4109 5510 4233
rect 5579 4205 5609 4233
rect 5563 4195 5629 4205
rect 5563 4161 5579 4195
rect 5613 4161 5629 4195
rect 5563 4151 5629 4161
rect 5480 4099 5649 4109
rect 5480 4079 5599 4099
rect 5583 4065 5599 4079
rect 5633 4065 5649 4099
rect 5583 4055 5649 4065
rect 5691 4085 5721 4221
rect 5879 4132 5909 4221
rect 5963 4206 5993 4221
rect 5963 4176 6026 4206
rect 5996 4153 6026 4176
rect 6427 4169 6821 4195
rect 5996 4137 6050 4153
rect 5879 4122 5954 4132
rect 5879 4088 5904 4122
rect 5938 4088 5954 4122
rect 5691 4069 5786 4085
rect 5480 4021 5541 4037
rect 5480 3987 5490 4021
rect 5524 3987 5541 4021
rect 5480 3971 5541 3987
rect 5511 3939 5541 3971
rect 5606 3939 5636 4055
rect 5691 4035 5742 4069
rect 5776 4035 5786 4069
rect 5691 4019 5786 4035
rect 5879 4078 5954 4088
rect 5996 4103 6006 4137
rect 6040 4103 6050 4137
rect 6645 4147 6821 4169
rect 5996 4087 6050 4103
rect 6427 4111 6603 4127
rect 5691 3939 5721 4019
rect 5879 3989 5909 4078
rect 5996 4034 6026 4087
rect 6427 4077 6443 4111
rect 6477 4077 6553 4111
rect 6587 4077 6603 4111
rect 6645 4113 6661 4147
rect 6695 4113 6771 4147
rect 6805 4113 6821 4147
rect 6645 4097 6821 4113
rect 6979 4153 7009 4175
rect 7167 4153 7197 4175
rect 7259 4153 7289 4175
rect 7343 4153 7373 4175
rect 7531 4169 7741 4195
rect 7900 4172 7930 4221
rect 7986 4172 8016 4221
rect 8072 4172 8102 4221
rect 8158 4172 8188 4221
rect 7657 4163 7741 4169
rect 6979 4137 7063 4153
rect 6979 4103 7019 4137
rect 7053 4103 7063 4137
rect 6979 4087 7063 4103
rect 7144 4137 7201 4153
rect 7144 4103 7157 4137
rect 7191 4103 7201 4137
rect 7144 4087 7201 4103
rect 7247 4137 7301 4153
rect 7247 4103 7257 4137
rect 7291 4103 7301 4137
rect 7247 4087 7301 4103
rect 7343 4137 7429 4153
rect 7343 4103 7385 4137
rect 7419 4103 7429 4137
rect 7657 4147 7799 4163
rect 6427 4055 6603 4077
rect 6983 4055 7013 4087
rect 7144 4055 7174 4087
rect 7252 4055 7282 4087
rect 7343 4083 7429 4103
rect 7473 4111 7615 4127
rect 7343 4055 7373 4083
rect 7473 4077 7489 4111
rect 7523 4077 7615 4111
rect 7657 4113 7749 4147
rect 7783 4113 7799 4147
rect 7657 4097 7799 4113
rect 7841 4137 8188 4172
rect 7841 4103 7857 4137
rect 7891 4103 8188 4137
rect 7473 4061 7615 4077
rect 7841 4070 8188 4103
rect 7531 4055 7615 4061
rect 7900 4055 7930 4070
rect 7986 4055 8016 4070
rect 8072 4055 8102 4070
rect 8158 4055 8188 4070
rect 8244 4162 8274 4221
rect 8330 4162 8360 4221
rect 8416 4162 8446 4221
rect 8502 4162 8532 4221
rect 8588 4162 8618 4221
rect 8674 4162 8704 4221
rect 8760 4162 8790 4221
rect 8846 4162 8876 4221
rect 8931 4162 8961 4221
rect 9017 4162 9047 4221
rect 9103 4162 9133 4221
rect 9189 4162 9219 4221
rect 9275 4162 9305 4221
rect 9361 4162 9391 4221
rect 9447 4162 9477 4221
rect 9533 4162 9563 4221
rect 9739 4169 10317 4195
rect 8244 4137 9563 4162
rect 8244 4103 8284 4137
rect 8318 4103 8352 4137
rect 8386 4103 8420 4137
rect 8454 4103 8488 4137
rect 8522 4103 8556 4137
rect 8590 4103 8624 4137
rect 8658 4103 8692 4137
rect 8726 4103 8760 4137
rect 8794 4103 8828 4137
rect 8862 4103 8896 4137
rect 8930 4103 8964 4137
rect 8998 4103 9032 4137
rect 9066 4103 9100 4137
rect 9134 4103 9168 4137
rect 9202 4103 9236 4137
rect 9270 4103 9304 4137
rect 9338 4103 9563 4137
rect 10045 4147 10317 4169
rect 8244 4087 9563 4103
rect 8244 4055 8274 4087
rect 8330 4055 8360 4087
rect 8416 4055 8446 4087
rect 8502 4055 8532 4087
rect 8588 4055 8618 4087
rect 8674 4055 8704 4087
rect 8760 4055 8790 4087
rect 8846 4055 8876 4087
rect 8931 4055 8961 4087
rect 9017 4055 9047 4087
rect 9103 4055 9133 4087
rect 9189 4055 9219 4087
rect 9275 4055 9305 4087
rect 9361 4055 9391 4087
rect 9447 4055 9477 4087
rect 9533 4055 9563 4087
rect 9739 4111 10003 4127
rect 9739 4077 9755 4111
rect 9789 4077 9854 4111
rect 9888 4077 9953 4111
rect 9987 4077 10003 4111
rect 10045 4113 10061 4147
rect 10095 4113 10164 4147
rect 10198 4113 10267 4147
rect 10301 4113 10317 4147
rect 10045 4097 10317 4113
rect 10567 4153 10597 4175
rect 10755 4153 10785 4175
rect 10847 4153 10877 4175
rect 10931 4153 10961 4175
rect 11119 4169 11329 4195
rect 11763 4206 11793 4221
rect 11245 4163 11329 4169
rect 11730 4176 11793 4206
rect 10567 4137 10651 4153
rect 10567 4103 10607 4137
rect 10641 4103 10651 4137
rect 10567 4087 10651 4103
rect 10732 4137 10789 4153
rect 10732 4103 10745 4137
rect 10779 4103 10789 4137
rect 10732 4087 10789 4103
rect 10835 4137 10889 4153
rect 10835 4103 10845 4137
rect 10879 4103 10889 4137
rect 10835 4087 10889 4103
rect 10931 4137 11017 4153
rect 10931 4103 10973 4137
rect 11007 4103 11017 4137
rect 11245 4147 11387 4163
rect 11730 4153 11760 4176
rect 9739 4055 10003 4077
rect 10571 4055 10601 4087
rect 10732 4055 10762 4087
rect 10840 4055 10870 4087
rect 10931 4083 11017 4103
rect 11061 4111 11203 4127
rect 10931 4055 10961 4083
rect 11061 4077 11077 4111
rect 11111 4077 11203 4111
rect 11245 4113 11337 4147
rect 11371 4113 11387 4147
rect 11245 4097 11387 4113
rect 11706 4137 11760 4153
rect 11706 4103 11716 4137
rect 11750 4103 11760 4137
rect 11847 4132 11877 4221
rect 11706 4087 11760 4103
rect 11061 4061 11203 4077
rect 11119 4055 11203 4061
rect 5963 4004 6026 4034
rect 6427 4029 6821 4055
rect 5963 3989 5993 4004
rect 4127 3829 4521 3855
rect 4689 3829 4719 3855
rect 4773 3829 4803 3855
rect 4983 3829 5013 3855
rect 5097 3829 5127 3855
rect 5181 3829 5211 3855
rect 5276 3829 5306 3855
rect 5408 3829 5438 3855
rect 5511 3829 5541 3855
rect 5606 3829 5636 3855
rect 5691 3829 5721 3855
rect 5879 3835 5909 3861
rect 5963 3835 5993 3861
rect 7531 4029 7741 4055
rect 9739 4029 10317 4055
rect 11119 4029 11329 4055
rect 11730 4034 11760 4087
rect 11802 4122 11877 4132
rect 11802 4088 11818 4122
rect 11852 4088 11877 4122
rect 11802 4078 11877 4088
rect 12035 4085 12065 4221
rect 12147 4205 12177 4233
rect 12127 4195 12193 4205
rect 12127 4161 12143 4195
rect 12177 4161 12193 4195
rect 12127 4151 12193 4161
rect 12246 4109 12276 4233
rect 12345 4193 12375 4221
rect 11730 4004 11793 4034
rect 11763 3989 11793 4004
rect 11847 3989 11877 4078
rect 11970 4069 12065 4085
rect 11970 4035 11980 4069
rect 12014 4035 12065 4069
rect 12107 4099 12276 4109
rect 12107 4065 12123 4099
rect 12157 4079 12276 4099
rect 12318 4183 12392 4193
rect 12318 4149 12342 4183
rect 12376 4149 12392 4183
rect 12565 4211 12595 4233
rect 12565 4195 12629 4211
rect 12464 4162 12494 4177
rect 12318 4139 12392 4149
rect 12157 4065 12173 4079
rect 12107 4055 12173 4065
rect 11970 4019 12065 4035
rect 12035 3939 12065 4019
rect 12120 3939 12150 4055
rect 12215 4021 12276 4037
rect 12215 3987 12232 4021
rect 12266 3987 12276 4021
rect 12215 3971 12276 3987
rect 12215 3939 12245 3971
rect 12318 3939 12348 4139
rect 12450 4132 12494 4162
rect 12565 4161 12585 4195
rect 12619 4161 12629 4195
rect 12565 4145 12629 4161
rect 12450 4097 12480 4132
rect 12671 4103 12701 4233
rect 12390 4087 12480 4097
rect 12390 4053 12406 4087
rect 12440 4053 12480 4087
rect 12390 4043 12480 4053
rect 12450 4005 12480 4043
rect 12532 4087 12701 4103
rect 12532 4053 12542 4087
rect 12576 4073 12701 4087
rect 12576 4053 12586 4073
rect 12532 4037 12586 4053
rect 12766 4037 12796 4221
rect 12955 4153 12985 4175
rect 13039 4153 13069 4175
rect 13235 4169 14181 4195
rect 14339 4169 15285 4195
rect 12843 4137 12985 4153
rect 12843 4103 12853 4137
rect 12887 4103 12985 4137
rect 12843 4087 12985 4103
rect 13027 4137 13081 4153
rect 13027 4103 13037 4137
rect 13071 4103 13081 4137
rect 13727 4147 14181 4169
rect 13027 4087 13081 4103
rect 13235 4111 13685 4127
rect 12953 4055 12983 4087
rect 13037 4055 13067 4087
rect 13235 4077 13507 4111
rect 13541 4077 13685 4111
rect 13727 4113 13871 4147
rect 13905 4113 14181 4147
rect 14831 4147 15285 4169
rect 13727 4097 14181 4113
rect 14339 4111 14789 4127
rect 13235 4055 13685 4077
rect 14339 4077 14611 4111
rect 14645 4077 14789 4111
rect 14831 4113 14975 4147
rect 15009 4113 15285 4147
rect 15535 4140 15565 4201
rect 15623 4186 15653 4201
rect 16951 4277 16981 4303
rect 17035 4277 17065 4303
rect 15623 4162 15659 4186
rect 15811 4169 16389 4195
rect 15629 4153 15659 4162
rect 14831 4097 15285 4113
rect 15531 4124 15585 4140
rect 14339 4055 14789 4077
rect 15531 4090 15541 4124
rect 15575 4090 15585 4124
rect 15531 4074 15585 4090
rect 15629 4137 15705 4153
rect 15629 4103 15661 4137
rect 15695 4103 15705 4137
rect 16117 4147 16389 4169
rect 16951 4153 16981 4193
rect 15629 4087 15705 4103
rect 15811 4111 16075 4127
rect 6427 3829 6821 3855
rect 6983 3829 7013 3855
rect 7144 3829 7174 3855
rect 7252 3829 7282 3855
rect 7343 3829 7373 3855
rect 7531 3829 7741 3855
rect 7900 3829 7930 3855
rect 7986 3829 8016 3855
rect 8072 3829 8102 3855
rect 8158 3829 8188 3855
rect 8244 3829 8274 3855
rect 8330 3829 8360 3855
rect 8416 3829 8446 3855
rect 8502 3829 8532 3855
rect 8588 3829 8618 3855
rect 8674 3829 8704 3855
rect 8760 3829 8790 3855
rect 8846 3829 8876 3855
rect 8931 3829 8961 3855
rect 9017 3829 9047 3855
rect 9103 3829 9133 3855
rect 9189 3829 9219 3855
rect 9275 3829 9305 3855
rect 9361 3829 9391 3855
rect 9447 3829 9477 3855
rect 9533 3829 9563 3855
rect 9739 3829 10317 3855
rect 10571 3829 10601 3855
rect 10732 3829 10762 3855
rect 10840 3829 10870 3855
rect 10931 3829 10961 3855
rect 11119 3829 11329 3855
rect 11763 3835 11793 3861
rect 11847 3835 11877 3861
rect 12545 3939 12575 4037
rect 12628 4021 12694 4031
rect 12628 3987 12644 4021
rect 12678 3987 12694 4021
rect 12628 3977 12694 3987
rect 12743 4021 12824 4037
rect 12743 3987 12780 4021
rect 12814 3987 12824 4021
rect 12629 3939 12659 3977
rect 12743 3971 12824 3987
rect 12743 3939 12773 3971
rect 13235 4029 14181 4055
rect 14339 4029 15285 4055
rect 15535 4013 15565 4074
rect 15629 4052 15659 4087
rect 15623 4028 15659 4052
rect 15811 4077 15827 4111
rect 15861 4077 15926 4111
rect 15960 4077 16025 4111
rect 16059 4077 16075 4111
rect 16117 4113 16133 4147
rect 16167 4113 16236 4147
rect 16270 4113 16339 4147
rect 16373 4113 16389 4147
rect 16117 4097 16389 4113
rect 16894 4137 16981 4153
rect 16894 4103 16910 4137
rect 16944 4103 16981 4137
rect 16894 4087 16981 4103
rect 15811 4055 16075 4077
rect 15811 4029 16389 4055
rect 15623 4013 15653 4028
rect 16951 3981 16981 4087
rect 17035 4153 17065 4193
rect 17143 4153 17173 4175
rect 17375 4169 18321 4195
rect 17035 4137 17101 4153
rect 17035 4103 17051 4137
rect 17085 4103 17101 4137
rect 17035 4087 17101 4103
rect 17143 4137 17209 4153
rect 17143 4103 17159 4137
rect 17193 4103 17209 4137
rect 17867 4147 18321 4169
rect 18663 4169 18781 4195
rect 18663 4167 18701 4169
rect 17143 4087 17209 4103
rect 17375 4111 17825 4127
rect 17035 3981 17065 4087
rect 17143 4055 17173 4087
rect 17375 4077 17647 4111
rect 17681 4077 17825 4111
rect 17867 4113 18011 4147
rect 18045 4113 18321 4147
rect 17867 4097 18321 4113
rect 18635 4151 18701 4167
rect 18635 4117 18651 4151
rect 18685 4117 18701 4151
rect 18635 4101 18701 4117
rect 18743 4111 18809 4127
rect 17375 4055 17825 4077
rect 18743 4077 18759 4111
rect 18793 4077 18809 4111
rect 18743 4061 18809 4077
rect 18743 4059 18781 4061
rect 16951 3871 16981 3897
rect 17035 3871 17065 3897
rect 17375 4029 18321 4055
rect 18663 4029 18781 4059
rect 12035 3829 12065 3855
rect 12120 3829 12150 3855
rect 12215 3829 12245 3855
rect 12318 3829 12348 3855
rect 12450 3829 12480 3855
rect 12545 3829 12575 3855
rect 12629 3829 12659 3855
rect 12743 3829 12773 3855
rect 12953 3829 12983 3855
rect 13037 3829 13067 3855
rect 13235 3829 14181 3855
rect 14339 3829 15285 3855
rect 15535 3829 15565 3855
rect 15623 3829 15653 3855
rect 15811 3829 16389 3855
rect 17143 3829 17173 3855
rect 17375 3829 18321 3855
rect 18663 3829 18781 3855
rect 1183 3761 1301 3787
rect 1459 3761 1853 3787
rect 2103 3755 2133 3781
rect 2187 3755 2217 3781
rect 2375 3761 2405 3787
rect 2460 3761 2490 3787
rect 2555 3761 2585 3787
rect 2658 3761 2688 3787
rect 2790 3761 2820 3787
rect 2885 3761 2915 3787
rect 2969 3761 2999 3787
rect 3083 3761 3113 3787
rect 3293 3761 3323 3787
rect 3377 3761 3407 3787
rect 2103 3612 2133 3627
rect 1183 3557 1301 3587
rect 1459 3561 1853 3587
rect 2070 3582 2133 3612
rect 1183 3555 1221 3557
rect 1155 3539 1221 3555
rect 1155 3505 1171 3539
rect 1205 3505 1221 3539
rect 1459 3539 1635 3561
rect 1155 3489 1221 3505
rect 1263 3499 1329 3515
rect 1263 3465 1279 3499
rect 1313 3465 1329 3499
rect 1459 3505 1475 3539
rect 1509 3505 1585 3539
rect 1619 3505 1635 3539
rect 2070 3529 2100 3582
rect 2187 3538 2217 3627
rect 2375 3597 2405 3677
rect 1459 3489 1635 3505
rect 1677 3503 1853 3519
rect 1263 3449 1329 3465
rect 1677 3469 1693 3503
rect 1727 3469 1803 3503
rect 1837 3469 1853 3503
rect 1263 3447 1301 3449
rect 1677 3447 1853 3469
rect 2046 3513 2100 3529
rect 2046 3479 2056 3513
rect 2090 3479 2100 3513
rect 2142 3528 2217 3538
rect 2310 3581 2405 3597
rect 2310 3547 2320 3581
rect 2354 3547 2405 3581
rect 2460 3561 2490 3677
rect 2555 3645 2585 3677
rect 2555 3629 2616 3645
rect 2555 3595 2572 3629
rect 2606 3595 2616 3629
rect 2555 3579 2616 3595
rect 2310 3531 2405 3547
rect 2142 3494 2158 3528
rect 2192 3494 2217 3528
rect 2142 3484 2217 3494
rect 2046 3463 2100 3479
rect 1183 3421 1301 3447
rect 1459 3421 1853 3447
rect 2070 3440 2100 3463
rect 2070 3410 2133 3440
rect 2103 3395 2133 3410
rect 2187 3395 2217 3484
rect 2375 3395 2405 3531
rect 2447 3551 2513 3561
rect 2447 3517 2463 3551
rect 2497 3537 2513 3551
rect 2497 3517 2616 3537
rect 2447 3507 2616 3517
rect 2467 3455 2533 3465
rect 2467 3421 2483 3455
rect 2517 3421 2533 3455
rect 2467 3411 2533 3421
rect 2487 3383 2517 3411
rect 2586 3383 2616 3507
rect 2658 3477 2688 3677
rect 2790 3573 2820 3611
rect 2885 3579 2915 3677
rect 2969 3639 2999 3677
rect 3083 3645 3113 3677
rect 2968 3629 3034 3639
rect 2968 3595 2984 3629
rect 3018 3595 3034 3629
rect 2968 3585 3034 3595
rect 3083 3629 3164 3645
rect 3083 3595 3120 3629
rect 3154 3595 3164 3629
rect 3083 3579 3164 3595
rect 2730 3563 2820 3573
rect 2730 3529 2746 3563
rect 2780 3529 2820 3563
rect 2730 3519 2820 3529
rect 2790 3484 2820 3519
rect 2872 3563 2926 3579
rect 2872 3529 2882 3563
rect 2916 3543 2926 3563
rect 2916 3529 3041 3543
rect 2872 3513 3041 3529
rect 2658 3467 2732 3477
rect 2658 3433 2682 3467
rect 2716 3433 2732 3467
rect 2790 3454 2834 3484
rect 2804 3439 2834 3454
rect 2905 3455 2969 3471
rect 2658 3423 2732 3433
rect 2685 3395 2715 3423
rect 2905 3421 2925 3455
rect 2959 3421 2969 3455
rect 2905 3405 2969 3421
rect 2905 3383 2935 3405
rect 3011 3383 3041 3513
rect 3106 3395 3136 3579
rect 4035 3755 4065 3781
rect 4119 3755 4149 3781
rect 4307 3761 4337 3787
rect 4392 3761 4422 3787
rect 4487 3761 4517 3787
rect 4590 3761 4620 3787
rect 4722 3761 4752 3787
rect 4817 3761 4847 3787
rect 4901 3761 4931 3787
rect 5015 3761 5045 3787
rect 5225 3761 5255 3787
rect 5309 3761 5339 3787
rect 5507 3761 6085 3787
rect 6339 3761 6369 3787
rect 6500 3761 6530 3787
rect 6608 3761 6638 3787
rect 6699 3761 6729 3787
rect 6887 3761 7097 3787
rect 4035 3612 4065 3627
rect 4002 3582 4065 3612
rect 3293 3529 3323 3561
rect 3377 3529 3407 3561
rect 4002 3529 4032 3582
rect 4119 3538 4149 3627
rect 4307 3597 4337 3677
rect 3183 3513 3325 3529
rect 3183 3479 3193 3513
rect 3227 3479 3325 3513
rect 3183 3463 3325 3479
rect 3367 3513 3421 3529
rect 3367 3479 3377 3513
rect 3411 3479 3421 3513
rect 3367 3463 3421 3479
rect 3978 3513 4032 3529
rect 3978 3479 3988 3513
rect 4022 3479 4032 3513
rect 4074 3528 4149 3538
rect 4242 3581 4337 3597
rect 4242 3547 4252 3581
rect 4286 3547 4337 3581
rect 4392 3561 4422 3677
rect 4487 3645 4517 3677
rect 4487 3629 4548 3645
rect 4487 3595 4504 3629
rect 4538 3595 4548 3629
rect 4487 3579 4548 3595
rect 4242 3531 4337 3547
rect 4074 3494 4090 3528
rect 4124 3494 4149 3528
rect 4074 3484 4149 3494
rect 3978 3463 4032 3479
rect 3295 3441 3325 3463
rect 3379 3441 3409 3463
rect 4002 3440 4032 3463
rect 4002 3410 4065 3440
rect 4035 3395 4065 3410
rect 4119 3395 4149 3484
rect 4307 3395 4337 3531
rect 4379 3551 4445 3561
rect 4379 3517 4395 3551
rect 4429 3537 4445 3551
rect 4429 3517 4548 3537
rect 4379 3507 4548 3517
rect 4399 3455 4465 3465
rect 4399 3421 4415 3455
rect 4449 3421 4465 3455
rect 4399 3411 4465 3421
rect 4419 3383 4449 3411
rect 4518 3383 4548 3507
rect 4590 3477 4620 3677
rect 4722 3573 4752 3611
rect 4817 3579 4847 3677
rect 4901 3639 4931 3677
rect 5015 3645 5045 3677
rect 4900 3629 4966 3639
rect 4900 3595 4916 3629
rect 4950 3595 4966 3629
rect 4900 3585 4966 3595
rect 5015 3629 5096 3645
rect 5015 3595 5052 3629
rect 5086 3595 5096 3629
rect 5015 3579 5096 3595
rect 4662 3563 4752 3573
rect 4662 3529 4678 3563
rect 4712 3529 4752 3563
rect 4662 3519 4752 3529
rect 4722 3484 4752 3519
rect 4804 3563 4858 3579
rect 4804 3529 4814 3563
rect 4848 3543 4858 3563
rect 4848 3529 4973 3543
rect 4804 3513 4973 3529
rect 4590 3467 4664 3477
rect 4590 3433 4614 3467
rect 4648 3433 4664 3467
rect 4722 3454 4766 3484
rect 4736 3439 4766 3454
rect 4837 3455 4901 3471
rect 4590 3423 4664 3433
rect 4617 3395 4647 3423
rect 4837 3421 4857 3455
rect 4891 3421 4901 3455
rect 4837 3405 4901 3421
rect 4837 3383 4867 3405
rect 4943 3383 4973 3513
rect 5038 3395 5068 3579
rect 5507 3561 6085 3587
rect 7255 3755 7285 3781
rect 7339 3755 7369 3781
rect 7527 3761 7557 3787
rect 7612 3761 7642 3787
rect 7707 3761 7737 3787
rect 7810 3761 7840 3787
rect 7942 3761 7972 3787
rect 8037 3761 8067 3787
rect 8121 3761 8151 3787
rect 8235 3761 8265 3787
rect 8445 3761 8475 3787
rect 8529 3761 8559 3787
rect 9003 3761 9581 3787
rect 7255 3612 7285 3627
rect 6887 3561 7097 3587
rect 7222 3582 7285 3612
rect 5225 3529 5255 3561
rect 5309 3529 5339 3561
rect 5507 3539 5771 3561
rect 5115 3513 5257 3529
rect 5115 3479 5125 3513
rect 5159 3479 5257 3513
rect 5115 3463 5257 3479
rect 5299 3513 5353 3529
rect 5299 3479 5309 3513
rect 5343 3479 5353 3513
rect 5507 3505 5523 3539
rect 5557 3505 5622 3539
rect 5656 3505 5721 3539
rect 5755 3505 5771 3539
rect 6339 3529 6369 3561
rect 6500 3529 6530 3561
rect 6608 3529 6638 3561
rect 6699 3533 6729 3561
rect 6887 3555 6971 3561
rect 6829 3539 6971 3555
rect 5507 3489 5771 3505
rect 5813 3503 6085 3519
rect 5299 3463 5353 3479
rect 5813 3469 5829 3503
rect 5863 3469 5932 3503
rect 5966 3469 6035 3503
rect 6069 3469 6085 3503
rect 5227 3441 5257 3463
rect 5311 3441 5341 3463
rect 5813 3447 6085 3469
rect 5507 3421 6085 3447
rect 6335 3513 6419 3529
rect 6335 3479 6375 3513
rect 6409 3479 6419 3513
rect 6335 3463 6419 3479
rect 6500 3513 6557 3529
rect 6500 3479 6513 3513
rect 6547 3479 6557 3513
rect 6500 3463 6557 3479
rect 6603 3513 6657 3529
rect 6603 3479 6613 3513
rect 6647 3479 6657 3513
rect 6603 3463 6657 3479
rect 6699 3513 6785 3533
rect 6699 3479 6741 3513
rect 6775 3479 6785 3513
rect 6829 3505 6845 3539
rect 6879 3505 6971 3539
rect 7222 3529 7252 3582
rect 7339 3538 7369 3627
rect 7527 3597 7557 3677
rect 6829 3489 6971 3505
rect 7013 3503 7155 3519
rect 6699 3463 6785 3479
rect 7013 3469 7105 3503
rect 7139 3469 7155 3503
rect 6335 3441 6365 3463
rect 6523 3441 6553 3463
rect 6615 3441 6645 3463
rect 6699 3441 6729 3463
rect 7013 3453 7155 3469
rect 7198 3513 7252 3529
rect 7198 3479 7208 3513
rect 7242 3479 7252 3513
rect 7294 3528 7369 3538
rect 7462 3581 7557 3597
rect 7462 3547 7472 3581
rect 7506 3547 7557 3581
rect 7612 3561 7642 3677
rect 7707 3645 7737 3677
rect 7707 3629 7768 3645
rect 7707 3595 7724 3629
rect 7758 3595 7768 3629
rect 7707 3579 7768 3595
rect 7462 3531 7557 3547
rect 7294 3494 7310 3528
rect 7344 3494 7369 3528
rect 7294 3484 7369 3494
rect 7198 3463 7252 3479
rect 7013 3447 7097 3453
rect 6887 3421 7097 3447
rect 7222 3440 7252 3463
rect 7222 3410 7285 3440
rect 7255 3395 7285 3410
rect 7339 3395 7369 3484
rect 7527 3395 7557 3531
rect 7599 3551 7665 3561
rect 7599 3517 7615 3551
rect 7649 3537 7665 3551
rect 7649 3517 7768 3537
rect 7599 3507 7768 3517
rect 7619 3455 7685 3465
rect 7619 3421 7635 3455
rect 7669 3421 7685 3455
rect 7619 3411 7685 3421
rect 7639 3383 7669 3411
rect 7738 3383 7768 3507
rect 7810 3477 7840 3677
rect 7942 3573 7972 3611
rect 8037 3579 8067 3677
rect 8121 3639 8151 3677
rect 8235 3645 8265 3677
rect 8120 3629 8186 3639
rect 8120 3595 8136 3629
rect 8170 3595 8186 3629
rect 8120 3585 8186 3595
rect 8235 3629 8316 3645
rect 8235 3595 8272 3629
rect 8306 3595 8316 3629
rect 8235 3579 8316 3595
rect 7882 3563 7972 3573
rect 7882 3529 7898 3563
rect 7932 3529 7972 3563
rect 7882 3519 7972 3529
rect 7942 3484 7972 3519
rect 8024 3563 8078 3579
rect 8024 3529 8034 3563
rect 8068 3543 8078 3563
rect 8068 3529 8193 3543
rect 8024 3513 8193 3529
rect 7810 3467 7884 3477
rect 7810 3433 7834 3467
rect 7868 3433 7884 3467
rect 7942 3454 7986 3484
rect 7956 3439 7986 3454
rect 8057 3455 8121 3471
rect 7810 3423 7884 3433
rect 7837 3395 7867 3423
rect 8057 3421 8077 3455
rect 8111 3421 8121 3455
rect 8057 3405 8121 3421
rect 8057 3383 8087 3405
rect 8163 3383 8193 3513
rect 8258 3395 8288 3579
rect 9831 3755 9861 3781
rect 9915 3755 9945 3781
rect 10103 3761 10133 3787
rect 10188 3761 10218 3787
rect 10283 3761 10313 3787
rect 10386 3761 10416 3787
rect 10518 3761 10548 3787
rect 10613 3761 10643 3787
rect 10697 3761 10727 3787
rect 10811 3761 10841 3787
rect 11021 3761 11051 3787
rect 11105 3761 11135 3787
rect 11303 3761 11697 3787
rect 9831 3612 9861 3627
rect 9003 3561 9581 3587
rect 9798 3582 9861 3612
rect 8445 3529 8475 3561
rect 8529 3529 8559 3561
rect 9003 3539 9267 3561
rect 8335 3513 8477 3529
rect 8335 3479 8345 3513
rect 8379 3479 8477 3513
rect 8335 3463 8477 3479
rect 8519 3513 8573 3529
rect 8519 3479 8529 3513
rect 8563 3479 8573 3513
rect 9003 3505 9019 3539
rect 9053 3505 9118 3539
rect 9152 3505 9217 3539
rect 9251 3505 9267 3539
rect 9798 3529 9828 3582
rect 9915 3538 9945 3627
rect 10103 3597 10133 3677
rect 9003 3489 9267 3505
rect 9309 3503 9581 3519
rect 8519 3463 8573 3479
rect 9309 3469 9325 3503
rect 9359 3469 9428 3503
rect 9462 3469 9531 3503
rect 9565 3469 9581 3503
rect 8447 3441 8477 3463
rect 8531 3441 8561 3463
rect 9309 3447 9581 3469
rect 9774 3513 9828 3529
rect 9774 3479 9784 3513
rect 9818 3479 9828 3513
rect 9870 3528 9945 3538
rect 10038 3581 10133 3597
rect 10038 3547 10048 3581
rect 10082 3547 10133 3581
rect 10188 3561 10218 3677
rect 10283 3645 10313 3677
rect 10283 3629 10344 3645
rect 10283 3595 10300 3629
rect 10334 3595 10344 3629
rect 10283 3579 10344 3595
rect 10038 3531 10133 3547
rect 9870 3494 9886 3528
rect 9920 3494 9945 3528
rect 9870 3484 9945 3494
rect 9774 3463 9828 3479
rect 9003 3421 9581 3447
rect 9798 3440 9828 3463
rect 9798 3410 9861 3440
rect 9831 3395 9861 3410
rect 9915 3395 9945 3484
rect 10103 3395 10133 3531
rect 10175 3551 10241 3561
rect 10175 3517 10191 3551
rect 10225 3537 10241 3551
rect 10225 3517 10344 3537
rect 10175 3507 10344 3517
rect 10195 3455 10261 3465
rect 10195 3421 10211 3455
rect 10245 3421 10261 3455
rect 10195 3411 10261 3421
rect 10215 3383 10245 3411
rect 10314 3383 10344 3507
rect 10386 3477 10416 3677
rect 10518 3573 10548 3611
rect 10613 3579 10643 3677
rect 10697 3639 10727 3677
rect 10811 3645 10841 3677
rect 10696 3629 10762 3639
rect 10696 3595 10712 3629
rect 10746 3595 10762 3629
rect 10696 3585 10762 3595
rect 10811 3629 10892 3645
rect 10811 3595 10848 3629
rect 10882 3595 10892 3629
rect 10811 3579 10892 3595
rect 10458 3563 10548 3573
rect 10458 3529 10474 3563
rect 10508 3529 10548 3563
rect 10458 3519 10548 3529
rect 10518 3484 10548 3519
rect 10600 3563 10654 3579
rect 10600 3529 10610 3563
rect 10644 3543 10654 3563
rect 10644 3529 10769 3543
rect 10600 3513 10769 3529
rect 10386 3467 10460 3477
rect 10386 3433 10410 3467
rect 10444 3433 10460 3467
rect 10518 3454 10562 3484
rect 10532 3439 10562 3454
rect 10633 3455 10697 3471
rect 10386 3423 10460 3433
rect 10413 3395 10443 3423
rect 10633 3421 10653 3455
rect 10687 3421 10697 3455
rect 10633 3405 10697 3421
rect 10633 3383 10663 3405
rect 10739 3383 10769 3513
rect 10834 3395 10864 3579
rect 11855 3755 11885 3781
rect 11939 3755 11969 3781
rect 12127 3761 12157 3787
rect 12212 3761 12242 3787
rect 12307 3761 12337 3787
rect 12410 3761 12440 3787
rect 12542 3761 12572 3787
rect 12637 3761 12667 3787
rect 12721 3761 12751 3787
rect 12835 3761 12865 3787
rect 13045 3761 13075 3787
rect 13129 3761 13159 3787
rect 13327 3761 13905 3787
rect 14155 3761 15101 3787
rect 15259 3761 15653 3787
rect 15811 3761 15841 3787
rect 15899 3761 15929 3787
rect 16087 3761 16297 3787
rect 16499 3761 16529 3787
rect 16915 3761 17125 3787
rect 17327 3761 17357 3787
rect 17743 3761 18321 3787
rect 18663 3761 18781 3787
rect 11855 3612 11885 3627
rect 11303 3561 11697 3587
rect 11822 3582 11885 3612
rect 11021 3529 11051 3561
rect 11105 3529 11135 3561
rect 11303 3539 11479 3561
rect 10911 3513 11053 3529
rect 10911 3479 10921 3513
rect 10955 3479 11053 3513
rect 10911 3463 11053 3479
rect 11095 3513 11149 3529
rect 11095 3479 11105 3513
rect 11139 3479 11149 3513
rect 11303 3505 11319 3539
rect 11353 3505 11429 3539
rect 11463 3505 11479 3539
rect 11822 3529 11852 3582
rect 11939 3538 11969 3627
rect 12127 3597 12157 3677
rect 11303 3489 11479 3505
rect 11521 3503 11697 3519
rect 11095 3463 11149 3479
rect 11521 3469 11537 3503
rect 11571 3469 11647 3503
rect 11681 3469 11697 3503
rect 11023 3441 11053 3463
rect 11107 3441 11137 3463
rect 11521 3447 11697 3469
rect 11798 3513 11852 3529
rect 11798 3479 11808 3513
rect 11842 3479 11852 3513
rect 11894 3528 11969 3538
rect 12062 3581 12157 3597
rect 12062 3547 12072 3581
rect 12106 3547 12157 3581
rect 12212 3561 12242 3677
rect 12307 3645 12337 3677
rect 12307 3629 12368 3645
rect 12307 3595 12324 3629
rect 12358 3595 12368 3629
rect 12307 3579 12368 3595
rect 12062 3531 12157 3547
rect 11894 3494 11910 3528
rect 11944 3494 11969 3528
rect 11894 3484 11969 3494
rect 11798 3463 11852 3479
rect 11303 3421 11697 3447
rect 11822 3440 11852 3463
rect 11822 3410 11885 3440
rect 11855 3395 11885 3410
rect 11939 3395 11969 3484
rect 12127 3395 12157 3531
rect 12199 3551 12265 3561
rect 12199 3517 12215 3551
rect 12249 3537 12265 3551
rect 12249 3517 12368 3537
rect 12199 3507 12368 3517
rect 12219 3455 12285 3465
rect 12219 3421 12235 3455
rect 12269 3421 12285 3455
rect 12219 3411 12285 3421
rect 12239 3383 12269 3411
rect 12338 3383 12368 3507
rect 12410 3477 12440 3677
rect 12542 3573 12572 3611
rect 12637 3579 12667 3677
rect 12721 3639 12751 3677
rect 12835 3645 12865 3677
rect 12720 3629 12786 3639
rect 12720 3595 12736 3629
rect 12770 3595 12786 3629
rect 12720 3585 12786 3595
rect 12835 3629 12916 3645
rect 12835 3595 12872 3629
rect 12906 3595 12916 3629
rect 12835 3579 12916 3595
rect 12482 3563 12572 3573
rect 12482 3529 12498 3563
rect 12532 3529 12572 3563
rect 12482 3519 12572 3529
rect 12542 3484 12572 3519
rect 12624 3563 12678 3579
rect 12624 3529 12634 3563
rect 12668 3543 12678 3563
rect 12668 3529 12793 3543
rect 12624 3513 12793 3529
rect 12410 3467 12484 3477
rect 12410 3433 12434 3467
rect 12468 3433 12484 3467
rect 12542 3454 12586 3484
rect 12556 3439 12586 3454
rect 12657 3455 12721 3471
rect 12410 3423 12484 3433
rect 12437 3395 12467 3423
rect 12657 3421 12677 3455
rect 12711 3421 12721 3455
rect 12657 3405 12721 3421
rect 12657 3383 12687 3405
rect 12763 3383 12793 3513
rect 12858 3395 12888 3579
rect 13327 3561 13905 3587
rect 14155 3561 15101 3587
rect 15259 3561 15653 3587
rect 13045 3529 13075 3561
rect 13129 3529 13159 3561
rect 13327 3539 13591 3561
rect 12935 3513 13077 3529
rect 12935 3479 12945 3513
rect 12979 3479 13077 3513
rect 12935 3463 13077 3479
rect 13119 3513 13173 3529
rect 13119 3479 13129 3513
rect 13163 3479 13173 3513
rect 13327 3505 13343 3539
rect 13377 3505 13442 3539
rect 13476 3505 13541 3539
rect 13575 3505 13591 3539
rect 14155 3539 14605 3561
rect 13327 3489 13591 3505
rect 13633 3503 13905 3519
rect 13119 3463 13173 3479
rect 13633 3469 13649 3503
rect 13683 3469 13752 3503
rect 13786 3469 13855 3503
rect 13889 3469 13905 3503
rect 14155 3505 14427 3539
rect 14461 3505 14605 3539
rect 15259 3539 15435 3561
rect 15811 3542 15841 3603
rect 15899 3588 15929 3603
rect 15899 3564 15935 3588
rect 14155 3489 14605 3505
rect 14647 3503 15101 3519
rect 13047 3441 13077 3463
rect 13131 3441 13161 3463
rect 13633 3447 13905 3469
rect 14647 3469 14791 3503
rect 14825 3469 15101 3503
rect 15259 3505 15275 3539
rect 15309 3505 15385 3539
rect 15419 3505 15435 3539
rect 15807 3526 15861 3542
rect 15259 3489 15435 3505
rect 15477 3503 15653 3519
rect 14647 3447 15101 3469
rect 15477 3469 15493 3503
rect 15527 3469 15603 3503
rect 15637 3469 15653 3503
rect 15807 3492 15817 3526
rect 15851 3492 15861 3526
rect 15807 3476 15861 3492
rect 15905 3529 15935 3564
rect 16087 3561 16297 3587
rect 16607 3719 16637 3745
rect 16691 3719 16721 3745
rect 16087 3555 16171 3561
rect 16029 3539 16171 3555
rect 15905 3513 15981 3529
rect 15905 3479 15937 3513
rect 15971 3479 15981 3513
rect 16029 3505 16045 3539
rect 16079 3505 16171 3539
rect 16499 3529 16529 3561
rect 16607 3529 16637 3635
rect 16029 3489 16171 3505
rect 16213 3503 16355 3519
rect 15477 3447 15653 3469
rect 13327 3421 13905 3447
rect 14155 3421 15101 3447
rect 15259 3421 15653 3447
rect 15811 3415 15841 3476
rect 15905 3463 15981 3479
rect 16213 3469 16305 3503
rect 16339 3469 16355 3503
rect 15905 3454 15935 3463
rect 15899 3430 15935 3454
rect 16213 3453 16355 3469
rect 16463 3513 16529 3529
rect 16463 3479 16479 3513
rect 16513 3479 16529 3513
rect 16463 3463 16529 3479
rect 16571 3513 16637 3529
rect 16571 3479 16587 3513
rect 16621 3479 16637 3513
rect 16571 3463 16637 3479
rect 16213 3447 16297 3453
rect 15899 3415 15929 3430
rect 16087 3421 16297 3447
rect 16499 3441 16529 3463
rect 16607 3423 16637 3463
rect 16691 3529 16721 3635
rect 16915 3561 17125 3587
rect 17435 3719 17465 3745
rect 17519 3719 17549 3745
rect 16915 3555 16999 3561
rect 16857 3539 16999 3555
rect 16691 3513 16778 3529
rect 16691 3479 16728 3513
rect 16762 3479 16778 3513
rect 16857 3505 16873 3539
rect 16907 3505 16999 3539
rect 17327 3529 17357 3561
rect 17435 3529 17465 3635
rect 16857 3489 16999 3505
rect 17041 3503 17183 3519
rect 16691 3463 16778 3479
rect 17041 3469 17133 3503
rect 17167 3469 17183 3503
rect 16691 3423 16721 3463
rect 17041 3453 17183 3469
rect 17291 3513 17357 3529
rect 17291 3479 17307 3513
rect 17341 3479 17357 3513
rect 17291 3463 17357 3479
rect 17399 3513 17465 3529
rect 17399 3479 17415 3513
rect 17449 3479 17465 3513
rect 17399 3463 17465 3479
rect 17041 3447 17125 3453
rect 16915 3421 17125 3447
rect 17327 3441 17357 3463
rect 16607 3313 16637 3339
rect 16691 3313 16721 3339
rect 17435 3423 17465 3463
rect 17519 3529 17549 3635
rect 17743 3561 18321 3587
rect 17743 3539 18007 3561
rect 18663 3557 18781 3587
rect 17519 3513 17606 3529
rect 17519 3479 17556 3513
rect 17590 3479 17606 3513
rect 17743 3505 17759 3539
rect 17793 3505 17858 3539
rect 17892 3505 17957 3539
rect 17991 3505 18007 3539
rect 18743 3555 18781 3557
rect 18743 3539 18809 3555
rect 17743 3489 18007 3505
rect 18049 3503 18321 3519
rect 17519 3463 17606 3479
rect 18049 3469 18065 3503
rect 18099 3469 18168 3503
rect 18202 3469 18271 3503
rect 18305 3469 18321 3503
rect 17519 3423 17549 3463
rect 18049 3447 18321 3469
rect 18635 3499 18701 3515
rect 18635 3465 18651 3499
rect 18685 3465 18701 3499
rect 18743 3505 18759 3539
rect 18793 3505 18809 3539
rect 18743 3489 18809 3505
rect 18635 3449 18701 3465
rect 17743 3421 18321 3447
rect 18663 3447 18701 3449
rect 18663 3421 18781 3447
rect 17435 3313 17465 3339
rect 17519 3313 17549 3339
rect 1183 3285 1301 3311
rect 1459 3285 1853 3311
rect 2103 3285 2133 3311
rect 2187 3285 2217 3311
rect 2375 3285 2405 3311
rect 2487 3285 2517 3311
rect 2586 3285 2616 3311
rect 2685 3285 2715 3311
rect 2804 3285 2834 3311
rect 2905 3285 2935 3311
rect 3011 3285 3041 3311
rect 3106 3285 3136 3311
rect 3295 3285 3325 3311
rect 3379 3285 3409 3311
rect 4035 3285 4065 3311
rect 4119 3285 4149 3311
rect 4307 3285 4337 3311
rect 4419 3285 4449 3311
rect 4518 3285 4548 3311
rect 4617 3285 4647 3311
rect 4736 3285 4766 3311
rect 4837 3285 4867 3311
rect 4943 3285 4973 3311
rect 5038 3285 5068 3311
rect 5227 3285 5257 3311
rect 5311 3285 5341 3311
rect 5507 3285 6085 3311
rect 6335 3285 6365 3311
rect 6523 3285 6553 3311
rect 6615 3285 6645 3311
rect 6699 3285 6729 3311
rect 6887 3285 7097 3311
rect 7255 3285 7285 3311
rect 7339 3285 7369 3311
rect 7527 3285 7557 3311
rect 7639 3285 7669 3311
rect 7738 3285 7768 3311
rect 7837 3285 7867 3311
rect 7956 3285 7986 3311
rect 8057 3285 8087 3311
rect 8163 3285 8193 3311
rect 8258 3285 8288 3311
rect 8447 3285 8477 3311
rect 8531 3285 8561 3311
rect 9003 3285 9581 3311
rect 9831 3285 9861 3311
rect 9915 3285 9945 3311
rect 10103 3285 10133 3311
rect 10215 3285 10245 3311
rect 10314 3285 10344 3311
rect 10413 3285 10443 3311
rect 10532 3285 10562 3311
rect 10633 3285 10663 3311
rect 10739 3285 10769 3311
rect 10834 3285 10864 3311
rect 11023 3285 11053 3311
rect 11107 3285 11137 3311
rect 11303 3285 11697 3311
rect 11855 3285 11885 3311
rect 11939 3285 11969 3311
rect 12127 3285 12157 3311
rect 12239 3285 12269 3311
rect 12338 3285 12368 3311
rect 12437 3285 12467 3311
rect 12556 3285 12586 3311
rect 12657 3285 12687 3311
rect 12763 3285 12793 3311
rect 12858 3285 12888 3311
rect 13047 3285 13077 3311
rect 13131 3285 13161 3311
rect 13327 3285 13905 3311
rect 14155 3285 15101 3311
rect 15259 3285 15653 3311
rect 15811 3285 15841 3311
rect 15899 3285 15929 3311
rect 16087 3285 16297 3311
rect 16499 3285 16529 3311
rect 16915 3285 17125 3311
rect 17327 3285 17357 3311
rect 17743 3285 18321 3311
rect 18663 3285 18781 3311
rect 1183 3217 1301 3243
rect 1459 3217 1669 3243
rect 1920 3217 1950 3243
rect 2015 3217 2045 3243
rect 2099 3217 2129 3243
rect 2287 3217 2497 3243
rect 2673 3217 2703 3243
rect 2759 3217 2789 3243
rect 2845 3217 2875 3243
rect 2931 3217 2961 3243
rect 3017 3217 3047 3243
rect 3103 3217 3133 3243
rect 3189 3217 3219 3243
rect 3275 3217 3305 3243
rect 3360 3217 3390 3243
rect 3446 3217 3476 3243
rect 3532 3217 3562 3243
rect 3618 3217 3648 3243
rect 3704 3217 3734 3243
rect 3790 3217 3820 3243
rect 3876 3217 3906 3243
rect 3962 3217 3992 3243
rect 4048 3217 4078 3243
rect 4134 3217 4164 3243
rect 4220 3217 4250 3243
rect 4306 3217 4336 3243
rect 4495 3217 5441 3243
rect 5599 3217 6177 3243
rect 6427 3217 7005 3243
rect 1183 3081 1301 3107
rect 1459 3081 1669 3107
rect 1263 3079 1301 3081
rect 1263 3063 1329 3079
rect 1155 3023 1221 3039
rect 1155 2989 1171 3023
rect 1205 2989 1221 3023
rect 1263 3029 1279 3063
rect 1313 3029 1329 3063
rect 1585 3075 1669 3081
rect 1920 3084 1950 3133
rect 2015 3115 2045 3133
rect 2099 3115 2129 3133
rect 1585 3059 1727 3075
rect 1920 3069 1973 3084
rect 1263 3013 1329 3029
rect 1401 3023 1543 3039
rect 1155 2973 1221 2989
rect 1401 2989 1417 3023
rect 1451 2989 1543 3023
rect 1585 3025 1677 3059
rect 1711 3025 1727 3059
rect 1585 3009 1727 3025
rect 1909 3049 1973 3069
rect 1909 3015 1929 3049
rect 1963 3015 1973 3049
rect 1401 2973 1543 2989
rect 1909 2985 1973 3015
rect 2015 3049 2129 3115
rect 2287 3081 2497 3107
rect 2015 3015 2033 3049
rect 2067 3015 2129 3049
rect 2413 3075 2497 3081
rect 2413 3059 2555 3075
rect 2015 2985 2129 3015
rect 1183 2971 1221 2973
rect 1183 2941 1301 2971
rect 1459 2967 1543 2973
rect 1920 2967 1950 2985
rect 2015 2967 2045 2985
rect 2099 2967 2129 2985
rect 2229 3023 2371 3039
rect 2229 2989 2245 3023
rect 2279 2989 2371 3023
rect 2413 3025 2505 3059
rect 2539 3025 2555 3059
rect 2413 3009 2555 3025
rect 2673 3074 2703 3133
rect 2759 3074 2789 3133
rect 2845 3074 2875 3133
rect 2931 3074 2961 3133
rect 3017 3074 3047 3133
rect 3103 3074 3133 3133
rect 3189 3074 3219 3133
rect 3275 3074 3305 3133
rect 3360 3074 3390 3133
rect 3446 3074 3476 3133
rect 3532 3074 3562 3133
rect 3618 3074 3648 3133
rect 3704 3074 3734 3133
rect 3790 3074 3820 3133
rect 3876 3074 3906 3133
rect 3962 3074 3992 3133
rect 2673 3049 3992 3074
rect 2673 3015 2898 3049
rect 2932 3015 2966 3049
rect 3000 3015 3034 3049
rect 3068 3015 3102 3049
rect 3136 3015 3170 3049
rect 3204 3015 3238 3049
rect 3272 3015 3306 3049
rect 3340 3015 3374 3049
rect 3408 3015 3442 3049
rect 3476 3015 3510 3049
rect 3544 3015 3578 3049
rect 3612 3015 3646 3049
rect 3680 3015 3714 3049
rect 3748 3015 3782 3049
rect 3816 3015 3850 3049
rect 3884 3015 3918 3049
rect 3952 3015 3992 3049
rect 2229 2973 2371 2989
rect 2287 2967 2371 2973
rect 2673 2999 3992 3015
rect 2673 2967 2703 2999
rect 2759 2967 2789 2999
rect 2845 2967 2875 2999
rect 2931 2967 2961 2999
rect 3017 2967 3047 2999
rect 3103 2967 3133 2999
rect 3189 2967 3219 2999
rect 3275 2967 3305 2999
rect 3360 2967 3390 2999
rect 3446 2967 3476 2999
rect 3532 2967 3562 2999
rect 3618 2967 3648 2999
rect 3704 2967 3734 2999
rect 3790 2967 3820 2999
rect 3876 2967 3906 2999
rect 3962 2967 3992 2999
rect 4048 3084 4078 3133
rect 4134 3084 4164 3133
rect 4220 3084 4250 3133
rect 4306 3084 4336 3133
rect 4048 3049 4395 3084
rect 4495 3081 5441 3107
rect 5599 3081 6177 3107
rect 7439 3217 7649 3243
rect 7808 3217 7838 3243
rect 7894 3217 7924 3243
rect 7980 3217 8010 3243
rect 8066 3217 8096 3243
rect 8152 3217 8182 3243
rect 8238 3217 8268 3243
rect 8324 3217 8354 3243
rect 8410 3217 8440 3243
rect 8496 3217 8526 3243
rect 8582 3217 8612 3243
rect 8668 3217 8698 3243
rect 8754 3217 8784 3243
rect 8839 3217 8869 3243
rect 8925 3217 8955 3243
rect 9011 3217 9041 3243
rect 9097 3217 9127 3243
rect 9183 3217 9213 3243
rect 9269 3217 9299 3243
rect 9355 3217 9385 3243
rect 9441 3217 9471 3243
rect 9647 3217 10593 3243
rect 10751 3217 11329 3243
rect 11763 3217 11793 3243
rect 11847 3217 11877 3243
rect 12035 3217 12065 3243
rect 12147 3217 12177 3243
rect 12246 3217 12276 3243
rect 12345 3217 12375 3243
rect 12464 3217 12494 3243
rect 12565 3217 12595 3243
rect 12671 3217 12701 3243
rect 12766 3217 12796 3243
rect 12955 3217 12985 3243
rect 13039 3217 13069 3243
rect 13235 3217 14181 3243
rect 14339 3217 15285 3243
rect 15443 3217 16389 3243
rect 16915 3217 16945 3243
rect 17003 3217 17033 3243
rect 17191 3217 18137 3243
rect 18295 3217 18505 3243
rect 18663 3217 18781 3243
rect 6427 3081 7005 3107
rect 7439 3081 7649 3107
rect 7808 3084 7838 3133
rect 7894 3084 7924 3133
rect 7980 3084 8010 3133
rect 8066 3084 8096 3133
rect 4048 3015 4345 3049
rect 4379 3015 4395 3049
rect 4987 3059 5441 3081
rect 4048 2982 4395 3015
rect 4495 3023 4945 3039
rect 4495 2989 4767 3023
rect 4801 2989 4945 3023
rect 4987 3025 5131 3059
rect 5165 3025 5441 3059
rect 5905 3059 6177 3081
rect 4987 3009 5441 3025
rect 5599 3023 5863 3039
rect 4048 2967 4078 2982
rect 4134 2967 4164 2982
rect 4220 2967 4250 2982
rect 4306 2967 4336 2982
rect 4495 2967 4945 2989
rect 5599 2989 5615 3023
rect 5649 2989 5714 3023
rect 5748 2989 5813 3023
rect 5847 2989 5863 3023
rect 5905 3025 5921 3059
rect 5955 3025 6024 3059
rect 6058 3025 6127 3059
rect 6161 3025 6177 3059
rect 6733 3059 7005 3081
rect 5905 3009 6177 3025
rect 6427 3023 6691 3039
rect 5599 2967 5863 2989
rect 6427 2989 6443 3023
rect 6477 2989 6542 3023
rect 6576 2989 6641 3023
rect 6675 2989 6691 3023
rect 6733 3025 6749 3059
rect 6783 3025 6852 3059
rect 6886 3025 6955 3059
rect 6989 3025 7005 3059
rect 7565 3075 7649 3081
rect 7565 3059 7707 3075
rect 6733 3009 7005 3025
rect 7381 3023 7523 3039
rect 6427 2967 6691 2989
rect 7381 2989 7397 3023
rect 7431 2989 7523 3023
rect 7565 3025 7657 3059
rect 7691 3025 7707 3059
rect 7565 3009 7707 3025
rect 7749 3049 8096 3084
rect 7749 3015 7765 3049
rect 7799 3015 8096 3049
rect 7381 2973 7523 2989
rect 7749 2982 8096 3015
rect 7439 2967 7523 2973
rect 7808 2967 7838 2982
rect 7894 2967 7924 2982
rect 7980 2967 8010 2982
rect 8066 2967 8096 2982
rect 8152 3074 8182 3133
rect 8238 3074 8268 3133
rect 8324 3074 8354 3133
rect 8410 3074 8440 3133
rect 8496 3074 8526 3133
rect 8582 3074 8612 3133
rect 8668 3074 8698 3133
rect 8754 3074 8784 3133
rect 8839 3074 8869 3133
rect 8925 3074 8955 3133
rect 9011 3074 9041 3133
rect 9097 3074 9127 3133
rect 9183 3074 9213 3133
rect 9269 3074 9299 3133
rect 9355 3074 9385 3133
rect 9441 3074 9471 3133
rect 9647 3081 10593 3107
rect 10751 3081 11329 3107
rect 11763 3118 11793 3133
rect 8152 3049 9471 3074
rect 8152 3015 8192 3049
rect 8226 3015 8260 3049
rect 8294 3015 8328 3049
rect 8362 3015 8396 3049
rect 8430 3015 8464 3049
rect 8498 3015 8532 3049
rect 8566 3015 8600 3049
rect 8634 3015 8668 3049
rect 8702 3015 8736 3049
rect 8770 3015 8804 3049
rect 8838 3015 8872 3049
rect 8906 3015 8940 3049
rect 8974 3015 9008 3049
rect 9042 3015 9076 3049
rect 9110 3015 9144 3049
rect 9178 3015 9212 3049
rect 9246 3015 9471 3049
rect 10139 3059 10593 3081
rect 8152 2999 9471 3015
rect 8152 2967 8182 2999
rect 8238 2967 8268 2999
rect 8324 2967 8354 2999
rect 8410 2967 8440 2999
rect 8496 2967 8526 2999
rect 8582 2967 8612 2999
rect 8668 2967 8698 2999
rect 8754 2967 8784 2999
rect 8839 2967 8869 2999
rect 8925 2967 8955 2999
rect 9011 2967 9041 2999
rect 9097 2967 9127 2999
rect 9183 2967 9213 2999
rect 9269 2967 9299 2999
rect 9355 2967 9385 2999
rect 9441 2967 9471 2999
rect 9647 3023 10097 3039
rect 9647 2989 9919 3023
rect 9953 2989 10097 3023
rect 10139 3025 10283 3059
rect 10317 3025 10593 3059
rect 11057 3059 11329 3081
rect 11730 3088 11793 3118
rect 11730 3065 11760 3088
rect 10139 3009 10593 3025
rect 10751 3023 11015 3039
rect 9647 2967 10097 2989
rect 10751 2989 10767 3023
rect 10801 2989 10866 3023
rect 10900 2989 10965 3023
rect 10999 2989 11015 3023
rect 11057 3025 11073 3059
rect 11107 3025 11176 3059
rect 11210 3025 11279 3059
rect 11313 3025 11329 3059
rect 11057 3009 11329 3025
rect 11706 3049 11760 3065
rect 11706 3015 11716 3049
rect 11750 3015 11760 3049
rect 11847 3044 11877 3133
rect 11706 2999 11760 3015
rect 10751 2967 11015 2989
rect 1459 2941 1669 2967
rect 2287 2941 2497 2967
rect 4495 2941 5441 2967
rect 5599 2941 6177 2967
rect 6427 2941 7005 2967
rect 7439 2941 7649 2967
rect 9647 2941 10593 2967
rect 10751 2941 11329 2967
rect 11730 2946 11760 2999
rect 11802 3034 11877 3044
rect 11802 3000 11818 3034
rect 11852 3000 11877 3034
rect 11802 2990 11877 3000
rect 12035 2997 12065 3133
rect 12147 3117 12177 3145
rect 12127 3107 12193 3117
rect 12127 3073 12143 3107
rect 12177 3073 12193 3107
rect 12127 3063 12193 3073
rect 12246 3021 12276 3145
rect 12345 3105 12375 3133
rect 11730 2916 11793 2946
rect 11763 2901 11793 2916
rect 11847 2901 11877 2990
rect 11970 2981 12065 2997
rect 11970 2947 11980 2981
rect 12014 2947 12065 2981
rect 12107 3011 12276 3021
rect 12107 2977 12123 3011
rect 12157 2991 12276 3011
rect 12318 3095 12392 3105
rect 12318 3061 12342 3095
rect 12376 3061 12392 3095
rect 12565 3123 12595 3145
rect 12565 3107 12629 3123
rect 12464 3074 12494 3089
rect 12318 3051 12392 3061
rect 12157 2977 12173 2991
rect 12107 2967 12173 2977
rect 11970 2931 12065 2947
rect 12035 2851 12065 2931
rect 12120 2851 12150 2967
rect 12215 2933 12276 2949
rect 12215 2899 12232 2933
rect 12266 2899 12276 2933
rect 12215 2883 12276 2899
rect 12215 2851 12245 2883
rect 12318 2851 12348 3051
rect 12450 3044 12494 3074
rect 12565 3073 12585 3107
rect 12619 3073 12629 3107
rect 12565 3057 12629 3073
rect 12450 3009 12480 3044
rect 12671 3015 12701 3145
rect 12390 2999 12480 3009
rect 12390 2965 12406 2999
rect 12440 2965 12480 2999
rect 12390 2955 12480 2965
rect 12450 2917 12480 2955
rect 12532 2999 12701 3015
rect 12532 2965 12542 2999
rect 12576 2985 12701 2999
rect 12576 2965 12586 2985
rect 12532 2949 12586 2965
rect 12766 2949 12796 3133
rect 12955 3065 12985 3087
rect 13039 3065 13069 3087
rect 13235 3081 14181 3107
rect 14339 3081 15285 3107
rect 15443 3081 16389 3107
rect 12843 3049 12985 3065
rect 12843 3015 12853 3049
rect 12887 3015 12985 3049
rect 12843 2999 12985 3015
rect 13027 3049 13081 3065
rect 13027 3015 13037 3049
rect 13071 3015 13081 3049
rect 13727 3059 14181 3081
rect 13027 2999 13081 3015
rect 13235 3023 13685 3039
rect 12953 2967 12983 2999
rect 13037 2967 13067 2999
rect 13235 2989 13507 3023
rect 13541 2989 13685 3023
rect 13727 3025 13871 3059
rect 13905 3025 14181 3059
rect 14831 3059 15285 3081
rect 13727 3009 14181 3025
rect 14339 3023 14789 3039
rect 13235 2967 13685 2989
rect 14339 2989 14611 3023
rect 14645 2989 14789 3023
rect 14831 3025 14975 3059
rect 15009 3025 15285 3059
rect 15935 3059 16389 3081
rect 14831 3009 15285 3025
rect 15443 3023 15893 3039
rect 14339 2967 14789 2989
rect 15443 2989 15715 3023
rect 15749 2989 15893 3023
rect 15935 3025 16079 3059
rect 16113 3025 16389 3059
rect 16915 3052 16945 3113
rect 17003 3098 17033 3113
rect 17003 3074 17039 3098
rect 17191 3081 18137 3107
rect 18295 3081 18505 3107
rect 17009 3065 17039 3074
rect 15935 3009 16389 3025
rect 16911 3036 16965 3052
rect 15443 2967 15893 2989
rect 16911 3002 16921 3036
rect 16955 3002 16965 3036
rect 16911 2986 16965 3002
rect 17009 3049 17085 3065
rect 17009 3015 17041 3049
rect 17075 3015 17085 3049
rect 17683 3059 18137 3081
rect 17009 2999 17085 3015
rect 17191 3023 17641 3039
rect 1183 2741 1301 2767
rect 1459 2741 1669 2767
rect 1920 2741 1950 2767
rect 2015 2741 2045 2767
rect 2099 2741 2129 2767
rect 2287 2741 2497 2767
rect 2673 2741 2703 2767
rect 2759 2741 2789 2767
rect 2845 2741 2875 2767
rect 2931 2741 2961 2767
rect 3017 2741 3047 2767
rect 3103 2741 3133 2767
rect 3189 2741 3219 2767
rect 3275 2741 3305 2767
rect 3360 2741 3390 2767
rect 3446 2741 3476 2767
rect 3532 2741 3562 2767
rect 3618 2741 3648 2767
rect 3704 2741 3734 2767
rect 3790 2741 3820 2767
rect 3876 2741 3906 2767
rect 3962 2741 3992 2767
rect 4048 2741 4078 2767
rect 4134 2741 4164 2767
rect 4220 2741 4250 2767
rect 4306 2741 4336 2767
rect 4495 2741 5441 2767
rect 5599 2741 6177 2767
rect 6427 2741 7005 2767
rect 7439 2741 7649 2767
rect 7808 2741 7838 2767
rect 7894 2741 7924 2767
rect 7980 2741 8010 2767
rect 8066 2741 8096 2767
rect 8152 2741 8182 2767
rect 8238 2741 8268 2767
rect 8324 2741 8354 2767
rect 8410 2741 8440 2767
rect 8496 2741 8526 2767
rect 8582 2741 8612 2767
rect 8668 2741 8698 2767
rect 8754 2741 8784 2767
rect 8839 2741 8869 2767
rect 8925 2741 8955 2767
rect 9011 2741 9041 2767
rect 9097 2741 9127 2767
rect 9183 2741 9213 2767
rect 9269 2741 9299 2767
rect 9355 2741 9385 2767
rect 9441 2741 9471 2767
rect 9647 2741 10593 2767
rect 10751 2741 11329 2767
rect 11763 2747 11793 2773
rect 11847 2747 11877 2773
rect 12545 2851 12575 2949
rect 12628 2933 12694 2943
rect 12628 2899 12644 2933
rect 12678 2899 12694 2933
rect 12628 2889 12694 2899
rect 12743 2933 12824 2949
rect 12743 2899 12780 2933
rect 12814 2899 12824 2933
rect 12629 2851 12659 2889
rect 12743 2883 12824 2899
rect 12743 2851 12773 2883
rect 13235 2941 14181 2967
rect 14339 2941 15285 2967
rect 15443 2941 16389 2967
rect 16915 2925 16945 2986
rect 17009 2964 17039 2999
rect 17003 2940 17039 2964
rect 17191 2989 17463 3023
rect 17497 2989 17641 3023
rect 17683 3025 17827 3059
rect 17861 3025 18137 3059
rect 18421 3075 18505 3081
rect 18663 3081 18781 3107
rect 18663 3079 18701 3081
rect 18421 3059 18563 3075
rect 17683 3009 18137 3025
rect 18237 3023 18379 3039
rect 17191 2967 17641 2989
rect 18237 2989 18253 3023
rect 18287 2989 18379 3023
rect 18421 3025 18513 3059
rect 18547 3025 18563 3059
rect 18421 3009 18563 3025
rect 18635 3063 18701 3079
rect 18635 3029 18651 3063
rect 18685 3029 18701 3063
rect 18635 3013 18701 3029
rect 18743 3023 18809 3039
rect 18237 2973 18379 2989
rect 18295 2967 18379 2973
rect 18743 2989 18759 3023
rect 18793 2989 18809 3023
rect 18743 2973 18809 2989
rect 18743 2971 18781 2973
rect 17191 2941 18137 2967
rect 18295 2941 18505 2967
rect 18663 2941 18781 2971
rect 17003 2925 17033 2940
rect 12035 2741 12065 2767
rect 12120 2741 12150 2767
rect 12215 2741 12245 2767
rect 12318 2741 12348 2767
rect 12450 2741 12480 2767
rect 12545 2741 12575 2767
rect 12629 2741 12659 2767
rect 12743 2741 12773 2767
rect 12953 2741 12983 2767
rect 13037 2741 13067 2767
rect 13235 2741 14181 2767
rect 14339 2741 15285 2767
rect 15443 2741 16389 2767
rect 16915 2741 16945 2767
rect 17003 2741 17033 2767
rect 17191 2741 18137 2767
rect 18295 2741 18505 2767
rect 18663 2741 18781 2767
rect 1183 2673 1301 2699
rect 1459 2673 1853 2699
rect 2113 2673 2143 2699
rect 2197 2673 2227 2699
rect 2407 2673 2437 2699
rect 2521 2673 2551 2699
rect 2605 2673 2635 2699
rect 2700 2673 2730 2699
rect 2832 2673 2862 2699
rect 2935 2673 2965 2699
rect 3030 2673 3060 2699
rect 3115 2673 3145 2699
rect 1183 2469 1301 2499
rect 1459 2473 1853 2499
rect 2407 2557 2437 2589
rect 2356 2541 2437 2557
rect 2521 2551 2551 2589
rect 2356 2507 2366 2541
rect 2400 2507 2437 2541
rect 2356 2491 2437 2507
rect 2486 2541 2552 2551
rect 2486 2507 2502 2541
rect 2536 2507 2552 2541
rect 2486 2497 2552 2507
rect 2605 2491 2635 2589
rect 3303 2667 3333 2693
rect 3387 2667 3417 2693
rect 4219 2673 4429 2699
rect 1183 2467 1221 2469
rect 1155 2451 1221 2467
rect 1155 2417 1171 2451
rect 1205 2417 1221 2451
rect 1459 2451 1635 2473
rect 1155 2401 1221 2417
rect 1263 2411 1329 2427
rect 1263 2377 1279 2411
rect 1313 2377 1329 2411
rect 1459 2417 1475 2451
rect 1509 2417 1585 2451
rect 1619 2417 1635 2451
rect 2113 2441 2143 2473
rect 2197 2441 2227 2473
rect 1459 2401 1635 2417
rect 1677 2415 1853 2431
rect 1263 2361 1329 2377
rect 1677 2381 1693 2415
rect 1727 2381 1803 2415
rect 1837 2381 1853 2415
rect 1263 2359 1301 2361
rect 1677 2359 1853 2381
rect 2099 2425 2153 2441
rect 2099 2391 2109 2425
rect 2143 2391 2153 2425
rect 2099 2375 2153 2391
rect 2195 2425 2337 2441
rect 2195 2391 2293 2425
rect 2327 2391 2337 2425
rect 2195 2375 2337 2391
rect 1183 2333 1301 2359
rect 1459 2333 1853 2359
rect 2111 2353 2141 2375
rect 2195 2353 2225 2375
rect 2384 2307 2414 2491
rect 2594 2475 2648 2491
rect 2594 2455 2604 2475
rect 2479 2441 2604 2455
rect 2638 2441 2648 2475
rect 2479 2425 2648 2441
rect 2700 2485 2730 2523
rect 2700 2475 2790 2485
rect 2700 2441 2740 2475
rect 2774 2441 2790 2475
rect 2700 2431 2790 2441
rect 2479 2295 2509 2425
rect 2700 2396 2730 2431
rect 2551 2367 2615 2383
rect 2551 2333 2561 2367
rect 2595 2333 2615 2367
rect 2686 2366 2730 2396
rect 2832 2389 2862 2589
rect 2935 2557 2965 2589
rect 2904 2541 2965 2557
rect 2904 2507 2914 2541
rect 2948 2507 2965 2541
rect 2904 2491 2965 2507
rect 3030 2473 3060 2589
rect 3115 2509 3145 2589
rect 3115 2493 3210 2509
rect 3007 2463 3073 2473
rect 3007 2449 3023 2463
rect 2788 2379 2862 2389
rect 2686 2351 2716 2366
rect 2551 2317 2615 2333
rect 2585 2295 2615 2317
rect 2788 2345 2804 2379
rect 2838 2345 2862 2379
rect 2788 2335 2862 2345
rect 2904 2429 3023 2449
rect 3057 2429 3073 2463
rect 2904 2419 3073 2429
rect 3115 2459 3166 2493
rect 3200 2459 3210 2493
rect 3115 2443 3210 2459
rect 3303 2450 3333 2539
rect 3387 2524 3417 2539
rect 3387 2494 3450 2524
rect 2805 2307 2835 2335
rect 2904 2295 2934 2419
rect 2987 2367 3053 2377
rect 2987 2333 3003 2367
rect 3037 2333 3053 2367
rect 2987 2323 3053 2333
rect 3003 2295 3033 2323
rect 3115 2307 3145 2443
rect 3303 2440 3378 2450
rect 3303 2406 3328 2440
rect 3362 2406 3378 2440
rect 3303 2396 3378 2406
rect 3420 2441 3450 2494
rect 4679 2667 4709 2693
rect 4763 2667 4793 2693
rect 4951 2673 4981 2699
rect 5036 2673 5066 2699
rect 5131 2673 5161 2699
rect 5234 2673 5264 2699
rect 5366 2673 5396 2699
rect 5461 2673 5491 2699
rect 5545 2673 5575 2699
rect 5659 2673 5689 2699
rect 5869 2673 5899 2699
rect 5953 2673 5983 2699
rect 6427 2673 7005 2699
rect 7265 2673 7295 2699
rect 7349 2673 7379 2699
rect 7559 2673 7589 2699
rect 7673 2673 7703 2699
rect 7757 2673 7787 2699
rect 7852 2673 7882 2699
rect 7984 2673 8014 2699
rect 8087 2673 8117 2699
rect 8182 2673 8212 2699
rect 8267 2673 8297 2699
rect 4679 2524 4709 2539
rect 4219 2473 4429 2499
rect 4646 2494 4709 2524
rect 4219 2467 4303 2473
rect 4161 2451 4303 2467
rect 3420 2425 3474 2441
rect 3303 2307 3333 2396
rect 3420 2391 3430 2425
rect 3464 2391 3474 2425
rect 4161 2417 4177 2451
rect 4211 2417 4303 2451
rect 4646 2441 4676 2494
rect 4763 2450 4793 2539
rect 4951 2509 4981 2589
rect 4161 2401 4303 2417
rect 4345 2415 4487 2431
rect 3420 2375 3474 2391
rect 4345 2381 4437 2415
rect 4471 2381 4487 2415
rect 3420 2352 3450 2375
rect 4345 2365 4487 2381
rect 4622 2425 4676 2441
rect 4622 2391 4632 2425
rect 4666 2391 4676 2425
rect 4718 2440 4793 2450
rect 4886 2493 4981 2509
rect 4886 2459 4896 2493
rect 4930 2459 4981 2493
rect 5036 2473 5066 2589
rect 5131 2557 5161 2589
rect 5131 2541 5192 2557
rect 5131 2507 5148 2541
rect 5182 2507 5192 2541
rect 5131 2491 5192 2507
rect 4886 2443 4981 2459
rect 4718 2406 4734 2440
rect 4768 2406 4793 2440
rect 4718 2396 4793 2406
rect 4622 2375 4676 2391
rect 4345 2359 4429 2365
rect 3387 2322 3450 2352
rect 3387 2307 3417 2322
rect 4219 2333 4429 2359
rect 4646 2352 4676 2375
rect 1183 2197 1301 2223
rect 1459 2197 1853 2223
rect 2111 2197 2141 2223
rect 2195 2197 2225 2223
rect 2384 2197 2414 2223
rect 2479 2197 2509 2223
rect 2585 2197 2615 2223
rect 2686 2197 2716 2223
rect 2805 2197 2835 2223
rect 2904 2197 2934 2223
rect 3003 2197 3033 2223
rect 3115 2197 3145 2223
rect 3303 2197 3333 2223
rect 3387 2197 3417 2223
rect 4646 2322 4709 2352
rect 4679 2307 4709 2322
rect 4763 2307 4793 2396
rect 4951 2307 4981 2443
rect 5023 2463 5089 2473
rect 5023 2429 5039 2463
rect 5073 2449 5089 2463
rect 5073 2429 5192 2449
rect 5023 2419 5192 2429
rect 5043 2367 5109 2377
rect 5043 2333 5059 2367
rect 5093 2333 5109 2367
rect 5043 2323 5109 2333
rect 5063 2295 5093 2323
rect 5162 2295 5192 2419
rect 5234 2389 5264 2589
rect 5366 2485 5396 2523
rect 5461 2491 5491 2589
rect 5545 2551 5575 2589
rect 5659 2557 5689 2589
rect 5544 2541 5610 2551
rect 5544 2507 5560 2541
rect 5594 2507 5610 2541
rect 5544 2497 5610 2507
rect 5659 2541 5740 2557
rect 5659 2507 5696 2541
rect 5730 2507 5740 2541
rect 5659 2491 5740 2507
rect 5306 2475 5396 2485
rect 5306 2441 5322 2475
rect 5356 2441 5396 2475
rect 5306 2431 5396 2441
rect 5366 2396 5396 2431
rect 5448 2475 5502 2491
rect 5448 2441 5458 2475
rect 5492 2455 5502 2475
rect 5492 2441 5617 2455
rect 5448 2425 5617 2441
rect 5234 2379 5308 2389
rect 5234 2345 5258 2379
rect 5292 2345 5308 2379
rect 5366 2366 5410 2396
rect 5380 2351 5410 2366
rect 5481 2367 5545 2383
rect 5234 2335 5308 2345
rect 5261 2307 5291 2335
rect 5481 2333 5501 2367
rect 5535 2333 5545 2367
rect 5481 2317 5545 2333
rect 5481 2295 5511 2317
rect 5587 2295 5617 2425
rect 5682 2307 5712 2491
rect 6427 2473 7005 2499
rect 7559 2557 7589 2589
rect 7508 2541 7589 2557
rect 7673 2551 7703 2589
rect 7508 2507 7518 2541
rect 7552 2507 7589 2541
rect 7508 2491 7589 2507
rect 7638 2541 7704 2551
rect 7638 2507 7654 2541
rect 7688 2507 7704 2541
rect 7638 2497 7704 2507
rect 7757 2491 7787 2589
rect 8455 2667 8485 2693
rect 8539 2667 8569 2693
rect 9003 2673 9581 2699
rect 5869 2441 5899 2473
rect 5953 2441 5983 2473
rect 6427 2451 6691 2473
rect 5759 2425 5901 2441
rect 5759 2391 5769 2425
rect 5803 2391 5901 2425
rect 5759 2375 5901 2391
rect 5943 2425 5997 2441
rect 5943 2391 5953 2425
rect 5987 2391 5997 2425
rect 6427 2417 6443 2451
rect 6477 2417 6542 2451
rect 6576 2417 6641 2451
rect 6675 2417 6691 2451
rect 7265 2441 7295 2473
rect 7349 2441 7379 2473
rect 6427 2401 6691 2417
rect 6733 2415 7005 2431
rect 5943 2375 5997 2391
rect 6733 2381 6749 2415
rect 6783 2381 6852 2415
rect 6886 2381 6955 2415
rect 6989 2381 7005 2415
rect 5871 2353 5901 2375
rect 5955 2353 5985 2375
rect 6733 2359 7005 2381
rect 7251 2425 7305 2441
rect 7251 2391 7261 2425
rect 7295 2391 7305 2425
rect 7251 2375 7305 2391
rect 7347 2425 7489 2441
rect 7347 2391 7445 2425
rect 7479 2391 7489 2425
rect 7347 2375 7489 2391
rect 6427 2333 7005 2359
rect 7263 2353 7293 2375
rect 7347 2353 7377 2375
rect 7536 2307 7566 2491
rect 7746 2475 7800 2491
rect 7746 2455 7756 2475
rect 7631 2441 7756 2455
rect 7790 2441 7800 2475
rect 7631 2425 7800 2441
rect 7852 2485 7882 2523
rect 7852 2475 7942 2485
rect 7852 2441 7892 2475
rect 7926 2441 7942 2475
rect 7852 2431 7942 2441
rect 7631 2295 7661 2425
rect 7852 2396 7882 2431
rect 7703 2367 7767 2383
rect 7703 2333 7713 2367
rect 7747 2333 7767 2367
rect 7838 2366 7882 2396
rect 7984 2389 8014 2589
rect 8087 2557 8117 2589
rect 8056 2541 8117 2557
rect 8056 2507 8066 2541
rect 8100 2507 8117 2541
rect 8056 2491 8117 2507
rect 8182 2473 8212 2589
rect 8267 2509 8297 2589
rect 8267 2493 8362 2509
rect 8159 2463 8225 2473
rect 8159 2449 8175 2463
rect 7940 2379 8014 2389
rect 7838 2351 7868 2366
rect 7703 2317 7767 2333
rect 7737 2295 7767 2317
rect 7940 2345 7956 2379
rect 7990 2345 8014 2379
rect 7940 2335 8014 2345
rect 8056 2429 8175 2449
rect 8209 2429 8225 2463
rect 8056 2419 8225 2429
rect 8267 2459 8318 2493
rect 8352 2459 8362 2493
rect 8267 2443 8362 2459
rect 8455 2450 8485 2539
rect 8539 2524 8569 2539
rect 8539 2494 8602 2524
rect 7957 2307 7987 2335
rect 8056 2295 8086 2419
rect 8139 2367 8205 2377
rect 8139 2333 8155 2367
rect 8189 2333 8205 2367
rect 8139 2323 8205 2333
rect 8155 2295 8185 2323
rect 8267 2307 8297 2443
rect 8455 2440 8530 2450
rect 8455 2406 8480 2440
rect 8514 2406 8530 2440
rect 8455 2396 8530 2406
rect 8572 2441 8602 2494
rect 9831 2667 9861 2693
rect 9915 2667 9945 2693
rect 10103 2673 10133 2699
rect 10188 2673 10218 2699
rect 10283 2673 10313 2699
rect 10386 2673 10416 2699
rect 10518 2673 10548 2699
rect 10613 2673 10643 2699
rect 10697 2673 10727 2699
rect 10811 2673 10841 2699
rect 11021 2673 11051 2699
rect 11105 2673 11135 2699
rect 11579 2673 11789 2699
rect 11957 2673 11987 2699
rect 12041 2673 12071 2699
rect 12251 2673 12281 2699
rect 12365 2673 12395 2699
rect 12449 2673 12479 2699
rect 12544 2673 12574 2699
rect 12676 2673 12706 2699
rect 12779 2673 12809 2699
rect 12874 2673 12904 2699
rect 12959 2673 12989 2699
rect 9831 2524 9861 2539
rect 9003 2473 9581 2499
rect 9798 2494 9861 2524
rect 9003 2451 9267 2473
rect 8572 2425 8626 2441
rect 8455 2307 8485 2396
rect 8572 2391 8582 2425
rect 8616 2391 8626 2425
rect 9003 2417 9019 2451
rect 9053 2417 9118 2451
rect 9152 2417 9217 2451
rect 9251 2417 9267 2451
rect 9798 2441 9828 2494
rect 9915 2450 9945 2539
rect 10103 2509 10133 2589
rect 9003 2401 9267 2417
rect 9309 2415 9581 2431
rect 8572 2375 8626 2391
rect 9309 2381 9325 2415
rect 9359 2381 9428 2415
rect 9462 2381 9531 2415
rect 9565 2381 9581 2415
rect 8572 2352 8602 2375
rect 9309 2359 9581 2381
rect 9774 2425 9828 2441
rect 9774 2391 9784 2425
rect 9818 2391 9828 2425
rect 9870 2440 9945 2450
rect 10038 2493 10133 2509
rect 10038 2459 10048 2493
rect 10082 2459 10133 2493
rect 10188 2473 10218 2589
rect 10283 2557 10313 2589
rect 10283 2541 10344 2557
rect 10283 2507 10300 2541
rect 10334 2507 10344 2541
rect 10283 2491 10344 2507
rect 10038 2443 10133 2459
rect 9870 2406 9886 2440
rect 9920 2406 9945 2440
rect 9870 2396 9945 2406
rect 9774 2375 9828 2391
rect 8539 2322 8602 2352
rect 8539 2307 8569 2322
rect 9003 2333 9581 2359
rect 9798 2352 9828 2375
rect 9798 2322 9861 2352
rect 9831 2307 9861 2322
rect 9915 2307 9945 2396
rect 10103 2307 10133 2443
rect 10175 2463 10241 2473
rect 10175 2429 10191 2463
rect 10225 2449 10241 2463
rect 10225 2429 10344 2449
rect 10175 2419 10344 2429
rect 10195 2367 10261 2377
rect 10195 2333 10211 2367
rect 10245 2333 10261 2367
rect 10195 2323 10261 2333
rect 10215 2295 10245 2323
rect 10314 2295 10344 2419
rect 10386 2389 10416 2589
rect 10518 2485 10548 2523
rect 10613 2491 10643 2589
rect 10697 2551 10727 2589
rect 10811 2557 10841 2589
rect 10696 2541 10762 2551
rect 10696 2507 10712 2541
rect 10746 2507 10762 2541
rect 10696 2497 10762 2507
rect 10811 2541 10892 2557
rect 10811 2507 10848 2541
rect 10882 2507 10892 2541
rect 10811 2491 10892 2507
rect 10458 2475 10548 2485
rect 10458 2441 10474 2475
rect 10508 2441 10548 2475
rect 10458 2431 10548 2441
rect 10518 2396 10548 2431
rect 10600 2475 10654 2491
rect 10600 2441 10610 2475
rect 10644 2455 10654 2475
rect 10644 2441 10769 2455
rect 10600 2425 10769 2441
rect 10386 2379 10460 2389
rect 10386 2345 10410 2379
rect 10444 2345 10460 2379
rect 10518 2366 10562 2396
rect 10532 2351 10562 2366
rect 10633 2367 10697 2383
rect 10386 2335 10460 2345
rect 10413 2307 10443 2335
rect 10633 2333 10653 2367
rect 10687 2333 10697 2367
rect 10633 2317 10697 2333
rect 10633 2295 10663 2317
rect 10739 2295 10769 2425
rect 10834 2307 10864 2491
rect 11579 2473 11789 2499
rect 12251 2557 12281 2589
rect 12200 2541 12281 2557
rect 12365 2551 12395 2589
rect 12200 2507 12210 2541
rect 12244 2507 12281 2541
rect 12200 2491 12281 2507
rect 12330 2541 12396 2551
rect 12330 2507 12346 2541
rect 12380 2507 12396 2541
rect 12330 2497 12396 2507
rect 12449 2491 12479 2589
rect 13147 2667 13177 2693
rect 13231 2667 13261 2693
rect 13419 2673 13813 2699
rect 11021 2441 11051 2473
rect 11105 2441 11135 2473
rect 11579 2467 11663 2473
rect 11521 2451 11663 2467
rect 10911 2425 11053 2441
rect 10911 2391 10921 2425
rect 10955 2391 11053 2425
rect 10911 2375 11053 2391
rect 11095 2425 11149 2441
rect 11095 2391 11105 2425
rect 11139 2391 11149 2425
rect 11521 2417 11537 2451
rect 11571 2417 11663 2451
rect 11957 2441 11987 2473
rect 12041 2441 12071 2473
rect 11521 2401 11663 2417
rect 11705 2415 11847 2431
rect 11095 2375 11149 2391
rect 11705 2381 11797 2415
rect 11831 2381 11847 2415
rect 11023 2353 11053 2375
rect 11107 2353 11137 2375
rect 11705 2365 11847 2381
rect 11943 2425 11997 2441
rect 11943 2391 11953 2425
rect 11987 2391 11997 2425
rect 11943 2375 11997 2391
rect 12039 2425 12181 2441
rect 12039 2391 12137 2425
rect 12171 2391 12181 2425
rect 12039 2375 12181 2391
rect 11705 2359 11789 2365
rect 11579 2333 11789 2359
rect 11955 2353 11985 2375
rect 12039 2353 12069 2375
rect 12228 2307 12258 2491
rect 12438 2475 12492 2491
rect 12438 2455 12448 2475
rect 12323 2441 12448 2455
rect 12482 2441 12492 2475
rect 12323 2425 12492 2441
rect 12544 2485 12574 2523
rect 12544 2475 12634 2485
rect 12544 2441 12584 2475
rect 12618 2441 12634 2475
rect 12544 2431 12634 2441
rect 12323 2295 12353 2425
rect 12544 2396 12574 2431
rect 12395 2367 12459 2383
rect 12395 2333 12405 2367
rect 12439 2333 12459 2367
rect 12530 2366 12574 2396
rect 12676 2389 12706 2589
rect 12779 2557 12809 2589
rect 12748 2541 12809 2557
rect 12748 2507 12758 2541
rect 12792 2507 12809 2541
rect 12748 2491 12809 2507
rect 12874 2473 12904 2589
rect 12959 2509 12989 2589
rect 12959 2493 13054 2509
rect 12851 2463 12917 2473
rect 12851 2449 12867 2463
rect 12632 2379 12706 2389
rect 12530 2351 12560 2366
rect 12395 2317 12459 2333
rect 12429 2295 12459 2317
rect 12632 2345 12648 2379
rect 12682 2345 12706 2379
rect 12632 2335 12706 2345
rect 12748 2429 12867 2449
rect 12901 2429 12917 2463
rect 12748 2419 12917 2429
rect 12959 2459 13010 2493
rect 13044 2459 13054 2493
rect 12959 2443 13054 2459
rect 13147 2450 13177 2539
rect 13231 2524 13261 2539
rect 13231 2494 13294 2524
rect 14281 2660 14377 2699
rect 12649 2307 12679 2335
rect 12748 2295 12778 2419
rect 12831 2367 12897 2377
rect 12831 2333 12847 2367
rect 12881 2333 12897 2367
rect 12831 2323 12897 2333
rect 12847 2295 12877 2323
rect 12959 2307 12989 2443
rect 13147 2440 13222 2450
rect 13147 2406 13172 2440
rect 13206 2406 13222 2440
rect 13147 2396 13222 2406
rect 13264 2441 13294 2494
rect 13419 2473 13813 2499
rect 14281 2626 14331 2660
rect 14365 2626 14377 2660
rect 14281 2592 14377 2626
rect 14281 2558 14331 2592
rect 14365 2558 14377 2592
rect 13419 2451 13595 2473
rect 13264 2425 13318 2441
rect 13147 2307 13177 2396
rect 13264 2391 13274 2425
rect 13308 2391 13318 2425
rect 13419 2417 13435 2451
rect 13469 2417 13545 2451
rect 13579 2417 13595 2451
rect 13419 2401 13595 2417
rect 13637 2415 13813 2431
rect 13264 2375 13318 2391
rect 13637 2381 13653 2415
rect 13687 2381 13763 2415
rect 13797 2381 13813 2415
rect 13264 2352 13294 2375
rect 13637 2359 13813 2381
rect 13231 2322 13294 2352
rect 13419 2333 13813 2359
rect 14281 2417 14377 2558
rect 13231 2307 13261 2322
rect 14281 2325 14377 2408
rect 14281 2291 14331 2325
rect 14365 2291 14377 2325
rect 14281 2257 14377 2291
rect 14281 2223 14331 2257
rect 14365 2223 14377 2257
rect 4219 2197 4429 2223
rect 4679 2197 4709 2223
rect 4763 2197 4793 2223
rect 4951 2197 4981 2223
rect 5063 2197 5093 2223
rect 5162 2197 5192 2223
rect 5261 2197 5291 2223
rect 5380 2197 5410 2223
rect 5481 2197 5511 2223
rect 5587 2197 5617 2223
rect 5682 2197 5712 2223
rect 5871 2197 5901 2223
rect 5955 2197 5985 2223
rect 6427 2197 7005 2223
rect 7263 2197 7293 2223
rect 7347 2197 7377 2223
rect 7536 2197 7566 2223
rect 7631 2197 7661 2223
rect 7737 2197 7767 2223
rect 7838 2197 7868 2223
rect 7957 2197 7987 2223
rect 8056 2197 8086 2223
rect 8155 2197 8185 2223
rect 8267 2197 8297 2223
rect 8455 2197 8485 2223
rect 8539 2197 8569 2223
rect 9003 2197 9581 2223
rect 9831 2197 9861 2223
rect 9915 2197 9945 2223
rect 10103 2197 10133 2223
rect 10215 2197 10245 2223
rect 10314 2197 10344 2223
rect 10413 2197 10443 2223
rect 10532 2197 10562 2223
rect 10633 2197 10663 2223
rect 10739 2197 10769 2223
rect 10834 2197 10864 2223
rect 11023 2197 11053 2223
rect 11107 2197 11137 2223
rect 11579 2197 11789 2223
rect 11955 2197 11985 2223
rect 12039 2197 12069 2223
rect 12228 2197 12258 2223
rect 12323 2197 12353 2223
rect 12429 2197 12459 2223
rect 12530 2197 12560 2223
rect 12649 2197 12679 2223
rect 12748 2197 12778 2223
rect 12847 2197 12877 2223
rect 12959 2197 12989 2223
rect 13147 2197 13177 2223
rect 13231 2197 13261 2223
rect 13419 2197 13813 2223
rect 14281 2197 14377 2223
rect 14419 2660 14515 2699
rect 14615 2673 15561 2699
rect 15719 2673 16297 2699
rect 16915 2673 16945 2699
rect 17003 2673 17033 2699
rect 17191 2673 17401 2699
rect 14419 2626 14431 2660
rect 14465 2626 14515 2660
rect 14419 2592 14515 2626
rect 14419 2558 14431 2592
rect 14465 2558 14515 2592
rect 14419 2417 14515 2558
rect 14419 2329 14515 2408
rect 14615 2473 15561 2499
rect 15719 2473 16297 2499
rect 14615 2451 15065 2473
rect 14615 2417 14887 2451
rect 14921 2417 15065 2451
rect 15719 2451 15983 2473
rect 16915 2454 16945 2515
rect 17003 2500 17033 2515
rect 17003 2476 17039 2500
rect 17559 2665 17589 2691
rect 17654 2673 17684 2699
rect 17738 2673 17768 2699
rect 17927 2673 18505 2699
rect 18663 2673 18781 2699
rect 14615 2401 15065 2417
rect 15107 2415 15561 2431
rect 15107 2381 15251 2415
rect 15285 2381 15561 2415
rect 15719 2417 15735 2451
rect 15769 2417 15834 2451
rect 15868 2417 15933 2451
rect 15967 2417 15983 2451
rect 16911 2438 16965 2454
rect 15719 2401 15983 2417
rect 16025 2415 16297 2431
rect 15107 2359 15561 2381
rect 16025 2381 16041 2415
rect 16075 2381 16144 2415
rect 16178 2381 16247 2415
rect 16281 2381 16297 2415
rect 16911 2404 16921 2438
rect 16955 2404 16965 2438
rect 16911 2388 16965 2404
rect 17009 2441 17039 2476
rect 17191 2473 17401 2499
rect 17191 2467 17275 2473
rect 17133 2451 17275 2467
rect 17009 2425 17085 2441
rect 17009 2391 17041 2425
rect 17075 2391 17085 2425
rect 17133 2417 17149 2451
rect 17183 2417 17275 2451
rect 17559 2441 17589 2537
rect 17927 2473 18505 2499
rect 17654 2441 17684 2473
rect 17738 2441 17768 2473
rect 17133 2401 17275 2417
rect 17317 2415 17459 2431
rect 16025 2359 16297 2381
rect 14615 2333 15561 2359
rect 15719 2333 16297 2359
rect 14419 2295 14431 2329
rect 14465 2295 14515 2329
rect 14419 2261 14515 2295
rect 14419 2227 14431 2261
rect 14465 2227 14515 2261
rect 14419 2197 14515 2227
rect 16915 2327 16945 2388
rect 17009 2375 17085 2391
rect 17317 2381 17409 2415
rect 17443 2381 17459 2415
rect 17009 2366 17039 2375
rect 17003 2342 17039 2366
rect 17317 2365 17459 2381
rect 17507 2425 17589 2441
rect 17507 2391 17517 2425
rect 17551 2391 17589 2425
rect 17507 2375 17589 2391
rect 17631 2425 17768 2441
rect 17631 2391 17641 2425
rect 17675 2391 17768 2425
rect 17927 2451 18191 2473
rect 18663 2469 18781 2499
rect 17927 2417 17943 2451
rect 17977 2417 18042 2451
rect 18076 2417 18141 2451
rect 18175 2417 18191 2451
rect 18743 2467 18781 2469
rect 18743 2451 18809 2467
rect 17927 2401 18191 2417
rect 18233 2415 18505 2431
rect 17631 2375 17768 2391
rect 17317 2359 17401 2365
rect 17003 2327 17033 2342
rect 17191 2333 17401 2359
rect 17559 2307 17589 2375
rect 17654 2353 17684 2375
rect 17738 2353 17768 2375
rect 18233 2381 18249 2415
rect 18283 2381 18352 2415
rect 18386 2381 18455 2415
rect 18489 2381 18505 2415
rect 18233 2359 18505 2381
rect 18635 2411 18701 2427
rect 18635 2377 18651 2411
rect 18685 2377 18701 2411
rect 18743 2417 18759 2451
rect 18793 2417 18809 2451
rect 18743 2401 18809 2417
rect 18635 2361 18701 2377
rect 17927 2333 18505 2359
rect 18663 2359 18701 2361
rect 18663 2333 18781 2359
rect 14615 2197 15561 2223
rect 15719 2197 16297 2223
rect 16915 2197 16945 2223
rect 17003 2197 17033 2223
rect 17191 2197 17401 2223
rect 17559 2197 17589 2223
rect 17654 2197 17684 2223
rect 17738 2197 17768 2223
rect 17927 2197 18505 2223
rect 18663 2197 18781 2223
<< polycont >>
rect 1171 7341 1205 7375
rect 1279 7381 1313 7415
rect 1737 7367 1771 7401
rect 1861 7367 1895 7401
rect 2283 7341 2317 7375
rect 2647 7377 2681 7411
rect 3131 7341 3165 7375
rect 3241 7341 3275 7375
rect 3349 7377 3383 7411
rect 3459 7377 3493 7411
rect 4129 7367 4163 7401
rect 4253 7367 4287 7401
rect 4675 7341 4709 7375
rect 5039 7377 5073 7411
rect 5785 7367 5819 7401
rect 5909 7367 5943 7401
rect 6047 7341 6081 7375
rect 6155 7381 6189 7415
rect 6699 7341 6733 7375
rect 7063 7377 7097 7411
rect 7489 7341 7523 7375
rect 7749 7377 7783 7411
rect 7857 7367 7891 7401
rect 7981 7367 8015 7401
rect 8283 7341 8317 7375
rect 8393 7341 8427 7375
rect 8501 7377 8535 7411
rect 8611 7377 8645 7411
rect 9019 7341 9053 7375
rect 9129 7341 9163 7375
rect 9237 7377 9271 7411
rect 9347 7377 9381 7411
rect 9697 7341 9731 7375
rect 9957 7377 9991 7411
rect 10117 7367 10151 7401
rect 10221 7367 10255 7401
rect 10491 7341 10525 7375
rect 10590 7341 10624 7375
rect 10689 7341 10723 7375
rect 10797 7377 10831 7411
rect 10900 7377 10934 7411
rect 11003 7377 11037 7411
rect 11199 7341 11233 7375
rect 11307 7381 11341 7415
rect 11595 7341 11629 7375
rect 11694 7341 11728 7375
rect 11793 7341 11827 7375
rect 11901 7377 11935 7411
rect 12004 7377 12038 7411
rect 12107 7377 12141 7411
rect 12273 7367 12307 7401
rect 12397 7367 12431 7401
rect 12955 7341 12989 7375
rect 13319 7377 13353 7411
rect 13775 7341 13809 7375
rect 13883 7381 13917 7415
rect 14113 7341 14147 7375
rect 14373 7377 14407 7411
rect 14481 7367 14515 7401
rect 14605 7367 14639 7401
rect 15163 7341 15197 7375
rect 15527 7377 15561 7411
rect 16011 7341 16045 7375
rect 16121 7341 16155 7375
rect 16229 7377 16263 7411
rect 16339 7377 16373 7411
rect 16873 7367 16907 7401
rect 16997 7367 17031 7401
rect 17299 7341 17333 7375
rect 17398 7341 17432 7375
rect 17497 7341 17531 7375
rect 17605 7377 17639 7411
rect 17708 7377 17742 7411
rect 17811 7377 17845 7411
rect 18069 7367 18103 7401
rect 18193 7367 18227 7401
rect 18651 7381 18685 7415
rect 18759 7341 18793 7375
rect 1171 6769 1205 6803
rect 1279 6729 1313 6763
rect 1731 6769 1765 6803
rect 2095 6733 2129 6767
rect 2835 6769 2869 6803
rect 3199 6733 3233 6767
rect 4123 6769 4157 6803
rect 4487 6733 4521 6767
rect 5227 6769 5261 6803
rect 5591 6733 5625 6767
rect 6331 6769 6365 6803
rect 6695 6733 6729 6767
rect 7435 6769 7469 6803
rect 7799 6733 7833 6767
rect 8283 6769 8317 6803
rect 8393 6769 8427 6803
rect 8501 6733 8535 6767
rect 8611 6733 8645 6767
rect 9275 6769 9309 6803
rect 9639 6733 9673 6767
rect 10379 6769 10413 6803
rect 10743 6733 10777 6767
rect 11483 6769 11517 6803
rect 11847 6733 11881 6767
rect 12587 6769 12621 6803
rect 12951 6733 12985 6767
rect 13435 6769 13469 6803
rect 13545 6769 13579 6803
rect 13653 6733 13687 6767
rect 13763 6733 13797 6767
rect 14427 6769 14461 6803
rect 14791 6733 14825 6767
rect 15531 6769 15565 6803
rect 15895 6733 15929 6767
rect 16635 6769 16669 6803
rect 16999 6733 17033 6767
rect 17739 6769 17773 6803
rect 18103 6733 18137 6767
rect 18651 6729 18685 6763
rect 18759 6769 18793 6803
rect 1171 6253 1205 6287
rect 1279 6293 1313 6327
rect 1731 6253 1765 6287
rect 2095 6289 2129 6323
rect 2835 6253 2869 6287
rect 3199 6289 3233 6323
rect 3939 6253 3973 6287
rect 4303 6289 4337 6323
rect 5043 6253 5077 6287
rect 5407 6289 5441 6323
rect 5833 6253 5867 6287
rect 6093 6289 6127 6323
rect 6699 6253 6733 6287
rect 7063 6289 7097 6323
rect 7803 6253 7837 6287
rect 8167 6289 8201 6323
rect 8907 6253 8941 6287
rect 9271 6289 9305 6323
rect 10011 6253 10045 6287
rect 10375 6289 10409 6323
rect 10859 6253 10893 6287
rect 10969 6253 11003 6287
rect 11077 6289 11111 6323
rect 11187 6289 11221 6323
rect 11851 6253 11885 6287
rect 12215 6289 12249 6323
rect 12955 6253 12989 6287
rect 13319 6289 13353 6323
rect 14059 6253 14093 6287
rect 14423 6289 14457 6323
rect 15163 6253 15197 6287
rect 15527 6289 15561 6323
rect 16011 6253 16045 6287
rect 16121 6253 16155 6287
rect 16229 6289 16263 6323
rect 16339 6289 16373 6323
rect 17003 6253 17037 6287
rect 17367 6289 17401 6323
rect 17851 6253 17885 6287
rect 17950 6253 17984 6287
rect 18049 6253 18083 6287
rect 18157 6289 18191 6323
rect 18260 6289 18294 6323
rect 18363 6289 18397 6323
rect 18651 6293 18685 6327
rect 18759 6253 18793 6287
rect 1171 5681 1205 5715
rect 1279 5641 1313 5675
rect 1475 5681 1509 5715
rect 1574 5681 1608 5715
rect 1673 5681 1707 5715
rect 1781 5645 1815 5679
rect 1884 5645 1918 5679
rect 1987 5645 2021 5679
rect 2245 5655 2279 5689
rect 2365 5668 2399 5702
rect 2579 5681 2613 5715
rect 2689 5681 2723 5715
rect 2797 5645 2831 5679
rect 2907 5645 2941 5679
rect 3121 5668 3155 5702
rect 3241 5655 3275 5689
rect 3349 5681 3383 5715
rect 3609 5645 3643 5679
rect 4123 5681 4157 5715
rect 4487 5645 4521 5679
rect 5227 5681 5261 5715
rect 5591 5645 5625 5679
rect 6075 5681 6109 5715
rect 6174 5681 6208 5715
rect 6273 5681 6307 5715
rect 6381 5645 6415 5679
rect 6484 5645 6518 5679
rect 6587 5645 6621 5679
rect 6802 5655 6836 5689
rect 6898 5655 6932 5689
rect 7207 5732 7241 5766
rect 7039 5619 7073 5653
rect 7375 5732 7409 5766
rect 7135 5619 7169 5653
rect 7297 5619 7331 5653
rect 7895 5681 7929 5715
rect 8259 5645 8293 5679
rect 9019 5681 9053 5715
rect 9118 5681 9152 5715
rect 9217 5681 9251 5715
rect 9325 5645 9359 5679
rect 9428 5645 9462 5679
rect 9531 5645 9565 5679
rect 9930 5655 9964 5689
rect 10026 5655 10060 5689
rect 10335 5732 10369 5766
rect 10167 5619 10201 5653
rect 10503 5732 10537 5766
rect 10263 5619 10297 5653
rect 10425 5619 10459 5653
rect 10709 5681 10743 5715
rect 10969 5645 11003 5679
rect 11143 5655 11177 5689
rect 11251 5655 11285 5689
rect 11392 5655 11426 5689
rect 11595 5681 11629 5715
rect 11694 5681 11728 5715
rect 11793 5681 11827 5715
rect 11901 5645 11935 5679
rect 12004 5645 12038 5679
rect 12107 5645 12141 5679
rect 12322 5655 12356 5689
rect 12418 5655 12452 5689
rect 12727 5732 12761 5766
rect 12559 5619 12593 5653
rect 12895 5732 12929 5766
rect 12655 5619 12689 5653
rect 12817 5619 12851 5653
rect 13159 5681 13193 5715
rect 13258 5681 13292 5715
rect 13357 5681 13391 5715
rect 13465 5645 13499 5679
rect 13568 5645 13602 5679
rect 13671 5645 13705 5679
rect 14346 5655 14380 5689
rect 14442 5655 14476 5689
rect 14751 5732 14785 5766
rect 14583 5619 14617 5653
rect 14919 5732 14953 5766
rect 14679 5619 14713 5653
rect 14841 5619 14875 5653
rect 15439 5681 15473 5715
rect 15803 5645 15837 5679
rect 16543 5681 16577 5715
rect 16907 5645 16941 5679
rect 17647 5681 17681 5715
rect 18011 5645 18045 5679
rect 18651 5641 18685 5675
rect 18759 5681 18793 5715
rect 1171 5165 1205 5199
rect 1279 5205 1313 5239
rect 1475 5165 1509 5199
rect 1585 5165 1619 5199
rect 1693 5201 1727 5235
rect 1803 5201 1837 5235
rect 2035 5191 2069 5225
rect 2143 5191 2177 5225
rect 2284 5191 2318 5225
rect 2429 5165 2463 5199
rect 2689 5201 2723 5235
rect 2955 5191 2989 5225
rect 3063 5191 3097 5225
rect 3204 5191 3238 5225
rect 3349 5165 3383 5199
rect 3609 5201 3643 5235
rect 3717 5191 3751 5225
rect 3841 5191 3875 5225
rect 4085 5165 4119 5199
rect 4345 5201 4379 5235
rect 4453 5191 4487 5225
rect 5043 5165 5077 5199
rect 5407 5201 5441 5235
rect 5881 5178 5915 5212
rect 6001 5191 6035 5225
rect 6415 5165 6449 5199
rect 6523 5205 6557 5239
rect 6710 5191 6744 5225
rect 6806 5191 6840 5225
rect 6947 5227 6981 5261
rect 7043 5227 7077 5261
rect 7205 5227 7239 5261
rect 7115 5114 7149 5148
rect 7489 5165 7523 5199
rect 7749 5201 7783 5235
rect 7906 5191 7940 5225
rect 8002 5191 8036 5225
rect 8143 5227 8177 5261
rect 8239 5227 8273 5261
rect 8401 5227 8435 5261
rect 7283 5114 7317 5148
rect 8311 5114 8345 5148
rect 8685 5165 8719 5199
rect 8945 5201 8979 5235
rect 9227 5191 9261 5225
rect 9365 5191 9399 5225
rect 9465 5191 9499 5225
rect 9593 5191 9627 5225
rect 8479 5114 8513 5148
rect 9755 5165 9789 5199
rect 9854 5165 9888 5199
rect 9953 5165 9987 5199
rect 10061 5201 10095 5235
rect 10164 5201 10198 5235
rect 10267 5201 10301 5235
rect 10482 5191 10516 5225
rect 10578 5191 10612 5225
rect 10719 5227 10753 5261
rect 10815 5227 10849 5261
rect 10977 5227 11011 5261
rect 10887 5114 10921 5148
rect 11055 5114 11089 5148
rect 11851 5165 11885 5199
rect 12215 5201 12249 5235
rect 12641 5165 12675 5199
rect 12901 5201 12935 5235
rect 13150 5191 13184 5225
rect 13246 5191 13280 5225
rect 13387 5227 13421 5261
rect 13483 5227 13517 5261
rect 13645 5227 13679 5261
rect 13555 5114 13589 5148
rect 13723 5114 13757 5148
rect 14243 5165 14277 5199
rect 14607 5201 14641 5235
rect 15347 5165 15381 5199
rect 15711 5201 15745 5235
rect 16137 5165 16171 5199
rect 16397 5201 16431 5235
rect 17003 5165 17037 5199
rect 17367 5201 17401 5235
rect 17851 5165 17885 5199
rect 17950 5165 17984 5199
rect 18049 5165 18083 5199
rect 18157 5201 18191 5235
rect 18260 5201 18294 5235
rect 18363 5201 18397 5235
rect 18651 5205 18685 5239
rect 18759 5165 18793 5199
rect 1171 4593 1205 4627
rect 1279 4553 1313 4587
rect 1475 4593 1509 4627
rect 1585 4593 1619 4627
rect 1693 4557 1727 4591
rect 1803 4557 1837 4591
rect 2056 4567 2090 4601
rect 2320 4635 2354 4669
rect 2572 4683 2606 4717
rect 2158 4582 2192 4616
rect 2463 4605 2497 4639
rect 2483 4509 2517 4543
rect 2984 4683 3018 4717
rect 3120 4683 3154 4717
rect 2746 4617 2780 4651
rect 2882 4617 2916 4651
rect 2682 4521 2716 4555
rect 2925 4509 2959 4543
rect 3193 4567 3227 4601
rect 3377 4567 3411 4601
rect 4059 4567 4093 4601
rect 4167 4567 4201 4601
rect 4308 4567 4342 4601
rect 4453 4593 4487 4627
rect 4713 4557 4747 4591
rect 4995 4567 5029 4601
rect 5133 4567 5167 4601
rect 5233 4567 5267 4601
rect 5361 4567 5395 4601
rect 5465 4593 5499 4627
rect 5725 4557 5759 4591
rect 5915 4567 5949 4601
rect 6053 4567 6087 4601
rect 6153 4567 6187 4601
rect 6281 4567 6315 4601
rect 6385 4593 6419 4627
rect 6645 4557 6679 4591
rect 6748 4567 6782 4601
rect 7012 4635 7046 4669
rect 7264 4683 7298 4717
rect 6850 4582 6884 4616
rect 7155 4605 7189 4639
rect 7175 4509 7209 4543
rect 7676 4683 7710 4717
rect 7812 4683 7846 4717
rect 7438 4617 7472 4651
rect 7574 4617 7608 4651
rect 7374 4521 7408 4555
rect 7617 4509 7651 4543
rect 7885 4567 7919 4601
rect 8069 4567 8103 4601
rect 8283 4593 8317 4627
rect 8393 4593 8427 4627
rect 10278 4683 10312 4717
rect 10414 4683 10448 4717
rect 8501 4557 8535 4591
rect 8611 4557 8645 4591
rect 9019 4593 9053 4627
rect 9118 4593 9152 4627
rect 9217 4593 9251 4627
rect 9325 4557 9359 4591
rect 9428 4557 9462 4591
rect 9531 4557 9565 4591
rect 9727 4593 9761 4627
rect 9835 4553 9869 4587
rect 10021 4567 10055 4601
rect 10205 4567 10239 4601
rect 10516 4617 10550 4651
rect 10652 4617 10686 4651
rect 10473 4509 10507 4543
rect 10826 4683 10860 4717
rect 10716 4521 10750 4555
rect 10935 4605 10969 4639
rect 11078 4635 11112 4669
rect 10915 4509 10949 4543
rect 11240 4582 11274 4616
rect 11342 4567 11376 4601
rect 11445 4593 11479 4627
rect 11705 4557 11739 4591
rect 11895 4567 11929 4601
rect 12033 4567 12067 4601
rect 12133 4567 12167 4601
rect 12261 4567 12295 4601
rect 12365 4593 12399 4627
rect 12625 4557 12659 4591
rect 12815 4567 12849 4601
rect 12953 4567 12987 4601
rect 13053 4567 13087 4601
rect 13181 4567 13215 4601
rect 13343 4593 13377 4627
rect 13442 4593 13476 4627
rect 13541 4593 13575 4627
rect 13649 4557 13683 4591
rect 13752 4557 13786 4591
rect 13855 4557 13889 4591
rect 14143 4593 14177 4627
rect 14251 4553 14285 4587
rect 14426 4567 14460 4601
rect 14567 4567 14601 4601
rect 14675 4567 14709 4601
rect 15163 4593 15197 4627
rect 15527 4557 15561 4591
rect 16267 4593 16301 4627
rect 16631 4557 16665 4591
rect 17371 4593 17405 4627
rect 17735 4557 17769 4591
rect 18161 4593 18195 4627
rect 18421 4557 18455 4591
rect 18651 4553 18685 4587
rect 18759 4593 18793 4627
rect 1171 4077 1205 4111
rect 1279 4117 1313 4151
rect 1475 4077 1509 4111
rect 1585 4077 1619 4111
rect 1693 4113 1727 4147
rect 1803 4113 1837 4147
rect 1969 4103 2003 4137
rect 2089 4090 2123 4124
rect 2245 4077 2279 4111
rect 2505 4113 2539 4147
rect 2661 4103 2695 4137
rect 2845 4103 2879 4137
rect 3113 4161 3147 4195
rect 3356 4149 3390 4183
rect 3156 4053 3190 4087
rect 3292 4053 3326 4087
rect 2918 3987 2952 4021
rect 3054 3987 3088 4021
rect 3555 4161 3589 4195
rect 3575 4065 3609 4099
rect 3880 4088 3914 4122
rect 3466 3987 3500 4021
rect 3718 4035 3752 4069
rect 3982 4103 4016 4137
rect 4143 4077 4177 4111
rect 4253 4077 4287 4111
rect 4361 4113 4395 4147
rect 4471 4113 4505 4147
rect 4685 4103 4719 4137
rect 4869 4103 4903 4137
rect 5137 4161 5171 4195
rect 5380 4149 5414 4183
rect 5180 4053 5214 4087
rect 5316 4053 5350 4087
rect 4942 3987 4976 4021
rect 5078 3987 5112 4021
rect 5579 4161 5613 4195
rect 5599 4065 5633 4099
rect 5904 4088 5938 4122
rect 5490 3987 5524 4021
rect 5742 4035 5776 4069
rect 6006 4103 6040 4137
rect 6443 4077 6477 4111
rect 6553 4077 6587 4111
rect 6661 4113 6695 4147
rect 6771 4113 6805 4147
rect 7019 4103 7053 4137
rect 7157 4103 7191 4137
rect 7257 4103 7291 4137
rect 7385 4103 7419 4137
rect 7489 4077 7523 4111
rect 7749 4113 7783 4147
rect 7857 4103 7891 4137
rect 8284 4103 8318 4137
rect 8352 4103 8386 4137
rect 8420 4103 8454 4137
rect 8488 4103 8522 4137
rect 8556 4103 8590 4137
rect 8624 4103 8658 4137
rect 8692 4103 8726 4137
rect 8760 4103 8794 4137
rect 8828 4103 8862 4137
rect 8896 4103 8930 4137
rect 8964 4103 8998 4137
rect 9032 4103 9066 4137
rect 9100 4103 9134 4137
rect 9168 4103 9202 4137
rect 9236 4103 9270 4137
rect 9304 4103 9338 4137
rect 9755 4077 9789 4111
rect 9854 4077 9888 4111
rect 9953 4077 9987 4111
rect 10061 4113 10095 4147
rect 10164 4113 10198 4147
rect 10267 4113 10301 4147
rect 10607 4103 10641 4137
rect 10745 4103 10779 4137
rect 10845 4103 10879 4137
rect 10973 4103 11007 4137
rect 11077 4077 11111 4111
rect 11337 4113 11371 4147
rect 11716 4103 11750 4137
rect 11818 4088 11852 4122
rect 12143 4161 12177 4195
rect 11980 4035 12014 4069
rect 12123 4065 12157 4099
rect 12342 4149 12376 4183
rect 12232 3987 12266 4021
rect 12585 4161 12619 4195
rect 12406 4053 12440 4087
rect 12542 4053 12576 4087
rect 12853 4103 12887 4137
rect 13037 4103 13071 4137
rect 13507 4077 13541 4111
rect 13871 4113 13905 4147
rect 14611 4077 14645 4111
rect 14975 4113 15009 4147
rect 15541 4090 15575 4124
rect 15661 4103 15695 4137
rect 12644 3987 12678 4021
rect 12780 3987 12814 4021
rect 15827 4077 15861 4111
rect 15926 4077 15960 4111
rect 16025 4077 16059 4111
rect 16133 4113 16167 4147
rect 16236 4113 16270 4147
rect 16339 4113 16373 4147
rect 16910 4103 16944 4137
rect 17051 4103 17085 4137
rect 17159 4103 17193 4137
rect 17647 4077 17681 4111
rect 18011 4113 18045 4147
rect 18651 4117 18685 4151
rect 18759 4077 18793 4111
rect 1171 3505 1205 3539
rect 1279 3465 1313 3499
rect 1475 3505 1509 3539
rect 1585 3505 1619 3539
rect 1693 3469 1727 3503
rect 1803 3469 1837 3503
rect 2056 3479 2090 3513
rect 2320 3547 2354 3581
rect 2572 3595 2606 3629
rect 2158 3494 2192 3528
rect 2463 3517 2497 3551
rect 2483 3421 2517 3455
rect 2984 3595 3018 3629
rect 3120 3595 3154 3629
rect 2746 3529 2780 3563
rect 2882 3529 2916 3563
rect 2682 3433 2716 3467
rect 2925 3421 2959 3455
rect 3193 3479 3227 3513
rect 3377 3479 3411 3513
rect 3988 3479 4022 3513
rect 4252 3547 4286 3581
rect 4504 3595 4538 3629
rect 4090 3494 4124 3528
rect 4395 3517 4429 3551
rect 4415 3421 4449 3455
rect 4916 3595 4950 3629
rect 5052 3595 5086 3629
rect 4678 3529 4712 3563
rect 4814 3529 4848 3563
rect 4614 3433 4648 3467
rect 4857 3421 4891 3455
rect 5125 3479 5159 3513
rect 5309 3479 5343 3513
rect 5523 3505 5557 3539
rect 5622 3505 5656 3539
rect 5721 3505 5755 3539
rect 5829 3469 5863 3503
rect 5932 3469 5966 3503
rect 6035 3469 6069 3503
rect 6375 3479 6409 3513
rect 6513 3479 6547 3513
rect 6613 3479 6647 3513
rect 6741 3479 6775 3513
rect 6845 3505 6879 3539
rect 7105 3469 7139 3503
rect 7208 3479 7242 3513
rect 7472 3547 7506 3581
rect 7724 3595 7758 3629
rect 7310 3494 7344 3528
rect 7615 3517 7649 3551
rect 7635 3421 7669 3455
rect 8136 3595 8170 3629
rect 8272 3595 8306 3629
rect 7898 3529 7932 3563
rect 8034 3529 8068 3563
rect 7834 3433 7868 3467
rect 8077 3421 8111 3455
rect 8345 3479 8379 3513
rect 8529 3479 8563 3513
rect 9019 3505 9053 3539
rect 9118 3505 9152 3539
rect 9217 3505 9251 3539
rect 9325 3469 9359 3503
rect 9428 3469 9462 3503
rect 9531 3469 9565 3503
rect 9784 3479 9818 3513
rect 10048 3547 10082 3581
rect 10300 3595 10334 3629
rect 9886 3494 9920 3528
rect 10191 3517 10225 3551
rect 10211 3421 10245 3455
rect 10712 3595 10746 3629
rect 10848 3595 10882 3629
rect 10474 3529 10508 3563
rect 10610 3529 10644 3563
rect 10410 3433 10444 3467
rect 10653 3421 10687 3455
rect 10921 3479 10955 3513
rect 11105 3479 11139 3513
rect 11319 3505 11353 3539
rect 11429 3505 11463 3539
rect 11537 3469 11571 3503
rect 11647 3469 11681 3503
rect 11808 3479 11842 3513
rect 12072 3547 12106 3581
rect 12324 3595 12358 3629
rect 11910 3494 11944 3528
rect 12215 3517 12249 3551
rect 12235 3421 12269 3455
rect 12736 3595 12770 3629
rect 12872 3595 12906 3629
rect 12498 3529 12532 3563
rect 12634 3529 12668 3563
rect 12434 3433 12468 3467
rect 12677 3421 12711 3455
rect 12945 3479 12979 3513
rect 13129 3479 13163 3513
rect 13343 3505 13377 3539
rect 13442 3505 13476 3539
rect 13541 3505 13575 3539
rect 13649 3469 13683 3503
rect 13752 3469 13786 3503
rect 13855 3469 13889 3503
rect 14427 3505 14461 3539
rect 14791 3469 14825 3503
rect 15275 3505 15309 3539
rect 15385 3505 15419 3539
rect 15493 3469 15527 3503
rect 15603 3469 15637 3503
rect 15817 3492 15851 3526
rect 15937 3479 15971 3513
rect 16045 3505 16079 3539
rect 16305 3469 16339 3503
rect 16479 3479 16513 3513
rect 16587 3479 16621 3513
rect 16728 3479 16762 3513
rect 16873 3505 16907 3539
rect 17133 3469 17167 3503
rect 17307 3479 17341 3513
rect 17415 3479 17449 3513
rect 17556 3479 17590 3513
rect 17759 3505 17793 3539
rect 17858 3505 17892 3539
rect 17957 3505 17991 3539
rect 18065 3469 18099 3503
rect 18168 3469 18202 3503
rect 18271 3469 18305 3503
rect 18651 3465 18685 3499
rect 18759 3505 18793 3539
rect 1171 2989 1205 3023
rect 1279 3029 1313 3063
rect 1417 2989 1451 3023
rect 1677 3025 1711 3059
rect 1929 3015 1963 3049
rect 2033 3015 2067 3049
rect 2245 2989 2279 3023
rect 2505 3025 2539 3059
rect 2898 3015 2932 3049
rect 2966 3015 3000 3049
rect 3034 3015 3068 3049
rect 3102 3015 3136 3049
rect 3170 3015 3204 3049
rect 3238 3015 3272 3049
rect 3306 3015 3340 3049
rect 3374 3015 3408 3049
rect 3442 3015 3476 3049
rect 3510 3015 3544 3049
rect 3578 3015 3612 3049
rect 3646 3015 3680 3049
rect 3714 3015 3748 3049
rect 3782 3015 3816 3049
rect 3850 3015 3884 3049
rect 3918 3015 3952 3049
rect 4345 3015 4379 3049
rect 4767 2989 4801 3023
rect 5131 3025 5165 3059
rect 5615 2989 5649 3023
rect 5714 2989 5748 3023
rect 5813 2989 5847 3023
rect 5921 3025 5955 3059
rect 6024 3025 6058 3059
rect 6127 3025 6161 3059
rect 6443 2989 6477 3023
rect 6542 2989 6576 3023
rect 6641 2989 6675 3023
rect 6749 3025 6783 3059
rect 6852 3025 6886 3059
rect 6955 3025 6989 3059
rect 7397 2989 7431 3023
rect 7657 3025 7691 3059
rect 7765 3015 7799 3049
rect 8192 3015 8226 3049
rect 8260 3015 8294 3049
rect 8328 3015 8362 3049
rect 8396 3015 8430 3049
rect 8464 3015 8498 3049
rect 8532 3015 8566 3049
rect 8600 3015 8634 3049
rect 8668 3015 8702 3049
rect 8736 3015 8770 3049
rect 8804 3015 8838 3049
rect 8872 3015 8906 3049
rect 8940 3015 8974 3049
rect 9008 3015 9042 3049
rect 9076 3015 9110 3049
rect 9144 3015 9178 3049
rect 9212 3015 9246 3049
rect 9919 2989 9953 3023
rect 10283 3025 10317 3059
rect 10767 2989 10801 3023
rect 10866 2989 10900 3023
rect 10965 2989 10999 3023
rect 11073 3025 11107 3059
rect 11176 3025 11210 3059
rect 11279 3025 11313 3059
rect 11716 3015 11750 3049
rect 11818 3000 11852 3034
rect 12143 3073 12177 3107
rect 11980 2947 12014 2981
rect 12123 2977 12157 3011
rect 12342 3061 12376 3095
rect 12232 2899 12266 2933
rect 12585 3073 12619 3107
rect 12406 2965 12440 2999
rect 12542 2965 12576 2999
rect 12853 3015 12887 3049
rect 13037 3015 13071 3049
rect 13507 2989 13541 3023
rect 13871 3025 13905 3059
rect 14611 2989 14645 3023
rect 14975 3025 15009 3059
rect 15715 2989 15749 3023
rect 16079 3025 16113 3059
rect 16921 3002 16955 3036
rect 17041 3015 17075 3049
rect 12644 2899 12678 2933
rect 12780 2899 12814 2933
rect 17463 2989 17497 3023
rect 17827 3025 17861 3059
rect 18253 2989 18287 3023
rect 18513 3025 18547 3059
rect 18651 3029 18685 3063
rect 18759 2989 18793 3023
rect 2366 2507 2400 2541
rect 2502 2507 2536 2541
rect 1171 2417 1205 2451
rect 1279 2377 1313 2411
rect 1475 2417 1509 2451
rect 1585 2417 1619 2451
rect 1693 2381 1727 2415
rect 1803 2381 1837 2415
rect 2109 2391 2143 2425
rect 2293 2391 2327 2425
rect 2604 2441 2638 2475
rect 2740 2441 2774 2475
rect 2561 2333 2595 2367
rect 2914 2507 2948 2541
rect 2804 2345 2838 2379
rect 3023 2429 3057 2463
rect 3166 2459 3200 2493
rect 3003 2333 3037 2367
rect 3328 2406 3362 2440
rect 3430 2391 3464 2425
rect 4177 2417 4211 2451
rect 4437 2381 4471 2415
rect 4632 2391 4666 2425
rect 4896 2459 4930 2493
rect 5148 2507 5182 2541
rect 4734 2406 4768 2440
rect 5039 2429 5073 2463
rect 5059 2333 5093 2367
rect 5560 2507 5594 2541
rect 5696 2507 5730 2541
rect 5322 2441 5356 2475
rect 5458 2441 5492 2475
rect 5258 2345 5292 2379
rect 5501 2333 5535 2367
rect 7518 2507 7552 2541
rect 7654 2507 7688 2541
rect 5769 2391 5803 2425
rect 5953 2391 5987 2425
rect 6443 2417 6477 2451
rect 6542 2417 6576 2451
rect 6641 2417 6675 2451
rect 6749 2381 6783 2415
rect 6852 2381 6886 2415
rect 6955 2381 6989 2415
rect 7261 2391 7295 2425
rect 7445 2391 7479 2425
rect 7756 2441 7790 2475
rect 7892 2441 7926 2475
rect 7713 2333 7747 2367
rect 8066 2507 8100 2541
rect 7956 2345 7990 2379
rect 8175 2429 8209 2463
rect 8318 2459 8352 2493
rect 8155 2333 8189 2367
rect 8480 2406 8514 2440
rect 8582 2391 8616 2425
rect 9019 2417 9053 2451
rect 9118 2417 9152 2451
rect 9217 2417 9251 2451
rect 9325 2381 9359 2415
rect 9428 2381 9462 2415
rect 9531 2381 9565 2415
rect 9784 2391 9818 2425
rect 10048 2459 10082 2493
rect 10300 2507 10334 2541
rect 9886 2406 9920 2440
rect 10191 2429 10225 2463
rect 10211 2333 10245 2367
rect 10712 2507 10746 2541
rect 10848 2507 10882 2541
rect 10474 2441 10508 2475
rect 10610 2441 10644 2475
rect 10410 2345 10444 2379
rect 10653 2333 10687 2367
rect 12210 2507 12244 2541
rect 12346 2507 12380 2541
rect 10921 2391 10955 2425
rect 11105 2391 11139 2425
rect 11537 2417 11571 2451
rect 11797 2381 11831 2415
rect 11953 2391 11987 2425
rect 12137 2391 12171 2425
rect 12448 2441 12482 2475
rect 12584 2441 12618 2475
rect 12405 2333 12439 2367
rect 12758 2507 12792 2541
rect 12648 2345 12682 2379
rect 12867 2429 12901 2463
rect 13010 2459 13044 2493
rect 12847 2333 12881 2367
rect 13172 2406 13206 2440
rect 14331 2626 14365 2660
rect 14331 2558 14365 2592
rect 13274 2391 13308 2425
rect 13435 2417 13469 2451
rect 13545 2417 13579 2451
rect 13653 2381 13687 2415
rect 13763 2381 13797 2415
rect 14331 2291 14365 2325
rect 14331 2223 14365 2257
rect 14431 2626 14465 2660
rect 14431 2558 14465 2592
rect 14887 2417 14921 2451
rect 15251 2381 15285 2415
rect 15735 2417 15769 2451
rect 15834 2417 15868 2451
rect 15933 2417 15967 2451
rect 16041 2381 16075 2415
rect 16144 2381 16178 2415
rect 16247 2381 16281 2415
rect 16921 2404 16955 2438
rect 17041 2391 17075 2425
rect 17149 2417 17183 2451
rect 14431 2295 14465 2329
rect 14431 2227 14465 2261
rect 17409 2381 17443 2415
rect 17517 2391 17551 2425
rect 17641 2391 17675 2425
rect 17943 2417 17977 2451
rect 18042 2417 18076 2451
rect 18141 2417 18175 2451
rect 18249 2381 18283 2415
rect 18352 2381 18386 2415
rect 18455 2381 18489 2415
rect 18651 2377 18685 2411
rect 18759 2417 18793 2451
<< rmp >>
rect 14281 2408 14377 2417
rect 14419 2408 14515 2417
<< ndiode >>
rect 9503 7559 9629 7577
rect 9503 7525 9511 7559
rect 9545 7525 9586 7559
rect 9620 7525 9629 7559
rect 9503 7491 9629 7525
rect 9503 7457 9511 7491
rect 9545 7457 9586 7491
rect 9620 7457 9629 7491
rect 9503 7439 9629 7457
rect 7203 3207 7329 3225
rect 7203 3173 7211 3207
rect 7245 3173 7286 3207
rect 7320 3173 7329 3207
rect 7203 3139 7329 3173
rect 7203 3105 7211 3139
rect 7245 3105 7286 3139
rect 7320 3105 7329 3139
rect 7203 3087 7329 3105
rect 3983 2335 4109 2353
rect 3983 2301 3991 2335
rect 4025 2301 4066 2335
rect 4100 2301 4109 2335
rect 3983 2267 4109 2301
rect 3983 2233 3991 2267
rect 4025 2233 4066 2267
rect 4100 2233 4109 2267
rect 3983 2215 4109 2233
<< ndiodec >>
rect 9511 7525 9545 7559
rect 9586 7525 9620 7559
rect 9511 7457 9545 7491
rect 9586 7457 9620 7491
rect 7211 3173 7245 3207
rect 7286 3173 7320 3207
rect 7211 3105 7245 3139
rect 7286 3105 7320 3139
rect 3991 2301 4025 2335
rect 4066 2301 4100 2335
rect 3991 2233 4025 2267
rect 4066 2233 4100 2267
<< locali >>
rect 1104 7599 1133 7633
rect 1167 7599 1225 7633
rect 1259 7599 1317 7633
rect 1351 7599 1409 7633
rect 1443 7599 1501 7633
rect 1535 7599 1593 7633
rect 1627 7599 1685 7633
rect 1719 7599 1777 7633
rect 1811 7599 1869 7633
rect 1903 7599 1961 7633
rect 1995 7599 2053 7633
rect 2087 7599 2145 7633
rect 2179 7599 2237 7633
rect 2271 7599 2329 7633
rect 2363 7599 2421 7633
rect 2455 7599 2513 7633
rect 2547 7599 2605 7633
rect 2639 7599 2697 7633
rect 2731 7599 2789 7633
rect 2823 7599 2881 7633
rect 2915 7599 2973 7633
rect 3007 7599 3065 7633
rect 3099 7599 3157 7633
rect 3191 7599 3249 7633
rect 3283 7599 3341 7633
rect 3375 7599 3433 7633
rect 3467 7599 3525 7633
rect 3559 7599 3617 7633
rect 3651 7599 3709 7633
rect 3743 7599 3801 7633
rect 3835 7599 3893 7633
rect 3927 7599 3985 7633
rect 4019 7599 4077 7633
rect 4111 7599 4169 7633
rect 4203 7599 4261 7633
rect 4295 7599 4353 7633
rect 4387 7599 4445 7633
rect 4479 7599 4537 7633
rect 4571 7599 4629 7633
rect 4663 7599 4721 7633
rect 4755 7599 4813 7633
rect 4847 7599 4905 7633
rect 4939 7599 4997 7633
rect 5031 7599 5089 7633
rect 5123 7599 5181 7633
rect 5215 7599 5273 7633
rect 5307 7599 5365 7633
rect 5399 7599 5457 7633
rect 5491 7599 5549 7633
rect 5583 7599 5641 7633
rect 5675 7599 5733 7633
rect 5767 7599 5825 7633
rect 5859 7599 5917 7633
rect 5951 7599 6009 7633
rect 6043 7599 6101 7633
rect 6135 7599 6193 7633
rect 6227 7599 6285 7633
rect 6319 7599 6377 7633
rect 6411 7599 6469 7633
rect 6503 7599 6561 7633
rect 6595 7599 6653 7633
rect 6687 7599 6745 7633
rect 6779 7599 6837 7633
rect 6871 7599 6929 7633
rect 6963 7599 7021 7633
rect 7055 7599 7113 7633
rect 7147 7599 7205 7633
rect 7239 7599 7297 7633
rect 7331 7599 7389 7633
rect 7423 7599 7481 7633
rect 7515 7599 7573 7633
rect 7607 7599 7665 7633
rect 7699 7599 7757 7633
rect 7791 7599 7849 7633
rect 7883 7599 7941 7633
rect 7975 7599 8033 7633
rect 8067 7599 8125 7633
rect 8159 7599 8217 7633
rect 8251 7599 8309 7633
rect 8343 7599 8401 7633
rect 8435 7599 8493 7633
rect 8527 7599 8585 7633
rect 8619 7599 8677 7633
rect 8711 7599 8769 7633
rect 8803 7599 8861 7633
rect 8895 7599 8953 7633
rect 8987 7599 9045 7633
rect 9079 7599 9137 7633
rect 9171 7599 9229 7633
rect 9263 7599 9321 7633
rect 9355 7599 9413 7633
rect 9447 7599 9505 7633
rect 9539 7599 9597 7633
rect 9631 7599 9689 7633
rect 9723 7599 9781 7633
rect 9815 7599 9873 7633
rect 9907 7599 9965 7633
rect 9999 7599 10057 7633
rect 10091 7599 10149 7633
rect 10183 7599 10241 7633
rect 10275 7599 10333 7633
rect 10367 7599 10425 7633
rect 10459 7599 10517 7633
rect 10551 7599 10609 7633
rect 10643 7599 10701 7633
rect 10735 7599 10793 7633
rect 10827 7599 10885 7633
rect 10919 7599 10977 7633
rect 11011 7599 11069 7633
rect 11103 7599 11161 7633
rect 11195 7599 11253 7633
rect 11287 7599 11345 7633
rect 11379 7599 11437 7633
rect 11471 7599 11529 7633
rect 11563 7599 11621 7633
rect 11655 7599 11713 7633
rect 11747 7599 11805 7633
rect 11839 7599 11897 7633
rect 11931 7599 11989 7633
rect 12023 7599 12081 7633
rect 12115 7599 12173 7633
rect 12207 7599 12265 7633
rect 12299 7599 12357 7633
rect 12391 7599 12449 7633
rect 12483 7599 12541 7633
rect 12575 7599 12633 7633
rect 12667 7599 12725 7633
rect 12759 7599 12817 7633
rect 12851 7599 12909 7633
rect 12943 7599 13001 7633
rect 13035 7599 13093 7633
rect 13127 7599 13185 7633
rect 13219 7599 13277 7633
rect 13311 7599 13369 7633
rect 13403 7599 13461 7633
rect 13495 7599 13553 7633
rect 13587 7599 13645 7633
rect 13679 7599 13737 7633
rect 13771 7599 13829 7633
rect 13863 7599 13921 7633
rect 13955 7599 14013 7633
rect 14047 7599 14105 7633
rect 14139 7599 14197 7633
rect 14231 7599 14289 7633
rect 14323 7599 14381 7633
rect 14415 7599 14473 7633
rect 14507 7599 14565 7633
rect 14599 7599 14657 7633
rect 14691 7599 14749 7633
rect 14783 7599 14841 7633
rect 14875 7599 14933 7633
rect 14967 7599 15025 7633
rect 15059 7599 15117 7633
rect 15151 7599 15209 7633
rect 15243 7599 15301 7633
rect 15335 7599 15393 7633
rect 15427 7599 15485 7633
rect 15519 7599 15577 7633
rect 15611 7599 15669 7633
rect 15703 7599 15761 7633
rect 15795 7599 15853 7633
rect 15887 7599 15945 7633
rect 15979 7599 16037 7633
rect 16071 7599 16129 7633
rect 16163 7599 16221 7633
rect 16255 7599 16313 7633
rect 16347 7599 16405 7633
rect 16439 7599 16497 7633
rect 16531 7599 16589 7633
rect 16623 7599 16681 7633
rect 16715 7599 16773 7633
rect 16807 7599 16865 7633
rect 16899 7599 16957 7633
rect 16991 7599 17049 7633
rect 17083 7599 17141 7633
rect 17175 7599 17233 7633
rect 17267 7599 17325 7633
rect 17359 7599 17417 7633
rect 17451 7599 17509 7633
rect 17543 7599 17601 7633
rect 17635 7599 17693 7633
rect 17727 7599 17785 7633
rect 17819 7599 17877 7633
rect 17911 7599 17969 7633
rect 18003 7599 18061 7633
rect 18095 7599 18153 7633
rect 18187 7599 18245 7633
rect 18279 7599 18337 7633
rect 18371 7599 18429 7633
rect 18463 7599 18521 7633
rect 18555 7599 18613 7633
rect 18647 7599 18705 7633
rect 18739 7599 18797 7633
rect 18831 7599 18860 7633
rect 1121 7536 1363 7599
rect 1121 7502 1139 7536
rect 1173 7502 1311 7536
rect 1345 7502 1363 7536
rect 1121 7449 1363 7502
rect 1582 7553 1634 7599
rect 1582 7519 1600 7553
rect 1582 7485 1634 7519
rect 1582 7451 1600 7485
rect 1121 7375 1225 7449
rect 1582 7431 1634 7451
rect 1669 7531 1720 7565
rect 1669 7527 1685 7531
rect 1669 7493 1684 7527
rect 1719 7497 1720 7531
rect 1754 7557 1820 7599
rect 1754 7523 1770 7557
rect 1804 7523 1820 7557
rect 1863 7544 1897 7565
rect 1718 7493 1720 7497
rect 1669 7450 1720 7493
rect 1863 7489 1897 7510
rect 1949 7538 3018 7599
rect 1949 7504 1967 7538
rect 2001 7504 2967 7538
rect 3001 7504 3018 7538
rect 1949 7490 3018 7504
rect 3053 7538 3571 7599
rect 3053 7504 3071 7538
rect 3105 7504 3519 7538
rect 3553 7504 3571 7538
rect 1754 7455 1897 7489
rect 1121 7341 1171 7375
rect 1205 7341 1225 7375
rect 1259 7381 1279 7415
rect 1313 7381 1363 7415
rect 1259 7307 1363 7381
rect 1121 7260 1363 7307
rect 1121 7226 1139 7260
rect 1173 7226 1311 7260
rect 1345 7226 1363 7260
rect 1121 7165 1363 7226
rect 1121 7131 1139 7165
rect 1173 7131 1311 7165
rect 1345 7131 1363 7165
rect 1121 7089 1363 7131
rect 1582 7301 1634 7319
rect 1582 7267 1600 7301
rect 1582 7233 1634 7267
rect 1582 7199 1600 7233
rect 1582 7165 1634 7199
rect 1582 7131 1600 7165
rect 1582 7089 1634 7131
rect 1669 7304 1703 7450
rect 1754 7417 1788 7455
rect 1737 7401 1788 7417
rect 1771 7367 1788 7401
rect 1737 7351 1788 7367
rect 1754 7309 1788 7351
rect 1844 7401 1915 7419
rect 1844 7367 1861 7401
rect 1895 7395 1915 7401
rect 1844 7361 1869 7367
rect 1903 7361 1915 7395
rect 1844 7345 1915 7361
rect 2266 7375 2334 7490
rect 3053 7445 3571 7504
rect 3697 7505 3755 7599
rect 3697 7471 3709 7505
rect 3743 7471 3755 7505
rect 3697 7454 3755 7471
rect 3974 7553 4026 7599
rect 3974 7519 3992 7553
rect 3974 7485 4026 7519
rect 3974 7451 3992 7485
rect 2266 7341 2283 7375
rect 2317 7341 2334 7375
rect 2266 7324 2334 7341
rect 2630 7411 2700 7426
rect 2630 7377 2647 7411
rect 2681 7377 2700 7411
rect 1669 7270 1720 7304
rect 1754 7275 1897 7309
rect 1669 7236 1684 7270
rect 1718 7236 1720 7270
rect 1863 7241 1897 7275
rect 1669 7189 1720 7236
rect 1669 7155 1684 7189
rect 1718 7155 1720 7189
rect 1669 7123 1720 7155
rect 1754 7207 1770 7241
rect 1804 7207 1820 7241
rect 1754 7173 1820 7207
rect 1754 7139 1770 7173
rect 1804 7139 1820 7173
rect 1754 7089 1820 7139
rect 1863 7173 1897 7207
rect 2630 7176 2700 7377
rect 3053 7375 3295 7445
rect 3974 7431 4026 7451
rect 4061 7531 4112 7565
rect 4061 7527 4077 7531
rect 4061 7493 4076 7527
rect 4111 7497 4112 7531
rect 4146 7557 4212 7599
rect 4146 7523 4162 7557
rect 4196 7523 4212 7557
rect 4255 7544 4289 7565
rect 4110 7493 4112 7497
rect 4061 7450 4112 7493
rect 4255 7489 4289 7510
rect 4341 7538 5410 7599
rect 4341 7504 4359 7538
rect 4393 7504 5359 7538
rect 5393 7504 5410 7538
rect 4341 7490 5410 7504
rect 5630 7553 5682 7599
rect 5630 7519 5648 7553
rect 4146 7455 4289 7489
rect 3053 7341 3131 7375
rect 3165 7341 3241 7375
rect 3275 7341 3295 7375
rect 3329 7377 3349 7411
rect 3383 7377 3459 7411
rect 3493 7377 3571 7411
rect 3329 7307 3571 7377
rect 3053 7267 3571 7307
rect 3053 7233 3071 7267
rect 3105 7233 3519 7267
rect 3553 7233 3571 7267
rect 1863 7123 1897 7139
rect 1949 7165 3018 7176
rect 1949 7131 1967 7165
rect 2001 7131 2967 7165
rect 3001 7131 3018 7165
rect 1949 7089 3018 7131
rect 3053 7165 3571 7233
rect 3053 7131 3071 7165
rect 3105 7131 3519 7165
rect 3553 7131 3571 7165
rect 3053 7089 3571 7131
rect 3697 7287 3755 7322
rect 3697 7253 3709 7287
rect 3743 7253 3755 7287
rect 3697 7194 3755 7253
rect 3697 7160 3709 7194
rect 3743 7160 3755 7194
rect 3697 7089 3755 7160
rect 3974 7301 4026 7319
rect 3974 7267 3992 7301
rect 3974 7233 4026 7267
rect 3974 7199 3992 7233
rect 3974 7165 4026 7199
rect 3974 7131 3992 7165
rect 3974 7089 4026 7131
rect 4061 7304 4095 7450
rect 4146 7417 4180 7455
rect 4129 7401 4180 7417
rect 4163 7367 4180 7401
rect 4129 7351 4180 7367
rect 4146 7309 4180 7351
rect 4236 7401 4307 7419
rect 4236 7367 4253 7401
rect 4287 7395 4307 7401
rect 4236 7361 4261 7367
rect 4295 7361 4307 7395
rect 4236 7345 4307 7361
rect 4658 7375 4726 7490
rect 5630 7485 5682 7519
rect 5630 7451 5648 7485
rect 5630 7431 5682 7451
rect 5717 7531 5768 7565
rect 5717 7527 5733 7531
rect 5717 7493 5732 7527
rect 5767 7497 5768 7531
rect 5802 7557 5868 7599
rect 5802 7523 5818 7557
rect 5852 7523 5868 7557
rect 5911 7544 5945 7565
rect 5766 7493 5768 7497
rect 5717 7450 5768 7493
rect 5911 7489 5945 7510
rect 5802 7455 5945 7489
rect 5997 7536 6239 7599
rect 5997 7502 6015 7536
rect 6049 7502 6187 7536
rect 6221 7502 6239 7536
rect 4658 7341 4675 7375
rect 4709 7341 4726 7375
rect 4658 7324 4726 7341
rect 5022 7411 5092 7426
rect 5022 7377 5039 7411
rect 5073 7377 5092 7411
rect 4061 7270 4112 7304
rect 4146 7275 4289 7309
rect 4061 7236 4076 7270
rect 4110 7236 4112 7270
rect 4255 7241 4289 7275
rect 4061 7189 4112 7236
rect 4061 7155 4076 7189
rect 4110 7155 4112 7189
rect 4061 7123 4112 7155
rect 4146 7207 4162 7241
rect 4196 7207 4212 7241
rect 4146 7173 4212 7207
rect 4146 7139 4162 7173
rect 4196 7139 4212 7173
rect 4146 7089 4212 7139
rect 4255 7173 4289 7207
rect 5022 7176 5092 7377
rect 5630 7301 5682 7319
rect 5630 7267 5648 7301
rect 5630 7233 5682 7267
rect 5630 7199 5648 7233
rect 4255 7123 4289 7139
rect 4341 7165 5410 7176
rect 4341 7131 4359 7165
rect 4393 7131 5359 7165
rect 5393 7131 5410 7165
rect 4341 7089 5410 7131
rect 5630 7165 5682 7199
rect 5630 7131 5648 7165
rect 5630 7089 5682 7131
rect 5717 7304 5751 7450
rect 5802 7417 5836 7455
rect 5997 7449 6239 7502
rect 6273 7505 6331 7599
rect 6273 7471 6285 7505
rect 6319 7471 6331 7505
rect 6365 7538 7434 7599
rect 6365 7504 6383 7538
rect 6417 7504 7383 7538
rect 7417 7504 7434 7538
rect 6365 7490 7434 7504
rect 7469 7531 7803 7599
rect 7469 7497 7487 7531
rect 7521 7497 7751 7531
rect 7785 7497 7803 7531
rect 6273 7454 6331 7471
rect 5785 7401 5836 7417
rect 5819 7367 5836 7401
rect 5785 7351 5836 7367
rect 5802 7309 5836 7351
rect 5892 7401 5963 7419
rect 5892 7367 5909 7401
rect 5943 7395 5963 7401
rect 5892 7361 5917 7367
rect 5951 7361 5963 7395
rect 5892 7345 5963 7361
rect 5997 7375 6101 7449
rect 5997 7341 6047 7375
rect 6081 7341 6101 7375
rect 6135 7381 6155 7415
rect 6189 7381 6239 7415
rect 5717 7270 5768 7304
rect 5802 7275 5945 7309
rect 6135 7307 6239 7381
rect 6682 7375 6750 7490
rect 7469 7445 7803 7497
rect 7855 7544 7889 7565
rect 7932 7557 7998 7599
rect 7932 7523 7948 7557
rect 7982 7523 7998 7557
rect 8032 7531 8083 7565
rect 7855 7489 7889 7510
rect 8032 7497 8033 7531
rect 8067 7527 8083 7531
rect 8032 7493 8034 7497
rect 8068 7493 8083 7527
rect 7855 7455 7998 7489
rect 6682 7341 6699 7375
rect 6733 7341 6750 7375
rect 6682 7324 6750 7341
rect 7046 7411 7116 7426
rect 7046 7377 7063 7411
rect 7097 7377 7116 7411
rect 5717 7236 5732 7270
rect 5766 7236 5768 7270
rect 5911 7241 5945 7275
rect 5717 7189 5768 7236
rect 5717 7155 5732 7189
rect 5766 7155 5768 7189
rect 5717 7123 5768 7155
rect 5802 7207 5818 7241
rect 5852 7207 5868 7241
rect 5802 7173 5868 7207
rect 5802 7139 5818 7173
rect 5852 7139 5868 7173
rect 5802 7089 5868 7139
rect 5911 7173 5945 7207
rect 5911 7123 5945 7139
rect 5997 7260 6239 7307
rect 5997 7226 6015 7260
rect 6049 7226 6187 7260
rect 6221 7226 6239 7260
rect 5997 7165 6239 7226
rect 5997 7131 6015 7165
rect 6049 7131 6187 7165
rect 6221 7131 6239 7165
rect 5997 7089 6239 7131
rect 6273 7287 6331 7322
rect 6273 7253 6285 7287
rect 6319 7253 6331 7287
rect 6273 7194 6331 7253
rect 6273 7160 6285 7194
rect 6319 7160 6331 7194
rect 7046 7176 7116 7377
rect 7469 7375 7619 7445
rect 7469 7341 7489 7375
rect 7523 7341 7619 7375
rect 7653 7377 7749 7411
rect 7783 7377 7803 7411
rect 7653 7307 7803 7377
rect 7837 7401 7908 7419
rect 7837 7395 7857 7401
rect 7837 7361 7849 7395
rect 7891 7367 7908 7401
rect 7883 7361 7908 7367
rect 7837 7345 7908 7361
rect 7964 7417 7998 7455
rect 8032 7450 8083 7493
rect 7964 7401 8015 7417
rect 7964 7367 7981 7401
rect 7964 7351 8015 7367
rect 7964 7309 7998 7351
rect 7469 7267 7803 7307
rect 7469 7233 7487 7267
rect 7521 7233 7751 7267
rect 7785 7233 7803 7267
rect 6273 7089 6331 7160
rect 6365 7165 7434 7176
rect 6365 7131 6383 7165
rect 6417 7131 7383 7165
rect 7417 7131 7434 7165
rect 6365 7089 7434 7131
rect 7469 7165 7803 7233
rect 7469 7131 7487 7165
rect 7521 7131 7751 7165
rect 7785 7131 7803 7165
rect 7469 7089 7803 7131
rect 7855 7275 7998 7309
rect 8049 7304 8083 7450
rect 8118 7553 8170 7599
rect 8152 7519 8170 7553
rect 8118 7485 8170 7519
rect 8152 7451 8170 7485
rect 8118 7431 8170 7451
rect 8205 7538 8723 7599
rect 8205 7504 8223 7538
rect 8257 7504 8671 7538
rect 8705 7504 8723 7538
rect 8205 7445 8723 7504
rect 8849 7505 8907 7599
rect 8849 7471 8861 7505
rect 8895 7471 8907 7505
rect 8849 7454 8907 7471
rect 8941 7538 9459 7599
rect 8941 7504 8959 7538
rect 8993 7504 9407 7538
rect 9441 7504 9459 7538
rect 8941 7445 9459 7504
rect 9493 7559 9643 7565
rect 9493 7525 9511 7559
rect 9545 7525 9586 7559
rect 9620 7525 9643 7559
rect 9493 7491 9643 7525
rect 9493 7457 9511 7491
rect 9545 7457 9586 7491
rect 9620 7463 9643 7491
rect 8205 7375 8447 7445
rect 8205 7341 8283 7375
rect 8317 7341 8393 7375
rect 8427 7341 8447 7375
rect 8481 7377 8501 7411
rect 8535 7377 8611 7411
rect 8645 7377 8723 7411
rect 7855 7241 7889 7275
rect 8032 7270 8083 7304
rect 7855 7173 7889 7207
rect 7855 7123 7889 7139
rect 7932 7207 7948 7241
rect 7982 7207 7998 7241
rect 7932 7173 7998 7207
rect 7932 7139 7948 7173
rect 7982 7139 7998 7173
rect 7932 7089 7998 7139
rect 8032 7236 8034 7270
rect 8068 7236 8083 7270
rect 8032 7189 8083 7236
rect 8032 7155 8034 7189
rect 8068 7155 8083 7189
rect 8032 7123 8083 7155
rect 8118 7301 8170 7319
rect 8481 7307 8723 7377
rect 8941 7375 9183 7445
rect 9493 7429 9597 7457
rect 9631 7429 9643 7463
rect 8941 7341 9019 7375
rect 9053 7341 9129 7375
rect 9163 7341 9183 7375
rect 9217 7377 9237 7411
rect 9271 7377 9347 7411
rect 9381 7377 9459 7411
rect 8152 7267 8170 7301
rect 8118 7233 8170 7267
rect 8152 7199 8170 7233
rect 8118 7165 8170 7199
rect 8152 7131 8170 7165
rect 8118 7089 8170 7131
rect 8205 7267 8723 7307
rect 8205 7233 8223 7267
rect 8257 7233 8671 7267
rect 8705 7233 8723 7267
rect 8205 7165 8723 7233
rect 8205 7131 8223 7165
rect 8257 7131 8671 7165
rect 8705 7131 8723 7165
rect 8205 7089 8723 7131
rect 8849 7287 8907 7322
rect 9217 7307 9459 7377
rect 8849 7253 8861 7287
rect 8895 7253 8907 7287
rect 8849 7194 8907 7253
rect 8849 7160 8861 7194
rect 8895 7160 8907 7194
rect 8849 7089 8907 7160
rect 8941 7267 9459 7307
rect 8941 7233 8959 7267
rect 8993 7233 9407 7267
rect 9441 7233 9459 7267
rect 8941 7165 9459 7233
rect 8941 7131 8959 7165
rect 8993 7131 9407 7165
rect 9441 7131 9459 7165
rect 8941 7089 9459 7131
rect 9493 7123 9643 7429
rect 9677 7531 10011 7599
rect 9677 7497 9695 7531
rect 9729 7497 9959 7531
rect 9993 7497 10011 7531
rect 9677 7445 10011 7497
rect 10045 7549 10097 7565
rect 10045 7515 10063 7549
rect 10045 7499 10097 7515
rect 10139 7553 10194 7599
rect 10139 7519 10149 7553
rect 10183 7519 10194 7553
rect 10139 7503 10194 7519
rect 10236 7549 10277 7565
rect 10236 7515 10243 7549
rect 10311 7553 10378 7599
rect 10311 7519 10327 7553
rect 10361 7519 10378 7553
rect 10413 7538 11115 7599
rect 9677 7375 9827 7445
rect 9677 7341 9697 7375
rect 9731 7341 9827 7375
rect 9861 7377 9957 7411
rect 9991 7377 10011 7411
rect 9861 7307 10011 7377
rect 9677 7267 10011 7307
rect 9677 7233 9695 7267
rect 9729 7233 9959 7267
rect 9993 7233 10011 7267
rect 9677 7165 10011 7233
rect 9677 7131 9695 7165
rect 9729 7131 9959 7165
rect 9993 7131 10011 7165
rect 9677 7089 10011 7131
rect 10045 7317 10079 7499
rect 10236 7485 10277 7515
rect 10413 7504 10431 7538
rect 10465 7504 11063 7538
rect 11097 7504 11115 7538
rect 10113 7463 10185 7467
rect 10113 7429 10149 7463
rect 10183 7429 10185 7463
rect 10236 7451 10373 7485
rect 10113 7401 10185 7429
rect 10113 7367 10117 7401
rect 10151 7367 10185 7401
rect 10113 7351 10185 7367
rect 10221 7401 10271 7417
rect 10255 7367 10271 7401
rect 10221 7317 10271 7367
rect 10045 7284 10271 7317
rect 10045 7250 10063 7284
rect 10097 7283 10271 7284
rect 10097 7250 10099 7283
rect 10045 7179 10099 7250
rect 10305 7259 10373 7451
rect 10413 7445 11115 7504
rect 11149 7536 11391 7599
rect 11149 7502 11167 7536
rect 11201 7502 11339 7536
rect 11373 7502 11391 7536
rect 11149 7449 11391 7502
rect 11425 7505 11483 7599
rect 11425 7471 11437 7505
rect 11471 7471 11483 7505
rect 11425 7454 11483 7471
rect 11517 7538 12219 7599
rect 11517 7504 11535 7538
rect 11569 7504 12167 7538
rect 12201 7504 12219 7538
rect 10413 7375 10743 7445
rect 10413 7341 10491 7375
rect 10525 7341 10590 7375
rect 10624 7341 10689 7375
rect 10723 7341 10743 7375
rect 10777 7377 10797 7411
rect 10831 7377 10900 7411
rect 10934 7377 11003 7411
rect 11037 7377 11115 7411
rect 10777 7307 11115 7377
rect 11149 7375 11253 7449
rect 11517 7445 12219 7504
rect 12271 7544 12305 7565
rect 12348 7557 12414 7599
rect 12348 7523 12364 7557
rect 12398 7523 12414 7557
rect 12448 7531 12499 7565
rect 12271 7489 12305 7510
rect 12448 7497 12449 7531
rect 12483 7527 12499 7531
rect 12448 7493 12450 7497
rect 12484 7493 12499 7527
rect 12271 7455 12414 7489
rect 11149 7341 11199 7375
rect 11233 7341 11253 7375
rect 11287 7381 11307 7415
rect 11341 7381 11391 7415
rect 11287 7307 11391 7381
rect 11517 7375 11847 7445
rect 11517 7341 11595 7375
rect 11629 7341 11694 7375
rect 11728 7341 11793 7375
rect 11827 7341 11847 7375
rect 11881 7377 11901 7411
rect 11935 7377 12004 7411
rect 12038 7377 12107 7411
rect 12141 7377 12219 7411
rect 10305 7245 10333 7259
rect 10045 7145 10063 7179
rect 10097 7145 10099 7179
rect 10045 7129 10099 7145
rect 10133 7211 10149 7245
rect 10183 7211 10199 7245
rect 10133 7177 10199 7211
rect 10133 7143 10149 7177
rect 10183 7143 10199 7177
rect 10133 7089 10199 7143
rect 10240 7225 10333 7245
rect 10367 7225 10373 7259
rect 10240 7210 10373 7225
rect 10413 7267 11115 7307
rect 10413 7233 10431 7267
rect 10465 7233 11063 7267
rect 11097 7233 11115 7267
rect 10240 7179 10277 7210
rect 10240 7145 10243 7179
rect 10240 7129 10277 7145
rect 10311 7140 10327 7174
rect 10361 7140 10378 7174
rect 10311 7089 10378 7140
rect 10413 7165 11115 7233
rect 10413 7131 10431 7165
rect 10465 7131 11063 7165
rect 11097 7131 11115 7165
rect 10413 7089 11115 7131
rect 11149 7260 11391 7307
rect 11149 7226 11167 7260
rect 11201 7226 11339 7260
rect 11373 7226 11391 7260
rect 11149 7165 11391 7226
rect 11149 7131 11167 7165
rect 11201 7131 11339 7165
rect 11373 7131 11391 7165
rect 11149 7089 11391 7131
rect 11425 7287 11483 7322
rect 11881 7307 12219 7377
rect 12253 7401 12324 7419
rect 12253 7395 12273 7401
rect 12253 7361 12265 7395
rect 12307 7367 12324 7401
rect 12299 7361 12324 7367
rect 12253 7345 12324 7361
rect 12380 7417 12414 7455
rect 12448 7450 12499 7493
rect 12380 7401 12431 7417
rect 12380 7367 12397 7401
rect 12380 7351 12431 7367
rect 12380 7309 12414 7351
rect 11425 7253 11437 7287
rect 11471 7253 11483 7287
rect 11425 7194 11483 7253
rect 11425 7160 11437 7194
rect 11471 7160 11483 7194
rect 11425 7089 11483 7160
rect 11517 7267 12219 7307
rect 11517 7233 11535 7267
rect 11569 7233 12167 7267
rect 12201 7233 12219 7267
rect 11517 7165 12219 7233
rect 11517 7131 11535 7165
rect 11569 7131 12167 7165
rect 12201 7131 12219 7165
rect 11517 7089 12219 7131
rect 12271 7275 12414 7309
rect 12465 7304 12499 7450
rect 12534 7553 12586 7599
rect 12568 7519 12586 7553
rect 12534 7485 12586 7519
rect 12621 7538 13690 7599
rect 12621 7504 12639 7538
rect 12673 7504 13639 7538
rect 13673 7504 13690 7538
rect 12621 7490 13690 7504
rect 13725 7536 13967 7599
rect 13725 7502 13743 7536
rect 13777 7502 13915 7536
rect 13949 7502 13967 7536
rect 12568 7451 12586 7485
rect 12534 7431 12586 7451
rect 12938 7375 13006 7490
rect 13725 7449 13967 7502
rect 14001 7505 14059 7599
rect 14001 7471 14013 7505
rect 14047 7471 14059 7505
rect 14001 7454 14059 7471
rect 14093 7531 14427 7599
rect 14093 7497 14111 7531
rect 14145 7497 14375 7531
rect 14409 7497 14427 7531
rect 12938 7341 12955 7375
rect 12989 7341 13006 7375
rect 12938 7324 13006 7341
rect 13302 7411 13372 7426
rect 13302 7377 13319 7411
rect 13353 7377 13372 7411
rect 12271 7241 12305 7275
rect 12448 7270 12499 7304
rect 12271 7173 12305 7207
rect 12271 7123 12305 7139
rect 12348 7207 12364 7241
rect 12398 7207 12414 7241
rect 12348 7173 12414 7207
rect 12348 7139 12364 7173
rect 12398 7139 12414 7173
rect 12348 7089 12414 7139
rect 12448 7236 12450 7270
rect 12484 7236 12499 7270
rect 12448 7189 12499 7236
rect 12448 7155 12450 7189
rect 12484 7155 12499 7189
rect 12448 7123 12499 7155
rect 12534 7301 12586 7319
rect 12568 7267 12586 7301
rect 12534 7233 12586 7267
rect 12568 7199 12586 7233
rect 12534 7165 12586 7199
rect 13302 7176 13372 7377
rect 13725 7375 13829 7449
rect 14093 7445 14427 7497
rect 14479 7544 14513 7565
rect 14556 7557 14622 7599
rect 14556 7523 14572 7557
rect 14606 7523 14622 7557
rect 14656 7531 14707 7565
rect 14479 7489 14513 7510
rect 14656 7497 14657 7531
rect 14691 7527 14707 7531
rect 14656 7493 14658 7497
rect 14692 7493 14707 7527
rect 14479 7455 14622 7489
rect 13725 7341 13775 7375
rect 13809 7341 13829 7375
rect 13863 7381 13883 7415
rect 13917 7381 13967 7415
rect 13863 7307 13967 7381
rect 14093 7375 14243 7445
rect 14093 7341 14113 7375
rect 14147 7341 14243 7375
rect 14277 7377 14373 7411
rect 14407 7377 14427 7411
rect 13725 7260 13967 7307
rect 13725 7226 13743 7260
rect 13777 7226 13915 7260
rect 13949 7226 13967 7260
rect 12568 7131 12586 7165
rect 12534 7089 12586 7131
rect 12621 7165 13690 7176
rect 12621 7131 12639 7165
rect 12673 7131 13639 7165
rect 13673 7131 13690 7165
rect 12621 7089 13690 7131
rect 13725 7165 13967 7226
rect 13725 7131 13743 7165
rect 13777 7131 13915 7165
rect 13949 7131 13967 7165
rect 13725 7089 13967 7131
rect 14001 7287 14059 7322
rect 14277 7307 14427 7377
rect 14461 7401 14532 7419
rect 14461 7395 14481 7401
rect 14461 7361 14473 7395
rect 14515 7367 14532 7401
rect 14507 7361 14532 7367
rect 14461 7345 14532 7361
rect 14588 7417 14622 7455
rect 14656 7450 14707 7493
rect 14588 7401 14639 7417
rect 14588 7367 14605 7401
rect 14588 7351 14639 7367
rect 14588 7309 14622 7351
rect 14001 7253 14013 7287
rect 14047 7253 14059 7287
rect 14001 7194 14059 7253
rect 14001 7160 14013 7194
rect 14047 7160 14059 7194
rect 14001 7089 14059 7160
rect 14093 7267 14427 7307
rect 14093 7233 14111 7267
rect 14145 7233 14375 7267
rect 14409 7233 14427 7267
rect 14093 7165 14427 7233
rect 14093 7131 14111 7165
rect 14145 7131 14375 7165
rect 14409 7131 14427 7165
rect 14093 7089 14427 7131
rect 14479 7275 14622 7309
rect 14673 7304 14707 7450
rect 14742 7553 14794 7599
rect 14776 7519 14794 7553
rect 14742 7485 14794 7519
rect 14829 7538 15898 7599
rect 14829 7504 14847 7538
rect 14881 7504 15847 7538
rect 15881 7504 15898 7538
rect 14829 7490 15898 7504
rect 15933 7538 16451 7599
rect 15933 7504 15951 7538
rect 15985 7504 16399 7538
rect 16433 7504 16451 7538
rect 14776 7451 14794 7485
rect 14742 7431 14794 7451
rect 15146 7375 15214 7490
rect 15933 7445 16451 7504
rect 16577 7505 16635 7599
rect 16577 7471 16589 7505
rect 16623 7471 16635 7505
rect 16577 7454 16635 7471
rect 16871 7544 16905 7565
rect 16948 7557 17014 7599
rect 16948 7523 16964 7557
rect 16998 7523 17014 7557
rect 17048 7531 17099 7565
rect 16871 7489 16905 7510
rect 17048 7497 17049 7531
rect 17083 7527 17099 7531
rect 17048 7493 17050 7497
rect 17084 7493 17099 7527
rect 16871 7455 17014 7489
rect 15146 7341 15163 7375
rect 15197 7341 15214 7375
rect 15146 7324 15214 7341
rect 15510 7411 15580 7426
rect 15510 7377 15527 7411
rect 15561 7377 15580 7411
rect 14479 7241 14513 7275
rect 14656 7270 14707 7304
rect 14479 7173 14513 7207
rect 14479 7123 14513 7139
rect 14556 7207 14572 7241
rect 14606 7207 14622 7241
rect 14556 7173 14622 7207
rect 14556 7139 14572 7173
rect 14606 7139 14622 7173
rect 14556 7089 14622 7139
rect 14656 7236 14658 7270
rect 14692 7236 14707 7270
rect 14656 7189 14707 7236
rect 14656 7155 14658 7189
rect 14692 7155 14707 7189
rect 14656 7123 14707 7155
rect 14742 7301 14794 7319
rect 14776 7267 14794 7301
rect 14742 7233 14794 7267
rect 14776 7199 14794 7233
rect 14742 7165 14794 7199
rect 15510 7176 15580 7377
rect 15933 7375 16175 7445
rect 15933 7341 16011 7375
rect 16045 7341 16121 7375
rect 16155 7341 16175 7375
rect 16209 7377 16229 7411
rect 16263 7377 16339 7411
rect 16373 7377 16451 7411
rect 16209 7307 16451 7377
rect 16853 7401 16924 7419
rect 16853 7395 16873 7401
rect 16853 7361 16865 7395
rect 16907 7367 16924 7401
rect 16899 7361 16924 7367
rect 16853 7345 16924 7361
rect 16980 7417 17014 7455
rect 17048 7450 17099 7493
rect 16980 7401 17031 7417
rect 16980 7367 16997 7401
rect 16980 7351 17031 7367
rect 15933 7267 16451 7307
rect 15933 7233 15951 7267
rect 15985 7233 16399 7267
rect 16433 7233 16451 7267
rect 14776 7131 14794 7165
rect 14742 7089 14794 7131
rect 14829 7165 15898 7176
rect 14829 7131 14847 7165
rect 14881 7131 15847 7165
rect 15881 7131 15898 7165
rect 14829 7089 15898 7131
rect 15933 7165 16451 7233
rect 15933 7131 15951 7165
rect 15985 7131 16399 7165
rect 16433 7131 16451 7165
rect 15933 7089 16451 7131
rect 16577 7287 16635 7322
rect 16980 7309 17014 7351
rect 16577 7253 16589 7287
rect 16623 7253 16635 7287
rect 16577 7194 16635 7253
rect 16577 7160 16589 7194
rect 16623 7160 16635 7194
rect 16577 7089 16635 7160
rect 16871 7275 17014 7309
rect 17065 7304 17099 7450
rect 17134 7553 17186 7599
rect 17168 7519 17186 7553
rect 17134 7485 17186 7519
rect 17168 7451 17186 7485
rect 17134 7431 17186 7451
rect 17221 7538 17923 7599
rect 17221 7504 17239 7538
rect 17273 7504 17871 7538
rect 17905 7504 17923 7538
rect 17221 7445 17923 7504
rect 18067 7544 18101 7565
rect 18144 7557 18210 7599
rect 18144 7523 18160 7557
rect 18194 7523 18210 7557
rect 18244 7531 18295 7565
rect 18067 7489 18101 7510
rect 18244 7497 18245 7531
rect 18279 7527 18295 7531
rect 18244 7493 18246 7497
rect 18280 7493 18295 7527
rect 18067 7455 18210 7489
rect 17221 7375 17551 7445
rect 17221 7341 17299 7375
rect 17333 7341 17398 7375
rect 17432 7341 17497 7375
rect 17531 7341 17551 7375
rect 17585 7377 17605 7411
rect 17639 7377 17708 7411
rect 17742 7377 17811 7411
rect 17845 7377 17923 7411
rect 16871 7241 16905 7275
rect 17048 7270 17099 7304
rect 16871 7173 16905 7207
rect 16871 7123 16905 7139
rect 16948 7207 16964 7241
rect 16998 7207 17014 7241
rect 16948 7173 17014 7207
rect 16948 7139 16964 7173
rect 16998 7139 17014 7173
rect 16948 7089 17014 7139
rect 17048 7236 17050 7270
rect 17084 7236 17099 7270
rect 17048 7189 17099 7236
rect 17048 7155 17050 7189
rect 17084 7155 17099 7189
rect 17048 7123 17099 7155
rect 17134 7301 17186 7319
rect 17585 7307 17923 7377
rect 18049 7401 18120 7419
rect 18049 7395 18069 7401
rect 18049 7361 18061 7395
rect 18103 7367 18120 7401
rect 18095 7361 18120 7367
rect 18049 7345 18120 7361
rect 18176 7417 18210 7455
rect 18244 7450 18295 7493
rect 18176 7401 18227 7417
rect 18176 7367 18193 7401
rect 18176 7351 18227 7367
rect 18176 7309 18210 7351
rect 17168 7267 17186 7301
rect 17134 7233 17186 7267
rect 17168 7199 17186 7233
rect 17134 7165 17186 7199
rect 17168 7131 17186 7165
rect 17134 7089 17186 7131
rect 17221 7267 17923 7307
rect 17221 7233 17239 7267
rect 17273 7233 17871 7267
rect 17905 7233 17923 7267
rect 17221 7165 17923 7233
rect 17221 7131 17239 7165
rect 17273 7131 17871 7165
rect 17905 7131 17923 7165
rect 17221 7089 17923 7131
rect 18067 7275 18210 7309
rect 18261 7304 18295 7450
rect 18330 7553 18382 7599
rect 18364 7519 18382 7553
rect 18330 7485 18382 7519
rect 18364 7451 18382 7485
rect 18330 7431 18382 7451
rect 18601 7536 18843 7599
rect 18601 7502 18619 7536
rect 18653 7502 18791 7536
rect 18825 7502 18843 7536
rect 18601 7449 18843 7502
rect 18601 7381 18651 7415
rect 18685 7381 18705 7415
rect 18067 7241 18101 7275
rect 18244 7270 18295 7304
rect 18067 7173 18101 7207
rect 18067 7123 18101 7139
rect 18144 7207 18160 7241
rect 18194 7207 18210 7241
rect 18144 7173 18210 7207
rect 18144 7139 18160 7173
rect 18194 7139 18210 7173
rect 18144 7089 18210 7139
rect 18244 7236 18246 7270
rect 18280 7236 18295 7270
rect 18244 7189 18295 7236
rect 18244 7155 18246 7189
rect 18280 7155 18295 7189
rect 18244 7123 18295 7155
rect 18330 7301 18382 7319
rect 18364 7267 18382 7301
rect 18330 7233 18382 7267
rect 18364 7199 18382 7233
rect 18330 7165 18382 7199
rect 18364 7131 18382 7165
rect 18330 7089 18382 7131
rect 18601 7307 18705 7381
rect 18739 7375 18843 7449
rect 18739 7341 18759 7375
rect 18793 7341 18843 7375
rect 18601 7260 18843 7307
rect 18601 7226 18619 7260
rect 18653 7226 18791 7260
rect 18825 7226 18843 7260
rect 18601 7165 18843 7226
rect 18601 7131 18619 7165
rect 18653 7131 18791 7165
rect 18825 7131 18843 7165
rect 18601 7089 18843 7131
rect 1104 7055 1133 7089
rect 1167 7055 1225 7089
rect 1259 7055 1317 7089
rect 1351 7055 1409 7089
rect 1443 7055 1501 7089
rect 1535 7055 1593 7089
rect 1627 7055 1685 7089
rect 1719 7055 1777 7089
rect 1811 7055 1869 7089
rect 1903 7055 1961 7089
rect 1995 7055 2053 7089
rect 2087 7055 2145 7089
rect 2179 7055 2237 7089
rect 2271 7055 2329 7089
rect 2363 7055 2421 7089
rect 2455 7055 2513 7089
rect 2547 7055 2605 7089
rect 2639 7055 2697 7089
rect 2731 7055 2789 7089
rect 2823 7055 2881 7089
rect 2915 7055 2973 7089
rect 3007 7055 3065 7089
rect 3099 7055 3157 7089
rect 3191 7055 3249 7089
rect 3283 7055 3341 7089
rect 3375 7055 3433 7089
rect 3467 7055 3525 7089
rect 3559 7055 3617 7089
rect 3651 7055 3709 7089
rect 3743 7055 3801 7089
rect 3835 7055 3893 7089
rect 3927 7055 3985 7089
rect 4019 7055 4077 7089
rect 4111 7055 4169 7089
rect 4203 7055 4261 7089
rect 4295 7055 4353 7089
rect 4387 7055 4445 7089
rect 4479 7055 4537 7089
rect 4571 7055 4629 7089
rect 4663 7055 4721 7089
rect 4755 7055 4813 7089
rect 4847 7055 4905 7089
rect 4939 7055 4997 7089
rect 5031 7055 5089 7089
rect 5123 7055 5181 7089
rect 5215 7055 5273 7089
rect 5307 7055 5365 7089
rect 5399 7055 5457 7089
rect 5491 7055 5549 7089
rect 5583 7055 5641 7089
rect 5675 7055 5733 7089
rect 5767 7055 5825 7089
rect 5859 7055 5917 7089
rect 5951 7055 6009 7089
rect 6043 7055 6101 7089
rect 6135 7055 6193 7089
rect 6227 7055 6285 7089
rect 6319 7055 6377 7089
rect 6411 7055 6469 7089
rect 6503 7055 6561 7089
rect 6595 7055 6653 7089
rect 6687 7055 6745 7089
rect 6779 7055 6837 7089
rect 6871 7055 6929 7089
rect 6963 7055 7021 7089
rect 7055 7055 7113 7089
rect 7147 7055 7205 7089
rect 7239 7055 7297 7089
rect 7331 7055 7389 7089
rect 7423 7055 7481 7089
rect 7515 7055 7573 7089
rect 7607 7055 7665 7089
rect 7699 7055 7757 7089
rect 7791 7055 7849 7089
rect 7883 7055 7941 7089
rect 7975 7055 8033 7089
rect 8067 7055 8125 7089
rect 8159 7055 8217 7089
rect 8251 7055 8309 7089
rect 8343 7055 8401 7089
rect 8435 7055 8493 7089
rect 8527 7055 8585 7089
rect 8619 7055 8677 7089
rect 8711 7055 8769 7089
rect 8803 7055 8861 7089
rect 8895 7055 8953 7089
rect 8987 7055 9045 7089
rect 9079 7055 9137 7089
rect 9171 7055 9229 7089
rect 9263 7055 9321 7089
rect 9355 7055 9413 7089
rect 9447 7055 9505 7089
rect 9539 7055 9597 7089
rect 9631 7055 9689 7089
rect 9723 7055 9781 7089
rect 9815 7055 9873 7089
rect 9907 7055 9965 7089
rect 9999 7055 10057 7089
rect 10091 7055 10149 7089
rect 10183 7055 10241 7089
rect 10275 7055 10333 7089
rect 10367 7055 10425 7089
rect 10459 7055 10517 7089
rect 10551 7055 10609 7089
rect 10643 7055 10701 7089
rect 10735 7055 10793 7089
rect 10827 7055 10885 7089
rect 10919 7055 10977 7089
rect 11011 7055 11069 7089
rect 11103 7055 11161 7089
rect 11195 7055 11253 7089
rect 11287 7055 11345 7089
rect 11379 7055 11437 7089
rect 11471 7055 11529 7089
rect 11563 7055 11621 7089
rect 11655 7055 11713 7089
rect 11747 7055 11805 7089
rect 11839 7055 11897 7089
rect 11931 7055 11989 7089
rect 12023 7055 12081 7089
rect 12115 7055 12173 7089
rect 12207 7055 12265 7089
rect 12299 7055 12357 7089
rect 12391 7055 12449 7089
rect 12483 7055 12541 7089
rect 12575 7055 12633 7089
rect 12667 7055 12725 7089
rect 12759 7055 12817 7089
rect 12851 7055 12909 7089
rect 12943 7055 13001 7089
rect 13035 7055 13093 7089
rect 13127 7055 13185 7089
rect 13219 7055 13277 7089
rect 13311 7055 13369 7089
rect 13403 7055 13461 7089
rect 13495 7055 13553 7089
rect 13587 7055 13645 7089
rect 13679 7055 13737 7089
rect 13771 7055 13829 7089
rect 13863 7055 13921 7089
rect 13955 7055 14013 7089
rect 14047 7055 14105 7089
rect 14139 7055 14197 7089
rect 14231 7055 14289 7089
rect 14323 7055 14381 7089
rect 14415 7055 14473 7089
rect 14507 7055 14565 7089
rect 14599 7055 14657 7089
rect 14691 7055 14749 7089
rect 14783 7055 14841 7089
rect 14875 7055 14933 7089
rect 14967 7055 15025 7089
rect 15059 7055 15117 7089
rect 15151 7055 15209 7089
rect 15243 7055 15301 7089
rect 15335 7055 15393 7089
rect 15427 7055 15485 7089
rect 15519 7055 15577 7089
rect 15611 7055 15669 7089
rect 15703 7055 15761 7089
rect 15795 7055 15853 7089
rect 15887 7055 15945 7089
rect 15979 7055 16037 7089
rect 16071 7055 16129 7089
rect 16163 7055 16221 7089
rect 16255 7055 16313 7089
rect 16347 7055 16405 7089
rect 16439 7055 16497 7089
rect 16531 7055 16589 7089
rect 16623 7055 16681 7089
rect 16715 7055 16773 7089
rect 16807 7055 16865 7089
rect 16899 7055 16957 7089
rect 16991 7055 17049 7089
rect 17083 7055 17141 7089
rect 17175 7055 17233 7089
rect 17267 7055 17325 7089
rect 17359 7055 17417 7089
rect 17451 7055 17509 7089
rect 17543 7055 17601 7089
rect 17635 7055 17693 7089
rect 17727 7055 17785 7089
rect 17819 7055 17877 7089
rect 17911 7055 17969 7089
rect 18003 7055 18061 7089
rect 18095 7055 18153 7089
rect 18187 7055 18245 7089
rect 18279 7055 18337 7089
rect 18371 7055 18429 7089
rect 18463 7055 18521 7089
rect 18555 7055 18613 7089
rect 18647 7055 18705 7089
rect 18739 7055 18797 7089
rect 18831 7055 18860 7089
rect 1121 7013 1363 7055
rect 1121 6979 1139 7013
rect 1173 6979 1311 7013
rect 1345 6979 1363 7013
rect 1121 6918 1363 6979
rect 1397 7013 2466 7055
rect 1397 6979 1415 7013
rect 1449 6979 2415 7013
rect 2449 6979 2466 7013
rect 1397 6968 2466 6979
rect 2501 7013 3570 7055
rect 2501 6979 2519 7013
rect 2553 6979 3519 7013
rect 3553 6979 3570 7013
rect 2501 6968 3570 6979
rect 3697 6984 3755 7055
rect 1121 6884 1139 6918
rect 1173 6884 1311 6918
rect 1345 6884 1363 6918
rect 1121 6837 1363 6884
rect 1121 6769 1171 6803
rect 1205 6769 1225 6803
rect 1121 6695 1225 6769
rect 1259 6763 1363 6837
rect 1259 6729 1279 6763
rect 1313 6729 1363 6763
rect 1714 6803 1782 6820
rect 1714 6769 1731 6803
rect 1765 6769 1782 6803
rect 1121 6642 1363 6695
rect 1714 6654 1782 6769
rect 2078 6767 2148 6968
rect 2078 6733 2095 6767
rect 2129 6733 2148 6767
rect 2078 6718 2148 6733
rect 2818 6803 2886 6820
rect 2818 6769 2835 6803
rect 2869 6769 2886 6803
rect 2818 6654 2886 6769
rect 3182 6767 3252 6968
rect 3697 6950 3709 6984
rect 3743 6950 3755 6984
rect 3789 7013 4858 7055
rect 3789 6979 3807 7013
rect 3841 6979 4807 7013
rect 4841 6979 4858 7013
rect 3789 6968 4858 6979
rect 4893 7013 5962 7055
rect 4893 6979 4911 7013
rect 4945 6979 5911 7013
rect 5945 6979 5962 7013
rect 4893 6968 5962 6979
rect 5997 7013 7066 7055
rect 5997 6979 6015 7013
rect 6049 6979 7015 7013
rect 7049 6979 7066 7013
rect 5997 6968 7066 6979
rect 7101 7013 8170 7055
rect 7101 6979 7119 7013
rect 7153 6979 8119 7013
rect 8153 6979 8170 7013
rect 7101 6968 8170 6979
rect 8205 7013 8723 7055
rect 8205 6979 8223 7013
rect 8257 6979 8671 7013
rect 8705 6979 8723 7013
rect 3697 6891 3755 6950
rect 3697 6857 3709 6891
rect 3743 6857 3755 6891
rect 3697 6822 3755 6857
rect 3182 6733 3199 6767
rect 3233 6733 3252 6767
rect 3182 6718 3252 6733
rect 4106 6803 4174 6820
rect 4106 6769 4123 6803
rect 4157 6769 4174 6803
rect 3697 6673 3755 6690
rect 1121 6608 1139 6642
rect 1173 6608 1311 6642
rect 1345 6608 1363 6642
rect 1121 6545 1363 6608
rect 1397 6640 2466 6654
rect 1397 6606 1415 6640
rect 1449 6606 2415 6640
rect 2449 6606 2466 6640
rect 1397 6545 2466 6606
rect 2501 6640 3570 6654
rect 2501 6606 2519 6640
rect 2553 6606 3519 6640
rect 3553 6606 3570 6640
rect 2501 6545 3570 6606
rect 3697 6639 3709 6673
rect 3743 6639 3755 6673
rect 4106 6654 4174 6769
rect 4470 6767 4540 6968
rect 4470 6733 4487 6767
rect 4521 6733 4540 6767
rect 4470 6718 4540 6733
rect 5210 6803 5278 6820
rect 5210 6769 5227 6803
rect 5261 6769 5278 6803
rect 5210 6654 5278 6769
rect 5574 6767 5644 6968
rect 5574 6733 5591 6767
rect 5625 6733 5644 6767
rect 5574 6718 5644 6733
rect 6314 6803 6382 6820
rect 6314 6769 6331 6803
rect 6365 6769 6382 6803
rect 6314 6654 6382 6769
rect 6678 6767 6748 6968
rect 6678 6733 6695 6767
rect 6729 6733 6748 6767
rect 6678 6718 6748 6733
rect 7418 6803 7486 6820
rect 7418 6769 7435 6803
rect 7469 6769 7486 6803
rect 7418 6654 7486 6769
rect 7782 6767 7852 6968
rect 8205 6911 8723 6979
rect 8205 6877 8223 6911
rect 8257 6877 8671 6911
rect 8705 6877 8723 6911
rect 8205 6837 8723 6877
rect 7782 6733 7799 6767
rect 7833 6733 7852 6767
rect 7782 6718 7852 6733
rect 8205 6769 8283 6803
rect 8317 6769 8393 6803
rect 8427 6769 8447 6803
rect 8205 6699 8447 6769
rect 8481 6767 8723 6837
rect 8849 6984 8907 7055
rect 8849 6950 8861 6984
rect 8895 6950 8907 6984
rect 8941 7013 10010 7055
rect 8941 6979 8959 7013
rect 8993 6979 9959 7013
rect 9993 6979 10010 7013
rect 8941 6968 10010 6979
rect 10045 7013 11114 7055
rect 10045 6979 10063 7013
rect 10097 6979 11063 7013
rect 11097 6979 11114 7013
rect 10045 6968 11114 6979
rect 11149 7013 12218 7055
rect 11149 6979 11167 7013
rect 11201 6979 12167 7013
rect 12201 6979 12218 7013
rect 11149 6968 12218 6979
rect 12253 7013 13322 7055
rect 12253 6979 12271 7013
rect 12305 6979 13271 7013
rect 13305 6979 13322 7013
rect 12253 6968 13322 6979
rect 13357 7013 13875 7055
rect 13357 6979 13375 7013
rect 13409 6979 13823 7013
rect 13857 6979 13875 7013
rect 8849 6891 8907 6950
rect 8849 6857 8861 6891
rect 8895 6857 8907 6891
rect 8849 6822 8907 6857
rect 8481 6733 8501 6767
rect 8535 6733 8611 6767
rect 8645 6733 8723 6767
rect 9258 6803 9326 6820
rect 9258 6769 9275 6803
rect 9309 6769 9326 6803
rect 3697 6545 3755 6639
rect 3789 6640 4858 6654
rect 3789 6606 3807 6640
rect 3841 6606 4807 6640
rect 4841 6606 4858 6640
rect 3789 6545 4858 6606
rect 4893 6640 5962 6654
rect 4893 6606 4911 6640
rect 4945 6606 5911 6640
rect 5945 6606 5962 6640
rect 4893 6545 5962 6606
rect 5997 6640 7066 6654
rect 5997 6606 6015 6640
rect 6049 6606 7015 6640
rect 7049 6606 7066 6640
rect 5997 6545 7066 6606
rect 7101 6640 8170 6654
rect 7101 6606 7119 6640
rect 7153 6606 8119 6640
rect 8153 6606 8170 6640
rect 7101 6545 8170 6606
rect 8205 6640 8723 6699
rect 8205 6606 8223 6640
rect 8257 6606 8671 6640
rect 8705 6606 8723 6640
rect 8205 6545 8723 6606
rect 8849 6673 8907 6690
rect 8849 6639 8861 6673
rect 8895 6639 8907 6673
rect 9258 6654 9326 6769
rect 9622 6767 9692 6968
rect 9622 6733 9639 6767
rect 9673 6733 9692 6767
rect 9622 6718 9692 6733
rect 10362 6803 10430 6820
rect 10362 6769 10379 6803
rect 10413 6769 10430 6803
rect 10362 6654 10430 6769
rect 10726 6767 10796 6968
rect 10726 6733 10743 6767
rect 10777 6733 10796 6767
rect 10726 6718 10796 6733
rect 11466 6803 11534 6820
rect 11466 6769 11483 6803
rect 11517 6769 11534 6803
rect 11466 6654 11534 6769
rect 11830 6767 11900 6968
rect 11830 6733 11847 6767
rect 11881 6733 11900 6767
rect 11830 6718 11900 6733
rect 12570 6803 12638 6820
rect 12570 6769 12587 6803
rect 12621 6769 12638 6803
rect 12570 6654 12638 6769
rect 12934 6767 13004 6968
rect 13357 6911 13875 6979
rect 13357 6877 13375 6911
rect 13409 6877 13823 6911
rect 13857 6877 13875 6911
rect 13357 6837 13875 6877
rect 12934 6733 12951 6767
rect 12985 6733 13004 6767
rect 12934 6718 13004 6733
rect 13357 6769 13435 6803
rect 13469 6769 13545 6803
rect 13579 6769 13599 6803
rect 13357 6699 13599 6769
rect 13633 6767 13875 6837
rect 14001 6984 14059 7055
rect 14001 6950 14013 6984
rect 14047 6950 14059 6984
rect 14093 7013 15162 7055
rect 14093 6979 14111 7013
rect 14145 6979 15111 7013
rect 15145 6979 15162 7013
rect 14093 6968 15162 6979
rect 15197 7013 16266 7055
rect 15197 6979 15215 7013
rect 15249 6979 16215 7013
rect 16249 6979 16266 7013
rect 15197 6968 16266 6979
rect 16301 7013 17370 7055
rect 16301 6979 16319 7013
rect 16353 6979 17319 7013
rect 17353 6979 17370 7013
rect 16301 6968 17370 6979
rect 17405 7013 18474 7055
rect 17405 6979 17423 7013
rect 17457 6979 18423 7013
rect 18457 6979 18474 7013
rect 17405 6968 18474 6979
rect 18601 7013 18843 7055
rect 18601 6979 18619 7013
rect 18653 6979 18791 7013
rect 18825 6979 18843 7013
rect 14001 6891 14059 6950
rect 14001 6857 14013 6891
rect 14047 6857 14059 6891
rect 14001 6822 14059 6857
rect 13633 6733 13653 6767
rect 13687 6733 13763 6767
rect 13797 6733 13875 6767
rect 14410 6803 14478 6820
rect 14410 6769 14427 6803
rect 14461 6769 14478 6803
rect 8849 6545 8907 6639
rect 8941 6640 10010 6654
rect 8941 6606 8959 6640
rect 8993 6606 9959 6640
rect 9993 6606 10010 6640
rect 8941 6545 10010 6606
rect 10045 6640 11114 6654
rect 10045 6606 10063 6640
rect 10097 6606 11063 6640
rect 11097 6606 11114 6640
rect 10045 6545 11114 6606
rect 11149 6640 12218 6654
rect 11149 6606 11167 6640
rect 11201 6606 12167 6640
rect 12201 6606 12218 6640
rect 11149 6545 12218 6606
rect 12253 6640 13322 6654
rect 12253 6606 12271 6640
rect 12305 6606 13271 6640
rect 13305 6606 13322 6640
rect 12253 6545 13322 6606
rect 13357 6640 13875 6699
rect 13357 6606 13375 6640
rect 13409 6606 13823 6640
rect 13857 6606 13875 6640
rect 13357 6545 13875 6606
rect 14001 6673 14059 6690
rect 14001 6639 14013 6673
rect 14047 6639 14059 6673
rect 14410 6654 14478 6769
rect 14774 6767 14844 6968
rect 14774 6733 14791 6767
rect 14825 6733 14844 6767
rect 14774 6718 14844 6733
rect 15514 6803 15582 6820
rect 15514 6769 15531 6803
rect 15565 6769 15582 6803
rect 15514 6654 15582 6769
rect 15878 6767 15948 6968
rect 15878 6733 15895 6767
rect 15929 6733 15948 6767
rect 15878 6718 15948 6733
rect 16618 6803 16686 6820
rect 16618 6769 16635 6803
rect 16669 6769 16686 6803
rect 16618 6654 16686 6769
rect 16982 6767 17052 6968
rect 16982 6733 16999 6767
rect 17033 6733 17052 6767
rect 16982 6718 17052 6733
rect 17722 6803 17790 6820
rect 17722 6769 17739 6803
rect 17773 6769 17790 6803
rect 17722 6654 17790 6769
rect 18086 6767 18156 6968
rect 18086 6733 18103 6767
rect 18137 6733 18156 6767
rect 18086 6718 18156 6733
rect 18601 6918 18843 6979
rect 18601 6884 18619 6918
rect 18653 6884 18791 6918
rect 18825 6884 18843 6918
rect 18601 6837 18843 6884
rect 18601 6763 18705 6837
rect 18601 6729 18651 6763
rect 18685 6729 18705 6763
rect 18739 6769 18759 6803
rect 18793 6769 18843 6803
rect 18739 6695 18843 6769
rect 14001 6545 14059 6639
rect 14093 6640 15162 6654
rect 14093 6606 14111 6640
rect 14145 6606 15111 6640
rect 15145 6606 15162 6640
rect 14093 6545 15162 6606
rect 15197 6640 16266 6654
rect 15197 6606 15215 6640
rect 15249 6606 16215 6640
rect 16249 6606 16266 6640
rect 15197 6545 16266 6606
rect 16301 6640 17370 6654
rect 16301 6606 16319 6640
rect 16353 6606 17319 6640
rect 17353 6606 17370 6640
rect 16301 6545 17370 6606
rect 17405 6640 18474 6654
rect 17405 6606 17423 6640
rect 17457 6606 18423 6640
rect 18457 6606 18474 6640
rect 17405 6545 18474 6606
rect 18601 6642 18843 6695
rect 18601 6608 18619 6642
rect 18653 6608 18791 6642
rect 18825 6608 18843 6642
rect 18601 6545 18843 6608
rect 1104 6511 1133 6545
rect 1167 6511 1225 6545
rect 1259 6511 1317 6545
rect 1351 6511 1409 6545
rect 1443 6511 1501 6545
rect 1535 6511 1593 6545
rect 1627 6511 1685 6545
rect 1719 6511 1777 6545
rect 1811 6511 1869 6545
rect 1903 6511 1961 6545
rect 1995 6511 2053 6545
rect 2087 6511 2145 6545
rect 2179 6511 2237 6545
rect 2271 6511 2329 6545
rect 2363 6511 2421 6545
rect 2455 6511 2513 6545
rect 2547 6511 2605 6545
rect 2639 6511 2697 6545
rect 2731 6511 2789 6545
rect 2823 6511 2881 6545
rect 2915 6511 2973 6545
rect 3007 6511 3065 6545
rect 3099 6511 3157 6545
rect 3191 6511 3249 6545
rect 3283 6511 3341 6545
rect 3375 6511 3433 6545
rect 3467 6511 3525 6545
rect 3559 6511 3617 6545
rect 3651 6511 3709 6545
rect 3743 6511 3801 6545
rect 3835 6511 3893 6545
rect 3927 6511 3985 6545
rect 4019 6511 4077 6545
rect 4111 6511 4169 6545
rect 4203 6511 4261 6545
rect 4295 6511 4353 6545
rect 4387 6511 4445 6545
rect 4479 6511 4537 6545
rect 4571 6511 4629 6545
rect 4663 6511 4721 6545
rect 4755 6511 4813 6545
rect 4847 6511 4905 6545
rect 4939 6511 4997 6545
rect 5031 6511 5089 6545
rect 5123 6511 5181 6545
rect 5215 6511 5273 6545
rect 5307 6511 5365 6545
rect 5399 6511 5457 6545
rect 5491 6511 5549 6545
rect 5583 6511 5641 6545
rect 5675 6511 5733 6545
rect 5767 6511 5825 6545
rect 5859 6511 5917 6545
rect 5951 6511 6009 6545
rect 6043 6511 6101 6545
rect 6135 6511 6193 6545
rect 6227 6511 6285 6545
rect 6319 6511 6377 6545
rect 6411 6511 6469 6545
rect 6503 6511 6561 6545
rect 6595 6511 6653 6545
rect 6687 6511 6745 6545
rect 6779 6511 6837 6545
rect 6871 6511 6929 6545
rect 6963 6511 7021 6545
rect 7055 6511 7113 6545
rect 7147 6511 7205 6545
rect 7239 6511 7297 6545
rect 7331 6511 7389 6545
rect 7423 6511 7481 6545
rect 7515 6511 7573 6545
rect 7607 6511 7665 6545
rect 7699 6511 7757 6545
rect 7791 6511 7849 6545
rect 7883 6511 7941 6545
rect 7975 6511 8033 6545
rect 8067 6511 8125 6545
rect 8159 6511 8217 6545
rect 8251 6511 8309 6545
rect 8343 6511 8401 6545
rect 8435 6511 8493 6545
rect 8527 6511 8585 6545
rect 8619 6511 8677 6545
rect 8711 6511 8769 6545
rect 8803 6511 8861 6545
rect 8895 6511 8953 6545
rect 8987 6511 9045 6545
rect 9079 6511 9137 6545
rect 9171 6511 9229 6545
rect 9263 6511 9321 6545
rect 9355 6511 9413 6545
rect 9447 6511 9505 6545
rect 9539 6511 9597 6545
rect 9631 6511 9689 6545
rect 9723 6511 9781 6545
rect 9815 6511 9873 6545
rect 9907 6511 9965 6545
rect 9999 6511 10057 6545
rect 10091 6511 10149 6545
rect 10183 6511 10241 6545
rect 10275 6511 10333 6545
rect 10367 6511 10425 6545
rect 10459 6511 10517 6545
rect 10551 6511 10609 6545
rect 10643 6511 10701 6545
rect 10735 6511 10793 6545
rect 10827 6511 10885 6545
rect 10919 6511 10977 6545
rect 11011 6511 11069 6545
rect 11103 6511 11161 6545
rect 11195 6511 11253 6545
rect 11287 6511 11345 6545
rect 11379 6511 11437 6545
rect 11471 6511 11529 6545
rect 11563 6511 11621 6545
rect 11655 6511 11713 6545
rect 11747 6511 11805 6545
rect 11839 6511 11897 6545
rect 11931 6511 11989 6545
rect 12023 6511 12081 6545
rect 12115 6511 12173 6545
rect 12207 6511 12265 6545
rect 12299 6511 12357 6545
rect 12391 6511 12449 6545
rect 12483 6511 12541 6545
rect 12575 6511 12633 6545
rect 12667 6511 12725 6545
rect 12759 6511 12817 6545
rect 12851 6511 12909 6545
rect 12943 6511 13001 6545
rect 13035 6511 13093 6545
rect 13127 6511 13185 6545
rect 13219 6511 13277 6545
rect 13311 6511 13369 6545
rect 13403 6511 13461 6545
rect 13495 6511 13553 6545
rect 13587 6511 13645 6545
rect 13679 6511 13737 6545
rect 13771 6511 13829 6545
rect 13863 6511 13921 6545
rect 13955 6511 14013 6545
rect 14047 6511 14105 6545
rect 14139 6511 14197 6545
rect 14231 6511 14289 6545
rect 14323 6511 14381 6545
rect 14415 6511 14473 6545
rect 14507 6511 14565 6545
rect 14599 6511 14657 6545
rect 14691 6511 14749 6545
rect 14783 6511 14841 6545
rect 14875 6511 14933 6545
rect 14967 6511 15025 6545
rect 15059 6511 15117 6545
rect 15151 6511 15209 6545
rect 15243 6511 15301 6545
rect 15335 6511 15393 6545
rect 15427 6511 15485 6545
rect 15519 6511 15577 6545
rect 15611 6511 15669 6545
rect 15703 6511 15761 6545
rect 15795 6511 15853 6545
rect 15887 6511 15945 6545
rect 15979 6511 16037 6545
rect 16071 6511 16129 6545
rect 16163 6511 16221 6545
rect 16255 6511 16313 6545
rect 16347 6511 16405 6545
rect 16439 6511 16497 6545
rect 16531 6511 16589 6545
rect 16623 6511 16681 6545
rect 16715 6511 16773 6545
rect 16807 6511 16865 6545
rect 16899 6511 16957 6545
rect 16991 6511 17049 6545
rect 17083 6511 17141 6545
rect 17175 6511 17233 6545
rect 17267 6511 17325 6545
rect 17359 6511 17417 6545
rect 17451 6511 17509 6545
rect 17543 6511 17601 6545
rect 17635 6511 17693 6545
rect 17727 6511 17785 6545
rect 17819 6511 17877 6545
rect 17911 6511 17969 6545
rect 18003 6511 18061 6545
rect 18095 6511 18153 6545
rect 18187 6511 18245 6545
rect 18279 6511 18337 6545
rect 18371 6511 18429 6545
rect 18463 6511 18521 6545
rect 18555 6511 18613 6545
rect 18647 6511 18705 6545
rect 18739 6511 18797 6545
rect 18831 6511 18860 6545
rect 1121 6448 1363 6511
rect 1121 6414 1139 6448
rect 1173 6414 1311 6448
rect 1345 6414 1363 6448
rect 1121 6361 1363 6414
rect 1397 6450 2466 6511
rect 1397 6416 1415 6450
rect 1449 6416 2415 6450
rect 2449 6416 2466 6450
rect 1397 6402 2466 6416
rect 2501 6450 3570 6511
rect 2501 6416 2519 6450
rect 2553 6416 3519 6450
rect 3553 6416 3570 6450
rect 2501 6402 3570 6416
rect 3605 6450 4674 6511
rect 3605 6416 3623 6450
rect 3657 6416 4623 6450
rect 4657 6416 4674 6450
rect 3605 6402 4674 6416
rect 4709 6450 5778 6511
rect 4709 6416 4727 6450
rect 4761 6416 5727 6450
rect 5761 6416 5778 6450
rect 4709 6402 5778 6416
rect 5813 6443 6147 6511
rect 5813 6409 5831 6443
rect 5865 6409 6095 6443
rect 6129 6409 6147 6443
rect 1121 6287 1225 6361
rect 1121 6253 1171 6287
rect 1205 6253 1225 6287
rect 1259 6293 1279 6327
rect 1313 6293 1363 6327
rect 1259 6219 1363 6293
rect 1714 6287 1782 6402
rect 1714 6253 1731 6287
rect 1765 6253 1782 6287
rect 1714 6236 1782 6253
rect 2078 6323 2148 6338
rect 2078 6289 2095 6323
rect 2129 6289 2148 6323
rect 1121 6172 1363 6219
rect 1121 6138 1139 6172
rect 1173 6138 1311 6172
rect 1345 6138 1363 6172
rect 1121 6077 1363 6138
rect 2078 6088 2148 6289
rect 2818 6287 2886 6402
rect 2818 6253 2835 6287
rect 2869 6253 2886 6287
rect 2818 6236 2886 6253
rect 3182 6323 3252 6338
rect 3182 6289 3199 6323
rect 3233 6289 3252 6323
rect 3182 6088 3252 6289
rect 3922 6287 3990 6402
rect 3922 6253 3939 6287
rect 3973 6253 3990 6287
rect 3922 6236 3990 6253
rect 4286 6323 4356 6338
rect 4286 6289 4303 6323
rect 4337 6289 4356 6323
rect 4286 6088 4356 6289
rect 5026 6287 5094 6402
rect 5813 6357 6147 6409
rect 6273 6417 6331 6511
rect 6273 6383 6285 6417
rect 6319 6383 6331 6417
rect 6365 6450 7434 6511
rect 6365 6416 6383 6450
rect 6417 6416 7383 6450
rect 7417 6416 7434 6450
rect 6365 6402 7434 6416
rect 7469 6450 8538 6511
rect 7469 6416 7487 6450
rect 7521 6416 8487 6450
rect 8521 6416 8538 6450
rect 7469 6402 8538 6416
rect 8573 6450 9642 6511
rect 8573 6416 8591 6450
rect 8625 6416 9591 6450
rect 9625 6416 9642 6450
rect 8573 6402 9642 6416
rect 9677 6450 10746 6511
rect 9677 6416 9695 6450
rect 9729 6416 10695 6450
rect 10729 6416 10746 6450
rect 9677 6402 10746 6416
rect 10781 6450 11299 6511
rect 10781 6416 10799 6450
rect 10833 6416 11247 6450
rect 11281 6416 11299 6450
rect 6273 6366 6331 6383
rect 5026 6253 5043 6287
rect 5077 6253 5094 6287
rect 5026 6236 5094 6253
rect 5390 6323 5460 6338
rect 5390 6289 5407 6323
rect 5441 6289 5460 6323
rect 5390 6088 5460 6289
rect 5813 6287 5963 6357
rect 5813 6253 5833 6287
rect 5867 6253 5963 6287
rect 5997 6289 6093 6323
rect 6127 6289 6147 6323
rect 5997 6219 6147 6289
rect 6682 6287 6750 6402
rect 6682 6253 6699 6287
rect 6733 6253 6750 6287
rect 6682 6236 6750 6253
rect 7046 6323 7116 6338
rect 7046 6289 7063 6323
rect 7097 6289 7116 6323
rect 5813 6179 6147 6219
rect 5813 6145 5831 6179
rect 5865 6145 6095 6179
rect 6129 6145 6147 6179
rect 1121 6043 1139 6077
rect 1173 6043 1311 6077
rect 1345 6043 1363 6077
rect 1121 6001 1363 6043
rect 1397 6077 2466 6088
rect 1397 6043 1415 6077
rect 1449 6043 2415 6077
rect 2449 6043 2466 6077
rect 1397 6001 2466 6043
rect 2501 6077 3570 6088
rect 2501 6043 2519 6077
rect 2553 6043 3519 6077
rect 3553 6043 3570 6077
rect 2501 6001 3570 6043
rect 3605 6077 4674 6088
rect 3605 6043 3623 6077
rect 3657 6043 4623 6077
rect 4657 6043 4674 6077
rect 3605 6001 4674 6043
rect 4709 6077 5778 6088
rect 4709 6043 4727 6077
rect 4761 6043 5727 6077
rect 5761 6043 5778 6077
rect 4709 6001 5778 6043
rect 5813 6077 6147 6145
rect 5813 6043 5831 6077
rect 5865 6043 6095 6077
rect 6129 6043 6147 6077
rect 5813 6001 6147 6043
rect 6273 6199 6331 6234
rect 6273 6165 6285 6199
rect 6319 6165 6331 6199
rect 6273 6106 6331 6165
rect 6273 6072 6285 6106
rect 6319 6072 6331 6106
rect 7046 6088 7116 6289
rect 7786 6287 7854 6402
rect 7786 6253 7803 6287
rect 7837 6253 7854 6287
rect 7786 6236 7854 6253
rect 8150 6323 8220 6338
rect 8150 6289 8167 6323
rect 8201 6289 8220 6323
rect 8150 6088 8220 6289
rect 8890 6287 8958 6402
rect 8890 6253 8907 6287
rect 8941 6253 8958 6287
rect 8890 6236 8958 6253
rect 9254 6323 9324 6338
rect 9254 6289 9271 6323
rect 9305 6289 9324 6323
rect 9254 6088 9324 6289
rect 9994 6287 10062 6402
rect 10781 6357 11299 6416
rect 11425 6417 11483 6511
rect 11425 6383 11437 6417
rect 11471 6383 11483 6417
rect 11517 6450 12586 6511
rect 11517 6416 11535 6450
rect 11569 6416 12535 6450
rect 12569 6416 12586 6450
rect 11517 6402 12586 6416
rect 12621 6450 13690 6511
rect 12621 6416 12639 6450
rect 12673 6416 13639 6450
rect 13673 6416 13690 6450
rect 12621 6402 13690 6416
rect 13725 6450 14794 6511
rect 13725 6416 13743 6450
rect 13777 6416 14743 6450
rect 14777 6416 14794 6450
rect 13725 6402 14794 6416
rect 14829 6450 15898 6511
rect 14829 6416 14847 6450
rect 14881 6416 15847 6450
rect 15881 6416 15898 6450
rect 14829 6402 15898 6416
rect 15933 6450 16451 6511
rect 15933 6416 15951 6450
rect 15985 6416 16399 6450
rect 16433 6416 16451 6450
rect 11425 6366 11483 6383
rect 9994 6253 10011 6287
rect 10045 6253 10062 6287
rect 9994 6236 10062 6253
rect 10358 6323 10428 6338
rect 10358 6289 10375 6323
rect 10409 6289 10428 6323
rect 10358 6088 10428 6289
rect 10781 6287 11023 6357
rect 10781 6253 10859 6287
rect 10893 6253 10969 6287
rect 11003 6253 11023 6287
rect 11057 6289 11077 6323
rect 11111 6289 11187 6323
rect 11221 6289 11299 6323
rect 11057 6219 11299 6289
rect 11834 6287 11902 6402
rect 11834 6253 11851 6287
rect 11885 6253 11902 6287
rect 11834 6236 11902 6253
rect 12198 6323 12268 6338
rect 12198 6289 12215 6323
rect 12249 6289 12268 6323
rect 10781 6179 11299 6219
rect 10781 6145 10799 6179
rect 10833 6145 11247 6179
rect 11281 6145 11299 6179
rect 6273 6001 6331 6072
rect 6365 6077 7434 6088
rect 6365 6043 6383 6077
rect 6417 6043 7383 6077
rect 7417 6043 7434 6077
rect 6365 6001 7434 6043
rect 7469 6077 8538 6088
rect 7469 6043 7487 6077
rect 7521 6043 8487 6077
rect 8521 6043 8538 6077
rect 7469 6001 8538 6043
rect 8573 6077 9642 6088
rect 8573 6043 8591 6077
rect 8625 6043 9591 6077
rect 9625 6043 9642 6077
rect 8573 6001 9642 6043
rect 9677 6077 10746 6088
rect 9677 6043 9695 6077
rect 9729 6043 10695 6077
rect 10729 6043 10746 6077
rect 9677 6001 10746 6043
rect 10781 6077 11299 6145
rect 10781 6043 10799 6077
rect 10833 6043 11247 6077
rect 11281 6043 11299 6077
rect 10781 6001 11299 6043
rect 11425 6199 11483 6234
rect 11425 6165 11437 6199
rect 11471 6165 11483 6199
rect 11425 6106 11483 6165
rect 11425 6072 11437 6106
rect 11471 6072 11483 6106
rect 12198 6088 12268 6289
rect 12938 6287 13006 6402
rect 12938 6253 12955 6287
rect 12989 6253 13006 6287
rect 12938 6236 13006 6253
rect 13302 6323 13372 6338
rect 13302 6289 13319 6323
rect 13353 6289 13372 6323
rect 13302 6088 13372 6289
rect 14042 6287 14110 6402
rect 14042 6253 14059 6287
rect 14093 6253 14110 6287
rect 14042 6236 14110 6253
rect 14406 6323 14476 6338
rect 14406 6289 14423 6323
rect 14457 6289 14476 6323
rect 14406 6088 14476 6289
rect 15146 6287 15214 6402
rect 15933 6357 16451 6416
rect 16577 6417 16635 6511
rect 16577 6383 16589 6417
rect 16623 6383 16635 6417
rect 16669 6450 17738 6511
rect 16669 6416 16687 6450
rect 16721 6416 17687 6450
rect 17721 6416 17738 6450
rect 16669 6402 17738 6416
rect 17773 6450 18475 6511
rect 17773 6416 17791 6450
rect 17825 6416 18423 6450
rect 18457 6416 18475 6450
rect 16577 6366 16635 6383
rect 15146 6253 15163 6287
rect 15197 6253 15214 6287
rect 15146 6236 15214 6253
rect 15510 6323 15580 6338
rect 15510 6289 15527 6323
rect 15561 6289 15580 6323
rect 15510 6088 15580 6289
rect 15933 6287 16175 6357
rect 15933 6253 16011 6287
rect 16045 6253 16121 6287
rect 16155 6253 16175 6287
rect 16209 6289 16229 6323
rect 16263 6289 16339 6323
rect 16373 6289 16451 6323
rect 16209 6219 16451 6289
rect 16986 6287 17054 6402
rect 17773 6357 18475 6416
rect 18601 6448 18843 6511
rect 18601 6414 18619 6448
rect 18653 6414 18791 6448
rect 18825 6414 18843 6448
rect 18601 6361 18843 6414
rect 16986 6253 17003 6287
rect 17037 6253 17054 6287
rect 16986 6236 17054 6253
rect 17350 6323 17420 6338
rect 17350 6289 17367 6323
rect 17401 6289 17420 6323
rect 15933 6179 16451 6219
rect 15933 6145 15951 6179
rect 15985 6145 16399 6179
rect 16433 6145 16451 6179
rect 11425 6001 11483 6072
rect 11517 6077 12586 6088
rect 11517 6043 11535 6077
rect 11569 6043 12535 6077
rect 12569 6043 12586 6077
rect 11517 6001 12586 6043
rect 12621 6077 13690 6088
rect 12621 6043 12639 6077
rect 12673 6043 13639 6077
rect 13673 6043 13690 6077
rect 12621 6001 13690 6043
rect 13725 6077 14794 6088
rect 13725 6043 13743 6077
rect 13777 6043 14743 6077
rect 14777 6043 14794 6077
rect 13725 6001 14794 6043
rect 14829 6077 15898 6088
rect 14829 6043 14847 6077
rect 14881 6043 15847 6077
rect 15881 6043 15898 6077
rect 14829 6001 15898 6043
rect 15933 6077 16451 6145
rect 15933 6043 15951 6077
rect 15985 6043 16399 6077
rect 16433 6043 16451 6077
rect 15933 6001 16451 6043
rect 16577 6199 16635 6234
rect 16577 6165 16589 6199
rect 16623 6165 16635 6199
rect 16577 6106 16635 6165
rect 16577 6072 16589 6106
rect 16623 6072 16635 6106
rect 17350 6088 17420 6289
rect 17773 6287 18103 6357
rect 17773 6253 17851 6287
rect 17885 6253 17950 6287
rect 17984 6253 18049 6287
rect 18083 6253 18103 6287
rect 18137 6289 18157 6323
rect 18191 6289 18260 6323
rect 18294 6289 18363 6323
rect 18397 6289 18475 6323
rect 18137 6219 18475 6289
rect 17773 6179 18475 6219
rect 17773 6145 17791 6179
rect 17825 6145 18423 6179
rect 18457 6145 18475 6179
rect 16577 6001 16635 6072
rect 16669 6077 17738 6088
rect 16669 6043 16687 6077
rect 16721 6043 17687 6077
rect 17721 6043 17738 6077
rect 16669 6001 17738 6043
rect 17773 6077 18475 6145
rect 17773 6043 17791 6077
rect 17825 6043 18423 6077
rect 18457 6043 18475 6077
rect 17773 6001 18475 6043
rect 18601 6293 18651 6327
rect 18685 6293 18705 6327
rect 18601 6219 18705 6293
rect 18739 6287 18843 6361
rect 18739 6253 18759 6287
rect 18793 6253 18843 6287
rect 18601 6172 18843 6219
rect 18601 6138 18619 6172
rect 18653 6138 18791 6172
rect 18825 6138 18843 6172
rect 18601 6077 18843 6138
rect 18601 6043 18619 6077
rect 18653 6043 18791 6077
rect 18825 6043 18843 6077
rect 18601 6001 18843 6043
rect 1104 5967 1133 6001
rect 1167 5967 1225 6001
rect 1259 5967 1317 6001
rect 1351 5967 1409 6001
rect 1443 5967 1501 6001
rect 1535 5967 1593 6001
rect 1627 5967 1685 6001
rect 1719 5967 1777 6001
rect 1811 5967 1869 6001
rect 1903 5967 1961 6001
rect 1995 5967 2053 6001
rect 2087 5967 2145 6001
rect 2179 5967 2237 6001
rect 2271 5967 2329 6001
rect 2363 5967 2421 6001
rect 2455 5967 2513 6001
rect 2547 5967 2605 6001
rect 2639 5967 2697 6001
rect 2731 5967 2789 6001
rect 2823 5967 2881 6001
rect 2915 5967 2973 6001
rect 3007 5967 3065 6001
rect 3099 5967 3157 6001
rect 3191 5967 3249 6001
rect 3283 5967 3341 6001
rect 3375 5967 3433 6001
rect 3467 5967 3525 6001
rect 3559 5967 3617 6001
rect 3651 5967 3709 6001
rect 3743 5967 3801 6001
rect 3835 5967 3893 6001
rect 3927 5967 3985 6001
rect 4019 5967 4077 6001
rect 4111 5967 4169 6001
rect 4203 5967 4261 6001
rect 4295 5967 4353 6001
rect 4387 5967 4445 6001
rect 4479 5967 4537 6001
rect 4571 5967 4629 6001
rect 4663 5967 4721 6001
rect 4755 5967 4813 6001
rect 4847 5967 4905 6001
rect 4939 5967 4997 6001
rect 5031 5967 5089 6001
rect 5123 5967 5181 6001
rect 5215 5967 5273 6001
rect 5307 5967 5365 6001
rect 5399 5967 5457 6001
rect 5491 5967 5549 6001
rect 5583 5967 5641 6001
rect 5675 5967 5733 6001
rect 5767 5967 5825 6001
rect 5859 5967 5917 6001
rect 5951 5967 6009 6001
rect 6043 5967 6101 6001
rect 6135 5967 6193 6001
rect 6227 5967 6285 6001
rect 6319 5967 6377 6001
rect 6411 5967 6469 6001
rect 6503 5967 6561 6001
rect 6595 5967 6653 6001
rect 6687 5967 6745 6001
rect 6779 5967 6837 6001
rect 6871 5967 6929 6001
rect 6963 5967 7021 6001
rect 7055 5967 7113 6001
rect 7147 5967 7205 6001
rect 7239 5967 7297 6001
rect 7331 5967 7389 6001
rect 7423 5967 7481 6001
rect 7515 5967 7573 6001
rect 7607 5967 7665 6001
rect 7699 5967 7757 6001
rect 7791 5967 7849 6001
rect 7883 5967 7941 6001
rect 7975 5967 8033 6001
rect 8067 5967 8125 6001
rect 8159 5967 8217 6001
rect 8251 5967 8309 6001
rect 8343 5967 8401 6001
rect 8435 5967 8493 6001
rect 8527 5967 8585 6001
rect 8619 5967 8677 6001
rect 8711 5967 8769 6001
rect 8803 5967 8861 6001
rect 8895 5967 8953 6001
rect 8987 5967 9045 6001
rect 9079 5967 9137 6001
rect 9171 5967 9229 6001
rect 9263 5967 9321 6001
rect 9355 5967 9413 6001
rect 9447 5967 9505 6001
rect 9539 5967 9597 6001
rect 9631 5967 9689 6001
rect 9723 5967 9781 6001
rect 9815 5967 9873 6001
rect 9907 5967 9965 6001
rect 9999 5967 10057 6001
rect 10091 5967 10149 6001
rect 10183 5967 10241 6001
rect 10275 5967 10333 6001
rect 10367 5967 10425 6001
rect 10459 5967 10517 6001
rect 10551 5967 10609 6001
rect 10643 5967 10701 6001
rect 10735 5967 10793 6001
rect 10827 5967 10885 6001
rect 10919 5967 10977 6001
rect 11011 5967 11069 6001
rect 11103 5967 11161 6001
rect 11195 5967 11253 6001
rect 11287 5967 11345 6001
rect 11379 5967 11437 6001
rect 11471 5967 11529 6001
rect 11563 5967 11621 6001
rect 11655 5967 11713 6001
rect 11747 5967 11805 6001
rect 11839 5967 11897 6001
rect 11931 5967 11989 6001
rect 12023 5967 12081 6001
rect 12115 5967 12173 6001
rect 12207 5967 12265 6001
rect 12299 5967 12357 6001
rect 12391 5967 12449 6001
rect 12483 5967 12541 6001
rect 12575 5967 12633 6001
rect 12667 5967 12725 6001
rect 12759 5967 12817 6001
rect 12851 5967 12909 6001
rect 12943 5967 13001 6001
rect 13035 5967 13093 6001
rect 13127 5967 13185 6001
rect 13219 5967 13277 6001
rect 13311 5967 13369 6001
rect 13403 5967 13461 6001
rect 13495 5967 13553 6001
rect 13587 5967 13645 6001
rect 13679 5967 13737 6001
rect 13771 5967 13829 6001
rect 13863 5967 13921 6001
rect 13955 5967 14013 6001
rect 14047 5967 14105 6001
rect 14139 5967 14197 6001
rect 14231 5967 14289 6001
rect 14323 5967 14381 6001
rect 14415 5967 14473 6001
rect 14507 5967 14565 6001
rect 14599 5967 14657 6001
rect 14691 5967 14749 6001
rect 14783 5967 14841 6001
rect 14875 5967 14933 6001
rect 14967 5967 15025 6001
rect 15059 5967 15117 6001
rect 15151 5967 15209 6001
rect 15243 5967 15301 6001
rect 15335 5967 15393 6001
rect 15427 5967 15485 6001
rect 15519 5967 15577 6001
rect 15611 5967 15669 6001
rect 15703 5967 15761 6001
rect 15795 5967 15853 6001
rect 15887 5967 15945 6001
rect 15979 5967 16037 6001
rect 16071 5967 16129 6001
rect 16163 5967 16221 6001
rect 16255 5967 16313 6001
rect 16347 5967 16405 6001
rect 16439 5967 16497 6001
rect 16531 5967 16589 6001
rect 16623 5967 16681 6001
rect 16715 5967 16773 6001
rect 16807 5967 16865 6001
rect 16899 5967 16957 6001
rect 16991 5967 17049 6001
rect 17083 5967 17141 6001
rect 17175 5967 17233 6001
rect 17267 5967 17325 6001
rect 17359 5967 17417 6001
rect 17451 5967 17509 6001
rect 17543 5967 17601 6001
rect 17635 5967 17693 6001
rect 17727 5967 17785 6001
rect 17819 5967 17877 6001
rect 17911 5967 17969 6001
rect 18003 5967 18061 6001
rect 18095 5967 18153 6001
rect 18187 5967 18245 6001
rect 18279 5967 18337 6001
rect 18371 5967 18429 6001
rect 18463 5967 18521 6001
rect 18555 5967 18613 6001
rect 18647 5967 18705 6001
rect 18739 5967 18797 6001
rect 18831 5967 18860 6001
rect 1121 5925 1363 5967
rect 1121 5891 1139 5925
rect 1173 5891 1311 5925
rect 1345 5891 1363 5925
rect 1121 5830 1363 5891
rect 1121 5796 1139 5830
rect 1173 5796 1311 5830
rect 1345 5796 1363 5830
rect 1121 5749 1363 5796
rect 1397 5925 2099 5967
rect 1397 5891 1415 5925
rect 1449 5891 2047 5925
rect 2081 5891 2099 5925
rect 1397 5823 2099 5891
rect 1397 5789 1415 5823
rect 1449 5789 2047 5823
rect 2081 5789 2099 5823
rect 1397 5749 2099 5789
rect 1121 5681 1171 5715
rect 1205 5681 1225 5715
rect 1121 5607 1225 5681
rect 1259 5675 1363 5749
rect 1259 5641 1279 5675
rect 1313 5641 1363 5675
rect 1397 5681 1475 5715
rect 1509 5681 1574 5715
rect 1608 5681 1673 5715
rect 1707 5681 1727 5715
rect 1397 5611 1727 5681
rect 1761 5679 2099 5749
rect 2243 5917 2277 5933
rect 2243 5849 2277 5883
rect 2313 5917 2379 5967
rect 2313 5883 2329 5917
rect 2363 5883 2379 5917
rect 2313 5849 2379 5883
rect 2313 5815 2329 5849
rect 2363 5815 2379 5849
rect 2413 5917 2467 5933
rect 2413 5883 2415 5917
rect 2449 5883 2467 5917
rect 2413 5836 2467 5883
rect 2243 5781 2277 5815
rect 2413 5802 2415 5836
rect 2449 5831 2467 5836
rect 2413 5797 2421 5802
rect 2455 5797 2467 5831
rect 2243 5747 2376 5781
rect 2413 5752 2467 5797
rect 2342 5718 2376 5747
rect 1761 5645 1781 5679
rect 1815 5645 1884 5679
rect 1918 5645 1987 5679
rect 2021 5645 2099 5679
rect 2229 5695 2295 5711
rect 2229 5661 2237 5695
rect 2271 5689 2295 5695
rect 2229 5655 2245 5661
rect 2279 5655 2295 5689
rect 2229 5637 2295 5655
rect 2342 5702 2399 5718
rect 2342 5668 2365 5702
rect 2342 5652 2399 5668
rect 1121 5554 1363 5607
rect 1121 5520 1139 5554
rect 1173 5520 1311 5554
rect 1345 5520 1363 5554
rect 1121 5457 1363 5520
rect 1397 5552 2099 5611
rect 2342 5601 2376 5652
rect 1397 5518 1415 5552
rect 1449 5518 2047 5552
rect 2081 5518 2099 5552
rect 1397 5457 2099 5518
rect 2243 5567 2376 5601
rect 2433 5592 2467 5752
rect 2501 5925 3019 5967
rect 2501 5891 2519 5925
rect 2553 5891 2967 5925
rect 3001 5891 3019 5925
rect 2501 5823 3019 5891
rect 2501 5789 2519 5823
rect 2553 5789 2967 5823
rect 3001 5789 3019 5823
rect 2501 5749 3019 5789
rect 2243 5546 2277 5567
rect 2415 5563 2467 5592
rect 2243 5491 2277 5512
rect 2313 5499 2329 5533
rect 2363 5499 2379 5533
rect 2313 5457 2379 5499
rect 2449 5529 2467 5563
rect 2415 5491 2467 5529
rect 2501 5681 2579 5715
rect 2613 5681 2689 5715
rect 2723 5681 2743 5715
rect 2501 5611 2743 5681
rect 2777 5679 3019 5749
rect 2777 5645 2797 5679
rect 2831 5645 2907 5679
rect 2941 5645 3019 5679
rect 3053 5917 3107 5933
rect 3053 5883 3071 5917
rect 3105 5883 3107 5917
rect 3053 5836 3107 5883
rect 3053 5802 3071 5836
rect 3105 5802 3107 5836
rect 3141 5917 3207 5967
rect 3141 5883 3157 5917
rect 3191 5883 3207 5917
rect 3141 5849 3207 5883
rect 3141 5815 3157 5849
rect 3191 5815 3207 5849
rect 3243 5917 3277 5933
rect 3243 5849 3277 5883
rect 3053 5752 3107 5802
rect 3243 5781 3277 5815
rect 2501 5552 3019 5611
rect 2501 5518 2519 5552
rect 2553 5518 2967 5552
rect 3001 5518 3019 5552
rect 2501 5457 3019 5518
rect 3053 5592 3087 5752
rect 3144 5747 3277 5781
rect 3329 5925 3663 5967
rect 3329 5891 3347 5925
rect 3381 5891 3611 5925
rect 3645 5891 3663 5925
rect 3329 5823 3663 5891
rect 3329 5789 3347 5823
rect 3381 5789 3611 5823
rect 3645 5789 3663 5823
rect 3329 5749 3663 5789
rect 3144 5718 3178 5747
rect 3121 5702 3178 5718
rect 3155 5668 3178 5702
rect 3121 5652 3178 5668
rect 3144 5601 3178 5652
rect 3225 5695 3291 5711
rect 3225 5689 3249 5695
rect 3225 5655 3241 5689
rect 3283 5661 3291 5695
rect 3275 5655 3291 5661
rect 3225 5637 3291 5655
rect 3329 5681 3349 5715
rect 3383 5681 3479 5715
rect 3329 5611 3479 5681
rect 3513 5679 3663 5749
rect 3697 5896 3755 5967
rect 3697 5862 3709 5896
rect 3743 5862 3755 5896
rect 3789 5925 4858 5967
rect 3789 5891 3807 5925
rect 3841 5891 4807 5925
rect 4841 5891 4858 5925
rect 3789 5880 4858 5891
rect 4893 5925 5962 5967
rect 4893 5891 4911 5925
rect 4945 5891 5911 5925
rect 5945 5891 5962 5925
rect 4893 5880 5962 5891
rect 5997 5925 6699 5967
rect 5997 5891 6015 5925
rect 6049 5891 6647 5925
rect 6681 5891 6699 5925
rect 3697 5803 3755 5862
rect 3697 5769 3709 5803
rect 3743 5769 3755 5803
rect 3697 5734 3755 5769
rect 3513 5645 3609 5679
rect 3643 5645 3663 5679
rect 4106 5715 4174 5732
rect 4106 5681 4123 5715
rect 4157 5681 4174 5715
rect 3053 5563 3105 5592
rect 3144 5567 3277 5601
rect 3053 5559 3071 5563
rect 3053 5525 3065 5559
rect 3243 5546 3277 5567
rect 3099 5525 3105 5529
rect 3053 5491 3105 5525
rect 3141 5499 3157 5533
rect 3191 5499 3207 5533
rect 3141 5457 3207 5499
rect 3243 5491 3277 5512
rect 3329 5559 3663 5611
rect 3329 5525 3347 5559
rect 3381 5525 3611 5559
rect 3645 5525 3663 5559
rect 3329 5457 3663 5525
rect 3697 5585 3755 5602
rect 3697 5551 3709 5585
rect 3743 5551 3755 5585
rect 4106 5566 4174 5681
rect 4470 5679 4540 5880
rect 4470 5645 4487 5679
rect 4521 5645 4540 5679
rect 4470 5630 4540 5645
rect 5210 5715 5278 5732
rect 5210 5681 5227 5715
rect 5261 5681 5278 5715
rect 5210 5566 5278 5681
rect 5574 5679 5644 5880
rect 5997 5823 6699 5891
rect 5997 5789 6015 5823
rect 6049 5789 6647 5823
rect 6681 5789 6699 5823
rect 5997 5749 6699 5789
rect 5574 5645 5591 5679
rect 5625 5645 5644 5679
rect 5574 5630 5644 5645
rect 5997 5681 6075 5715
rect 6109 5681 6174 5715
rect 6208 5681 6273 5715
rect 6307 5681 6327 5715
rect 5997 5611 6327 5681
rect 6361 5679 6699 5749
rect 6361 5645 6381 5679
rect 6415 5645 6484 5679
rect 6518 5645 6587 5679
rect 6621 5645 6699 5679
rect 6734 5925 6801 5933
rect 6734 5891 6751 5925
rect 6785 5891 6801 5925
rect 6734 5857 6801 5891
rect 6734 5823 6751 5857
rect 6785 5823 6801 5857
rect 6734 5789 6801 5823
rect 6734 5755 6751 5789
rect 6785 5755 6801 5789
rect 6734 5739 6801 5755
rect 6835 5925 6869 5967
rect 6835 5857 6869 5891
rect 6835 5789 6869 5823
rect 6835 5739 6869 5755
rect 6903 5899 7309 5933
rect 3697 5457 3755 5551
rect 3789 5552 4858 5566
rect 3789 5518 3807 5552
rect 3841 5518 4807 5552
rect 4841 5518 4858 5552
rect 3789 5457 4858 5518
rect 4893 5552 5962 5566
rect 4893 5518 4911 5552
rect 4945 5518 5911 5552
rect 5945 5518 5962 5552
rect 4893 5457 5962 5518
rect 5997 5552 6699 5611
rect 5997 5518 6015 5552
rect 6049 5518 6647 5552
rect 6681 5518 6699 5552
rect 5997 5457 6699 5518
rect 6734 5605 6768 5739
rect 6903 5705 6937 5899
rect 6802 5689 6853 5705
rect 6836 5655 6853 5689
rect 6802 5639 6853 5655
rect 6898 5689 6937 5705
rect 6932 5655 6937 5689
rect 6898 5639 6937 5655
rect 6971 5831 7071 5865
rect 7105 5831 7146 5865
rect 7180 5831 7196 5865
rect 6819 5605 6853 5639
rect 6971 5605 7005 5831
rect 6734 5559 6785 5605
rect 6819 5571 7005 5605
rect 7039 5766 7241 5797
rect 7039 5763 7207 5766
rect 7039 5653 7073 5763
rect 7203 5732 7207 5763
rect 7039 5603 7073 5619
rect 7114 5653 7169 5723
rect 7114 5619 7135 5653
rect 6734 5525 6745 5559
rect 6779 5552 6785 5559
rect 6970 5564 7005 5571
rect 6970 5548 7076 5564
rect 7114 5559 7169 5619
rect 6734 5518 6751 5525
rect 6734 5491 6785 5518
rect 6819 5533 6885 5537
rect 6819 5499 6835 5533
rect 6869 5499 6885 5533
rect 6819 5457 6885 5499
rect 6970 5514 7042 5548
rect 7147 5525 7169 5559
rect 6970 5491 7076 5514
rect 7114 5491 7169 5525
rect 7203 5627 7241 5732
rect 7275 5766 7309 5899
rect 7343 5865 7377 5967
rect 7561 5925 8630 5967
rect 7343 5815 7377 5831
rect 7424 5865 7527 5897
rect 7561 5891 7579 5925
rect 7613 5891 8579 5925
rect 8613 5891 8630 5925
rect 7561 5880 8630 5891
rect 8849 5896 8907 5967
rect 7424 5831 7429 5865
rect 7463 5831 7527 5865
rect 7424 5815 7527 5831
rect 7275 5763 7375 5766
rect 7275 5729 7297 5763
rect 7331 5732 7375 5763
rect 7409 5732 7425 5766
rect 7331 5729 7425 5732
rect 7275 5728 7425 5729
rect 7459 5653 7527 5815
rect 7203 5593 7205 5627
rect 7239 5593 7241 5627
rect 7281 5619 7297 5653
rect 7331 5619 7527 5653
rect 7878 5715 7946 5732
rect 7878 5681 7895 5715
rect 7929 5681 7946 5715
rect 7203 5491 7241 5593
rect 7277 5548 7379 5564
rect 7311 5514 7345 5548
rect 7277 5457 7379 5514
rect 7423 5548 7472 5619
rect 7878 5566 7946 5681
rect 8242 5679 8312 5880
rect 8849 5862 8861 5896
rect 8895 5862 8907 5896
rect 8849 5803 8907 5862
rect 8849 5769 8861 5803
rect 8895 5769 8907 5803
rect 8849 5734 8907 5769
rect 8941 5925 9643 5967
rect 8941 5891 8959 5925
rect 8993 5891 9591 5925
rect 9625 5891 9643 5925
rect 8941 5823 9643 5891
rect 8941 5789 8959 5823
rect 8993 5789 9591 5823
rect 9625 5789 9643 5823
rect 8941 5749 9643 5789
rect 8242 5645 8259 5679
rect 8293 5645 8312 5679
rect 8242 5630 8312 5645
rect 8941 5681 9019 5715
rect 9053 5681 9118 5715
rect 9152 5681 9217 5715
rect 9251 5681 9271 5715
rect 8941 5611 9271 5681
rect 9305 5679 9643 5749
rect 9305 5645 9325 5679
rect 9359 5645 9428 5679
rect 9462 5645 9531 5679
rect 9565 5645 9643 5679
rect 9862 5925 9929 5933
rect 9862 5891 9879 5925
rect 9913 5891 9929 5925
rect 9862 5857 9929 5891
rect 9862 5823 9879 5857
rect 9913 5823 9929 5857
rect 9862 5789 9929 5823
rect 9862 5755 9879 5789
rect 9913 5755 9929 5789
rect 9862 5739 9929 5755
rect 9963 5925 9997 5967
rect 9963 5857 9997 5891
rect 9963 5789 9997 5823
rect 9963 5739 9997 5755
rect 10031 5899 10437 5933
rect 8849 5585 8907 5602
rect 7423 5514 7429 5548
rect 7463 5514 7472 5548
rect 7423 5498 7472 5514
rect 7561 5552 8630 5566
rect 7561 5518 7579 5552
rect 7613 5518 8579 5552
rect 8613 5518 8630 5552
rect 7561 5457 8630 5518
rect 8849 5551 8861 5585
rect 8895 5551 8907 5585
rect 8849 5457 8907 5551
rect 8941 5552 9643 5611
rect 8941 5518 8959 5552
rect 8993 5518 9591 5552
rect 9625 5518 9643 5552
rect 8941 5457 9643 5518
rect 9862 5605 9896 5739
rect 10031 5705 10065 5899
rect 9930 5689 9981 5705
rect 9964 5655 9981 5689
rect 9930 5639 9981 5655
rect 10026 5689 10065 5705
rect 10060 5655 10065 5689
rect 10026 5639 10065 5655
rect 10099 5831 10199 5865
rect 10233 5831 10274 5865
rect 10308 5831 10324 5865
rect 9947 5605 9981 5639
rect 10099 5605 10133 5831
rect 9862 5559 9913 5605
rect 9947 5571 10133 5605
rect 10167 5766 10369 5797
rect 10167 5763 10335 5766
rect 10167 5653 10201 5763
rect 10331 5732 10335 5763
rect 10242 5695 10297 5723
rect 10275 5661 10297 5695
rect 10167 5603 10201 5619
rect 10242 5653 10297 5661
rect 10242 5619 10263 5653
rect 9862 5525 9873 5559
rect 9907 5552 9913 5559
rect 10098 5564 10133 5571
rect 10098 5548 10204 5564
rect 9862 5518 9879 5525
rect 9862 5491 9913 5518
rect 9947 5533 10013 5537
rect 9947 5499 9963 5533
rect 9997 5499 10013 5533
rect 9947 5457 10013 5499
rect 10098 5514 10170 5548
rect 10098 5491 10204 5514
rect 10242 5491 10297 5619
rect 10331 5627 10369 5732
rect 10403 5766 10437 5899
rect 10471 5865 10505 5967
rect 10689 5925 11023 5967
rect 10471 5815 10505 5831
rect 10552 5865 10655 5897
rect 10552 5831 10557 5865
rect 10591 5831 10655 5865
rect 10552 5815 10655 5831
rect 10403 5763 10503 5766
rect 10403 5729 10425 5763
rect 10459 5732 10503 5763
rect 10537 5732 10553 5766
rect 10459 5729 10553 5732
rect 10403 5728 10553 5729
rect 10587 5653 10655 5815
rect 10689 5891 10707 5925
rect 10741 5891 10971 5925
rect 11005 5891 11023 5925
rect 10689 5823 11023 5891
rect 10689 5789 10707 5823
rect 10741 5789 10971 5823
rect 11005 5789 11023 5823
rect 10689 5749 11023 5789
rect 10331 5593 10333 5627
rect 10367 5593 10369 5627
rect 10409 5619 10425 5653
rect 10459 5619 10655 5653
rect 10689 5681 10709 5715
rect 10743 5681 10839 5715
rect 10331 5491 10369 5593
rect 10405 5548 10507 5564
rect 10439 5514 10473 5548
rect 10405 5457 10507 5514
rect 10551 5548 10600 5619
rect 10551 5514 10557 5548
rect 10591 5514 10600 5548
rect 10551 5498 10600 5514
rect 10689 5611 10839 5681
rect 10873 5679 11023 5749
rect 10873 5645 10969 5679
rect 11003 5645 11023 5679
rect 11057 5925 11149 5933
rect 11057 5891 11099 5925
rect 11133 5891 11149 5925
rect 11057 5857 11149 5891
rect 11057 5823 11099 5857
rect 11133 5823 11149 5857
rect 11187 5925 11253 5967
rect 11187 5891 11203 5925
rect 11237 5891 11253 5925
rect 11187 5857 11253 5891
rect 11187 5823 11203 5857
rect 11237 5823 11253 5857
rect 11293 5883 11353 5899
rect 11293 5849 11311 5883
rect 11345 5849 11353 5883
rect 10689 5559 11023 5611
rect 10689 5525 10707 5559
rect 10741 5525 10971 5559
rect 11005 5525 11023 5559
rect 10689 5457 11023 5525
rect 11057 5559 11107 5823
rect 11293 5789 11353 5849
rect 11387 5883 11443 5967
rect 11387 5849 11395 5883
rect 11429 5849 11443 5883
rect 11387 5833 11443 5849
rect 11517 5925 12219 5967
rect 11517 5891 11535 5925
rect 11569 5891 12167 5925
rect 12201 5891 12219 5925
rect 11165 5755 11353 5789
rect 11517 5823 12219 5891
rect 11517 5789 11535 5823
rect 11569 5789 12167 5823
rect 12201 5789 12219 5823
rect 11427 5763 11480 5777
rect 11165 5705 11199 5755
rect 11427 5729 11437 5763
rect 11471 5729 11480 5763
rect 11517 5749 12219 5789
rect 11427 5705 11480 5729
rect 11141 5689 11199 5705
rect 11141 5655 11143 5689
rect 11177 5655 11199 5689
rect 11233 5695 11301 5705
rect 11233 5689 11253 5695
rect 11233 5655 11251 5689
rect 11287 5661 11301 5695
rect 11285 5655 11301 5661
rect 11345 5689 11480 5705
rect 11345 5655 11392 5689
rect 11426 5655 11480 5689
rect 11517 5681 11595 5715
rect 11629 5681 11694 5715
rect 11728 5681 11793 5715
rect 11827 5681 11847 5715
rect 11141 5639 11199 5655
rect 11165 5621 11199 5639
rect 11165 5583 11443 5621
rect 11057 5525 11069 5559
rect 11103 5549 11107 5559
rect 11377 5561 11443 5583
rect 11103 5533 11169 5549
rect 11103 5525 11119 5533
rect 11057 5499 11119 5525
rect 11153 5499 11169 5533
rect 11057 5491 11169 5499
rect 11203 5533 11253 5549
rect 11237 5499 11253 5533
rect 11377 5527 11395 5561
rect 11429 5527 11443 5561
rect 11377 5511 11443 5527
rect 11517 5611 11847 5681
rect 11881 5679 12219 5749
rect 11881 5645 11901 5679
rect 11935 5645 12004 5679
rect 12038 5645 12107 5679
rect 12141 5645 12219 5679
rect 12254 5925 12321 5933
rect 12254 5891 12271 5925
rect 12305 5891 12321 5925
rect 12254 5857 12321 5891
rect 12254 5831 12271 5857
rect 12254 5797 12265 5831
rect 12305 5823 12321 5857
rect 12299 5797 12321 5823
rect 12254 5789 12321 5797
rect 12254 5755 12271 5789
rect 12305 5755 12321 5789
rect 12254 5739 12321 5755
rect 12355 5925 12389 5967
rect 12355 5857 12389 5891
rect 12355 5789 12389 5823
rect 12355 5739 12389 5755
rect 12423 5899 12829 5933
rect 11517 5552 12219 5611
rect 11517 5518 11535 5552
rect 11569 5518 12167 5552
rect 12201 5518 12219 5552
rect 11203 5457 11253 5499
rect 11517 5457 12219 5518
rect 12254 5605 12288 5739
rect 12423 5705 12457 5899
rect 12322 5689 12373 5705
rect 12356 5655 12373 5689
rect 12322 5639 12373 5655
rect 12418 5689 12457 5705
rect 12452 5655 12457 5689
rect 12418 5639 12457 5655
rect 12491 5831 12591 5865
rect 12625 5831 12666 5865
rect 12700 5831 12716 5865
rect 12339 5605 12373 5639
rect 12491 5605 12525 5831
rect 12254 5552 12305 5605
rect 12339 5571 12525 5605
rect 12559 5766 12761 5797
rect 12559 5763 12727 5766
rect 12559 5653 12593 5763
rect 12723 5732 12727 5763
rect 12559 5603 12593 5619
rect 12634 5653 12689 5723
rect 12634 5619 12655 5653
rect 12254 5518 12271 5552
rect 12490 5564 12525 5571
rect 12490 5548 12596 5564
rect 12634 5559 12689 5619
rect 12254 5491 12305 5518
rect 12339 5533 12405 5537
rect 12339 5499 12355 5533
rect 12389 5499 12405 5533
rect 12339 5457 12405 5499
rect 12490 5514 12562 5548
rect 12667 5525 12689 5559
rect 12490 5491 12596 5514
rect 12634 5491 12689 5525
rect 12723 5627 12761 5732
rect 12795 5766 12829 5899
rect 12863 5865 12897 5967
rect 13081 5925 13783 5967
rect 12863 5815 12897 5831
rect 12944 5865 13047 5897
rect 12944 5831 12949 5865
rect 12983 5831 13047 5865
rect 12944 5815 13047 5831
rect 12795 5763 12895 5766
rect 12795 5729 12817 5763
rect 12851 5732 12895 5763
rect 12929 5732 12945 5766
rect 12851 5729 12945 5732
rect 12795 5728 12945 5729
rect 12979 5653 13047 5815
rect 13081 5891 13099 5925
rect 13133 5891 13731 5925
rect 13765 5891 13783 5925
rect 13081 5823 13783 5891
rect 13081 5789 13099 5823
rect 13133 5789 13731 5823
rect 13765 5789 13783 5823
rect 13081 5749 13783 5789
rect 12723 5593 12725 5627
rect 12759 5593 12761 5627
rect 12801 5619 12817 5653
rect 12851 5619 13047 5653
rect 13081 5681 13159 5715
rect 13193 5681 13258 5715
rect 13292 5681 13357 5715
rect 13391 5681 13411 5715
rect 12723 5491 12761 5593
rect 12797 5548 12899 5564
rect 12831 5514 12865 5548
rect 12797 5457 12899 5514
rect 12943 5548 12992 5619
rect 12943 5514 12949 5548
rect 12983 5514 12992 5548
rect 12943 5498 12992 5514
rect 13081 5611 13411 5681
rect 13445 5679 13783 5749
rect 14001 5896 14059 5967
rect 14001 5862 14013 5896
rect 14047 5862 14059 5896
rect 14001 5803 14059 5862
rect 14001 5769 14013 5803
rect 14047 5769 14059 5803
rect 14001 5734 14059 5769
rect 14278 5925 14345 5933
rect 14278 5891 14295 5925
rect 14329 5891 14345 5925
rect 14278 5857 14345 5891
rect 14278 5823 14295 5857
rect 14329 5823 14345 5857
rect 14278 5789 14345 5823
rect 14278 5755 14295 5789
rect 14329 5755 14345 5789
rect 14278 5739 14345 5755
rect 14379 5925 14413 5967
rect 14379 5857 14413 5891
rect 14379 5789 14413 5823
rect 14379 5739 14413 5755
rect 14447 5899 14853 5933
rect 13445 5645 13465 5679
rect 13499 5645 13568 5679
rect 13602 5645 13671 5679
rect 13705 5645 13783 5679
rect 13081 5552 13783 5611
rect 14278 5605 14312 5739
rect 14447 5705 14481 5899
rect 14346 5689 14397 5705
rect 14380 5655 14397 5689
rect 14346 5639 14397 5655
rect 14442 5689 14481 5705
rect 14476 5655 14481 5689
rect 14442 5639 14481 5655
rect 14515 5831 14615 5865
rect 14649 5831 14690 5865
rect 14724 5831 14740 5865
rect 14363 5605 14397 5639
rect 14515 5605 14549 5831
rect 13081 5518 13099 5552
rect 13133 5518 13731 5552
rect 13765 5518 13783 5552
rect 13081 5457 13783 5518
rect 14001 5585 14059 5602
rect 14001 5551 14013 5585
rect 14047 5551 14059 5585
rect 14001 5457 14059 5551
rect 14278 5559 14329 5605
rect 14363 5571 14549 5605
rect 14583 5766 14785 5797
rect 14583 5763 14751 5766
rect 14583 5653 14617 5763
rect 14747 5732 14751 5763
rect 14583 5603 14617 5619
rect 14658 5653 14713 5723
rect 14658 5619 14679 5653
rect 14278 5525 14289 5559
rect 14323 5552 14329 5559
rect 14514 5564 14549 5571
rect 14514 5548 14620 5564
rect 14658 5559 14713 5619
rect 14278 5518 14295 5525
rect 14278 5491 14329 5518
rect 14363 5533 14429 5537
rect 14363 5499 14379 5533
rect 14413 5499 14429 5533
rect 14363 5457 14429 5499
rect 14514 5514 14586 5548
rect 14691 5525 14713 5559
rect 14514 5491 14620 5514
rect 14658 5491 14713 5525
rect 14747 5627 14785 5732
rect 14819 5766 14853 5899
rect 14887 5865 14921 5967
rect 15105 5925 16174 5967
rect 14887 5815 14921 5831
rect 14968 5865 15071 5897
rect 15105 5891 15123 5925
rect 15157 5891 16123 5925
rect 16157 5891 16174 5925
rect 15105 5880 16174 5891
rect 16209 5925 17278 5967
rect 16209 5891 16227 5925
rect 16261 5891 17227 5925
rect 17261 5891 17278 5925
rect 16209 5880 17278 5891
rect 17313 5925 18382 5967
rect 17313 5891 17331 5925
rect 17365 5891 18331 5925
rect 18365 5891 18382 5925
rect 17313 5880 18382 5891
rect 18601 5925 18843 5967
rect 18601 5891 18619 5925
rect 18653 5891 18791 5925
rect 18825 5891 18843 5925
rect 14968 5831 14973 5865
rect 15007 5831 15071 5865
rect 14968 5815 15071 5831
rect 14819 5763 14919 5766
rect 14819 5729 14841 5763
rect 14875 5732 14919 5763
rect 14953 5732 14969 5766
rect 14875 5729 14969 5732
rect 14819 5728 14969 5729
rect 15003 5653 15071 5815
rect 14747 5593 14749 5627
rect 14783 5593 14785 5627
rect 14825 5619 14841 5653
rect 14875 5619 15071 5653
rect 15422 5715 15490 5732
rect 15422 5681 15439 5715
rect 15473 5681 15490 5715
rect 14747 5491 14785 5593
rect 14821 5548 14923 5564
rect 14855 5514 14889 5548
rect 14821 5457 14923 5514
rect 14967 5548 15016 5619
rect 15422 5566 15490 5681
rect 15786 5679 15856 5880
rect 15786 5645 15803 5679
rect 15837 5645 15856 5679
rect 15786 5630 15856 5645
rect 16526 5715 16594 5732
rect 16526 5681 16543 5715
rect 16577 5681 16594 5715
rect 16526 5566 16594 5681
rect 16890 5679 16960 5880
rect 16890 5645 16907 5679
rect 16941 5645 16960 5679
rect 16890 5630 16960 5645
rect 17630 5715 17698 5732
rect 17630 5681 17647 5715
rect 17681 5681 17698 5715
rect 17630 5566 17698 5681
rect 17994 5679 18064 5880
rect 17994 5645 18011 5679
rect 18045 5645 18064 5679
rect 17994 5630 18064 5645
rect 18601 5830 18843 5891
rect 18601 5796 18619 5830
rect 18653 5796 18791 5830
rect 18825 5796 18843 5830
rect 18601 5749 18843 5796
rect 18601 5675 18705 5749
rect 18601 5641 18651 5675
rect 18685 5641 18705 5675
rect 18739 5681 18759 5715
rect 18793 5681 18843 5715
rect 18739 5607 18843 5681
rect 14967 5514 14973 5548
rect 15007 5514 15016 5548
rect 14967 5498 15016 5514
rect 15105 5552 16174 5566
rect 15105 5518 15123 5552
rect 15157 5518 16123 5552
rect 16157 5518 16174 5552
rect 15105 5457 16174 5518
rect 16209 5552 17278 5566
rect 16209 5518 16227 5552
rect 16261 5518 17227 5552
rect 17261 5518 17278 5552
rect 16209 5457 17278 5518
rect 17313 5552 18382 5566
rect 17313 5518 17331 5552
rect 17365 5518 18331 5552
rect 18365 5518 18382 5552
rect 17313 5457 18382 5518
rect 18601 5554 18843 5607
rect 18601 5520 18619 5554
rect 18653 5520 18791 5554
rect 18825 5520 18843 5554
rect 18601 5457 18843 5520
rect 1104 5423 1133 5457
rect 1167 5423 1225 5457
rect 1259 5423 1317 5457
rect 1351 5423 1409 5457
rect 1443 5423 1501 5457
rect 1535 5423 1593 5457
rect 1627 5423 1685 5457
rect 1719 5423 1777 5457
rect 1811 5423 1869 5457
rect 1903 5423 1961 5457
rect 1995 5423 2053 5457
rect 2087 5423 2145 5457
rect 2179 5423 2237 5457
rect 2271 5423 2329 5457
rect 2363 5423 2421 5457
rect 2455 5423 2513 5457
rect 2547 5423 2605 5457
rect 2639 5423 2697 5457
rect 2731 5423 2789 5457
rect 2823 5423 2881 5457
rect 2915 5423 2973 5457
rect 3007 5423 3065 5457
rect 3099 5423 3157 5457
rect 3191 5423 3249 5457
rect 3283 5423 3341 5457
rect 3375 5423 3433 5457
rect 3467 5423 3525 5457
rect 3559 5423 3617 5457
rect 3651 5423 3709 5457
rect 3743 5423 3801 5457
rect 3835 5423 3893 5457
rect 3927 5423 3985 5457
rect 4019 5423 4077 5457
rect 4111 5423 4169 5457
rect 4203 5423 4261 5457
rect 4295 5423 4353 5457
rect 4387 5423 4445 5457
rect 4479 5423 4537 5457
rect 4571 5423 4629 5457
rect 4663 5423 4721 5457
rect 4755 5423 4813 5457
rect 4847 5423 4905 5457
rect 4939 5423 4997 5457
rect 5031 5423 5089 5457
rect 5123 5423 5181 5457
rect 5215 5423 5273 5457
rect 5307 5423 5365 5457
rect 5399 5423 5457 5457
rect 5491 5423 5549 5457
rect 5583 5423 5641 5457
rect 5675 5423 5733 5457
rect 5767 5423 5825 5457
rect 5859 5423 5917 5457
rect 5951 5423 6009 5457
rect 6043 5423 6101 5457
rect 6135 5423 6193 5457
rect 6227 5423 6285 5457
rect 6319 5423 6377 5457
rect 6411 5423 6469 5457
rect 6503 5423 6561 5457
rect 6595 5423 6653 5457
rect 6687 5423 6745 5457
rect 6779 5423 6837 5457
rect 6871 5423 6929 5457
rect 6963 5423 7021 5457
rect 7055 5423 7113 5457
rect 7147 5423 7205 5457
rect 7239 5423 7297 5457
rect 7331 5423 7389 5457
rect 7423 5423 7481 5457
rect 7515 5423 7573 5457
rect 7607 5423 7665 5457
rect 7699 5423 7757 5457
rect 7791 5423 7849 5457
rect 7883 5423 7941 5457
rect 7975 5423 8033 5457
rect 8067 5423 8125 5457
rect 8159 5423 8217 5457
rect 8251 5423 8309 5457
rect 8343 5423 8401 5457
rect 8435 5423 8493 5457
rect 8527 5423 8585 5457
rect 8619 5423 8677 5457
rect 8711 5423 8769 5457
rect 8803 5423 8861 5457
rect 8895 5423 8953 5457
rect 8987 5423 9045 5457
rect 9079 5423 9137 5457
rect 9171 5423 9229 5457
rect 9263 5423 9321 5457
rect 9355 5423 9413 5457
rect 9447 5423 9505 5457
rect 9539 5423 9597 5457
rect 9631 5423 9689 5457
rect 9723 5423 9781 5457
rect 9815 5423 9873 5457
rect 9907 5423 9965 5457
rect 9999 5423 10057 5457
rect 10091 5423 10149 5457
rect 10183 5423 10241 5457
rect 10275 5423 10333 5457
rect 10367 5423 10425 5457
rect 10459 5423 10517 5457
rect 10551 5423 10609 5457
rect 10643 5423 10701 5457
rect 10735 5423 10793 5457
rect 10827 5423 10885 5457
rect 10919 5423 10977 5457
rect 11011 5423 11069 5457
rect 11103 5423 11161 5457
rect 11195 5423 11253 5457
rect 11287 5423 11345 5457
rect 11379 5423 11437 5457
rect 11471 5423 11529 5457
rect 11563 5423 11621 5457
rect 11655 5423 11713 5457
rect 11747 5423 11805 5457
rect 11839 5423 11897 5457
rect 11931 5423 11989 5457
rect 12023 5423 12081 5457
rect 12115 5423 12173 5457
rect 12207 5423 12265 5457
rect 12299 5423 12357 5457
rect 12391 5423 12449 5457
rect 12483 5423 12541 5457
rect 12575 5423 12633 5457
rect 12667 5423 12725 5457
rect 12759 5423 12817 5457
rect 12851 5423 12909 5457
rect 12943 5423 13001 5457
rect 13035 5423 13093 5457
rect 13127 5423 13185 5457
rect 13219 5423 13277 5457
rect 13311 5423 13369 5457
rect 13403 5423 13461 5457
rect 13495 5423 13553 5457
rect 13587 5423 13645 5457
rect 13679 5423 13737 5457
rect 13771 5423 13829 5457
rect 13863 5423 13921 5457
rect 13955 5423 14013 5457
rect 14047 5423 14105 5457
rect 14139 5423 14197 5457
rect 14231 5423 14289 5457
rect 14323 5423 14381 5457
rect 14415 5423 14473 5457
rect 14507 5423 14565 5457
rect 14599 5423 14657 5457
rect 14691 5423 14749 5457
rect 14783 5423 14841 5457
rect 14875 5423 14933 5457
rect 14967 5423 15025 5457
rect 15059 5423 15117 5457
rect 15151 5423 15209 5457
rect 15243 5423 15301 5457
rect 15335 5423 15393 5457
rect 15427 5423 15485 5457
rect 15519 5423 15577 5457
rect 15611 5423 15669 5457
rect 15703 5423 15761 5457
rect 15795 5423 15853 5457
rect 15887 5423 15945 5457
rect 15979 5423 16037 5457
rect 16071 5423 16129 5457
rect 16163 5423 16221 5457
rect 16255 5423 16313 5457
rect 16347 5423 16405 5457
rect 16439 5423 16497 5457
rect 16531 5423 16589 5457
rect 16623 5423 16681 5457
rect 16715 5423 16773 5457
rect 16807 5423 16865 5457
rect 16899 5423 16957 5457
rect 16991 5423 17049 5457
rect 17083 5423 17141 5457
rect 17175 5423 17233 5457
rect 17267 5423 17325 5457
rect 17359 5423 17417 5457
rect 17451 5423 17509 5457
rect 17543 5423 17601 5457
rect 17635 5423 17693 5457
rect 17727 5423 17785 5457
rect 17819 5423 17877 5457
rect 17911 5423 17969 5457
rect 18003 5423 18061 5457
rect 18095 5423 18153 5457
rect 18187 5423 18245 5457
rect 18279 5423 18337 5457
rect 18371 5423 18429 5457
rect 18463 5423 18521 5457
rect 18555 5423 18613 5457
rect 18647 5423 18705 5457
rect 18739 5423 18797 5457
rect 18831 5423 18860 5457
rect 1121 5360 1363 5423
rect 1121 5326 1139 5360
rect 1173 5326 1311 5360
rect 1345 5326 1363 5360
rect 1121 5273 1363 5326
rect 1397 5362 1915 5423
rect 1397 5328 1415 5362
rect 1449 5328 1863 5362
rect 1897 5328 1915 5362
rect 1121 5199 1225 5273
rect 1397 5269 1915 5328
rect 1949 5381 2061 5389
rect 1949 5347 2011 5381
rect 2045 5347 2061 5381
rect 1949 5331 2061 5347
rect 2095 5381 2145 5423
rect 2129 5347 2145 5381
rect 2095 5331 2145 5347
rect 2269 5353 2335 5369
rect 1121 5165 1171 5199
rect 1205 5165 1225 5199
rect 1259 5205 1279 5239
rect 1313 5205 1363 5239
rect 1259 5131 1363 5205
rect 1397 5199 1639 5269
rect 1397 5165 1475 5199
rect 1509 5165 1585 5199
rect 1619 5165 1639 5199
rect 1673 5201 1693 5235
rect 1727 5201 1803 5235
rect 1837 5201 1915 5235
rect 1673 5131 1915 5201
rect 1121 5084 1363 5131
rect 1121 5050 1139 5084
rect 1173 5050 1311 5084
rect 1345 5050 1363 5084
rect 1121 4989 1363 5050
rect 1121 4955 1139 4989
rect 1173 4955 1311 4989
rect 1345 4955 1363 4989
rect 1121 4913 1363 4955
rect 1397 5091 1915 5131
rect 1397 5057 1415 5091
rect 1449 5057 1863 5091
rect 1897 5057 1915 5091
rect 1397 4989 1915 5057
rect 1397 4955 1415 4989
rect 1449 4955 1863 4989
rect 1897 4955 1915 4989
rect 1397 4913 1915 4955
rect 1949 5057 1999 5331
rect 2269 5319 2287 5353
rect 2321 5319 2335 5353
rect 2269 5297 2335 5319
rect 2057 5259 2335 5297
rect 2409 5355 2743 5423
rect 2409 5321 2427 5355
rect 2461 5321 2691 5355
rect 2725 5321 2743 5355
rect 2409 5269 2743 5321
rect 2869 5381 2981 5389
rect 2869 5355 2931 5381
rect 2869 5321 2881 5355
rect 2915 5347 2931 5355
rect 2965 5347 2981 5381
rect 2915 5331 2981 5347
rect 3015 5381 3065 5423
rect 3049 5347 3065 5381
rect 3015 5331 3065 5347
rect 3189 5353 3255 5369
rect 2915 5321 2919 5331
rect 2057 5241 2091 5259
rect 2033 5225 2091 5241
rect 2033 5191 2035 5225
rect 2069 5191 2091 5225
rect 2033 5175 2091 5191
rect 2125 5191 2143 5225
rect 2177 5219 2193 5225
rect 2125 5185 2145 5191
rect 2179 5185 2193 5219
rect 2125 5175 2193 5185
rect 2237 5191 2284 5225
rect 2318 5191 2372 5225
rect 2237 5175 2372 5191
rect 2057 5125 2091 5175
rect 2319 5151 2372 5175
rect 2409 5199 2559 5269
rect 2409 5165 2429 5199
rect 2463 5165 2559 5199
rect 2593 5201 2689 5235
rect 2723 5201 2743 5235
rect 2057 5091 2245 5125
rect 2319 5117 2329 5151
rect 2363 5117 2372 5151
rect 2593 5131 2743 5201
rect 2319 5103 2372 5117
rect 1949 5023 1991 5057
rect 2025 5023 2041 5057
rect 1949 5015 2041 5023
rect 1949 4981 1961 5015
rect 1995 4989 2041 5015
rect 1949 4955 1991 4981
rect 2025 4955 2041 4989
rect 1949 4947 2041 4955
rect 2079 5023 2095 5057
rect 2129 5023 2145 5057
rect 2079 4989 2145 5023
rect 2079 4955 2095 4989
rect 2129 4955 2145 4989
rect 2185 5031 2245 5091
rect 2409 5091 2743 5131
rect 2409 5057 2427 5091
rect 2461 5057 2691 5091
rect 2725 5057 2743 5091
rect 2185 4997 2203 5031
rect 2237 4997 2245 5031
rect 2185 4981 2245 4997
rect 2279 5031 2335 5047
rect 2279 4997 2287 5031
rect 2321 4997 2335 5031
rect 2079 4913 2145 4955
rect 2279 4913 2335 4997
rect 2409 4989 2743 5057
rect 2409 4955 2427 4989
rect 2461 4955 2691 4989
rect 2725 4955 2743 4989
rect 2409 4913 2743 4955
rect 2869 5057 2919 5321
rect 3189 5319 3207 5353
rect 3241 5319 3255 5353
rect 3189 5297 3255 5319
rect 2977 5259 3255 5297
rect 3329 5355 3663 5423
rect 3329 5321 3347 5355
rect 3381 5321 3611 5355
rect 3645 5321 3663 5355
rect 3329 5269 3663 5321
rect 3715 5368 3749 5389
rect 3792 5381 3858 5423
rect 3792 5347 3808 5381
rect 3842 5347 3858 5381
rect 3892 5355 3943 5389
rect 3715 5313 3749 5334
rect 3892 5321 3893 5355
rect 3927 5351 3943 5355
rect 3892 5317 3894 5321
rect 3928 5317 3943 5351
rect 3715 5279 3858 5313
rect 2977 5241 3011 5259
rect 2953 5225 3011 5241
rect 2953 5191 2955 5225
rect 2989 5191 3011 5225
rect 2953 5175 3011 5191
rect 3045 5191 3063 5225
rect 3097 5219 3113 5225
rect 3045 5185 3065 5191
rect 3099 5185 3113 5219
rect 3045 5175 3113 5185
rect 3157 5191 3204 5225
rect 3238 5219 3292 5225
rect 3238 5191 3249 5219
rect 3157 5185 3249 5191
rect 3283 5185 3292 5219
rect 3157 5175 3292 5185
rect 2977 5125 3011 5175
rect 2977 5091 3165 5125
rect 3239 5103 3292 5175
rect 3329 5199 3479 5269
rect 3329 5165 3349 5199
rect 3383 5165 3479 5199
rect 3513 5201 3609 5235
rect 3643 5201 3663 5235
rect 3513 5131 3663 5201
rect 3697 5225 3768 5243
rect 3697 5219 3717 5225
rect 3697 5185 3709 5219
rect 3751 5191 3768 5225
rect 3743 5185 3768 5191
rect 3697 5169 3768 5185
rect 3824 5241 3858 5279
rect 3892 5274 3943 5317
rect 3824 5225 3875 5241
rect 3824 5191 3841 5225
rect 3824 5175 3875 5191
rect 3824 5133 3858 5175
rect 2869 5023 2911 5057
rect 2945 5023 2961 5057
rect 2869 4989 2961 5023
rect 2869 4955 2911 4989
rect 2945 4955 2961 4989
rect 2869 4947 2961 4955
rect 2999 5023 3015 5057
rect 3049 5023 3065 5057
rect 2999 4989 3065 5023
rect 2999 4955 3015 4989
rect 3049 4955 3065 4989
rect 3105 5031 3165 5091
rect 3329 5091 3663 5131
rect 3329 5057 3347 5091
rect 3381 5057 3611 5091
rect 3645 5057 3663 5091
rect 3105 4997 3123 5031
rect 3157 4997 3165 5031
rect 3105 4981 3165 4997
rect 3199 5031 3255 5047
rect 3199 4997 3207 5031
rect 3241 4997 3255 5031
rect 2999 4913 3065 4955
rect 3199 4913 3255 4997
rect 3329 4989 3663 5057
rect 3329 4955 3347 4989
rect 3381 4955 3611 4989
rect 3645 4955 3663 4989
rect 3329 4913 3663 4955
rect 3715 5099 3858 5133
rect 3909 5128 3943 5274
rect 3978 5377 4030 5423
rect 4012 5343 4030 5377
rect 3978 5309 4030 5343
rect 4012 5275 4030 5309
rect 3978 5255 4030 5275
rect 4065 5355 4399 5423
rect 4065 5321 4083 5355
rect 4117 5321 4347 5355
rect 4381 5321 4399 5355
rect 4065 5269 4399 5321
rect 4441 5381 4487 5423
rect 4441 5347 4453 5381
rect 4441 5309 4487 5347
rect 4441 5275 4453 5309
rect 4065 5199 4215 5269
rect 4441 5259 4487 5275
rect 4521 5381 4587 5389
rect 4521 5347 4537 5381
rect 4571 5347 4587 5381
rect 4521 5309 4587 5347
rect 4521 5275 4537 5309
rect 4571 5275 4587 5309
rect 4521 5263 4587 5275
rect 4065 5165 4085 5199
rect 4119 5165 4215 5199
rect 4249 5201 4345 5235
rect 4379 5201 4399 5235
rect 3715 5065 3749 5099
rect 3892 5094 3943 5128
rect 3715 4997 3749 5031
rect 3715 4947 3749 4963
rect 3792 5031 3808 5065
rect 3842 5031 3858 5065
rect 3792 4997 3858 5031
rect 3792 4963 3808 4997
rect 3842 4963 3858 4997
rect 3792 4913 3858 4963
rect 3892 5060 3894 5094
rect 3928 5060 3943 5094
rect 3892 5013 3943 5060
rect 3892 4979 3894 5013
rect 3928 4979 3943 5013
rect 3892 4947 3943 4979
rect 3978 5125 4030 5143
rect 4249 5131 4399 5201
rect 4437 5219 4453 5225
rect 4437 5185 4445 5219
rect 4487 5191 4503 5225
rect 4479 5185 4503 5191
rect 4437 5175 4503 5185
rect 4537 5143 4587 5263
rect 4621 5381 4663 5423
rect 4655 5347 4663 5381
rect 4621 5309 4663 5347
rect 4709 5362 5778 5423
rect 4709 5328 4727 5362
rect 4761 5328 5727 5362
rect 5761 5328 5778 5362
rect 4709 5314 5778 5328
rect 5813 5351 5865 5389
rect 5813 5317 5831 5351
rect 5901 5381 5967 5423
rect 5901 5347 5917 5381
rect 5951 5347 5967 5381
rect 6003 5368 6037 5389
rect 4655 5275 4663 5309
rect 4621 5259 4663 5275
rect 5026 5199 5094 5314
rect 5813 5288 5865 5317
rect 6003 5313 6037 5334
rect 5026 5165 5043 5199
rect 5077 5165 5094 5199
rect 5026 5148 5094 5165
rect 5390 5235 5460 5250
rect 5390 5201 5407 5235
rect 5441 5201 5460 5235
rect 4012 5091 4030 5125
rect 3978 5057 4030 5091
rect 4012 5023 4030 5057
rect 3978 4989 4030 5023
rect 4012 4955 4030 4989
rect 3978 4913 4030 4955
rect 4065 5091 4399 5131
rect 4065 5057 4083 5091
rect 4117 5057 4347 5091
rect 4381 5057 4399 5091
rect 4065 4989 4399 5057
rect 4065 4955 4083 4989
rect 4117 4955 4347 4989
rect 4381 4955 4399 4989
rect 4065 4913 4399 4955
rect 4441 5125 4487 5141
rect 4441 5091 4453 5125
rect 4441 5057 4487 5091
rect 4441 5023 4453 5057
rect 4441 4989 4487 5023
rect 4441 4955 4453 4989
rect 4441 4913 4487 4955
rect 4521 5125 4587 5143
rect 4521 5091 4537 5125
rect 4571 5091 4587 5125
rect 4521 5057 4587 5091
rect 4521 5023 4537 5057
rect 4571 5023 4587 5057
rect 4521 5015 4587 5023
rect 4521 4955 4537 5015
rect 4571 4955 4587 5015
rect 4521 4947 4587 4955
rect 4621 5125 4663 5141
rect 4655 5091 4663 5125
rect 4621 5057 4663 5091
rect 4655 5023 4663 5057
rect 4621 4989 4663 5023
rect 5390 5000 5460 5201
rect 5813 5128 5847 5288
rect 5904 5279 6037 5313
rect 6273 5329 6331 5423
rect 6273 5295 6285 5329
rect 6319 5295 6331 5329
rect 5904 5228 5938 5279
rect 6273 5278 6331 5295
rect 6365 5360 6607 5423
rect 6365 5326 6383 5360
rect 6417 5326 6555 5360
rect 6589 5326 6607 5360
rect 6365 5273 6607 5326
rect 6642 5362 6693 5389
rect 6642 5328 6659 5362
rect 6727 5381 6793 5423
rect 6727 5347 6743 5381
rect 6777 5347 6793 5381
rect 6727 5343 6793 5347
rect 6878 5366 6984 5389
rect 6642 5275 6693 5328
rect 6878 5332 6950 5366
rect 7022 5355 7077 5389
rect 6878 5316 6984 5332
rect 7055 5321 7077 5355
rect 6878 5309 6913 5316
rect 6727 5275 6913 5309
rect 5881 5212 5938 5228
rect 5915 5178 5938 5212
rect 5881 5162 5938 5178
rect 5985 5225 6051 5243
rect 5985 5191 6001 5225
rect 6035 5219 6051 5225
rect 5985 5185 6009 5191
rect 6043 5185 6051 5219
rect 5985 5169 6051 5185
rect 6365 5199 6469 5273
rect 6365 5165 6415 5199
rect 6449 5165 6469 5199
rect 6503 5205 6523 5239
rect 6557 5205 6607 5239
rect 5904 5133 5938 5162
rect 5813 5078 5867 5128
rect 5904 5099 6037 5133
rect 5813 5044 5831 5078
rect 5865 5044 5867 5078
rect 6003 5065 6037 5099
rect 5813 5015 5867 5044
rect 4655 4955 4663 4989
rect 4621 4913 4663 4955
rect 4709 4989 5778 5000
rect 4709 4955 4727 4989
rect 4761 4955 5727 4989
rect 5761 4955 5778 4989
rect 4709 4913 5778 4955
rect 5813 4981 5825 5015
rect 5859 4997 5867 5015
rect 5813 4963 5831 4981
rect 5865 4963 5867 4997
rect 5813 4947 5867 4963
rect 5901 5031 5917 5065
rect 5951 5031 5967 5065
rect 5901 4997 5967 5031
rect 5901 4963 5917 4997
rect 5951 4963 5967 4997
rect 5901 4913 5967 4963
rect 6003 4997 6037 5031
rect 6003 4947 6037 4963
rect 6273 5111 6331 5146
rect 6503 5131 6607 5205
rect 6273 5077 6285 5111
rect 6319 5077 6331 5111
rect 6273 5018 6331 5077
rect 6273 4984 6285 5018
rect 6319 4984 6331 5018
rect 6273 4913 6331 4984
rect 6365 5084 6607 5131
rect 6365 5050 6383 5084
rect 6417 5050 6555 5084
rect 6589 5050 6607 5084
rect 6365 4989 6607 5050
rect 6365 4955 6383 4989
rect 6417 4955 6555 4989
rect 6589 4955 6607 4989
rect 6365 4913 6607 4955
rect 6642 5141 6676 5275
rect 6727 5241 6761 5275
rect 6710 5225 6761 5241
rect 6744 5191 6761 5225
rect 6710 5175 6761 5191
rect 6806 5225 6845 5241
rect 6840 5191 6845 5225
rect 6806 5175 6845 5191
rect 6642 5125 6709 5141
rect 6642 5091 6659 5125
rect 6693 5091 6709 5125
rect 6642 5057 6709 5091
rect 6642 5023 6659 5057
rect 6693 5023 6709 5057
rect 6642 5015 6709 5023
rect 6642 4981 6653 5015
rect 6687 4989 6709 5015
rect 6642 4955 6659 4981
rect 6693 4955 6709 4989
rect 6642 4947 6709 4955
rect 6743 5125 6777 5141
rect 6743 5057 6777 5091
rect 6743 4989 6777 5023
rect 6743 4913 6777 4955
rect 6811 4981 6845 5175
rect 6879 5049 6913 5275
rect 6947 5261 6981 5277
rect 6947 5117 6981 5227
rect 7022 5261 7077 5321
rect 7022 5227 7043 5261
rect 7022 5157 7077 5227
rect 7111 5355 7149 5389
rect 7111 5321 7113 5355
rect 7147 5321 7149 5355
rect 7111 5148 7149 5321
rect 7185 5366 7287 5423
rect 7219 5332 7253 5366
rect 7185 5316 7287 5332
rect 7331 5366 7380 5382
rect 7331 5332 7337 5366
rect 7371 5332 7380 5366
rect 7331 5261 7380 5332
rect 7469 5355 7803 5423
rect 7469 5321 7487 5355
rect 7521 5321 7751 5355
rect 7785 5321 7803 5355
rect 7469 5269 7803 5321
rect 7838 5362 7889 5389
rect 7838 5328 7855 5362
rect 7923 5381 7989 5423
rect 7923 5347 7939 5381
rect 7973 5347 7989 5381
rect 7923 5343 7989 5347
rect 8074 5366 8180 5389
rect 7838 5275 7889 5328
rect 8074 5332 8146 5366
rect 8074 5316 8180 5332
rect 8074 5309 8109 5316
rect 7923 5275 8109 5309
rect 7189 5227 7205 5261
rect 7239 5227 7435 5261
rect 7111 5117 7115 5148
rect 6947 5114 7115 5117
rect 6947 5083 7149 5114
rect 7183 5151 7333 5152
rect 7183 5148 7297 5151
rect 7183 5114 7283 5148
rect 7331 5117 7333 5151
rect 7317 5114 7333 5117
rect 6879 5015 6979 5049
rect 7013 5015 7054 5049
rect 7088 5015 7104 5049
rect 7183 4981 7217 5114
rect 7367 5065 7435 5227
rect 7469 5199 7619 5269
rect 7469 5165 7489 5199
rect 7523 5165 7619 5199
rect 7653 5201 7749 5235
rect 7783 5201 7803 5235
rect 7653 5131 7803 5201
rect 6811 4947 7217 4981
rect 7251 5049 7285 5065
rect 7251 4913 7285 5015
rect 7332 5049 7435 5065
rect 7332 5015 7337 5049
rect 7371 5015 7435 5049
rect 7332 4983 7435 5015
rect 7469 5091 7803 5131
rect 7469 5057 7487 5091
rect 7521 5057 7751 5091
rect 7785 5057 7803 5091
rect 7469 4989 7803 5057
rect 7469 4955 7487 4989
rect 7521 4955 7751 4989
rect 7785 4955 7803 4989
rect 7469 4913 7803 4955
rect 7838 5141 7872 5275
rect 7923 5241 7957 5275
rect 7906 5225 7957 5241
rect 7940 5191 7957 5225
rect 7906 5175 7957 5191
rect 8002 5225 8041 5241
rect 8036 5191 8041 5225
rect 8002 5175 8041 5191
rect 7838 5125 7905 5141
rect 7838 5091 7855 5125
rect 7889 5091 7905 5125
rect 7838 5057 7905 5091
rect 7838 5023 7855 5057
rect 7889 5023 7905 5057
rect 7838 5015 7905 5023
rect 7838 4981 7849 5015
rect 7883 4989 7905 5015
rect 7838 4955 7855 4981
rect 7889 4955 7905 4989
rect 7838 4947 7905 4955
rect 7939 5125 7973 5141
rect 7939 5057 7973 5091
rect 7939 4989 7973 5023
rect 7939 4913 7973 4955
rect 8007 4981 8041 5175
rect 8075 5049 8109 5275
rect 8143 5261 8177 5277
rect 8143 5117 8177 5227
rect 8218 5261 8273 5389
rect 8218 5227 8239 5261
rect 8218 5219 8273 5227
rect 8251 5185 8273 5219
rect 8218 5157 8273 5185
rect 8307 5355 8345 5389
rect 8307 5321 8309 5355
rect 8343 5321 8345 5355
rect 8307 5148 8345 5321
rect 8381 5366 8483 5423
rect 8415 5332 8449 5366
rect 8381 5316 8483 5332
rect 8527 5366 8576 5382
rect 8527 5332 8533 5366
rect 8567 5332 8576 5366
rect 8527 5261 8576 5332
rect 8665 5355 8999 5423
rect 8665 5321 8683 5355
rect 8717 5321 8947 5355
rect 8981 5321 8999 5355
rect 8665 5269 8999 5321
rect 9125 5378 9193 5389
rect 9125 5344 9143 5378
rect 9177 5344 9193 5378
rect 9125 5310 9193 5344
rect 9227 5381 9261 5423
rect 9227 5331 9261 5347
rect 9309 5377 9381 5389
rect 9309 5343 9331 5377
rect 9365 5343 9381 5377
rect 9309 5336 9381 5343
rect 9507 5381 9541 5423
rect 9309 5335 9380 5336
rect 9309 5333 9379 5335
rect 9309 5332 9378 5333
rect 9125 5276 9143 5310
rect 9177 5276 9193 5310
rect 9309 5330 9377 5332
rect 9507 5331 9541 5347
rect 9575 5377 9643 5389
rect 9575 5343 9591 5377
rect 9625 5343 9643 5377
rect 9309 5329 9376 5330
rect 9309 5327 9374 5329
rect 9309 5325 9372 5327
rect 9309 5309 9369 5325
rect 9309 5297 9331 5309
rect 8385 5227 8401 5261
rect 8435 5227 8631 5261
rect 8307 5117 8311 5148
rect 8143 5114 8311 5117
rect 8143 5083 8345 5114
rect 8379 5151 8529 5152
rect 8379 5117 8401 5151
rect 8435 5148 8529 5151
rect 8435 5117 8479 5148
rect 8379 5114 8479 5117
rect 8513 5114 8529 5148
rect 8075 5015 8175 5049
rect 8209 5015 8250 5049
rect 8284 5015 8300 5049
rect 8379 4981 8413 5114
rect 8563 5065 8631 5227
rect 8665 5199 8815 5269
rect 8665 5165 8685 5199
rect 8719 5165 8815 5199
rect 8849 5201 8945 5235
rect 8979 5201 8999 5235
rect 8849 5131 8999 5201
rect 8007 4947 8413 4981
rect 8447 5049 8481 5065
rect 8447 4913 8481 5015
rect 8528 5049 8631 5065
rect 8528 5015 8533 5049
rect 8567 5015 8631 5049
rect 8528 4983 8631 5015
rect 8665 5091 8999 5131
rect 8665 5057 8683 5091
rect 8717 5057 8947 5091
rect 8981 5057 8999 5091
rect 8665 4989 8999 5057
rect 8665 4955 8683 4989
rect 8717 4955 8947 4989
rect 8981 4955 8999 4989
rect 8665 4913 8999 4955
rect 9125 5234 9193 5276
rect 9227 5275 9331 5297
rect 9365 5275 9369 5309
rect 9227 5259 9369 5275
rect 9407 5279 9423 5313
rect 9457 5297 9473 5313
rect 9575 5309 9643 5343
rect 9575 5297 9591 5309
rect 9457 5279 9591 5297
rect 9407 5275 9591 5279
rect 9625 5275 9643 5309
rect 9407 5259 9643 5275
rect 9677 5362 10379 5423
rect 9677 5328 9695 5362
rect 9729 5328 10327 5362
rect 10361 5328 10379 5362
rect 9677 5269 10379 5328
rect 10414 5362 10465 5389
rect 10414 5328 10431 5362
rect 10499 5381 10565 5423
rect 10499 5347 10515 5381
rect 10549 5347 10565 5381
rect 10499 5343 10565 5347
rect 10650 5366 10756 5389
rect 10414 5275 10465 5328
rect 10650 5332 10722 5366
rect 10650 5316 10756 5332
rect 10650 5309 10685 5316
rect 10499 5275 10685 5309
rect 9125 5133 9181 5234
rect 9125 5099 9147 5133
rect 9227 5225 9284 5259
rect 9261 5191 9284 5225
rect 9227 5145 9284 5191
rect 9321 5219 9365 5225
rect 9355 5191 9365 5219
rect 9399 5191 9415 5225
rect 9355 5185 9415 5191
rect 9449 5191 9465 5225
rect 9499 5221 9515 5225
rect 9499 5219 9539 5221
rect 9499 5191 9505 5219
rect 9449 5185 9505 5191
rect 9577 5191 9593 5225
rect 9627 5191 9643 5225
rect 9577 5185 9643 5191
rect 9321 5179 9415 5185
rect 9227 5125 9457 5145
rect 9227 5102 9407 5125
rect 9125 5065 9181 5099
rect 9391 5091 9407 5102
rect 9441 5091 9457 5125
rect 9125 5031 9147 5065
rect 9125 5015 9181 5031
rect 9125 4981 9137 5015
rect 9171 4997 9181 5015
rect 9125 4963 9147 4981
rect 9125 4947 9181 4963
rect 9215 5057 9357 5068
rect 9215 5023 9233 5057
rect 9267 5023 9307 5057
rect 9341 5023 9357 5057
rect 9215 4989 9357 5023
rect 9215 4955 9233 4989
rect 9267 4955 9307 4989
rect 9341 4955 9357 4989
rect 9215 4913 9357 4955
rect 9391 5057 9457 5091
rect 9391 5023 9407 5057
rect 9441 5023 9457 5057
rect 9391 4989 9457 5023
rect 9391 4955 9407 4989
rect 9441 4955 9457 4989
rect 9496 4962 9539 5185
rect 9597 5151 9643 5185
rect 9677 5199 10007 5269
rect 9677 5165 9755 5199
rect 9789 5165 9854 5199
rect 9888 5165 9953 5199
rect 9987 5165 10007 5199
rect 10041 5201 10061 5235
rect 10095 5201 10164 5235
rect 10198 5201 10267 5235
rect 10301 5201 10379 5235
rect 9631 5117 9643 5151
rect 10041 5131 10379 5201
rect 9677 5091 10379 5131
rect 9677 5057 9695 5091
rect 9729 5057 10327 5091
rect 10361 5057 10379 5091
rect 9575 5023 9591 5057
rect 9625 5023 9641 5057
rect 9575 4989 9641 5023
rect 9391 4947 9457 4955
rect 9575 4955 9591 4989
rect 9625 4955 9641 4989
rect 9575 4913 9641 4955
rect 9677 4989 10379 5057
rect 9677 4955 9695 4989
rect 9729 4955 10327 4989
rect 10361 4955 10379 4989
rect 9677 4913 10379 4955
rect 10414 5141 10448 5275
rect 10499 5241 10533 5275
rect 10482 5225 10533 5241
rect 10516 5191 10533 5225
rect 10482 5175 10533 5191
rect 10578 5225 10617 5241
rect 10612 5191 10617 5225
rect 10578 5175 10617 5191
rect 10414 5125 10481 5141
rect 10414 5091 10431 5125
rect 10465 5091 10481 5125
rect 10414 5057 10481 5091
rect 10414 5023 10431 5057
rect 10465 5023 10481 5057
rect 10414 5015 10481 5023
rect 10414 4981 10425 5015
rect 10459 4989 10481 5015
rect 10414 4955 10431 4981
rect 10465 4955 10481 4989
rect 10414 4947 10481 4955
rect 10515 5125 10549 5141
rect 10515 5057 10549 5091
rect 10515 4989 10549 5023
rect 10515 4913 10549 4955
rect 10583 4981 10617 5175
rect 10651 5049 10685 5275
rect 10719 5261 10753 5277
rect 10719 5117 10753 5227
rect 10794 5261 10849 5389
rect 10794 5227 10815 5261
rect 10794 5219 10849 5227
rect 10827 5185 10849 5219
rect 10794 5157 10849 5185
rect 10883 5355 10921 5389
rect 10883 5321 10885 5355
rect 10919 5321 10921 5355
rect 10883 5148 10921 5321
rect 10957 5366 11059 5423
rect 10991 5332 11025 5366
rect 10957 5316 11059 5332
rect 11103 5366 11152 5382
rect 11103 5332 11109 5366
rect 11143 5332 11152 5366
rect 11103 5261 11152 5332
rect 11425 5329 11483 5423
rect 11425 5295 11437 5329
rect 11471 5295 11483 5329
rect 11517 5362 12586 5423
rect 11517 5328 11535 5362
rect 11569 5328 12535 5362
rect 12569 5328 12586 5362
rect 11517 5314 12586 5328
rect 12621 5355 12955 5423
rect 12621 5321 12639 5355
rect 12673 5321 12903 5355
rect 12937 5321 12955 5355
rect 11425 5278 11483 5295
rect 10961 5227 10977 5261
rect 11011 5227 11207 5261
rect 10883 5117 10887 5148
rect 10719 5114 10887 5117
rect 10719 5083 10921 5114
rect 10955 5151 11105 5152
rect 10955 5117 10977 5151
rect 11011 5148 11105 5151
rect 11011 5117 11055 5148
rect 10955 5114 11055 5117
rect 11089 5114 11105 5148
rect 10651 5015 10751 5049
rect 10785 5015 10826 5049
rect 10860 5015 10876 5049
rect 10955 4981 10989 5114
rect 11139 5065 11207 5227
rect 11834 5199 11902 5314
rect 12621 5269 12955 5321
rect 13082 5362 13133 5389
rect 13082 5328 13099 5362
rect 13167 5381 13233 5423
rect 13167 5347 13183 5381
rect 13217 5347 13233 5381
rect 13167 5343 13233 5347
rect 13318 5366 13424 5389
rect 13082 5275 13133 5328
rect 13318 5332 13390 5366
rect 13462 5355 13517 5389
rect 13318 5316 13424 5332
rect 13495 5321 13517 5355
rect 13318 5309 13353 5316
rect 13167 5275 13353 5309
rect 11834 5165 11851 5199
rect 11885 5165 11902 5199
rect 11834 5148 11902 5165
rect 12198 5235 12268 5250
rect 12198 5201 12215 5235
rect 12249 5201 12268 5235
rect 10583 4947 10989 4981
rect 11023 5049 11057 5065
rect 11023 4913 11057 5015
rect 11104 5049 11207 5065
rect 11104 5015 11109 5049
rect 11143 5015 11207 5049
rect 11104 4983 11207 5015
rect 11425 5111 11483 5146
rect 11425 5077 11437 5111
rect 11471 5077 11483 5111
rect 11425 5018 11483 5077
rect 11425 4984 11437 5018
rect 11471 4984 11483 5018
rect 12198 5000 12268 5201
rect 12621 5199 12771 5269
rect 12621 5165 12641 5199
rect 12675 5165 12771 5199
rect 12805 5201 12901 5235
rect 12935 5201 12955 5235
rect 12805 5131 12955 5201
rect 12621 5091 12955 5131
rect 12621 5057 12639 5091
rect 12673 5057 12903 5091
rect 12937 5057 12955 5091
rect 11425 4913 11483 4984
rect 11517 4989 12586 5000
rect 11517 4955 11535 4989
rect 11569 4955 12535 4989
rect 12569 4955 12586 4989
rect 11517 4913 12586 4955
rect 12621 4989 12955 5057
rect 12621 4955 12639 4989
rect 12673 4955 12903 4989
rect 12937 4955 12955 4989
rect 12621 4913 12955 4955
rect 13082 5141 13116 5275
rect 13167 5241 13201 5275
rect 13150 5225 13201 5241
rect 13184 5191 13201 5225
rect 13150 5175 13201 5191
rect 13246 5225 13285 5241
rect 13280 5191 13285 5225
rect 13246 5175 13285 5191
rect 13082 5125 13149 5141
rect 13082 5091 13099 5125
rect 13133 5091 13149 5125
rect 13082 5057 13149 5091
rect 13082 5023 13099 5057
rect 13133 5023 13149 5057
rect 13082 5015 13149 5023
rect 13082 4981 13093 5015
rect 13127 4989 13149 5015
rect 13082 4955 13099 4981
rect 13133 4955 13149 4989
rect 13082 4947 13149 4955
rect 13183 5125 13217 5141
rect 13183 5057 13217 5091
rect 13183 4989 13217 5023
rect 13183 4913 13217 4955
rect 13251 4981 13285 5175
rect 13319 5049 13353 5275
rect 13387 5261 13421 5277
rect 13387 5117 13421 5227
rect 13462 5261 13517 5321
rect 13462 5227 13483 5261
rect 13462 5157 13517 5227
rect 13551 5355 13589 5389
rect 13551 5321 13553 5355
rect 13587 5321 13589 5355
rect 13551 5148 13589 5321
rect 13625 5366 13727 5423
rect 13659 5332 13693 5366
rect 13625 5316 13727 5332
rect 13771 5366 13820 5382
rect 13771 5332 13777 5366
rect 13811 5332 13820 5366
rect 13771 5261 13820 5332
rect 13909 5362 14978 5423
rect 13909 5328 13927 5362
rect 13961 5328 14927 5362
rect 14961 5328 14978 5362
rect 13909 5314 14978 5328
rect 15013 5362 16082 5423
rect 15013 5328 15031 5362
rect 15065 5328 16031 5362
rect 16065 5328 16082 5362
rect 15013 5314 16082 5328
rect 16117 5355 16451 5423
rect 16117 5321 16135 5355
rect 16169 5321 16399 5355
rect 16433 5321 16451 5355
rect 13629 5227 13645 5261
rect 13679 5227 13875 5261
rect 13551 5117 13555 5148
rect 13387 5114 13555 5117
rect 13387 5083 13589 5114
rect 13623 5151 13773 5152
rect 13623 5117 13645 5151
rect 13679 5148 13773 5151
rect 13679 5117 13723 5148
rect 13623 5114 13723 5117
rect 13757 5114 13773 5148
rect 13319 5015 13419 5049
rect 13453 5015 13494 5049
rect 13528 5015 13544 5049
rect 13623 4981 13657 5114
rect 13807 5065 13875 5227
rect 14226 5199 14294 5314
rect 14226 5165 14243 5199
rect 14277 5165 14294 5199
rect 14226 5148 14294 5165
rect 14590 5235 14660 5250
rect 14590 5201 14607 5235
rect 14641 5201 14660 5235
rect 13251 4947 13657 4981
rect 13691 5049 13725 5065
rect 13691 4913 13725 5015
rect 13772 5049 13875 5065
rect 13772 5015 13777 5049
rect 13811 5015 13875 5049
rect 13772 4983 13875 5015
rect 14590 5000 14660 5201
rect 15330 5199 15398 5314
rect 16117 5269 16451 5321
rect 16577 5329 16635 5423
rect 16577 5295 16589 5329
rect 16623 5295 16635 5329
rect 16669 5362 17738 5423
rect 16669 5328 16687 5362
rect 16721 5328 17687 5362
rect 17721 5328 17738 5362
rect 16669 5314 17738 5328
rect 17773 5362 18475 5423
rect 17773 5328 17791 5362
rect 17825 5328 18423 5362
rect 18457 5328 18475 5362
rect 16577 5278 16635 5295
rect 15330 5165 15347 5199
rect 15381 5165 15398 5199
rect 15330 5148 15398 5165
rect 15694 5235 15764 5250
rect 15694 5201 15711 5235
rect 15745 5201 15764 5235
rect 15694 5000 15764 5201
rect 16117 5199 16267 5269
rect 16117 5165 16137 5199
rect 16171 5165 16267 5199
rect 16301 5201 16397 5235
rect 16431 5201 16451 5235
rect 16301 5131 16451 5201
rect 16986 5199 17054 5314
rect 17773 5269 18475 5328
rect 18601 5360 18843 5423
rect 18601 5326 18619 5360
rect 18653 5326 18791 5360
rect 18825 5326 18843 5360
rect 18601 5273 18843 5326
rect 16986 5165 17003 5199
rect 17037 5165 17054 5199
rect 16986 5148 17054 5165
rect 17350 5235 17420 5250
rect 17350 5201 17367 5235
rect 17401 5201 17420 5235
rect 16117 5091 16451 5131
rect 16117 5057 16135 5091
rect 16169 5057 16399 5091
rect 16433 5057 16451 5091
rect 13909 4989 14978 5000
rect 13909 4955 13927 4989
rect 13961 4955 14927 4989
rect 14961 4955 14978 4989
rect 13909 4913 14978 4955
rect 15013 4989 16082 5000
rect 15013 4955 15031 4989
rect 15065 4955 16031 4989
rect 16065 4955 16082 4989
rect 15013 4913 16082 4955
rect 16117 4989 16451 5057
rect 16117 4955 16135 4989
rect 16169 4955 16399 4989
rect 16433 4955 16451 4989
rect 16117 4913 16451 4955
rect 16577 5111 16635 5146
rect 16577 5077 16589 5111
rect 16623 5077 16635 5111
rect 16577 5018 16635 5077
rect 16577 4984 16589 5018
rect 16623 4984 16635 5018
rect 17350 5000 17420 5201
rect 17773 5199 18103 5269
rect 17773 5165 17851 5199
rect 17885 5165 17950 5199
rect 17984 5165 18049 5199
rect 18083 5165 18103 5199
rect 18137 5201 18157 5235
rect 18191 5201 18260 5235
rect 18294 5201 18363 5235
rect 18397 5201 18475 5235
rect 18137 5131 18475 5201
rect 17773 5091 18475 5131
rect 17773 5057 17791 5091
rect 17825 5057 18423 5091
rect 18457 5057 18475 5091
rect 16577 4913 16635 4984
rect 16669 4989 17738 5000
rect 16669 4955 16687 4989
rect 16721 4955 17687 4989
rect 17721 4955 17738 4989
rect 16669 4913 17738 4955
rect 17773 4989 18475 5057
rect 17773 4955 17791 4989
rect 17825 4955 18423 4989
rect 18457 4955 18475 4989
rect 17773 4913 18475 4955
rect 18601 5205 18651 5239
rect 18685 5205 18705 5239
rect 18601 5131 18705 5205
rect 18739 5199 18843 5273
rect 18739 5165 18759 5199
rect 18793 5165 18843 5199
rect 18601 5084 18843 5131
rect 18601 5050 18619 5084
rect 18653 5050 18791 5084
rect 18825 5050 18843 5084
rect 18601 4989 18843 5050
rect 18601 4955 18619 4989
rect 18653 4955 18791 4989
rect 18825 4955 18843 4989
rect 18601 4913 18843 4955
rect 1104 4879 1133 4913
rect 1167 4879 1225 4913
rect 1259 4879 1317 4913
rect 1351 4879 1409 4913
rect 1443 4879 1501 4913
rect 1535 4879 1593 4913
rect 1627 4879 1685 4913
rect 1719 4879 1777 4913
rect 1811 4879 1869 4913
rect 1903 4879 1961 4913
rect 1995 4879 2053 4913
rect 2087 4879 2145 4913
rect 2179 4879 2237 4913
rect 2271 4879 2329 4913
rect 2363 4879 2421 4913
rect 2455 4879 2513 4913
rect 2547 4879 2605 4913
rect 2639 4879 2697 4913
rect 2731 4879 2789 4913
rect 2823 4879 2881 4913
rect 2915 4879 2973 4913
rect 3007 4879 3065 4913
rect 3099 4879 3157 4913
rect 3191 4879 3249 4913
rect 3283 4879 3341 4913
rect 3375 4879 3433 4913
rect 3467 4879 3525 4913
rect 3559 4879 3617 4913
rect 3651 4879 3709 4913
rect 3743 4879 3801 4913
rect 3835 4879 3893 4913
rect 3927 4879 3985 4913
rect 4019 4879 4077 4913
rect 4111 4879 4169 4913
rect 4203 4879 4261 4913
rect 4295 4879 4353 4913
rect 4387 4879 4445 4913
rect 4479 4879 4537 4913
rect 4571 4879 4629 4913
rect 4663 4879 4721 4913
rect 4755 4879 4813 4913
rect 4847 4879 4905 4913
rect 4939 4879 4997 4913
rect 5031 4879 5089 4913
rect 5123 4879 5181 4913
rect 5215 4879 5273 4913
rect 5307 4879 5365 4913
rect 5399 4879 5457 4913
rect 5491 4879 5549 4913
rect 5583 4879 5641 4913
rect 5675 4879 5733 4913
rect 5767 4879 5825 4913
rect 5859 4879 5917 4913
rect 5951 4879 6009 4913
rect 6043 4879 6101 4913
rect 6135 4879 6193 4913
rect 6227 4879 6285 4913
rect 6319 4879 6377 4913
rect 6411 4879 6469 4913
rect 6503 4879 6561 4913
rect 6595 4879 6653 4913
rect 6687 4879 6745 4913
rect 6779 4879 6837 4913
rect 6871 4879 6929 4913
rect 6963 4879 7021 4913
rect 7055 4879 7113 4913
rect 7147 4879 7205 4913
rect 7239 4879 7297 4913
rect 7331 4879 7389 4913
rect 7423 4879 7481 4913
rect 7515 4879 7573 4913
rect 7607 4879 7665 4913
rect 7699 4879 7757 4913
rect 7791 4879 7849 4913
rect 7883 4879 7941 4913
rect 7975 4879 8033 4913
rect 8067 4879 8125 4913
rect 8159 4879 8217 4913
rect 8251 4879 8309 4913
rect 8343 4879 8401 4913
rect 8435 4879 8493 4913
rect 8527 4879 8585 4913
rect 8619 4879 8677 4913
rect 8711 4879 8769 4913
rect 8803 4879 8861 4913
rect 8895 4879 8953 4913
rect 8987 4879 9045 4913
rect 9079 4879 9137 4913
rect 9171 4879 9229 4913
rect 9263 4879 9321 4913
rect 9355 4879 9413 4913
rect 9447 4879 9505 4913
rect 9539 4879 9597 4913
rect 9631 4879 9689 4913
rect 9723 4879 9781 4913
rect 9815 4879 9873 4913
rect 9907 4879 9965 4913
rect 9999 4879 10057 4913
rect 10091 4879 10149 4913
rect 10183 4879 10241 4913
rect 10275 4879 10333 4913
rect 10367 4879 10425 4913
rect 10459 4879 10517 4913
rect 10551 4879 10609 4913
rect 10643 4879 10701 4913
rect 10735 4879 10793 4913
rect 10827 4879 10885 4913
rect 10919 4879 10977 4913
rect 11011 4879 11069 4913
rect 11103 4879 11161 4913
rect 11195 4879 11253 4913
rect 11287 4879 11345 4913
rect 11379 4879 11437 4913
rect 11471 4879 11529 4913
rect 11563 4879 11621 4913
rect 11655 4879 11713 4913
rect 11747 4879 11805 4913
rect 11839 4879 11897 4913
rect 11931 4879 11989 4913
rect 12023 4879 12081 4913
rect 12115 4879 12173 4913
rect 12207 4879 12265 4913
rect 12299 4879 12357 4913
rect 12391 4879 12449 4913
rect 12483 4879 12541 4913
rect 12575 4879 12633 4913
rect 12667 4879 12725 4913
rect 12759 4879 12817 4913
rect 12851 4879 12909 4913
rect 12943 4879 13001 4913
rect 13035 4879 13093 4913
rect 13127 4879 13185 4913
rect 13219 4879 13277 4913
rect 13311 4879 13369 4913
rect 13403 4879 13461 4913
rect 13495 4879 13553 4913
rect 13587 4879 13645 4913
rect 13679 4879 13737 4913
rect 13771 4879 13829 4913
rect 13863 4879 13921 4913
rect 13955 4879 14013 4913
rect 14047 4879 14105 4913
rect 14139 4879 14197 4913
rect 14231 4879 14289 4913
rect 14323 4879 14381 4913
rect 14415 4879 14473 4913
rect 14507 4879 14565 4913
rect 14599 4879 14657 4913
rect 14691 4879 14749 4913
rect 14783 4879 14841 4913
rect 14875 4879 14933 4913
rect 14967 4879 15025 4913
rect 15059 4879 15117 4913
rect 15151 4879 15209 4913
rect 15243 4879 15301 4913
rect 15335 4879 15393 4913
rect 15427 4879 15485 4913
rect 15519 4879 15577 4913
rect 15611 4879 15669 4913
rect 15703 4879 15761 4913
rect 15795 4879 15853 4913
rect 15887 4879 15945 4913
rect 15979 4879 16037 4913
rect 16071 4879 16129 4913
rect 16163 4879 16221 4913
rect 16255 4879 16313 4913
rect 16347 4879 16405 4913
rect 16439 4879 16497 4913
rect 16531 4879 16589 4913
rect 16623 4879 16681 4913
rect 16715 4879 16773 4913
rect 16807 4879 16865 4913
rect 16899 4879 16957 4913
rect 16991 4879 17049 4913
rect 17083 4879 17141 4913
rect 17175 4879 17233 4913
rect 17267 4879 17325 4913
rect 17359 4879 17417 4913
rect 17451 4879 17509 4913
rect 17543 4879 17601 4913
rect 17635 4879 17693 4913
rect 17727 4879 17785 4913
rect 17819 4879 17877 4913
rect 17911 4879 17969 4913
rect 18003 4879 18061 4913
rect 18095 4879 18153 4913
rect 18187 4879 18245 4913
rect 18279 4879 18337 4913
rect 18371 4879 18429 4913
rect 18463 4879 18521 4913
rect 18555 4879 18613 4913
rect 18647 4879 18705 4913
rect 18739 4879 18797 4913
rect 18831 4879 18860 4913
rect 1121 4837 1363 4879
rect 1121 4803 1139 4837
rect 1173 4803 1311 4837
rect 1345 4803 1363 4837
rect 1121 4742 1363 4803
rect 1121 4708 1139 4742
rect 1173 4708 1311 4742
rect 1345 4708 1363 4742
rect 1121 4661 1363 4708
rect 1397 4837 1915 4879
rect 1397 4803 1415 4837
rect 1449 4803 1863 4837
rect 1897 4803 1915 4837
rect 1397 4735 1915 4803
rect 1397 4701 1415 4735
rect 1449 4701 1863 4735
rect 1897 4701 1915 4735
rect 2059 4829 2093 4845
rect 2059 4761 2093 4795
rect 2127 4813 2193 4879
rect 2127 4779 2143 4813
rect 2177 4779 2193 4813
rect 2227 4829 2264 4845
rect 2261 4795 2264 4829
rect 2227 4761 2264 4795
rect 2312 4837 2365 4879
rect 2312 4803 2331 4837
rect 2312 4787 2365 4803
rect 2399 4829 2449 4845
rect 2399 4795 2415 4829
rect 2746 4837 2780 4879
rect 2093 4743 2192 4745
rect 2093 4727 2150 4743
rect 2059 4711 2150 4727
rect 1397 4661 1915 4701
rect 2146 4709 2150 4711
rect 2184 4709 2192 4743
rect 1121 4593 1171 4627
rect 1205 4593 1225 4627
rect 1121 4519 1225 4593
rect 1259 4587 1363 4661
rect 1259 4553 1279 4587
rect 1313 4553 1363 4587
rect 1397 4593 1475 4627
rect 1509 4593 1585 4627
rect 1619 4593 1639 4627
rect 1397 4523 1639 4593
rect 1673 4591 1915 4661
rect 1673 4557 1693 4591
rect 1727 4557 1803 4591
rect 1837 4557 1915 4591
rect 2042 4607 2112 4677
rect 2042 4573 2053 4607
rect 2087 4601 2112 4607
rect 2042 4567 2056 4573
rect 2090 4567 2112 4601
rect 2042 4547 2112 4567
rect 2146 4616 2192 4709
rect 2146 4582 2158 4616
rect 1121 4466 1363 4519
rect 1121 4432 1139 4466
rect 1173 4432 1311 4466
rect 1345 4432 1363 4466
rect 1121 4369 1363 4432
rect 1397 4464 1915 4523
rect 2146 4513 2192 4582
rect 1397 4430 1415 4464
rect 1449 4430 1863 4464
rect 1897 4430 1915 4464
rect 1397 4369 1915 4430
rect 2059 4479 2192 4513
rect 2261 4727 2264 4761
rect 2399 4760 2449 4795
rect 2491 4790 2507 4824
rect 2541 4790 2712 4824
rect 2227 4675 2264 4727
rect 2388 4734 2449 4760
rect 2538 4743 2644 4756
rect 2227 4641 2229 4675
rect 2263 4641 2264 4675
rect 2059 4471 2093 4479
rect 2227 4471 2264 4641
rect 2298 4669 2354 4685
rect 2298 4635 2320 4669
rect 2298 4607 2354 4635
rect 2298 4573 2320 4607
rect 2298 4495 2354 4573
rect 2388 4513 2422 4734
rect 2538 4709 2570 4743
rect 2604 4717 2644 4743
rect 2456 4675 2504 4696
rect 2456 4641 2467 4675
rect 2501 4641 2504 4675
rect 2456 4639 2504 4641
rect 2456 4605 2463 4639
rect 2497 4605 2504 4639
rect 2456 4577 2504 4605
rect 2538 4543 2572 4709
rect 2606 4683 2644 4717
rect 2678 4667 2712 4790
rect 2746 4769 2780 4803
rect 2746 4719 2780 4735
rect 2814 4829 2864 4845
rect 2814 4795 2830 4829
rect 3122 4829 3185 4879
rect 2814 4779 2864 4795
rect 2909 4785 2925 4819
rect 2959 4785 3086 4819
rect 2678 4651 2780 4667
rect 2678 4649 2746 4651
rect 2388 4487 2433 4513
rect 2467 4509 2483 4543
rect 2517 4509 2572 4543
rect 2467 4499 2572 4509
rect 2606 4617 2746 4649
rect 2606 4615 2780 4617
rect 2059 4421 2093 4437
rect 2127 4411 2143 4445
rect 2177 4411 2193 4445
rect 2261 4437 2264 4471
rect 2227 4421 2264 4437
rect 2315 4445 2365 4461
rect 2127 4369 2193 4411
rect 2315 4411 2331 4445
rect 2399 4459 2433 4487
rect 2606 4459 2640 4615
rect 2746 4601 2780 4615
rect 2682 4565 2722 4571
rect 2814 4565 2848 4779
rect 2882 4743 2920 4745
rect 2882 4709 2884 4743
rect 2918 4709 2920 4743
rect 2882 4651 2920 4709
rect 2916 4617 2920 4651
rect 2882 4601 2920 4617
rect 2954 4717 3018 4751
rect 2954 4683 2984 4717
rect 2954 4675 3018 4683
rect 2954 4641 2971 4675
rect 3005 4641 3018 4675
rect 2682 4555 2848 4565
rect 2954 4559 3018 4641
rect 2716 4521 2848 4555
rect 2682 4505 2848 4521
rect 2399 4425 2416 4459
rect 2450 4425 2466 4459
rect 2505 4425 2527 4459
rect 2561 4425 2640 4459
rect 2704 4453 2778 4469
rect 2315 4369 2365 4411
rect 2704 4419 2726 4453
rect 2760 4419 2778 4453
rect 2814 4459 2848 4505
rect 2925 4543 3018 4559
rect 2959 4509 3018 4543
rect 2925 4493 3018 4509
rect 3052 4617 3086 4785
rect 3122 4795 3124 4829
rect 3158 4795 3185 4829
rect 3122 4779 3185 4795
rect 3231 4837 3299 4845
rect 3231 4803 3247 4837
rect 3281 4803 3299 4837
rect 3231 4766 3299 4803
rect 3231 4733 3247 4766
rect 3120 4732 3247 4733
rect 3281 4732 3299 4766
rect 3120 4717 3299 4732
rect 3154 4695 3299 4717
rect 3154 4683 3247 4695
rect 3120 4661 3247 4683
rect 3281 4661 3299 4695
rect 3333 4807 3367 4879
rect 3333 4727 3367 4773
rect 3333 4677 3367 4693
rect 3401 4831 3467 4836
rect 3401 4797 3417 4831
rect 3451 4797 3467 4831
rect 3401 4763 3467 4797
rect 3401 4729 3417 4763
rect 3451 4729 3467 4763
rect 3401 4695 3467 4729
rect 3120 4658 3299 4661
rect 3261 4617 3299 4658
rect 3401 4661 3417 4695
rect 3451 4667 3467 4695
rect 3697 4808 3755 4879
rect 3697 4774 3709 4808
rect 3743 4774 3755 4808
rect 3697 4715 3755 4774
rect 3697 4681 3709 4715
rect 3743 4681 3755 4715
rect 3451 4661 3479 4667
rect 3401 4651 3479 4661
rect 3436 4641 3479 4651
rect 3697 4646 3755 4681
rect 3973 4837 4065 4845
rect 3973 4811 4015 4837
rect 3973 4777 3985 4811
rect 4049 4803 4065 4837
rect 4019 4777 4065 4803
rect 3973 4769 4065 4777
rect 3973 4735 4015 4769
rect 4049 4735 4065 4769
rect 4103 4837 4169 4879
rect 4103 4803 4119 4837
rect 4153 4803 4169 4837
rect 4103 4769 4169 4803
rect 4103 4735 4119 4769
rect 4153 4735 4169 4769
rect 4209 4795 4269 4811
rect 4209 4761 4227 4795
rect 4261 4761 4269 4795
rect 3052 4601 3227 4617
rect 3052 4567 3193 4601
rect 3052 4551 3227 4567
rect 3261 4601 3411 4617
rect 3261 4567 3377 4601
rect 3261 4551 3411 4567
rect 3052 4459 3086 4551
rect 3261 4517 3301 4551
rect 3445 4525 3479 4641
rect 3434 4517 3479 4525
rect 3235 4514 3301 4517
rect 3235 4480 3251 4514
rect 3285 4480 3301 4514
rect 3403 4516 3479 4517
rect 2814 4425 2845 4459
rect 2879 4425 2895 4459
rect 2929 4425 2948 4459
rect 2982 4425 3086 4459
rect 3141 4459 3183 4475
rect 3141 4425 3146 4459
rect 3180 4425 3183 4459
rect 2704 4369 2778 4419
rect 3141 4369 3183 4425
rect 3235 4446 3301 4480
rect 3235 4412 3251 4446
rect 3285 4412 3301 4446
rect 3335 4475 3369 4491
rect 3335 4369 3369 4441
rect 3403 4482 3419 4516
rect 3453 4500 3479 4516
rect 3453 4482 3469 4500
rect 3403 4471 3469 4482
rect 3403 4448 3433 4471
rect 3403 4414 3419 4448
rect 3467 4437 3469 4471
rect 3453 4414 3469 4437
rect 3403 4413 3469 4414
rect 3697 4497 3755 4514
rect 3697 4463 3709 4497
rect 3743 4463 3755 4497
rect 3697 4369 3755 4463
rect 3973 4461 4023 4735
rect 4209 4701 4269 4761
rect 4303 4795 4359 4879
rect 4303 4761 4311 4795
rect 4345 4761 4359 4795
rect 4303 4745 4359 4761
rect 4433 4837 4767 4879
rect 4433 4803 4451 4837
rect 4485 4803 4715 4837
rect 4749 4803 4767 4837
rect 4081 4667 4269 4701
rect 4433 4735 4767 4803
rect 4433 4701 4451 4735
rect 4485 4701 4715 4735
rect 4749 4701 4767 4735
rect 4343 4675 4396 4689
rect 4081 4617 4115 4667
rect 4343 4641 4353 4675
rect 4387 4641 4396 4675
rect 4433 4661 4767 4701
rect 4343 4617 4396 4641
rect 4057 4601 4115 4617
rect 4057 4567 4059 4601
rect 4093 4567 4115 4601
rect 4149 4607 4217 4617
rect 4149 4601 4169 4607
rect 4149 4567 4167 4601
rect 4203 4573 4217 4607
rect 4201 4567 4217 4573
rect 4261 4601 4396 4617
rect 4261 4567 4308 4601
rect 4342 4567 4396 4601
rect 4433 4593 4453 4627
rect 4487 4593 4583 4627
rect 4057 4551 4115 4567
rect 4081 4533 4115 4551
rect 4081 4495 4359 4533
rect 4293 4473 4359 4495
rect 3973 4445 4085 4461
rect 3973 4411 4035 4445
rect 4069 4411 4085 4445
rect 3973 4403 4085 4411
rect 4119 4445 4169 4461
rect 4153 4411 4169 4445
rect 4293 4439 4311 4473
rect 4345 4439 4359 4473
rect 4293 4423 4359 4439
rect 4433 4523 4583 4593
rect 4617 4591 4767 4661
rect 4617 4557 4713 4591
rect 4747 4557 4767 4591
rect 4893 4829 4949 4845
rect 4893 4795 4915 4829
rect 4893 4761 4949 4795
rect 4893 4727 4915 4761
rect 4893 4693 4949 4727
rect 4983 4837 5125 4879
rect 4983 4803 5001 4837
rect 5035 4803 5075 4837
rect 5109 4803 5125 4837
rect 4983 4769 5125 4803
rect 4983 4735 5001 4769
rect 5035 4735 5075 4769
rect 5109 4735 5125 4769
rect 4983 4724 5125 4735
rect 5159 4837 5225 4845
rect 5159 4803 5175 4837
rect 5209 4803 5225 4837
rect 5343 4837 5409 4879
rect 5159 4769 5225 4803
rect 5159 4735 5175 4769
rect 5209 4735 5225 4769
rect 4893 4659 4915 4693
rect 5159 4701 5225 4735
rect 5159 4690 5175 4701
rect 4893 4558 4949 4659
rect 4995 4667 5175 4690
rect 5209 4667 5225 4701
rect 4995 4647 5225 4667
rect 5264 4811 5307 4830
rect 5264 4777 5273 4811
rect 4995 4601 5052 4647
rect 5029 4567 5052 4601
rect 5089 4607 5183 4613
rect 5264 4607 5307 4777
rect 5343 4803 5359 4837
rect 5393 4803 5409 4837
rect 5343 4769 5409 4803
rect 5343 4735 5359 4769
rect 5393 4735 5409 4769
rect 5445 4837 5779 4879
rect 5445 4803 5463 4837
rect 5497 4803 5727 4837
rect 5761 4803 5779 4837
rect 5445 4735 5779 4803
rect 5445 4701 5463 4735
rect 5497 4701 5727 4735
rect 5761 4701 5779 4735
rect 5365 4641 5377 4675
rect 5445 4661 5779 4701
rect 5365 4607 5411 4641
rect 5123 4601 5183 4607
rect 5123 4573 5133 4601
rect 5089 4567 5133 4573
rect 5167 4567 5183 4601
rect 5217 4601 5307 4607
rect 5217 4567 5233 4601
rect 5267 4571 5307 4601
rect 5345 4601 5411 4607
rect 5267 4567 5283 4571
rect 5345 4567 5361 4601
rect 5395 4567 5411 4601
rect 5445 4593 5465 4627
rect 5499 4593 5595 4627
rect 4433 4471 4767 4523
rect 4433 4437 4451 4471
rect 4485 4437 4715 4471
rect 4749 4437 4767 4471
rect 4119 4369 4169 4411
rect 4433 4369 4767 4437
rect 4893 4516 4961 4558
rect 4893 4482 4911 4516
rect 4945 4482 4961 4516
rect 4995 4533 5052 4567
rect 4995 4517 5137 4533
rect 4995 4495 5099 4517
rect 4893 4471 4961 4482
rect 4893 4437 4905 4471
rect 4939 4448 4961 4471
rect 5077 4483 5099 4495
rect 5133 4483 5137 4517
rect 5077 4467 5137 4483
rect 5175 4517 5411 4533
rect 5175 4513 5359 4517
rect 5175 4479 5191 4513
rect 5225 4495 5359 4513
rect 5225 4479 5241 4495
rect 5343 4483 5359 4495
rect 5393 4483 5411 4517
rect 5077 4465 5140 4467
rect 5077 4463 5142 4465
rect 5077 4462 5144 4463
rect 4893 4414 4911 4437
rect 4945 4414 4961 4448
rect 4893 4403 4961 4414
rect 4995 4445 5029 4461
rect 4995 4369 5029 4411
rect 5077 4460 5145 4462
rect 5077 4459 5146 4460
rect 5077 4457 5147 4459
rect 5077 4456 5148 4457
rect 5077 4449 5149 4456
rect 5077 4415 5099 4449
rect 5133 4415 5149 4449
rect 5077 4403 5149 4415
rect 5275 4445 5309 4461
rect 5275 4369 5309 4411
rect 5343 4449 5411 4483
rect 5343 4415 5359 4449
rect 5393 4415 5411 4449
rect 5343 4403 5411 4415
rect 5445 4523 5595 4593
rect 5629 4591 5779 4661
rect 5629 4557 5725 4591
rect 5759 4557 5779 4591
rect 5813 4829 5869 4845
rect 5813 4795 5835 4829
rect 5813 4761 5869 4795
rect 5813 4727 5835 4761
rect 5813 4693 5869 4727
rect 5903 4837 6045 4879
rect 5903 4803 5921 4837
rect 5955 4803 5995 4837
rect 6029 4803 6045 4837
rect 5903 4769 6045 4803
rect 5903 4735 5921 4769
rect 5955 4735 5995 4769
rect 6029 4735 6045 4769
rect 5903 4724 6045 4735
rect 6079 4837 6145 4845
rect 6079 4803 6095 4837
rect 6129 4803 6145 4837
rect 6263 4837 6329 4879
rect 6079 4769 6145 4803
rect 6079 4735 6095 4769
rect 6129 4735 6145 4769
rect 5813 4659 5835 4693
rect 6079 4701 6145 4735
rect 6079 4690 6095 4701
rect 5813 4558 5869 4659
rect 5915 4667 6095 4690
rect 6129 4667 6145 4701
rect 5915 4647 6145 4667
rect 6184 4811 6227 4830
rect 6184 4777 6193 4811
rect 5915 4601 5972 4647
rect 5949 4567 5972 4601
rect 6009 4607 6103 4613
rect 6184 4607 6227 4777
rect 6263 4803 6279 4837
rect 6313 4803 6329 4837
rect 6263 4769 6329 4803
rect 6263 4735 6279 4769
rect 6313 4735 6329 4769
rect 6365 4837 6699 4879
rect 6365 4803 6383 4837
rect 6417 4803 6647 4837
rect 6681 4803 6699 4837
rect 6365 4735 6699 4803
rect 6365 4701 6383 4735
rect 6417 4701 6647 4735
rect 6681 4701 6699 4735
rect 6751 4829 6785 4845
rect 6751 4761 6785 4795
rect 6819 4813 6885 4879
rect 6819 4779 6835 4813
rect 6869 4779 6885 4813
rect 6919 4829 6956 4845
rect 6953 4795 6956 4829
rect 6919 4761 6956 4795
rect 7004 4837 7057 4879
rect 7004 4803 7023 4837
rect 7004 4787 7057 4803
rect 7091 4829 7141 4845
rect 7091 4795 7107 4829
rect 7438 4837 7472 4879
rect 6785 4743 6884 4745
rect 6785 4727 6842 4743
rect 6751 4711 6842 4727
rect 6319 4641 6331 4675
rect 6365 4661 6699 4701
rect 6838 4709 6842 4711
rect 6876 4709 6884 4743
rect 6285 4607 6331 4641
rect 6043 4601 6103 4607
rect 6043 4573 6053 4601
rect 6009 4567 6053 4573
rect 6087 4567 6103 4601
rect 6137 4601 6227 4607
rect 6137 4567 6153 4601
rect 6187 4571 6227 4601
rect 6265 4601 6331 4607
rect 6187 4567 6203 4571
rect 6265 4567 6281 4601
rect 6315 4567 6331 4601
rect 6365 4593 6385 4627
rect 6419 4593 6515 4627
rect 5445 4471 5779 4523
rect 5445 4437 5463 4471
rect 5497 4437 5727 4471
rect 5761 4437 5779 4471
rect 5445 4369 5779 4437
rect 5813 4516 5881 4558
rect 5813 4482 5831 4516
rect 5865 4482 5881 4516
rect 5915 4533 5972 4567
rect 5915 4517 6057 4533
rect 5915 4495 6019 4517
rect 5813 4471 5881 4482
rect 5813 4437 5825 4471
rect 5859 4448 5881 4471
rect 5997 4483 6019 4495
rect 6053 4483 6057 4517
rect 5997 4467 6057 4483
rect 6095 4517 6331 4533
rect 6095 4513 6279 4517
rect 6095 4479 6111 4513
rect 6145 4495 6279 4513
rect 6145 4479 6161 4495
rect 6263 4483 6279 4495
rect 6313 4483 6331 4517
rect 5997 4465 6060 4467
rect 5997 4463 6062 4465
rect 5997 4462 6064 4463
rect 5813 4414 5831 4437
rect 5865 4414 5881 4448
rect 5813 4403 5881 4414
rect 5915 4445 5949 4461
rect 5915 4369 5949 4411
rect 5997 4460 6065 4462
rect 5997 4459 6066 4460
rect 5997 4457 6067 4459
rect 5997 4456 6068 4457
rect 5997 4449 6069 4456
rect 5997 4415 6019 4449
rect 6053 4415 6069 4449
rect 5997 4403 6069 4415
rect 6195 4445 6229 4461
rect 6195 4369 6229 4411
rect 6263 4449 6331 4483
rect 6263 4415 6279 4449
rect 6313 4415 6331 4449
rect 6263 4403 6331 4415
rect 6365 4523 6515 4593
rect 6549 4591 6699 4661
rect 6549 4557 6645 4591
rect 6679 4557 6699 4591
rect 6734 4607 6804 4677
rect 6734 4573 6745 4607
rect 6779 4601 6804 4607
rect 6734 4567 6748 4573
rect 6782 4567 6804 4601
rect 6734 4547 6804 4567
rect 6838 4616 6884 4709
rect 6838 4582 6850 4616
rect 6365 4471 6699 4523
rect 6838 4513 6884 4582
rect 6365 4437 6383 4471
rect 6417 4437 6647 4471
rect 6681 4437 6699 4471
rect 6365 4369 6699 4437
rect 6751 4479 6884 4513
rect 6953 4727 6956 4761
rect 7091 4760 7141 4795
rect 7183 4790 7199 4824
rect 7233 4790 7404 4824
rect 6919 4675 6956 4727
rect 7080 4734 7141 4760
rect 7230 4743 7336 4756
rect 6919 4641 6921 4675
rect 6955 4641 6956 4675
rect 6751 4471 6785 4479
rect 6919 4471 6956 4641
rect 6990 4669 7046 4685
rect 6990 4635 7012 4669
rect 6990 4607 7046 4635
rect 6990 4573 7012 4607
rect 6990 4495 7046 4573
rect 7080 4513 7114 4734
rect 7230 4709 7262 4743
rect 7296 4717 7336 4743
rect 7148 4675 7196 4696
rect 7148 4641 7159 4675
rect 7193 4641 7196 4675
rect 7148 4639 7196 4641
rect 7148 4605 7155 4639
rect 7189 4605 7196 4639
rect 7148 4577 7196 4605
rect 7230 4543 7264 4709
rect 7298 4683 7336 4717
rect 7370 4667 7404 4790
rect 7438 4769 7472 4803
rect 7438 4719 7472 4735
rect 7506 4829 7556 4845
rect 7506 4795 7522 4829
rect 7814 4829 7877 4879
rect 7506 4779 7556 4795
rect 7601 4785 7617 4819
rect 7651 4785 7778 4819
rect 7370 4651 7472 4667
rect 7370 4649 7438 4651
rect 7080 4487 7125 4513
rect 7159 4509 7175 4543
rect 7209 4509 7264 4543
rect 7159 4499 7264 4509
rect 7298 4617 7438 4649
rect 7298 4615 7472 4617
rect 6751 4421 6785 4437
rect 6819 4411 6835 4445
rect 6869 4411 6885 4445
rect 6953 4437 6956 4471
rect 6919 4421 6956 4437
rect 7007 4445 7057 4461
rect 6819 4369 6885 4411
rect 7007 4411 7023 4445
rect 7091 4459 7125 4487
rect 7298 4459 7332 4615
rect 7438 4601 7472 4615
rect 7374 4565 7414 4571
rect 7506 4565 7540 4779
rect 7574 4743 7612 4745
rect 7574 4709 7576 4743
rect 7610 4709 7612 4743
rect 7574 4651 7612 4709
rect 7608 4617 7612 4651
rect 7574 4601 7612 4617
rect 7646 4717 7710 4751
rect 7646 4683 7676 4717
rect 7646 4675 7710 4683
rect 7646 4641 7663 4675
rect 7697 4641 7710 4675
rect 7374 4555 7540 4565
rect 7646 4559 7710 4641
rect 7408 4521 7540 4555
rect 7374 4505 7540 4521
rect 7091 4425 7108 4459
rect 7142 4425 7158 4459
rect 7197 4425 7219 4459
rect 7253 4425 7332 4459
rect 7396 4453 7470 4469
rect 7007 4369 7057 4411
rect 7396 4419 7418 4453
rect 7452 4419 7470 4453
rect 7506 4459 7540 4505
rect 7617 4543 7710 4559
rect 7651 4509 7710 4543
rect 7617 4493 7710 4509
rect 7744 4617 7778 4785
rect 7814 4795 7816 4829
rect 7850 4795 7877 4829
rect 7814 4779 7877 4795
rect 7923 4837 7991 4845
rect 7923 4803 7939 4837
rect 7973 4803 7991 4837
rect 7923 4766 7991 4803
rect 7923 4733 7939 4766
rect 7812 4732 7939 4733
rect 7973 4732 7991 4766
rect 7812 4717 7991 4732
rect 7846 4695 7991 4717
rect 7846 4683 7939 4695
rect 7812 4661 7939 4683
rect 7973 4661 7991 4695
rect 8025 4807 8059 4879
rect 8205 4837 8723 4879
rect 8025 4727 8059 4773
rect 8025 4677 8059 4693
rect 8093 4831 8159 4836
rect 8093 4797 8109 4831
rect 8143 4797 8159 4831
rect 8093 4763 8159 4797
rect 8093 4729 8109 4763
rect 8143 4729 8159 4763
rect 8093 4695 8159 4729
rect 7812 4658 7991 4661
rect 7953 4617 7991 4658
rect 8093 4661 8109 4695
rect 8143 4667 8159 4695
rect 8205 4803 8223 4837
rect 8257 4803 8671 4837
rect 8705 4803 8723 4837
rect 8205 4735 8723 4803
rect 8205 4701 8223 4735
rect 8257 4701 8671 4735
rect 8705 4701 8723 4735
rect 8143 4661 8171 4667
rect 8205 4661 8723 4701
rect 8093 4651 8171 4661
rect 8128 4641 8171 4651
rect 7744 4601 7919 4617
rect 7744 4567 7885 4601
rect 7744 4551 7919 4567
rect 7953 4601 8103 4617
rect 7953 4567 8069 4601
rect 7953 4551 8103 4567
rect 7744 4459 7778 4551
rect 7953 4517 7993 4551
rect 8137 4525 8171 4641
rect 8126 4517 8171 4525
rect 7927 4514 7993 4517
rect 7927 4480 7943 4514
rect 7977 4480 7993 4514
rect 8095 4516 8171 4517
rect 7506 4425 7537 4459
rect 7571 4425 7587 4459
rect 7621 4425 7640 4459
rect 7674 4425 7778 4459
rect 7833 4459 7875 4475
rect 7833 4425 7838 4459
rect 7872 4425 7875 4459
rect 7396 4369 7470 4419
rect 7833 4369 7875 4425
rect 7927 4446 7993 4480
rect 7927 4412 7943 4446
rect 7977 4412 7993 4446
rect 8027 4475 8061 4491
rect 8027 4369 8061 4441
rect 8095 4482 8111 4516
rect 8145 4500 8171 4516
rect 8205 4593 8283 4627
rect 8317 4593 8393 4627
rect 8427 4593 8447 4627
rect 8205 4523 8447 4593
rect 8481 4591 8723 4661
rect 8849 4808 8907 4879
rect 8849 4774 8861 4808
rect 8895 4774 8907 4808
rect 8849 4715 8907 4774
rect 8849 4681 8861 4715
rect 8895 4681 8907 4715
rect 8849 4646 8907 4681
rect 8941 4837 9643 4879
rect 8941 4803 8959 4837
rect 8993 4803 9591 4837
rect 9625 4803 9643 4837
rect 8941 4735 9643 4803
rect 8941 4701 8959 4735
rect 8993 4701 9591 4735
rect 9625 4701 9643 4735
rect 8941 4661 9643 4701
rect 9677 4837 9919 4879
rect 9677 4803 9695 4837
rect 9729 4803 9867 4837
rect 9901 4803 9919 4837
rect 9677 4742 9919 4803
rect 9677 4708 9695 4742
rect 9729 4708 9867 4742
rect 9901 4708 9919 4742
rect 9677 4661 9919 4708
rect 9965 4831 10031 4836
rect 9965 4811 9981 4831
rect 10015 4797 10031 4831
rect 9999 4777 10031 4797
rect 9965 4763 10031 4777
rect 9965 4729 9981 4763
rect 10015 4729 10031 4763
rect 9965 4695 10031 4729
rect 9965 4667 9981 4695
rect 8481 4557 8501 4591
rect 8535 4557 8611 4591
rect 8645 4557 8723 4591
rect 8941 4593 9019 4627
rect 9053 4593 9118 4627
rect 9152 4593 9217 4627
rect 9251 4593 9271 4627
rect 8941 4523 9271 4593
rect 9305 4591 9643 4661
rect 9305 4557 9325 4591
rect 9359 4557 9428 4591
rect 9462 4557 9531 4591
rect 9565 4557 9643 4591
rect 9677 4593 9727 4627
rect 9761 4593 9781 4627
rect 8145 4482 8161 4500
rect 8095 4471 8161 4482
rect 8095 4448 8125 4471
rect 8095 4414 8111 4448
rect 8159 4437 8161 4471
rect 8145 4414 8161 4437
rect 8095 4413 8161 4414
rect 8205 4464 8723 4523
rect 8205 4430 8223 4464
rect 8257 4430 8671 4464
rect 8705 4430 8723 4464
rect 8205 4369 8723 4430
rect 8849 4497 8907 4514
rect 8849 4463 8861 4497
rect 8895 4463 8907 4497
rect 8849 4369 8907 4463
rect 8941 4464 9643 4523
rect 8941 4430 8959 4464
rect 8993 4430 9591 4464
rect 9625 4430 9643 4464
rect 8941 4369 9643 4430
rect 9677 4519 9781 4593
rect 9815 4587 9919 4661
rect 9815 4553 9835 4587
rect 9869 4553 9919 4587
rect 9953 4661 9981 4667
rect 10015 4661 10031 4695
rect 10065 4807 10099 4879
rect 10065 4727 10099 4773
rect 10065 4677 10099 4693
rect 10133 4837 10201 4845
rect 10133 4803 10151 4837
rect 10185 4803 10201 4837
rect 10133 4766 10201 4803
rect 10247 4829 10310 4879
rect 10247 4795 10274 4829
rect 10308 4795 10310 4829
rect 10568 4829 10618 4845
rect 10247 4779 10310 4795
rect 10346 4785 10473 4819
rect 10507 4785 10523 4819
rect 10602 4795 10618 4829
rect 10133 4732 10151 4766
rect 10185 4733 10201 4766
rect 10185 4732 10312 4733
rect 10133 4717 10312 4732
rect 10133 4695 10278 4717
rect 9953 4651 10031 4661
rect 10133 4661 10151 4695
rect 10185 4683 10278 4695
rect 10185 4661 10312 4683
rect 10133 4658 10312 4661
rect 9953 4641 9996 4651
rect 9953 4525 9987 4641
rect 10133 4617 10171 4658
rect 10346 4617 10380 4785
rect 10568 4779 10618 4795
rect 10021 4601 10171 4617
rect 10055 4567 10171 4601
rect 10021 4551 10171 4567
rect 10205 4601 10380 4617
rect 10239 4567 10380 4601
rect 10205 4551 10380 4567
rect 9677 4466 9919 4519
rect 9953 4517 9998 4525
rect 10131 4517 10171 4551
rect 9953 4516 10029 4517
rect 9953 4500 9979 4516
rect 9677 4432 9695 4466
rect 9729 4432 9867 4466
rect 9901 4432 9919 4466
rect 9677 4369 9919 4432
rect 9963 4482 9979 4500
rect 10013 4482 10029 4516
rect 10131 4514 10197 4517
rect 9963 4448 10029 4482
rect 9963 4414 9979 4448
rect 10013 4414 10029 4448
rect 9963 4413 10029 4414
rect 10063 4475 10097 4491
rect 10063 4369 10097 4441
rect 10131 4480 10147 4514
rect 10181 4480 10197 4514
rect 10131 4446 10197 4480
rect 10131 4412 10147 4446
rect 10181 4412 10197 4446
rect 10249 4459 10291 4475
rect 10249 4425 10252 4459
rect 10286 4425 10291 4459
rect 10346 4459 10380 4551
rect 10414 4717 10478 4751
rect 10448 4683 10478 4717
rect 10414 4675 10478 4683
rect 10414 4641 10427 4675
rect 10461 4641 10478 4675
rect 10414 4559 10478 4641
rect 10512 4743 10550 4745
rect 10512 4709 10514 4743
rect 10548 4709 10550 4743
rect 10512 4651 10550 4709
rect 10512 4617 10516 4651
rect 10512 4601 10550 4617
rect 10584 4565 10618 4779
rect 10652 4837 10686 4879
rect 10983 4829 11033 4845
rect 10652 4769 10686 4803
rect 10652 4719 10686 4735
rect 10720 4790 10891 4824
rect 10925 4790 10941 4824
rect 11017 4795 11033 4829
rect 10720 4667 10754 4790
rect 10983 4760 11033 4795
rect 11067 4837 11120 4879
rect 11101 4803 11120 4837
rect 11067 4787 11120 4803
rect 11168 4829 11205 4845
rect 11168 4795 11171 4829
rect 11168 4761 11205 4795
rect 11239 4813 11305 4879
rect 11239 4779 11255 4813
rect 11289 4779 11305 4813
rect 11339 4829 11373 4845
rect 10788 4743 10894 4756
rect 10788 4717 10828 4743
rect 10788 4683 10826 4717
rect 10862 4709 10894 4743
rect 10983 4734 11044 4760
rect 10652 4651 10754 4667
rect 10686 4649 10754 4651
rect 10686 4617 10826 4649
rect 10652 4615 10826 4617
rect 10652 4601 10686 4615
rect 10710 4565 10750 4571
rect 10414 4543 10507 4559
rect 10414 4509 10473 4543
rect 10414 4493 10507 4509
rect 10584 4555 10750 4565
rect 10584 4521 10716 4555
rect 10584 4505 10750 4521
rect 10584 4459 10618 4505
rect 10346 4425 10450 4459
rect 10484 4425 10503 4459
rect 10537 4425 10553 4459
rect 10587 4425 10618 4459
rect 10654 4453 10728 4469
rect 10249 4369 10291 4425
rect 10654 4419 10672 4453
rect 10706 4419 10728 4453
rect 10792 4459 10826 4615
rect 10860 4543 10894 4709
rect 10928 4675 10976 4696
rect 10928 4641 10931 4675
rect 10965 4641 10976 4675
rect 10928 4639 10976 4641
rect 10928 4605 10935 4639
rect 10969 4605 10976 4639
rect 10928 4577 10976 4605
rect 10860 4509 10915 4543
rect 10949 4509 10965 4543
rect 11010 4513 11044 4734
rect 11168 4727 11171 4761
rect 11339 4761 11373 4795
rect 10860 4499 10965 4509
rect 10999 4487 11044 4513
rect 11078 4669 11134 4685
rect 11112 4635 11134 4669
rect 11078 4539 11134 4635
rect 11078 4505 11100 4539
rect 11078 4495 11134 4505
rect 11168 4675 11205 4727
rect 11168 4641 11169 4675
rect 11203 4641 11205 4675
rect 10999 4459 11033 4487
rect 11168 4471 11205 4641
rect 11240 4743 11339 4745
rect 11240 4709 11248 4743
rect 11282 4727 11339 4743
rect 11282 4711 11373 4727
rect 11425 4837 11759 4879
rect 11425 4803 11443 4837
rect 11477 4803 11707 4837
rect 11741 4803 11759 4837
rect 11425 4735 11759 4803
rect 11282 4709 11286 4711
rect 11240 4616 11286 4709
rect 11425 4701 11443 4735
rect 11477 4701 11707 4735
rect 11741 4701 11759 4735
rect 11274 4582 11286 4616
rect 11240 4513 11286 4582
rect 11320 4607 11390 4677
rect 11425 4661 11759 4701
rect 11320 4601 11345 4607
rect 11320 4567 11342 4601
rect 11379 4573 11390 4607
rect 11376 4567 11390 4573
rect 11320 4547 11390 4567
rect 11425 4593 11445 4627
rect 11479 4593 11575 4627
rect 11425 4523 11575 4593
rect 11609 4591 11759 4661
rect 11609 4557 11705 4591
rect 11739 4557 11759 4591
rect 11793 4829 11849 4845
rect 11793 4795 11815 4829
rect 11793 4761 11849 4795
rect 11793 4727 11815 4761
rect 11793 4693 11849 4727
rect 11883 4837 12025 4879
rect 11883 4803 11901 4837
rect 11935 4803 11975 4837
rect 12009 4803 12025 4837
rect 11883 4769 12025 4803
rect 11883 4735 11901 4769
rect 11935 4735 11975 4769
rect 12009 4735 12025 4769
rect 11883 4724 12025 4735
rect 12059 4837 12125 4845
rect 12059 4803 12075 4837
rect 12109 4803 12125 4837
rect 12243 4837 12309 4879
rect 12059 4769 12125 4803
rect 12059 4735 12075 4769
rect 12109 4735 12125 4769
rect 11793 4659 11815 4693
rect 12059 4701 12125 4735
rect 12059 4690 12075 4701
rect 11793 4558 11849 4659
rect 11895 4667 12075 4690
rect 12109 4667 12125 4701
rect 11895 4647 12125 4667
rect 12164 4811 12207 4830
rect 12164 4777 12173 4811
rect 11895 4601 11952 4647
rect 11929 4567 11952 4601
rect 11989 4607 12083 4613
rect 12164 4607 12207 4777
rect 12243 4803 12259 4837
rect 12293 4803 12309 4837
rect 12243 4769 12309 4803
rect 12243 4735 12259 4769
rect 12293 4735 12309 4769
rect 12345 4837 12679 4879
rect 12345 4803 12363 4837
rect 12397 4803 12627 4837
rect 12661 4803 12679 4837
rect 12345 4735 12679 4803
rect 12345 4701 12363 4735
rect 12397 4701 12627 4735
rect 12661 4701 12679 4735
rect 12299 4641 12311 4675
rect 12345 4661 12679 4701
rect 12265 4607 12311 4641
rect 12023 4601 12083 4607
rect 12023 4573 12033 4601
rect 11989 4567 12033 4573
rect 12067 4567 12083 4601
rect 12117 4601 12207 4607
rect 12117 4567 12133 4601
rect 12167 4571 12207 4601
rect 12245 4601 12311 4607
rect 12167 4567 12183 4571
rect 12245 4567 12261 4601
rect 12295 4567 12311 4601
rect 12345 4593 12365 4627
rect 12399 4593 12495 4627
rect 11240 4479 11373 4513
rect 10792 4425 10871 4459
rect 10905 4425 10927 4459
rect 10966 4425 10982 4459
rect 11016 4425 11033 4459
rect 11067 4445 11117 4461
rect 10654 4369 10728 4419
rect 11101 4411 11117 4445
rect 11168 4437 11171 4471
rect 11339 4471 11373 4479
rect 11168 4421 11205 4437
rect 11067 4369 11117 4411
rect 11239 4411 11255 4445
rect 11289 4411 11305 4445
rect 11339 4421 11373 4437
rect 11425 4471 11759 4523
rect 11425 4437 11443 4471
rect 11477 4437 11707 4471
rect 11741 4437 11759 4471
rect 11239 4369 11305 4411
rect 11425 4369 11759 4437
rect 11793 4516 11861 4558
rect 11793 4482 11811 4516
rect 11845 4482 11861 4516
rect 11895 4533 11952 4567
rect 11895 4517 12037 4533
rect 11895 4495 11999 4517
rect 11793 4471 11861 4482
rect 11793 4437 11805 4471
rect 11839 4448 11861 4471
rect 11977 4483 11999 4495
rect 12033 4483 12037 4517
rect 11977 4467 12037 4483
rect 12075 4517 12311 4533
rect 12075 4513 12259 4517
rect 12075 4479 12091 4513
rect 12125 4495 12259 4513
rect 12125 4479 12141 4495
rect 12243 4483 12259 4495
rect 12293 4483 12311 4517
rect 11977 4465 12040 4467
rect 11977 4463 12042 4465
rect 11977 4462 12044 4463
rect 11793 4414 11811 4437
rect 11845 4414 11861 4448
rect 11793 4403 11861 4414
rect 11895 4445 11929 4461
rect 11895 4369 11929 4411
rect 11977 4460 12045 4462
rect 11977 4459 12046 4460
rect 11977 4457 12047 4459
rect 11977 4456 12048 4457
rect 11977 4449 12049 4456
rect 11977 4415 11999 4449
rect 12033 4415 12049 4449
rect 11977 4403 12049 4415
rect 12175 4445 12209 4461
rect 12175 4369 12209 4411
rect 12243 4449 12311 4483
rect 12243 4415 12259 4449
rect 12293 4415 12311 4449
rect 12243 4403 12311 4415
rect 12345 4523 12495 4593
rect 12529 4591 12679 4661
rect 12529 4557 12625 4591
rect 12659 4557 12679 4591
rect 12713 4829 12769 4845
rect 12713 4795 12735 4829
rect 12713 4761 12769 4795
rect 12713 4727 12735 4761
rect 12713 4693 12769 4727
rect 12803 4837 12945 4879
rect 12803 4803 12821 4837
rect 12855 4803 12895 4837
rect 12929 4803 12945 4837
rect 12803 4769 12945 4803
rect 12803 4735 12821 4769
rect 12855 4735 12895 4769
rect 12929 4735 12945 4769
rect 12803 4724 12945 4735
rect 12979 4837 13045 4845
rect 12979 4803 12995 4837
rect 13029 4803 13045 4837
rect 13163 4837 13229 4879
rect 12979 4769 13045 4803
rect 12979 4735 12995 4769
rect 13029 4735 13045 4769
rect 12713 4659 12735 4693
rect 12979 4701 13045 4735
rect 12979 4690 12995 4701
rect 12713 4558 12769 4659
rect 12815 4667 12995 4690
rect 13029 4667 13045 4701
rect 12815 4647 13045 4667
rect 13084 4675 13127 4830
rect 13163 4803 13179 4837
rect 13213 4803 13229 4837
rect 13163 4769 13229 4803
rect 13163 4735 13179 4769
rect 13213 4735 13229 4769
rect 13265 4837 13967 4879
rect 13265 4803 13283 4837
rect 13317 4803 13915 4837
rect 13949 4803 13967 4837
rect 13265 4735 13967 4803
rect 13265 4701 13283 4735
rect 13317 4701 13915 4735
rect 13949 4701 13967 4735
rect 12815 4601 12872 4647
rect 13084 4641 13093 4675
rect 12849 4567 12872 4601
rect 12909 4607 13003 4613
rect 13084 4607 13127 4641
rect 13185 4607 13231 4675
rect 13265 4661 13967 4701
rect 12943 4601 13003 4607
rect 12943 4573 12953 4601
rect 12909 4567 12953 4573
rect 12987 4567 13003 4601
rect 13037 4601 13127 4607
rect 13037 4567 13053 4601
rect 13087 4571 13127 4601
rect 13165 4601 13185 4607
rect 13087 4567 13103 4571
rect 13165 4567 13181 4601
rect 13219 4573 13231 4607
rect 13215 4567 13231 4573
rect 13265 4593 13343 4627
rect 13377 4593 13442 4627
rect 13476 4593 13541 4627
rect 13575 4593 13595 4627
rect 12345 4471 12679 4523
rect 12345 4437 12363 4471
rect 12397 4437 12627 4471
rect 12661 4437 12679 4471
rect 12345 4369 12679 4437
rect 12713 4516 12781 4558
rect 12713 4482 12731 4516
rect 12765 4482 12781 4516
rect 12815 4533 12872 4567
rect 12815 4517 12957 4533
rect 12815 4495 12919 4517
rect 12713 4471 12781 4482
rect 12713 4437 12725 4471
rect 12759 4448 12781 4471
rect 12897 4483 12919 4495
rect 12953 4483 12957 4517
rect 12897 4467 12957 4483
rect 12995 4517 13231 4533
rect 12995 4513 13179 4517
rect 12995 4479 13011 4513
rect 13045 4495 13179 4513
rect 13045 4479 13061 4495
rect 13163 4483 13179 4495
rect 13213 4483 13231 4517
rect 12897 4465 12960 4467
rect 12897 4463 12962 4465
rect 12897 4462 12964 4463
rect 12713 4414 12731 4437
rect 12765 4414 12781 4448
rect 12713 4403 12781 4414
rect 12815 4445 12849 4461
rect 12815 4369 12849 4411
rect 12897 4460 12965 4462
rect 12897 4459 12966 4460
rect 12897 4457 12967 4459
rect 12897 4456 12968 4457
rect 12897 4449 12969 4456
rect 12897 4415 12919 4449
rect 12953 4415 12969 4449
rect 12897 4403 12969 4415
rect 13095 4445 13129 4461
rect 13095 4369 13129 4411
rect 13163 4449 13231 4483
rect 13163 4415 13179 4449
rect 13213 4415 13231 4449
rect 13163 4403 13231 4415
rect 13265 4523 13595 4593
rect 13629 4591 13967 4661
rect 14001 4808 14059 4879
rect 14001 4774 14013 4808
rect 14047 4774 14059 4808
rect 14001 4715 14059 4774
rect 14001 4681 14013 4715
rect 14047 4681 14059 4715
rect 14001 4646 14059 4681
rect 14093 4837 14335 4879
rect 14093 4803 14111 4837
rect 14145 4803 14283 4837
rect 14317 4803 14335 4837
rect 14093 4742 14335 4803
rect 14409 4795 14465 4879
rect 14599 4837 14665 4879
rect 14409 4761 14423 4795
rect 14457 4761 14465 4795
rect 14409 4745 14465 4761
rect 14499 4795 14559 4811
rect 14499 4761 14507 4795
rect 14541 4761 14559 4795
rect 14093 4708 14111 4742
rect 14145 4708 14283 4742
rect 14317 4708 14335 4742
rect 14093 4661 14335 4708
rect 14499 4701 14559 4761
rect 14599 4803 14615 4837
rect 14649 4803 14665 4837
rect 14599 4769 14665 4803
rect 14599 4735 14615 4769
rect 14649 4735 14665 4769
rect 14703 4837 14795 4845
rect 14703 4803 14719 4837
rect 14753 4803 14795 4837
rect 14703 4769 14795 4803
rect 14829 4837 15898 4879
rect 14829 4803 14847 4837
rect 14881 4803 15847 4837
rect 15881 4803 15898 4837
rect 14829 4792 15898 4803
rect 15933 4837 17002 4879
rect 15933 4803 15951 4837
rect 15985 4803 16951 4837
rect 16985 4803 17002 4837
rect 15933 4792 17002 4803
rect 17037 4837 18106 4879
rect 17037 4803 17055 4837
rect 17089 4803 18055 4837
rect 18089 4803 18106 4837
rect 17037 4792 18106 4803
rect 18141 4837 18475 4879
rect 18141 4803 18159 4837
rect 18193 4803 18423 4837
rect 18457 4803 18475 4837
rect 14703 4735 14719 4769
rect 14753 4735 14795 4769
rect 13629 4557 13649 4591
rect 13683 4557 13752 4591
rect 13786 4557 13855 4591
rect 13889 4557 13967 4591
rect 14093 4593 14143 4627
rect 14177 4593 14197 4627
rect 13265 4464 13967 4523
rect 14093 4519 14197 4593
rect 14231 4587 14335 4661
rect 14231 4553 14251 4587
rect 14285 4553 14335 4587
rect 14372 4617 14425 4689
rect 14499 4667 14687 4701
rect 14653 4617 14687 4667
rect 14372 4607 14507 4617
rect 14372 4573 14381 4607
rect 14415 4601 14507 4607
rect 14415 4573 14426 4601
rect 14372 4567 14426 4573
rect 14460 4567 14507 4601
rect 14551 4607 14619 4617
rect 14551 4573 14565 4607
rect 14599 4601 14619 4607
rect 14551 4567 14567 4573
rect 14601 4567 14619 4601
rect 14653 4601 14711 4617
rect 14653 4567 14675 4601
rect 14709 4567 14711 4601
rect 14653 4551 14711 4567
rect 14653 4533 14687 4551
rect 13265 4430 13283 4464
rect 13317 4430 13915 4464
rect 13949 4430 13967 4464
rect 13265 4369 13967 4430
rect 14001 4497 14059 4514
rect 14001 4463 14013 4497
rect 14047 4463 14059 4497
rect 14001 4369 14059 4463
rect 14093 4466 14335 4519
rect 14093 4432 14111 4466
rect 14145 4432 14283 4466
rect 14317 4432 14335 4466
rect 14093 4369 14335 4432
rect 14409 4495 14687 4533
rect 14409 4473 14475 4495
rect 14409 4439 14423 4473
rect 14457 4439 14475 4473
rect 14745 4471 14795 4735
rect 15146 4627 15214 4644
rect 15146 4593 15163 4627
rect 15197 4593 15214 4627
rect 15146 4478 15214 4593
rect 15510 4591 15580 4792
rect 15510 4557 15527 4591
rect 15561 4557 15580 4591
rect 15510 4542 15580 4557
rect 16250 4627 16318 4644
rect 16250 4593 16267 4627
rect 16301 4593 16318 4627
rect 16250 4478 16318 4593
rect 16614 4591 16684 4792
rect 16614 4557 16631 4591
rect 16665 4557 16684 4591
rect 16614 4542 16684 4557
rect 17354 4627 17422 4644
rect 17354 4593 17371 4627
rect 17405 4593 17422 4627
rect 17354 4478 17422 4593
rect 17718 4591 17788 4792
rect 18141 4735 18475 4803
rect 18141 4701 18159 4735
rect 18193 4701 18423 4735
rect 18457 4701 18475 4735
rect 18141 4661 18475 4701
rect 17718 4557 17735 4591
rect 17769 4557 17788 4591
rect 17718 4542 17788 4557
rect 18141 4593 18161 4627
rect 18195 4593 18291 4627
rect 18141 4523 18291 4593
rect 18325 4591 18475 4661
rect 18325 4557 18421 4591
rect 18455 4557 18475 4591
rect 18601 4837 18843 4879
rect 18601 4803 18619 4837
rect 18653 4803 18791 4837
rect 18825 4803 18843 4837
rect 18601 4742 18843 4803
rect 18601 4708 18619 4742
rect 18653 4708 18791 4742
rect 18825 4708 18843 4742
rect 18601 4661 18843 4708
rect 18601 4587 18705 4661
rect 18601 4553 18651 4587
rect 18685 4553 18705 4587
rect 18739 4593 18759 4627
rect 18793 4593 18843 4627
rect 14745 4461 14749 4471
rect 14409 4423 14475 4439
rect 14599 4445 14649 4461
rect 14599 4411 14615 4445
rect 14599 4369 14649 4411
rect 14683 4445 14749 4461
rect 14683 4411 14699 4445
rect 14733 4437 14749 4445
rect 14783 4437 14795 4471
rect 14733 4411 14795 4437
rect 14683 4403 14795 4411
rect 14829 4464 15898 4478
rect 14829 4430 14847 4464
rect 14881 4430 15847 4464
rect 15881 4430 15898 4464
rect 14829 4369 15898 4430
rect 15933 4464 17002 4478
rect 15933 4430 15951 4464
rect 15985 4430 16951 4464
rect 16985 4430 17002 4464
rect 15933 4369 17002 4430
rect 17037 4464 18106 4478
rect 17037 4430 17055 4464
rect 17089 4430 18055 4464
rect 18089 4430 18106 4464
rect 17037 4369 18106 4430
rect 18141 4471 18475 4523
rect 18739 4519 18843 4593
rect 18141 4437 18159 4471
rect 18193 4437 18423 4471
rect 18457 4437 18475 4471
rect 18141 4369 18475 4437
rect 18601 4466 18843 4519
rect 18601 4432 18619 4466
rect 18653 4432 18791 4466
rect 18825 4432 18843 4466
rect 18601 4369 18843 4432
rect 1104 4335 1133 4369
rect 1167 4335 1225 4369
rect 1259 4335 1317 4369
rect 1351 4335 1409 4369
rect 1443 4335 1501 4369
rect 1535 4335 1593 4369
rect 1627 4335 1685 4369
rect 1719 4335 1777 4369
rect 1811 4335 1869 4369
rect 1903 4335 1961 4369
rect 1995 4335 2053 4369
rect 2087 4335 2145 4369
rect 2179 4335 2237 4369
rect 2271 4335 2329 4369
rect 2363 4335 2421 4369
rect 2455 4335 2513 4369
rect 2547 4335 2605 4369
rect 2639 4335 2697 4369
rect 2731 4335 2789 4369
rect 2823 4335 2881 4369
rect 2915 4335 2973 4369
rect 3007 4335 3065 4369
rect 3099 4335 3157 4369
rect 3191 4335 3249 4369
rect 3283 4335 3341 4369
rect 3375 4335 3433 4369
rect 3467 4335 3525 4369
rect 3559 4335 3617 4369
rect 3651 4335 3709 4369
rect 3743 4335 3801 4369
rect 3835 4335 3893 4369
rect 3927 4335 3985 4369
rect 4019 4335 4077 4369
rect 4111 4335 4169 4369
rect 4203 4335 4261 4369
rect 4295 4335 4353 4369
rect 4387 4335 4445 4369
rect 4479 4335 4537 4369
rect 4571 4335 4629 4369
rect 4663 4335 4721 4369
rect 4755 4335 4813 4369
rect 4847 4335 4905 4369
rect 4939 4335 4997 4369
rect 5031 4335 5089 4369
rect 5123 4335 5181 4369
rect 5215 4335 5273 4369
rect 5307 4335 5365 4369
rect 5399 4335 5457 4369
rect 5491 4335 5549 4369
rect 5583 4335 5641 4369
rect 5675 4335 5733 4369
rect 5767 4335 5825 4369
rect 5859 4335 5917 4369
rect 5951 4335 6009 4369
rect 6043 4335 6101 4369
rect 6135 4335 6193 4369
rect 6227 4335 6285 4369
rect 6319 4335 6377 4369
rect 6411 4335 6469 4369
rect 6503 4335 6561 4369
rect 6595 4335 6653 4369
rect 6687 4335 6745 4369
rect 6779 4335 6837 4369
rect 6871 4335 6929 4369
rect 6963 4335 7021 4369
rect 7055 4335 7113 4369
rect 7147 4335 7205 4369
rect 7239 4335 7297 4369
rect 7331 4335 7389 4369
rect 7423 4335 7481 4369
rect 7515 4335 7573 4369
rect 7607 4335 7665 4369
rect 7699 4335 7757 4369
rect 7791 4335 7849 4369
rect 7883 4335 7941 4369
rect 7975 4335 8033 4369
rect 8067 4335 8125 4369
rect 8159 4335 8217 4369
rect 8251 4335 8309 4369
rect 8343 4335 8401 4369
rect 8435 4335 8493 4369
rect 8527 4335 8585 4369
rect 8619 4335 8677 4369
rect 8711 4335 8769 4369
rect 8803 4335 8861 4369
rect 8895 4335 8953 4369
rect 8987 4335 9045 4369
rect 9079 4335 9137 4369
rect 9171 4335 9229 4369
rect 9263 4335 9321 4369
rect 9355 4335 9413 4369
rect 9447 4335 9505 4369
rect 9539 4335 9597 4369
rect 9631 4335 9689 4369
rect 9723 4335 9781 4369
rect 9815 4335 9873 4369
rect 9907 4335 9965 4369
rect 9999 4335 10057 4369
rect 10091 4335 10149 4369
rect 10183 4335 10241 4369
rect 10275 4335 10333 4369
rect 10367 4335 10425 4369
rect 10459 4335 10517 4369
rect 10551 4335 10609 4369
rect 10643 4335 10701 4369
rect 10735 4335 10793 4369
rect 10827 4335 10885 4369
rect 10919 4335 10977 4369
rect 11011 4335 11069 4369
rect 11103 4335 11161 4369
rect 11195 4335 11253 4369
rect 11287 4335 11345 4369
rect 11379 4335 11437 4369
rect 11471 4335 11529 4369
rect 11563 4335 11621 4369
rect 11655 4335 11713 4369
rect 11747 4335 11805 4369
rect 11839 4335 11897 4369
rect 11931 4335 11989 4369
rect 12023 4335 12081 4369
rect 12115 4335 12173 4369
rect 12207 4335 12265 4369
rect 12299 4335 12357 4369
rect 12391 4335 12449 4369
rect 12483 4335 12541 4369
rect 12575 4335 12633 4369
rect 12667 4335 12725 4369
rect 12759 4335 12817 4369
rect 12851 4335 12909 4369
rect 12943 4335 13001 4369
rect 13035 4335 13093 4369
rect 13127 4335 13185 4369
rect 13219 4335 13277 4369
rect 13311 4335 13369 4369
rect 13403 4335 13461 4369
rect 13495 4335 13553 4369
rect 13587 4335 13645 4369
rect 13679 4335 13737 4369
rect 13771 4335 13829 4369
rect 13863 4335 13921 4369
rect 13955 4335 14013 4369
rect 14047 4335 14105 4369
rect 14139 4335 14197 4369
rect 14231 4335 14289 4369
rect 14323 4335 14381 4369
rect 14415 4335 14473 4369
rect 14507 4335 14565 4369
rect 14599 4335 14657 4369
rect 14691 4335 14749 4369
rect 14783 4335 14841 4369
rect 14875 4335 14933 4369
rect 14967 4335 15025 4369
rect 15059 4335 15117 4369
rect 15151 4335 15209 4369
rect 15243 4335 15301 4369
rect 15335 4335 15393 4369
rect 15427 4335 15485 4369
rect 15519 4335 15577 4369
rect 15611 4335 15669 4369
rect 15703 4335 15761 4369
rect 15795 4335 15853 4369
rect 15887 4335 15945 4369
rect 15979 4335 16037 4369
rect 16071 4335 16129 4369
rect 16163 4335 16221 4369
rect 16255 4335 16313 4369
rect 16347 4335 16405 4369
rect 16439 4335 16497 4369
rect 16531 4335 16589 4369
rect 16623 4335 16681 4369
rect 16715 4335 16773 4369
rect 16807 4335 16865 4369
rect 16899 4335 16957 4369
rect 16991 4335 17049 4369
rect 17083 4335 17141 4369
rect 17175 4335 17233 4369
rect 17267 4335 17325 4369
rect 17359 4335 17417 4369
rect 17451 4335 17509 4369
rect 17543 4335 17601 4369
rect 17635 4335 17693 4369
rect 17727 4335 17785 4369
rect 17819 4335 17877 4369
rect 17911 4335 17969 4369
rect 18003 4335 18061 4369
rect 18095 4335 18153 4369
rect 18187 4335 18245 4369
rect 18279 4335 18337 4369
rect 18371 4335 18429 4369
rect 18463 4335 18521 4369
rect 18555 4335 18613 4369
rect 18647 4335 18705 4369
rect 18739 4335 18797 4369
rect 18831 4335 18860 4369
rect 1121 4272 1363 4335
rect 1121 4238 1139 4272
rect 1173 4238 1311 4272
rect 1345 4238 1363 4272
rect 1121 4185 1363 4238
rect 1397 4274 1915 4335
rect 1397 4240 1415 4274
rect 1449 4240 1863 4274
rect 1897 4240 1915 4274
rect 1121 4111 1225 4185
rect 1397 4181 1915 4240
rect 1967 4280 2001 4301
rect 2037 4293 2103 4335
rect 2037 4259 2053 4293
rect 2087 4259 2103 4293
rect 2139 4263 2191 4301
rect 1967 4225 2001 4246
rect 2173 4229 2191 4263
rect 1967 4191 2100 4225
rect 2139 4200 2191 4229
rect 1121 4077 1171 4111
rect 1205 4077 1225 4111
rect 1259 4117 1279 4151
rect 1313 4117 1363 4151
rect 1259 4043 1363 4117
rect 1397 4111 1639 4181
rect 1397 4077 1475 4111
rect 1509 4077 1585 4111
rect 1619 4077 1639 4111
rect 1673 4113 1693 4147
rect 1727 4113 1803 4147
rect 1837 4113 1915 4147
rect 1673 4043 1915 4113
rect 1953 4137 2019 4155
rect 1953 4131 1969 4137
rect 1953 4097 1961 4131
rect 2003 4103 2019 4137
rect 1995 4097 2019 4103
rect 1953 4081 2019 4097
rect 2066 4140 2100 4191
rect 2066 4124 2123 4140
rect 2066 4090 2089 4124
rect 2066 4074 2123 4090
rect 2066 4045 2100 4074
rect 1121 3996 1363 4043
rect 1121 3962 1139 3996
rect 1173 3962 1311 3996
rect 1345 3962 1363 3996
rect 1121 3901 1363 3962
rect 1121 3867 1139 3901
rect 1173 3867 1311 3901
rect 1345 3867 1363 3901
rect 1121 3825 1363 3867
rect 1397 4003 1915 4043
rect 1397 3969 1415 4003
rect 1449 3969 1863 4003
rect 1897 3969 1915 4003
rect 1397 3901 1915 3969
rect 1397 3867 1415 3901
rect 1449 3867 1863 3901
rect 1897 3867 1915 3901
rect 1397 3825 1915 3867
rect 1967 4011 2100 4045
rect 2157 4040 2191 4200
rect 2225 4267 2559 4335
rect 2225 4233 2243 4267
rect 2277 4233 2507 4267
rect 2541 4233 2559 4267
rect 2225 4181 2559 4233
rect 2603 4290 2669 4291
rect 2603 4267 2619 4290
rect 2603 4233 2605 4267
rect 2653 4256 2669 4290
rect 2639 4233 2669 4256
rect 2603 4222 2669 4233
rect 2603 4204 2619 4222
rect 2593 4188 2619 4204
rect 2653 4188 2669 4222
rect 2703 4263 2737 4335
rect 2703 4213 2737 4229
rect 2771 4258 2787 4292
rect 2821 4258 2837 4292
rect 2771 4224 2837 4258
rect 2889 4279 2931 4335
rect 3294 4285 3368 4335
rect 2889 4245 2892 4279
rect 2926 4245 2931 4279
rect 2889 4229 2931 4245
rect 2986 4245 3090 4279
rect 3124 4245 3143 4279
rect 3177 4245 3193 4279
rect 3227 4245 3258 4279
rect 2593 4187 2669 4188
rect 2771 4190 2787 4224
rect 2821 4190 2837 4224
rect 2771 4187 2837 4190
rect 2225 4111 2375 4181
rect 2593 4179 2638 4187
rect 2225 4077 2245 4111
rect 2279 4077 2375 4111
rect 2409 4113 2505 4147
rect 2539 4113 2559 4147
rect 2409 4043 2559 4113
rect 1967 3977 2001 4011
rect 2137 3995 2191 4040
rect 2137 3990 2145 3995
rect 1967 3909 2001 3943
rect 1967 3859 2001 3875
rect 2037 3943 2053 3977
rect 2087 3943 2103 3977
rect 2037 3909 2103 3943
rect 2037 3875 2053 3909
rect 2087 3875 2103 3909
rect 2037 3825 2103 3875
rect 2137 3956 2139 3990
rect 2179 3961 2191 3995
rect 2173 3956 2191 3961
rect 2137 3909 2191 3956
rect 2137 3875 2139 3909
rect 2173 3875 2191 3909
rect 2137 3859 2191 3875
rect 2225 4003 2559 4043
rect 2593 4063 2627 4179
rect 2771 4153 2811 4187
rect 2986 4153 3020 4245
rect 2661 4137 2811 4153
rect 2695 4103 2811 4137
rect 2661 4087 2811 4103
rect 2845 4137 3020 4153
rect 2879 4103 3020 4137
rect 2845 4087 3020 4103
rect 2593 4053 2636 4063
rect 2593 4043 2671 4053
rect 2593 4037 2621 4043
rect 2225 3969 2243 4003
rect 2277 3969 2507 4003
rect 2541 3969 2559 4003
rect 2225 3901 2559 3969
rect 2225 3867 2243 3901
rect 2277 3867 2507 3901
rect 2541 3867 2559 3901
rect 2605 4009 2621 4037
rect 2655 4009 2671 4043
rect 2773 4046 2811 4087
rect 2773 4043 2952 4046
rect 2605 3975 2671 4009
rect 2605 3941 2621 3975
rect 2655 3941 2671 3975
rect 2605 3907 2671 3941
rect 2605 3873 2621 3907
rect 2655 3873 2671 3907
rect 2605 3868 2671 3873
rect 2705 4011 2739 4027
rect 2705 3931 2739 3977
rect 2225 3825 2559 3867
rect 2705 3825 2739 3897
rect 2773 4009 2791 4043
rect 2825 4021 2952 4043
rect 2825 4009 2918 4021
rect 2773 3987 2918 4009
rect 2773 3972 2952 3987
rect 2773 3938 2791 3972
rect 2825 3971 2952 3972
rect 2825 3938 2841 3971
rect 2773 3901 2841 3938
rect 2773 3867 2791 3901
rect 2825 3867 2841 3901
rect 2773 3859 2841 3867
rect 2887 3909 2950 3925
rect 2887 3875 2914 3909
rect 2948 3875 2950 3909
rect 2986 3919 3020 4087
rect 3054 4195 3147 4211
rect 3054 4161 3113 4195
rect 3054 4145 3147 4161
rect 3224 4199 3258 4245
rect 3294 4251 3312 4285
rect 3346 4251 3368 4285
rect 3707 4293 3757 4335
rect 3294 4235 3368 4251
rect 3432 4245 3511 4279
rect 3545 4245 3567 4279
rect 3606 4245 3622 4279
rect 3656 4245 3673 4279
rect 3224 4183 3390 4199
rect 3224 4149 3356 4183
rect 3054 4063 3118 4145
rect 3224 4139 3390 4149
rect 3054 4029 3067 4063
rect 3101 4029 3118 4063
rect 3054 4021 3118 4029
rect 3088 3987 3118 4021
rect 3054 3953 3118 3987
rect 3152 4087 3190 4103
rect 3152 4053 3156 4087
rect 3152 3995 3190 4053
rect 3152 3961 3154 3995
rect 3188 3961 3190 3995
rect 3152 3959 3190 3961
rect 3224 3925 3258 4139
rect 3350 4133 3390 4139
rect 3292 4089 3326 4103
rect 3432 4089 3466 4245
rect 3639 4217 3673 4245
rect 3741 4259 3757 4293
rect 3879 4293 3945 4335
rect 3707 4243 3757 4259
rect 3808 4267 3845 4283
rect 3808 4233 3811 4267
rect 3879 4259 3895 4293
rect 3929 4259 3945 4293
rect 3979 4267 4013 4283
rect 3292 4087 3466 4089
rect 3326 4055 3466 4087
rect 3500 4195 3605 4205
rect 3500 4161 3555 4195
rect 3589 4161 3605 4195
rect 3639 4191 3684 4217
rect 3326 4053 3394 4055
rect 3292 4037 3394 4053
rect 2986 3885 3113 3919
rect 3147 3885 3163 3919
rect 3208 3909 3258 3925
rect 2887 3825 2950 3875
rect 3242 3875 3258 3909
rect 3208 3859 3258 3875
rect 3292 3969 3326 3985
rect 3292 3901 3326 3935
rect 3360 3914 3394 4037
rect 3428 3987 3466 4021
rect 3500 3995 3534 4161
rect 3568 4099 3616 4127
rect 3568 4065 3575 4099
rect 3609 4065 3616 4099
rect 3568 4063 3616 4065
rect 3568 4029 3571 4063
rect 3605 4029 3616 4063
rect 3568 4008 3616 4029
rect 3428 3961 3468 3987
rect 3502 3961 3534 3995
rect 3650 3970 3684 4191
rect 3718 4131 3774 4209
rect 3718 4097 3729 4131
rect 3763 4097 3774 4131
rect 3718 4069 3774 4097
rect 3752 4035 3774 4069
rect 3718 4019 3774 4035
rect 3808 4063 3845 4233
rect 3979 4225 4013 4233
rect 3808 4029 3809 4063
rect 3843 4029 3845 4063
rect 3428 3948 3534 3961
rect 3623 3944 3684 3970
rect 3808 3977 3845 4029
rect 3360 3880 3531 3914
rect 3565 3880 3581 3914
rect 3623 3909 3673 3944
rect 3808 3943 3811 3977
rect 3880 4191 4013 4225
rect 4065 4274 4583 4335
rect 4065 4240 4083 4274
rect 4117 4240 4531 4274
rect 4565 4240 4583 4274
rect 3880 4122 3926 4191
rect 4065 4181 4583 4240
rect 4627 4290 4693 4291
rect 4627 4267 4643 4290
rect 4627 4233 4629 4267
rect 4677 4256 4693 4290
rect 4663 4233 4693 4256
rect 4627 4222 4693 4233
rect 4627 4204 4643 4222
rect 4617 4188 4643 4204
rect 4677 4188 4693 4222
rect 4727 4263 4761 4335
rect 4727 4213 4761 4229
rect 4795 4258 4811 4292
rect 4845 4258 4861 4292
rect 4795 4224 4861 4258
rect 4913 4279 4955 4335
rect 5318 4285 5392 4335
rect 4913 4245 4916 4279
rect 4950 4245 4955 4279
rect 4913 4229 4955 4245
rect 5010 4245 5114 4279
rect 5148 4245 5167 4279
rect 5201 4245 5217 4279
rect 5251 4245 5282 4279
rect 4617 4187 4693 4188
rect 4795 4190 4811 4224
rect 4845 4190 4861 4224
rect 4795 4187 4861 4190
rect 3914 4088 3926 4122
rect 3880 3995 3926 4088
rect 3960 4137 4030 4157
rect 3960 4103 3982 4137
rect 4016 4131 4030 4137
rect 3960 4097 3985 4103
rect 4019 4097 4030 4131
rect 3960 4027 4030 4097
rect 4065 4111 4307 4181
rect 4617 4179 4662 4187
rect 4065 4077 4143 4111
rect 4177 4077 4253 4111
rect 4287 4077 4307 4111
rect 4341 4113 4361 4147
rect 4395 4113 4471 4147
rect 4505 4113 4583 4147
rect 4341 4043 4583 4113
rect 3880 3961 3888 3995
rect 3922 3993 3926 3995
rect 4065 4003 4583 4043
rect 4617 4063 4651 4179
rect 4795 4153 4835 4187
rect 5010 4153 5044 4245
rect 4685 4137 4835 4153
rect 4719 4103 4835 4137
rect 4685 4087 4835 4103
rect 4869 4137 5044 4153
rect 4903 4103 5044 4137
rect 4869 4087 5044 4103
rect 4617 4053 4660 4063
rect 4617 4043 4695 4053
rect 4617 4037 4645 4043
rect 3922 3977 4013 3993
rect 3922 3961 3979 3977
rect 3880 3959 3979 3961
rect 3292 3825 3326 3867
rect 3657 3875 3673 3909
rect 3623 3859 3673 3875
rect 3707 3901 3760 3917
rect 3741 3867 3760 3901
rect 3707 3825 3760 3867
rect 3808 3909 3845 3943
rect 3808 3875 3811 3909
rect 3808 3859 3845 3875
rect 3879 3891 3895 3925
rect 3929 3891 3945 3925
rect 3879 3825 3945 3891
rect 3979 3909 4013 3943
rect 3979 3859 4013 3875
rect 4065 3969 4083 4003
rect 4117 3969 4531 4003
rect 4565 3969 4583 4003
rect 4065 3901 4583 3969
rect 4065 3867 4083 3901
rect 4117 3867 4531 3901
rect 4565 3867 4583 3901
rect 4629 4009 4645 4037
rect 4679 4009 4695 4043
rect 4797 4046 4835 4087
rect 4797 4043 4976 4046
rect 4629 3975 4695 4009
rect 4629 3941 4645 3975
rect 4679 3941 4695 3975
rect 4629 3907 4695 3941
rect 4629 3873 4645 3907
rect 4679 3873 4695 3907
rect 4629 3868 4695 3873
rect 4729 4011 4763 4027
rect 4729 3931 4763 3977
rect 4065 3825 4583 3867
rect 4729 3825 4763 3897
rect 4797 4009 4815 4043
rect 4849 4021 4976 4043
rect 4849 4009 4942 4021
rect 4797 3987 4942 4009
rect 4797 3972 4976 3987
rect 4797 3938 4815 3972
rect 4849 3971 4976 3972
rect 4849 3938 4865 3971
rect 4797 3901 4865 3938
rect 4797 3867 4815 3901
rect 4849 3867 4865 3901
rect 4797 3859 4865 3867
rect 4911 3909 4974 3925
rect 4911 3875 4938 3909
rect 4972 3875 4974 3909
rect 5010 3919 5044 4087
rect 5078 4195 5171 4211
rect 5078 4161 5137 4195
rect 5078 4145 5171 4161
rect 5248 4199 5282 4245
rect 5318 4251 5336 4285
rect 5370 4251 5392 4285
rect 5731 4293 5781 4335
rect 5318 4235 5392 4251
rect 5456 4245 5535 4279
rect 5569 4245 5591 4279
rect 5630 4245 5646 4279
rect 5680 4245 5697 4279
rect 5248 4183 5414 4199
rect 5248 4149 5380 4183
rect 5078 4063 5142 4145
rect 5248 4139 5414 4149
rect 5078 4029 5091 4063
rect 5125 4029 5142 4063
rect 5078 4021 5142 4029
rect 5112 3987 5142 4021
rect 5078 3953 5142 3987
rect 5176 4087 5214 4103
rect 5176 4053 5180 4087
rect 5176 3995 5214 4053
rect 5176 3961 5178 3995
rect 5212 3961 5214 3995
rect 5176 3959 5214 3961
rect 5248 3925 5282 4139
rect 5374 4133 5414 4139
rect 5316 4089 5350 4103
rect 5456 4089 5490 4245
rect 5663 4217 5697 4245
rect 5765 4259 5781 4293
rect 5903 4293 5969 4335
rect 5731 4243 5781 4259
rect 5832 4267 5869 4283
rect 5832 4233 5835 4267
rect 5903 4259 5919 4293
rect 5953 4259 5969 4293
rect 6003 4267 6037 4283
rect 5316 4087 5490 4089
rect 5350 4055 5490 4087
rect 5524 4195 5629 4205
rect 5524 4161 5579 4195
rect 5613 4161 5629 4195
rect 5663 4191 5708 4217
rect 5350 4053 5418 4055
rect 5316 4037 5418 4053
rect 5010 3885 5137 3919
rect 5171 3885 5187 3919
rect 5232 3909 5282 3925
rect 4911 3825 4974 3875
rect 5266 3875 5282 3909
rect 5232 3859 5282 3875
rect 5316 3969 5350 3985
rect 5316 3901 5350 3935
rect 5384 3914 5418 4037
rect 5452 3987 5490 4021
rect 5524 3995 5558 4161
rect 5592 4099 5640 4127
rect 5592 4065 5599 4099
rect 5633 4065 5640 4099
rect 5592 4063 5640 4065
rect 5592 4029 5595 4063
rect 5629 4029 5640 4063
rect 5592 4008 5640 4029
rect 5452 3961 5492 3987
rect 5526 3961 5558 3995
rect 5674 3970 5708 4191
rect 5742 4131 5798 4209
rect 5776 4097 5798 4131
rect 5742 4069 5798 4097
rect 5776 4035 5798 4069
rect 5742 4019 5798 4035
rect 5832 4063 5869 4233
rect 6003 4225 6037 4233
rect 5832 4029 5833 4063
rect 5867 4029 5869 4063
rect 5452 3948 5558 3961
rect 5647 3944 5708 3970
rect 5832 3977 5869 4029
rect 5384 3880 5555 3914
rect 5589 3880 5605 3914
rect 5647 3909 5697 3944
rect 5832 3943 5835 3977
rect 5904 4191 6037 4225
rect 6273 4241 6331 4335
rect 6273 4207 6285 4241
rect 6319 4207 6331 4241
rect 5904 4122 5950 4191
rect 6273 4190 6331 4207
rect 6365 4274 6883 4335
rect 6365 4240 6383 4274
rect 6417 4240 6831 4274
rect 6865 4240 6883 4274
rect 6365 4181 6883 4240
rect 6917 4290 6985 4301
rect 6917 4256 6935 4290
rect 6969 4256 6985 4290
rect 6917 4222 6985 4256
rect 7019 4293 7053 4335
rect 7019 4243 7053 4259
rect 7101 4289 7173 4301
rect 7101 4255 7123 4289
rect 7157 4255 7173 4289
rect 7101 4248 7173 4255
rect 7299 4293 7333 4335
rect 7101 4247 7172 4248
rect 7101 4245 7171 4247
rect 7101 4244 7170 4245
rect 6917 4188 6935 4222
rect 6969 4188 6985 4222
rect 7101 4242 7169 4244
rect 7299 4243 7333 4259
rect 7367 4289 7435 4301
rect 7367 4255 7383 4289
rect 7417 4255 7435 4289
rect 7101 4241 7168 4242
rect 7101 4239 7166 4241
rect 7101 4237 7164 4239
rect 7101 4221 7161 4237
rect 7101 4209 7123 4221
rect 5938 4088 5950 4122
rect 5904 3995 5950 4088
rect 5984 4137 6054 4157
rect 5984 4103 6006 4137
rect 6040 4131 6054 4137
rect 5984 4097 6009 4103
rect 6043 4097 6054 4131
rect 5984 4027 6054 4097
rect 6365 4111 6607 4181
rect 6365 4077 6443 4111
rect 6477 4077 6553 4111
rect 6587 4077 6607 4111
rect 6641 4113 6661 4147
rect 6695 4113 6771 4147
rect 6805 4113 6883 4147
rect 5904 3961 5912 3995
rect 5946 3993 5950 3995
rect 6273 4023 6331 4058
rect 6641 4043 6883 4113
rect 5946 3977 6037 3993
rect 5946 3961 6003 3977
rect 5904 3959 6003 3961
rect 5316 3825 5350 3867
rect 5681 3875 5697 3909
rect 5647 3859 5697 3875
rect 5731 3901 5784 3917
rect 5765 3867 5784 3901
rect 5731 3825 5784 3867
rect 5832 3909 5869 3943
rect 5832 3875 5835 3909
rect 5832 3859 5869 3875
rect 5903 3891 5919 3925
rect 5953 3891 5969 3925
rect 5903 3825 5969 3891
rect 6003 3909 6037 3943
rect 6003 3859 6037 3875
rect 6273 3989 6285 4023
rect 6319 3989 6331 4023
rect 6273 3930 6331 3989
rect 6273 3896 6285 3930
rect 6319 3896 6331 3930
rect 6273 3825 6331 3896
rect 6365 4003 6883 4043
rect 6365 3969 6383 4003
rect 6417 3969 6831 4003
rect 6865 3969 6883 4003
rect 6365 3901 6883 3969
rect 6365 3867 6383 3901
rect 6417 3867 6831 3901
rect 6865 3867 6883 3901
rect 6365 3825 6883 3867
rect 6917 4146 6985 4188
rect 7019 4187 7123 4209
rect 7157 4187 7161 4221
rect 7019 4171 7161 4187
rect 7199 4191 7215 4225
rect 7249 4209 7265 4225
rect 7367 4221 7435 4255
rect 7367 4209 7383 4221
rect 7249 4191 7383 4209
rect 7199 4187 7383 4191
rect 7417 4187 7435 4221
rect 7199 4171 7435 4187
rect 7469 4267 7803 4335
rect 7469 4233 7487 4267
rect 7521 4233 7751 4267
rect 7785 4233 7803 4267
rect 7837 4293 7898 4335
rect 7837 4259 7855 4293
rect 7889 4259 7898 4293
rect 7837 4233 7898 4259
rect 7934 4280 7984 4299
rect 7934 4246 7941 4280
rect 7975 4246 7984 4280
rect 7469 4181 7803 4233
rect 6917 4045 6973 4146
rect 6917 4011 6939 4045
rect 7019 4137 7076 4171
rect 7053 4103 7076 4137
rect 7019 4057 7076 4103
rect 7113 4131 7157 4137
rect 7147 4103 7157 4131
rect 7191 4103 7207 4137
rect 7147 4097 7207 4103
rect 7241 4103 7257 4137
rect 7291 4133 7307 4137
rect 7291 4131 7331 4133
rect 7291 4103 7297 4131
rect 7241 4097 7297 4103
rect 7369 4103 7385 4137
rect 7419 4103 7435 4137
rect 7369 4097 7435 4103
rect 7113 4091 7207 4097
rect 7019 4037 7249 4057
rect 7019 4014 7199 4037
rect 6917 3977 6973 4011
rect 7183 4003 7199 4014
rect 7233 4003 7249 4037
rect 6917 3943 6939 3977
rect 6917 3927 6973 3943
rect 6917 3893 6929 3927
rect 6963 3909 6973 3927
rect 6917 3875 6939 3893
rect 6917 3859 6973 3875
rect 7007 3969 7149 3980
rect 7007 3935 7025 3969
rect 7059 3935 7099 3969
rect 7133 3935 7149 3969
rect 7007 3901 7149 3935
rect 7007 3867 7025 3901
rect 7059 3867 7099 3901
rect 7133 3867 7149 3901
rect 7007 3825 7149 3867
rect 7183 3969 7249 4003
rect 7183 3935 7199 3969
rect 7233 3935 7249 3969
rect 7183 3901 7249 3935
rect 7183 3867 7199 3901
rect 7233 3867 7249 3901
rect 7288 3874 7331 4097
rect 7389 4063 7435 4097
rect 7469 4111 7619 4181
rect 7837 4165 7849 4199
rect 7883 4165 7900 4199
rect 7469 4077 7489 4111
rect 7523 4077 7619 4111
rect 7653 4113 7749 4147
rect 7783 4113 7803 4147
rect 7423 4029 7435 4063
rect 7653 4043 7803 4113
rect 7837 4137 7900 4165
rect 7837 4103 7857 4137
rect 7891 4103 7900 4137
rect 7837 4087 7900 4103
rect 7934 4137 7984 4246
rect 8018 4280 8070 4335
rect 8018 4246 8027 4280
rect 8061 4246 8070 4280
rect 8018 4230 8070 4246
rect 8106 4280 8156 4299
rect 8106 4246 8113 4280
rect 8147 4246 8156 4280
rect 8106 4137 8156 4246
rect 8190 4280 8242 4335
rect 8190 4246 8199 4280
rect 8233 4246 8242 4280
rect 8190 4223 8242 4246
rect 8276 4280 8328 4296
rect 8276 4246 8285 4280
rect 8319 4246 8328 4280
rect 8276 4205 8328 4246
rect 8362 4289 8414 4335
rect 8362 4255 8371 4289
rect 8405 4255 8414 4289
rect 8362 4239 8414 4255
rect 8448 4280 8500 4296
rect 8448 4246 8457 4280
rect 8491 4246 8500 4280
rect 8448 4205 8500 4246
rect 8534 4289 8586 4335
rect 8534 4255 8543 4289
rect 8577 4255 8586 4289
rect 8534 4239 8586 4255
rect 8620 4280 8672 4296
rect 8620 4246 8629 4280
rect 8663 4246 8672 4280
rect 8620 4205 8672 4246
rect 8706 4289 8755 4335
rect 8706 4255 8715 4289
rect 8749 4255 8755 4289
rect 8706 4239 8755 4255
rect 8789 4280 8844 4296
rect 8789 4246 8801 4280
rect 8835 4246 8844 4280
rect 8789 4205 8844 4246
rect 8878 4289 8927 4335
rect 8878 4255 8887 4289
rect 8921 4255 8927 4289
rect 8878 4239 8927 4255
rect 8961 4280 9013 4296
rect 8961 4246 8972 4280
rect 9006 4246 9013 4280
rect 8961 4205 9013 4246
rect 9049 4289 9099 4335
rect 9049 4255 9058 4289
rect 9092 4255 9099 4289
rect 9049 4239 9099 4255
rect 9133 4280 9185 4296
rect 9133 4246 9144 4280
rect 9178 4246 9185 4280
rect 9133 4205 9185 4246
rect 9221 4289 9271 4335
rect 9221 4255 9230 4289
rect 9264 4255 9271 4289
rect 9221 4239 9271 4255
rect 9305 4280 9357 4296
rect 9305 4246 9316 4280
rect 9350 4246 9357 4280
rect 9305 4205 9357 4246
rect 9393 4289 9445 4335
rect 9393 4255 9402 4289
rect 9436 4255 9445 4289
rect 9393 4239 9445 4255
rect 9479 4280 9531 4296
rect 9479 4246 9488 4280
rect 9522 4246 9531 4280
rect 9479 4205 9531 4246
rect 9565 4289 9625 4335
rect 9565 4255 9574 4289
rect 9608 4255 9625 4289
rect 9565 4239 9625 4255
rect 9677 4274 10379 4335
rect 9677 4240 9695 4274
rect 9729 4240 10327 4274
rect 10361 4240 10379 4274
rect 8276 4171 9625 4205
rect 7934 4103 8284 4137
rect 8318 4103 8352 4137
rect 8386 4103 8420 4137
rect 8454 4103 8488 4137
rect 8522 4103 8556 4137
rect 8590 4103 8624 4137
rect 8658 4103 8692 4137
rect 8726 4103 8760 4137
rect 8794 4103 8828 4137
rect 8862 4103 8896 4137
rect 8930 4103 8964 4137
rect 8998 4103 9032 4137
rect 9066 4103 9100 4137
rect 9134 4103 9168 4137
rect 9202 4103 9236 4137
rect 9270 4103 9304 4137
rect 9338 4103 9358 4137
rect 7934 4087 9358 4103
rect 7469 4003 7803 4043
rect 7469 3969 7487 4003
rect 7521 3969 7751 4003
rect 7785 3969 7803 4003
rect 7367 3935 7383 3969
rect 7417 3935 7433 3969
rect 7367 3901 7433 3935
rect 7183 3859 7249 3867
rect 7367 3867 7383 3901
rect 7417 3867 7433 3901
rect 7367 3825 7433 3867
rect 7469 3901 7803 3969
rect 7469 3867 7487 3901
rect 7521 3867 7751 3901
rect 7785 3867 7803 3901
rect 7469 3825 7803 3867
rect 7839 3969 7898 3987
rect 7839 3935 7855 3969
rect 7889 3935 7898 3969
rect 7839 3901 7898 3935
rect 7839 3867 7855 3901
rect 7889 3867 7898 3901
rect 7839 3825 7898 3867
rect 7934 3977 7983 4087
rect 7934 3943 7941 3977
rect 7975 3943 7983 3977
rect 7934 3909 7983 3943
rect 7934 3875 7941 3909
rect 7975 3875 7983 3909
rect 7934 3859 7983 3875
rect 8018 3969 8070 3987
rect 8018 3935 8027 3969
rect 8061 3935 8070 3969
rect 8018 3901 8070 3935
rect 8018 3867 8027 3901
rect 8061 3867 8070 3901
rect 8018 3825 8070 3867
rect 8106 3985 8156 4087
rect 9392 4063 9625 4171
rect 9677 4181 10379 4240
rect 10505 4290 10573 4301
rect 10505 4256 10523 4290
rect 10557 4256 10573 4290
rect 10505 4222 10573 4256
rect 10607 4293 10641 4335
rect 10607 4243 10641 4259
rect 10689 4289 10761 4301
rect 10689 4255 10711 4289
rect 10745 4255 10761 4289
rect 10689 4248 10761 4255
rect 10887 4293 10921 4335
rect 10689 4247 10760 4248
rect 10689 4245 10759 4247
rect 10689 4244 10758 4245
rect 10505 4188 10523 4222
rect 10557 4188 10573 4222
rect 10689 4242 10757 4244
rect 10887 4243 10921 4259
rect 10955 4289 11023 4301
rect 10955 4255 10971 4289
rect 11005 4255 11023 4289
rect 10689 4241 10756 4242
rect 10689 4239 10754 4241
rect 10689 4237 10752 4239
rect 10689 4221 10749 4237
rect 10689 4209 10711 4221
rect 9677 4111 10007 4181
rect 9677 4077 9755 4111
rect 9789 4077 9854 4111
rect 9888 4077 9953 4111
rect 9987 4077 10007 4111
rect 10041 4113 10061 4147
rect 10095 4113 10164 4147
rect 10198 4113 10267 4147
rect 10301 4113 10379 4147
rect 9392 4053 9597 4063
rect 8276 4031 9597 4053
rect 8276 3997 8285 4031
rect 8319 4005 8457 4031
rect 8319 3997 8328 4005
rect 8106 3951 8113 3985
rect 8147 3951 8156 3985
rect 8106 3917 8156 3951
rect 8106 3883 8113 3917
rect 8147 3883 8156 3917
rect 8106 3860 8156 3883
rect 8190 3969 8242 3985
rect 8190 3935 8199 3969
rect 8233 3935 8242 3969
rect 8190 3901 8242 3935
rect 8190 3867 8199 3901
rect 8233 3867 8242 3901
rect 8190 3826 8242 3867
rect 8276 3945 8328 3997
rect 8448 3997 8457 4005
rect 8491 4005 8629 4031
rect 8491 3997 8500 4005
rect 8276 3911 8285 3945
rect 8319 3911 8328 3945
rect 8276 3860 8328 3911
rect 8362 3925 8414 3971
rect 8362 3891 8371 3925
rect 8405 3891 8414 3925
rect 8362 3826 8414 3891
rect 8448 3945 8500 3997
rect 8620 3997 8629 4005
rect 8663 4005 8801 4031
rect 8663 3997 8672 4005
rect 8448 3911 8457 3945
rect 8491 3911 8500 3945
rect 8448 3860 8500 3911
rect 8534 3925 8586 3971
rect 8534 3891 8543 3925
rect 8577 3891 8586 3925
rect 8534 3826 8586 3891
rect 8620 3945 8672 3997
rect 8792 3997 8801 4005
rect 8835 4005 8972 4031
rect 8835 3997 8844 4005
rect 8620 3911 8629 3945
rect 8663 3911 8672 3945
rect 8620 3860 8672 3911
rect 8706 3925 8758 3971
rect 8706 3891 8715 3925
rect 8749 3891 8758 3925
rect 8706 3826 8758 3891
rect 8792 3945 8844 3997
rect 8961 3997 8972 4005
rect 9006 4005 9144 4031
rect 9006 3997 9013 4005
rect 8792 3911 8801 3945
rect 8835 3911 8844 3945
rect 8792 3860 8844 3911
rect 8878 3925 8927 3971
rect 8878 3891 8887 3925
rect 8921 3891 8927 3925
rect 8878 3826 8927 3891
rect 8961 3945 9013 3997
rect 9133 3997 9144 4005
rect 9178 4005 9316 4031
rect 9178 3997 9185 4005
rect 8961 3911 8972 3945
rect 9006 3911 9013 3945
rect 8961 3860 9013 3911
rect 9050 3925 9099 3971
rect 9050 3891 9058 3925
rect 9092 3891 9099 3925
rect 9050 3826 9099 3891
rect 9133 3945 9185 3997
rect 9305 3997 9316 4005
rect 9350 4008 9488 4031
rect 9350 3997 9357 4008
rect 9133 3911 9144 3945
rect 9178 3911 9185 3945
rect 9133 3860 9185 3911
rect 9222 3925 9271 3971
rect 9222 3891 9230 3925
rect 9264 3891 9271 3925
rect 9222 3826 9271 3891
rect 9305 3945 9357 3997
rect 9479 3997 9488 4008
rect 9522 4029 9597 4031
rect 10041 4043 10379 4113
rect 9522 4008 9625 4029
rect 9522 3997 9537 4008
rect 9305 3911 9316 3945
rect 9350 3911 9357 3945
rect 9305 3860 9357 3911
rect 9394 3925 9445 3971
rect 9394 3891 9402 3925
rect 9436 3891 9445 3925
rect 9394 3826 9445 3891
rect 9479 3945 9537 3997
rect 9677 4003 10379 4043
rect 9479 3911 9488 3945
rect 9522 3911 9537 3945
rect 9479 3860 9537 3911
rect 9571 3925 9625 3974
rect 9571 3891 9574 3925
rect 9608 3891 9625 3925
rect 8190 3825 9445 3826
rect 9571 3825 9625 3891
rect 9677 3969 9695 4003
rect 9729 3969 10327 4003
rect 10361 3969 10379 4003
rect 9677 3901 10379 3969
rect 9677 3867 9695 3901
rect 9729 3867 10327 3901
rect 10361 3867 10379 3901
rect 9677 3825 10379 3867
rect 10505 4146 10573 4188
rect 10607 4187 10711 4209
rect 10745 4187 10749 4221
rect 10607 4171 10749 4187
rect 10787 4191 10803 4225
rect 10837 4209 10853 4225
rect 10955 4221 11023 4255
rect 10955 4209 10971 4221
rect 10837 4191 10971 4209
rect 10787 4187 10971 4191
rect 11005 4187 11023 4221
rect 10787 4171 11023 4187
rect 11057 4267 11391 4335
rect 11057 4233 11075 4267
rect 11109 4233 11339 4267
rect 11373 4233 11391 4267
rect 11057 4181 11391 4233
rect 11425 4241 11483 4335
rect 11787 4293 11853 4335
rect 11425 4207 11437 4241
rect 11471 4207 11483 4241
rect 11425 4190 11483 4207
rect 11719 4267 11753 4283
rect 11787 4259 11803 4293
rect 11837 4259 11853 4293
rect 11975 4293 12025 4335
rect 11887 4267 11924 4283
rect 11719 4225 11753 4233
rect 11921 4233 11924 4267
rect 11975 4259 11991 4293
rect 12364 4285 12438 4335
rect 11975 4243 12025 4259
rect 12059 4245 12076 4279
rect 12110 4245 12126 4279
rect 12165 4245 12187 4279
rect 12221 4245 12300 4279
rect 11719 4191 11852 4225
rect 10505 4045 10561 4146
rect 10505 4011 10527 4045
rect 10607 4137 10664 4171
rect 10641 4103 10664 4137
rect 10607 4057 10664 4103
rect 10701 4131 10745 4137
rect 10735 4103 10745 4131
rect 10779 4103 10795 4137
rect 10735 4097 10795 4103
rect 10829 4103 10845 4137
rect 10879 4133 10895 4137
rect 10879 4103 10919 4133
rect 10829 4097 10919 4103
rect 10957 4103 10973 4137
rect 11007 4103 11023 4137
rect 10957 4097 11023 4103
rect 10701 4091 10795 4097
rect 10607 4037 10837 4057
rect 10607 4014 10787 4037
rect 10505 3977 10561 4011
rect 10771 4003 10787 4014
rect 10821 4003 10837 4037
rect 10505 3943 10527 3977
rect 10505 3927 10561 3943
rect 10505 3893 10517 3927
rect 10551 3909 10561 3927
rect 10505 3875 10527 3893
rect 10505 3859 10561 3875
rect 10595 3969 10737 3980
rect 10595 3935 10613 3969
rect 10647 3935 10687 3969
rect 10721 3935 10737 3969
rect 10595 3901 10737 3935
rect 10595 3867 10613 3901
rect 10647 3867 10687 3901
rect 10721 3867 10737 3901
rect 10595 3825 10737 3867
rect 10771 3969 10837 4003
rect 10771 3935 10787 3969
rect 10821 3935 10837 3969
rect 10771 3901 10837 3935
rect 10771 3867 10787 3901
rect 10821 3867 10837 3901
rect 10876 3995 10919 4097
rect 10977 4063 11023 4097
rect 11057 4111 11207 4181
rect 11057 4077 11077 4111
rect 11111 4077 11207 4111
rect 11241 4113 11337 4147
rect 11371 4113 11391 4147
rect 11011 4029 11023 4063
rect 11241 4043 11391 4113
rect 11702 4137 11772 4157
rect 11702 4131 11716 4137
rect 11702 4097 11713 4131
rect 11750 4103 11772 4137
rect 11747 4097 11772 4103
rect 10876 3961 10885 3995
rect 11057 4003 11391 4043
rect 11057 3969 11075 4003
rect 11109 3969 11339 4003
rect 11373 3969 11391 4003
rect 10876 3874 10919 3961
rect 10955 3935 10971 3969
rect 11005 3935 11021 3969
rect 10955 3901 11021 3935
rect 10771 3859 10837 3867
rect 10955 3867 10971 3901
rect 11005 3867 11021 3901
rect 10955 3825 11021 3867
rect 11057 3901 11391 3969
rect 11057 3867 11075 3901
rect 11109 3867 11339 3901
rect 11373 3867 11391 3901
rect 11057 3825 11391 3867
rect 11425 4023 11483 4058
rect 11702 4027 11772 4097
rect 11806 4122 11852 4191
rect 11806 4088 11818 4122
rect 11425 3989 11437 4023
rect 11471 3989 11483 4023
rect 11806 3995 11852 4088
rect 11806 3993 11810 3995
rect 11425 3930 11483 3989
rect 11425 3896 11437 3930
rect 11471 3896 11483 3930
rect 11425 3825 11483 3896
rect 11719 3977 11810 3993
rect 11753 3961 11810 3977
rect 11844 3961 11852 3995
rect 11753 3959 11852 3961
rect 11887 4063 11924 4233
rect 12059 4217 12093 4245
rect 11887 4029 11889 4063
rect 11923 4029 11924 4063
rect 11887 3977 11924 4029
rect 11958 4199 12014 4209
rect 11958 4165 11980 4199
rect 11958 4069 12014 4165
rect 11958 4035 11980 4069
rect 11958 4019 12014 4035
rect 12048 4191 12093 4217
rect 12127 4195 12232 4205
rect 11719 3909 11753 3943
rect 11921 3943 11924 3977
rect 12048 3970 12082 4191
rect 12127 4161 12143 4195
rect 12177 4161 12232 4195
rect 12116 4099 12164 4127
rect 12116 4065 12123 4099
rect 12157 4065 12164 4099
rect 12116 4063 12164 4065
rect 12116 4029 12127 4063
rect 12161 4029 12164 4063
rect 12116 4008 12164 4029
rect 12198 3995 12232 4161
rect 12266 4089 12300 4245
rect 12364 4251 12386 4285
rect 12420 4251 12438 4285
rect 12801 4279 12843 4335
rect 12364 4235 12438 4251
rect 12474 4245 12505 4279
rect 12539 4245 12555 4279
rect 12589 4245 12608 4279
rect 12642 4245 12746 4279
rect 12474 4199 12508 4245
rect 12342 4183 12508 4199
rect 12376 4149 12508 4183
rect 12342 4139 12508 4149
rect 12585 4195 12678 4211
rect 12619 4161 12678 4195
rect 12585 4145 12678 4161
rect 12342 4133 12382 4139
rect 12406 4089 12440 4103
rect 12266 4087 12440 4089
rect 12266 4055 12406 4087
rect 12338 4053 12406 4055
rect 12338 4037 12440 4053
rect 12048 3944 12109 3970
rect 12198 3961 12230 3995
rect 12266 3987 12304 4021
rect 12264 3961 12304 3987
rect 12198 3948 12304 3961
rect 11719 3859 11753 3875
rect 11787 3891 11803 3925
rect 11837 3891 11853 3925
rect 11787 3825 11853 3891
rect 11887 3909 11924 3943
rect 11921 3875 11924 3909
rect 11887 3859 11924 3875
rect 11972 3901 12025 3917
rect 11972 3867 11991 3901
rect 11972 3825 12025 3867
rect 12059 3909 12109 3944
rect 12338 3914 12372 4037
rect 12059 3875 12075 3909
rect 12151 3880 12167 3914
rect 12201 3880 12372 3914
rect 12406 3969 12440 3985
rect 12406 3901 12440 3935
rect 12059 3859 12109 3875
rect 12406 3825 12440 3867
rect 12474 3925 12508 4139
rect 12542 4087 12580 4103
rect 12576 4053 12580 4087
rect 12542 3995 12580 4053
rect 12542 3961 12544 3995
rect 12578 3961 12580 3995
rect 12542 3959 12580 3961
rect 12614 4063 12678 4145
rect 12614 4029 12631 4063
rect 12665 4029 12678 4063
rect 12614 4021 12678 4029
rect 12614 3987 12644 4021
rect 12614 3953 12678 3987
rect 12712 4153 12746 4245
rect 12801 4245 12806 4279
rect 12840 4245 12843 4279
rect 12801 4229 12843 4245
rect 12895 4258 12911 4292
rect 12945 4258 12961 4292
rect 12895 4224 12961 4258
rect 12895 4190 12911 4224
rect 12945 4190 12961 4224
rect 12995 4263 13029 4335
rect 12995 4213 13029 4229
rect 13063 4290 13129 4291
rect 13063 4256 13079 4290
rect 13113 4267 13129 4290
rect 13063 4233 13093 4256
rect 13127 4233 13129 4267
rect 13063 4222 13129 4233
rect 13173 4274 14242 4335
rect 13173 4240 13191 4274
rect 13225 4240 14191 4274
rect 14225 4240 14242 4274
rect 13173 4226 14242 4240
rect 14277 4274 15346 4335
rect 14277 4240 14295 4274
rect 14329 4240 15295 4274
rect 15329 4240 15346 4274
rect 14277 4226 15346 4240
rect 15473 4263 15525 4301
rect 15473 4229 15491 4263
rect 15561 4293 15627 4335
rect 15561 4259 15577 4293
rect 15611 4259 15627 4293
rect 15663 4280 15697 4301
rect 12895 4187 12961 4190
rect 13063 4188 13079 4222
rect 13113 4204 13129 4222
rect 13113 4188 13139 4204
rect 13063 4187 13139 4188
rect 12921 4153 12961 4187
rect 13094 4179 13139 4187
rect 12712 4137 12887 4153
rect 12712 4103 12853 4137
rect 12712 4087 12887 4103
rect 12921 4137 13071 4153
rect 12921 4103 13037 4137
rect 12921 4087 13071 4103
rect 12474 3909 12524 3925
rect 12712 3919 12746 4087
rect 12921 4046 12959 4087
rect 13105 4063 13139 4179
rect 13096 4053 13139 4063
rect 13490 4111 13558 4226
rect 13490 4077 13507 4111
rect 13541 4077 13558 4111
rect 13490 4060 13558 4077
rect 13854 4147 13924 4162
rect 13854 4113 13871 4147
rect 13905 4113 13924 4147
rect 12780 4043 12959 4046
rect 12780 4021 12907 4043
rect 12814 4009 12907 4021
rect 12941 4009 12959 4043
rect 13061 4043 13139 4053
rect 12814 3987 12959 4009
rect 12780 3972 12959 3987
rect 12780 3971 12907 3972
rect 12891 3938 12907 3971
rect 12941 3938 12959 3972
rect 12474 3875 12490 3909
rect 12569 3885 12585 3919
rect 12619 3885 12746 3919
rect 12782 3909 12845 3925
rect 12474 3859 12524 3875
rect 12782 3875 12784 3909
rect 12818 3875 12845 3909
rect 12782 3825 12845 3875
rect 12891 3901 12959 3938
rect 12891 3867 12907 3901
rect 12941 3867 12959 3901
rect 12891 3859 12959 3867
rect 12993 4011 13027 4027
rect 12993 3931 13027 3977
rect 12993 3825 13027 3897
rect 13061 4009 13077 4043
rect 13111 4037 13139 4043
rect 13111 4009 13127 4037
rect 13061 3975 13127 4009
rect 13061 3941 13077 3975
rect 13111 3941 13127 3975
rect 13061 3907 13127 3941
rect 13854 3912 13924 4113
rect 14594 4111 14662 4226
rect 15473 4200 15525 4229
rect 15663 4225 15697 4246
rect 14594 4077 14611 4111
rect 14645 4077 14662 4111
rect 14594 4060 14662 4077
rect 14958 4147 15028 4162
rect 14958 4113 14975 4147
rect 15009 4113 15028 4147
rect 14958 3912 15028 4113
rect 15473 4040 15507 4200
rect 15564 4191 15697 4225
rect 15749 4274 16451 4335
rect 15749 4240 15767 4274
rect 15801 4240 16399 4274
rect 16433 4240 16451 4274
rect 15564 4140 15598 4191
rect 15749 4181 16451 4240
rect 16577 4241 16635 4335
rect 17083 4293 17133 4335
rect 16577 4207 16589 4241
rect 16623 4207 16635 4241
rect 16577 4190 16635 4207
rect 16893 4265 16959 4281
rect 16893 4231 16907 4265
rect 16941 4231 16959 4265
rect 17083 4259 17099 4293
rect 17083 4243 17133 4259
rect 17167 4293 17279 4301
rect 17167 4259 17183 4293
rect 17217 4259 17279 4293
rect 17167 4243 17279 4259
rect 16893 4209 16959 4231
rect 15541 4124 15598 4140
rect 15575 4090 15598 4124
rect 15541 4074 15598 4090
rect 15645 4137 15711 4155
rect 15645 4103 15661 4137
rect 15695 4131 15711 4137
rect 15645 4097 15669 4103
rect 15703 4097 15711 4131
rect 15645 4081 15711 4097
rect 15749 4111 16079 4181
rect 16893 4171 17171 4209
rect 17137 4153 17171 4171
rect 15749 4077 15827 4111
rect 15861 4077 15926 4111
rect 15960 4077 16025 4111
rect 16059 4077 16079 4111
rect 16113 4113 16133 4147
rect 16167 4113 16236 4147
rect 16270 4113 16339 4147
rect 16373 4113 16451 4147
rect 17137 4137 17195 4153
rect 15564 4045 15598 4074
rect 15473 3990 15527 4040
rect 15564 4011 15697 4045
rect 16113 4043 16451 4113
rect 16856 4103 16910 4137
rect 16944 4103 16991 4137
rect 16856 4087 16991 4103
rect 17035 4131 17051 4137
rect 17035 4097 17049 4131
rect 17085 4103 17103 4137
rect 17083 4097 17103 4103
rect 17035 4087 17103 4097
rect 17137 4103 17159 4137
rect 17193 4103 17195 4137
rect 17137 4087 17195 4103
rect 16856 4063 16909 4087
rect 15473 3956 15491 3990
rect 15525 3956 15527 3990
rect 15663 3977 15697 4011
rect 15473 3927 15527 3956
rect 13061 3873 13077 3907
rect 13111 3873 13127 3907
rect 13061 3868 13127 3873
rect 13173 3901 14242 3912
rect 13173 3867 13191 3901
rect 13225 3867 14191 3901
rect 14225 3867 14242 3901
rect 13173 3825 14242 3867
rect 14277 3901 15346 3912
rect 14277 3867 14295 3901
rect 14329 3867 15295 3901
rect 15329 3867 15346 3901
rect 14277 3825 15346 3867
rect 15473 3893 15485 3927
rect 15519 3909 15527 3927
rect 15473 3875 15491 3893
rect 15525 3875 15527 3909
rect 15473 3859 15527 3875
rect 15561 3943 15577 3977
rect 15611 3943 15627 3977
rect 15561 3909 15627 3943
rect 15561 3875 15577 3909
rect 15611 3875 15627 3909
rect 15561 3825 15627 3875
rect 15663 3909 15697 3943
rect 15663 3859 15697 3875
rect 15749 4003 16451 4043
rect 15749 3969 15767 4003
rect 15801 3969 16399 4003
rect 16433 3969 16451 4003
rect 15749 3901 16451 3969
rect 15749 3867 15767 3901
rect 15801 3867 16399 3901
rect 16433 3867 16451 3901
rect 15749 3825 16451 3867
rect 16577 4023 16635 4058
rect 16577 3989 16589 4023
rect 16623 3989 16635 4023
rect 16856 4029 16865 4063
rect 16899 4029 16909 4063
rect 17137 4037 17171 4087
rect 16856 4015 16909 4029
rect 16577 3930 16635 3989
rect 16983 4003 17171 4037
rect 16577 3896 16589 3930
rect 16623 3896 16635 3930
rect 16577 3825 16635 3896
rect 16893 3943 16949 3959
rect 16893 3909 16907 3943
rect 16941 3909 16949 3943
rect 16893 3825 16949 3909
rect 16983 3943 17043 4003
rect 17229 3969 17279 4243
rect 17313 4274 18382 4335
rect 17313 4240 17331 4274
rect 17365 4240 18331 4274
rect 18365 4240 18382 4274
rect 17313 4226 18382 4240
rect 18601 4272 18843 4335
rect 18601 4238 18619 4272
rect 18653 4238 18791 4272
rect 18825 4238 18843 4272
rect 17630 4111 17698 4226
rect 18601 4185 18843 4238
rect 17630 4077 17647 4111
rect 17681 4077 17698 4111
rect 17630 4060 17698 4077
rect 17994 4147 18064 4162
rect 17994 4113 18011 4147
rect 18045 4113 18064 4147
rect 16983 3909 16991 3943
rect 17025 3909 17043 3943
rect 16983 3893 17043 3909
rect 17083 3935 17099 3969
rect 17133 3935 17149 3969
rect 17083 3901 17149 3935
rect 17083 3867 17099 3901
rect 17133 3867 17149 3901
rect 17083 3825 17149 3867
rect 17187 3935 17203 3969
rect 17237 3935 17279 3969
rect 17187 3927 17279 3935
rect 17187 3901 17233 3927
rect 17187 3867 17203 3901
rect 17267 3893 17279 3927
rect 17994 3912 18064 4113
rect 18601 4117 18651 4151
rect 18685 4117 18705 4151
rect 18601 4043 18705 4117
rect 18739 4111 18843 4185
rect 18739 4077 18759 4111
rect 18793 4077 18843 4111
rect 18601 3996 18843 4043
rect 18601 3962 18619 3996
rect 18653 3962 18791 3996
rect 18825 3962 18843 3996
rect 17237 3867 17279 3893
rect 17187 3859 17279 3867
rect 17313 3901 18382 3912
rect 17313 3867 17331 3901
rect 17365 3867 18331 3901
rect 18365 3867 18382 3901
rect 17313 3825 18382 3867
rect 18601 3901 18843 3962
rect 18601 3867 18619 3901
rect 18653 3867 18791 3901
rect 18825 3867 18843 3901
rect 18601 3825 18843 3867
rect 1104 3791 1133 3825
rect 1167 3791 1225 3825
rect 1259 3791 1317 3825
rect 1351 3791 1409 3825
rect 1443 3791 1501 3825
rect 1535 3791 1593 3825
rect 1627 3791 1685 3825
rect 1719 3791 1777 3825
rect 1811 3791 1869 3825
rect 1903 3791 1961 3825
rect 1995 3791 2053 3825
rect 2087 3791 2145 3825
rect 2179 3791 2237 3825
rect 2271 3791 2329 3825
rect 2363 3791 2421 3825
rect 2455 3791 2513 3825
rect 2547 3791 2605 3825
rect 2639 3791 2697 3825
rect 2731 3791 2789 3825
rect 2823 3791 2881 3825
rect 2915 3791 2973 3825
rect 3007 3791 3065 3825
rect 3099 3791 3157 3825
rect 3191 3791 3249 3825
rect 3283 3791 3341 3825
rect 3375 3791 3433 3825
rect 3467 3791 3525 3825
rect 3559 3791 3617 3825
rect 3651 3791 3709 3825
rect 3743 3791 3801 3825
rect 3835 3791 3893 3825
rect 3927 3791 3985 3825
rect 4019 3791 4077 3825
rect 4111 3791 4169 3825
rect 4203 3791 4261 3825
rect 4295 3791 4353 3825
rect 4387 3791 4445 3825
rect 4479 3791 4537 3825
rect 4571 3791 4629 3825
rect 4663 3791 4721 3825
rect 4755 3791 4813 3825
rect 4847 3791 4905 3825
rect 4939 3791 4997 3825
rect 5031 3791 5089 3825
rect 5123 3791 5181 3825
rect 5215 3791 5273 3825
rect 5307 3791 5365 3825
rect 5399 3791 5457 3825
rect 5491 3791 5549 3825
rect 5583 3791 5641 3825
rect 5675 3791 5733 3825
rect 5767 3791 5825 3825
rect 5859 3791 5917 3825
rect 5951 3791 6009 3825
rect 6043 3791 6101 3825
rect 6135 3791 6193 3825
rect 6227 3791 6285 3825
rect 6319 3791 6377 3825
rect 6411 3791 6469 3825
rect 6503 3791 6561 3825
rect 6595 3791 6653 3825
rect 6687 3791 6745 3825
rect 6779 3791 6837 3825
rect 6871 3791 6929 3825
rect 6963 3791 7021 3825
rect 7055 3791 7113 3825
rect 7147 3791 7205 3825
rect 7239 3791 7297 3825
rect 7331 3791 7389 3825
rect 7423 3791 7481 3825
rect 7515 3791 7573 3825
rect 7607 3791 7665 3825
rect 7699 3791 7757 3825
rect 7791 3791 7849 3825
rect 7883 3791 7941 3825
rect 7975 3791 8033 3825
rect 8067 3791 8125 3825
rect 8159 3791 8217 3825
rect 8251 3791 8309 3825
rect 8343 3791 8401 3825
rect 8435 3791 8493 3825
rect 8527 3791 8585 3825
rect 8619 3791 8677 3825
rect 8711 3791 8769 3825
rect 8803 3791 8861 3825
rect 8895 3791 8953 3825
rect 8987 3791 9045 3825
rect 9079 3791 9137 3825
rect 9171 3791 9229 3825
rect 9263 3791 9321 3825
rect 9355 3791 9413 3825
rect 9447 3791 9505 3825
rect 9539 3791 9597 3825
rect 9631 3791 9689 3825
rect 9723 3791 9781 3825
rect 9815 3791 9873 3825
rect 9907 3791 9965 3825
rect 9999 3791 10057 3825
rect 10091 3791 10149 3825
rect 10183 3791 10241 3825
rect 10275 3791 10333 3825
rect 10367 3791 10425 3825
rect 10459 3791 10517 3825
rect 10551 3791 10609 3825
rect 10643 3791 10701 3825
rect 10735 3791 10793 3825
rect 10827 3791 10885 3825
rect 10919 3791 10977 3825
rect 11011 3791 11069 3825
rect 11103 3791 11161 3825
rect 11195 3791 11253 3825
rect 11287 3791 11345 3825
rect 11379 3791 11437 3825
rect 11471 3791 11529 3825
rect 11563 3791 11621 3825
rect 11655 3791 11713 3825
rect 11747 3791 11805 3825
rect 11839 3791 11897 3825
rect 11931 3791 11989 3825
rect 12023 3791 12081 3825
rect 12115 3791 12173 3825
rect 12207 3791 12265 3825
rect 12299 3791 12357 3825
rect 12391 3791 12449 3825
rect 12483 3791 12541 3825
rect 12575 3791 12633 3825
rect 12667 3791 12725 3825
rect 12759 3791 12817 3825
rect 12851 3791 12909 3825
rect 12943 3791 13001 3825
rect 13035 3791 13093 3825
rect 13127 3791 13185 3825
rect 13219 3791 13277 3825
rect 13311 3791 13369 3825
rect 13403 3791 13461 3825
rect 13495 3791 13553 3825
rect 13587 3791 13645 3825
rect 13679 3791 13737 3825
rect 13771 3791 13829 3825
rect 13863 3791 13921 3825
rect 13955 3791 14013 3825
rect 14047 3791 14105 3825
rect 14139 3791 14197 3825
rect 14231 3791 14289 3825
rect 14323 3791 14381 3825
rect 14415 3791 14473 3825
rect 14507 3791 14565 3825
rect 14599 3791 14657 3825
rect 14691 3791 14749 3825
rect 14783 3791 14841 3825
rect 14875 3791 14933 3825
rect 14967 3791 15025 3825
rect 15059 3791 15117 3825
rect 15151 3791 15209 3825
rect 15243 3791 15301 3825
rect 15335 3791 15393 3825
rect 15427 3791 15485 3825
rect 15519 3791 15577 3825
rect 15611 3791 15669 3825
rect 15703 3791 15761 3825
rect 15795 3791 15853 3825
rect 15887 3791 15945 3825
rect 15979 3791 16037 3825
rect 16071 3791 16129 3825
rect 16163 3791 16221 3825
rect 16255 3791 16313 3825
rect 16347 3791 16405 3825
rect 16439 3791 16497 3825
rect 16531 3791 16589 3825
rect 16623 3791 16681 3825
rect 16715 3791 16773 3825
rect 16807 3791 16865 3825
rect 16899 3791 16957 3825
rect 16991 3791 17049 3825
rect 17083 3791 17141 3825
rect 17175 3791 17233 3825
rect 17267 3791 17325 3825
rect 17359 3791 17417 3825
rect 17451 3791 17509 3825
rect 17543 3791 17601 3825
rect 17635 3791 17693 3825
rect 17727 3791 17785 3825
rect 17819 3791 17877 3825
rect 17911 3791 17969 3825
rect 18003 3791 18061 3825
rect 18095 3791 18153 3825
rect 18187 3791 18245 3825
rect 18279 3791 18337 3825
rect 18371 3791 18429 3825
rect 18463 3791 18521 3825
rect 18555 3791 18613 3825
rect 18647 3791 18705 3825
rect 18739 3791 18797 3825
rect 18831 3791 18860 3825
rect 1121 3749 1363 3791
rect 1121 3715 1139 3749
rect 1173 3715 1311 3749
rect 1345 3715 1363 3749
rect 1121 3654 1363 3715
rect 1121 3620 1139 3654
rect 1173 3620 1311 3654
rect 1345 3620 1363 3654
rect 1121 3573 1363 3620
rect 1397 3749 1915 3791
rect 1397 3715 1415 3749
rect 1449 3715 1863 3749
rect 1897 3715 1915 3749
rect 1397 3647 1915 3715
rect 1397 3613 1415 3647
rect 1449 3613 1863 3647
rect 1897 3613 1915 3647
rect 2059 3741 2093 3757
rect 2059 3673 2093 3707
rect 2127 3725 2193 3791
rect 2127 3691 2143 3725
rect 2177 3691 2193 3725
rect 2227 3741 2264 3757
rect 2261 3707 2264 3741
rect 2227 3673 2264 3707
rect 2312 3749 2365 3791
rect 2312 3715 2331 3749
rect 2312 3699 2365 3715
rect 2399 3741 2449 3757
rect 2399 3707 2415 3741
rect 2746 3749 2780 3791
rect 2093 3655 2192 3657
rect 2093 3639 2150 3655
rect 2059 3623 2150 3639
rect 1397 3573 1915 3613
rect 2146 3621 2150 3623
rect 2184 3621 2192 3655
rect 1121 3505 1171 3539
rect 1205 3505 1225 3539
rect 1121 3431 1225 3505
rect 1259 3499 1363 3573
rect 1259 3465 1279 3499
rect 1313 3465 1363 3499
rect 1397 3505 1475 3539
rect 1509 3505 1585 3539
rect 1619 3505 1639 3539
rect 1397 3435 1639 3505
rect 1673 3503 1915 3573
rect 1673 3469 1693 3503
rect 1727 3469 1803 3503
rect 1837 3469 1915 3503
rect 2042 3519 2112 3589
rect 2042 3485 2053 3519
rect 2087 3513 2112 3519
rect 2042 3479 2056 3485
rect 2090 3479 2112 3513
rect 2042 3459 2112 3479
rect 2146 3528 2192 3621
rect 2146 3494 2158 3528
rect 1121 3378 1363 3431
rect 1121 3344 1139 3378
rect 1173 3344 1311 3378
rect 1345 3344 1363 3378
rect 1121 3281 1363 3344
rect 1397 3376 1915 3435
rect 2146 3425 2192 3494
rect 1397 3342 1415 3376
rect 1449 3342 1863 3376
rect 1897 3342 1915 3376
rect 1397 3281 1915 3342
rect 2059 3391 2192 3425
rect 2261 3639 2264 3673
rect 2399 3672 2449 3707
rect 2491 3702 2507 3736
rect 2541 3702 2712 3736
rect 2227 3587 2264 3639
rect 2388 3646 2449 3672
rect 2538 3655 2644 3668
rect 2227 3553 2229 3587
rect 2263 3553 2264 3587
rect 2059 3383 2093 3391
rect 2227 3383 2264 3553
rect 2298 3581 2354 3597
rect 2298 3547 2320 3581
rect 2298 3451 2354 3547
rect 2298 3417 2320 3451
rect 2298 3407 2354 3417
rect 2388 3425 2422 3646
rect 2538 3621 2570 3655
rect 2604 3629 2644 3655
rect 2456 3587 2504 3608
rect 2456 3553 2467 3587
rect 2501 3553 2504 3587
rect 2456 3551 2504 3553
rect 2456 3517 2463 3551
rect 2497 3517 2504 3551
rect 2456 3489 2504 3517
rect 2538 3455 2572 3621
rect 2606 3595 2644 3629
rect 2678 3579 2712 3702
rect 2746 3681 2780 3715
rect 2746 3631 2780 3647
rect 2814 3741 2864 3757
rect 2814 3707 2830 3741
rect 3122 3741 3185 3791
rect 2814 3691 2864 3707
rect 2909 3697 2925 3731
rect 2959 3697 3086 3731
rect 2678 3563 2780 3579
rect 2678 3561 2746 3563
rect 2388 3399 2433 3425
rect 2467 3421 2483 3455
rect 2517 3421 2572 3455
rect 2467 3411 2572 3421
rect 2606 3529 2746 3561
rect 2606 3527 2780 3529
rect 2059 3333 2093 3349
rect 2127 3323 2143 3357
rect 2177 3323 2193 3357
rect 2261 3349 2264 3383
rect 2227 3333 2264 3349
rect 2315 3357 2365 3373
rect 2127 3281 2193 3323
rect 2315 3323 2331 3357
rect 2399 3371 2433 3399
rect 2606 3371 2640 3527
rect 2746 3513 2780 3527
rect 2682 3477 2722 3483
rect 2814 3477 2848 3691
rect 2882 3655 2920 3657
rect 2882 3621 2884 3655
rect 2918 3621 2920 3655
rect 2882 3563 2920 3621
rect 2916 3529 2920 3563
rect 2882 3513 2920 3529
rect 2954 3629 3018 3663
rect 2954 3595 2984 3629
rect 2954 3587 3018 3595
rect 2954 3553 2971 3587
rect 3005 3553 3018 3587
rect 2682 3467 2848 3477
rect 2954 3471 3018 3553
rect 2716 3433 2848 3467
rect 2682 3417 2848 3433
rect 2399 3337 2416 3371
rect 2450 3337 2466 3371
rect 2505 3337 2527 3371
rect 2561 3337 2640 3371
rect 2704 3365 2778 3381
rect 2315 3281 2365 3323
rect 2704 3331 2726 3365
rect 2760 3331 2778 3365
rect 2814 3371 2848 3417
rect 2925 3455 3018 3471
rect 2959 3421 3018 3455
rect 2925 3405 3018 3421
rect 3052 3529 3086 3697
rect 3122 3707 3124 3741
rect 3158 3707 3185 3741
rect 3122 3691 3185 3707
rect 3231 3749 3299 3757
rect 3231 3715 3247 3749
rect 3281 3715 3299 3749
rect 3231 3678 3299 3715
rect 3231 3645 3247 3678
rect 3120 3644 3247 3645
rect 3281 3644 3299 3678
rect 3120 3629 3299 3644
rect 3154 3607 3299 3629
rect 3154 3595 3247 3607
rect 3120 3573 3247 3595
rect 3281 3573 3299 3607
rect 3333 3719 3367 3791
rect 3333 3639 3367 3685
rect 3333 3589 3367 3605
rect 3401 3743 3467 3748
rect 3401 3709 3417 3743
rect 3451 3723 3467 3743
rect 3401 3689 3433 3709
rect 3401 3675 3467 3689
rect 3401 3641 3417 3675
rect 3451 3641 3467 3675
rect 3401 3607 3467 3641
rect 3120 3570 3299 3573
rect 3261 3529 3299 3570
rect 3401 3573 3417 3607
rect 3451 3579 3467 3607
rect 3697 3720 3755 3791
rect 3697 3686 3709 3720
rect 3743 3686 3755 3720
rect 3697 3627 3755 3686
rect 3697 3593 3709 3627
rect 3743 3593 3755 3627
rect 3991 3741 4025 3757
rect 3991 3673 4025 3707
rect 4059 3725 4125 3791
rect 4059 3691 4075 3725
rect 4109 3691 4125 3725
rect 4159 3741 4196 3757
rect 4193 3707 4196 3741
rect 4159 3673 4196 3707
rect 4244 3749 4297 3791
rect 4244 3715 4263 3749
rect 4244 3699 4297 3715
rect 4331 3741 4381 3757
rect 4331 3707 4347 3741
rect 4678 3749 4712 3791
rect 4025 3655 4124 3657
rect 4025 3639 4082 3655
rect 3991 3623 4082 3639
rect 3451 3573 3479 3579
rect 3401 3563 3479 3573
rect 3436 3553 3479 3563
rect 3697 3558 3755 3593
rect 4078 3621 4082 3623
rect 4116 3621 4124 3655
rect 3974 3587 4044 3589
rect 3052 3513 3227 3529
rect 3052 3479 3193 3513
rect 3052 3463 3227 3479
rect 3261 3513 3411 3529
rect 3261 3479 3377 3513
rect 3261 3463 3411 3479
rect 3052 3371 3086 3463
rect 3261 3429 3301 3463
rect 3445 3437 3479 3553
rect 3974 3553 3985 3587
rect 4019 3553 4044 3587
rect 3974 3513 4044 3553
rect 3974 3479 3988 3513
rect 4022 3479 4044 3513
rect 3974 3459 4044 3479
rect 4078 3528 4124 3621
rect 4078 3494 4090 3528
rect 3434 3429 3479 3437
rect 3235 3426 3301 3429
rect 3235 3392 3251 3426
rect 3285 3392 3301 3426
rect 3403 3428 3479 3429
rect 2814 3337 2845 3371
rect 2879 3337 2895 3371
rect 2929 3337 2948 3371
rect 2982 3337 3086 3371
rect 3141 3371 3183 3387
rect 3141 3337 3146 3371
rect 3180 3337 3183 3371
rect 2704 3281 2778 3331
rect 3141 3281 3183 3337
rect 3235 3358 3301 3392
rect 3235 3324 3251 3358
rect 3285 3324 3301 3358
rect 3335 3387 3369 3403
rect 3335 3281 3369 3353
rect 3403 3394 3419 3428
rect 3453 3412 3479 3428
rect 3453 3394 3469 3412
rect 3403 3360 3469 3394
rect 3403 3326 3419 3360
rect 3453 3326 3469 3360
rect 3403 3325 3469 3326
rect 3697 3409 3755 3426
rect 4078 3425 4124 3494
rect 3697 3375 3709 3409
rect 3743 3375 3755 3409
rect 3697 3281 3755 3375
rect 3991 3391 4124 3425
rect 4193 3639 4196 3673
rect 4331 3672 4381 3707
rect 4423 3702 4439 3736
rect 4473 3702 4644 3736
rect 4159 3587 4196 3639
rect 4320 3646 4381 3672
rect 4470 3655 4576 3668
rect 4159 3553 4161 3587
rect 4195 3553 4196 3587
rect 3991 3383 4025 3391
rect 4159 3383 4196 3553
rect 4230 3581 4286 3597
rect 4230 3547 4252 3581
rect 4230 3519 4286 3547
rect 4230 3485 4252 3519
rect 4230 3407 4286 3485
rect 4320 3425 4354 3646
rect 4470 3621 4502 3655
rect 4536 3629 4576 3655
rect 4388 3587 4436 3608
rect 4388 3553 4399 3587
rect 4433 3553 4436 3587
rect 4388 3551 4436 3553
rect 4388 3517 4395 3551
rect 4429 3517 4436 3551
rect 4388 3489 4436 3517
rect 4470 3455 4504 3621
rect 4538 3595 4576 3629
rect 4610 3579 4644 3702
rect 4678 3681 4712 3715
rect 4678 3631 4712 3647
rect 4746 3741 4796 3757
rect 4746 3707 4762 3741
rect 5054 3741 5117 3791
rect 4746 3691 4796 3707
rect 4841 3697 4857 3731
rect 4891 3697 5018 3731
rect 4610 3563 4712 3579
rect 4610 3561 4678 3563
rect 4320 3399 4365 3425
rect 4399 3421 4415 3455
rect 4449 3421 4504 3455
rect 4399 3411 4504 3421
rect 4538 3529 4678 3561
rect 4538 3527 4712 3529
rect 3991 3333 4025 3349
rect 4059 3323 4075 3357
rect 4109 3323 4125 3357
rect 4193 3349 4196 3383
rect 4159 3333 4196 3349
rect 4247 3357 4297 3373
rect 4059 3281 4125 3323
rect 4247 3323 4263 3357
rect 4331 3371 4365 3399
rect 4538 3371 4572 3527
rect 4678 3513 4712 3527
rect 4614 3477 4654 3483
rect 4746 3477 4780 3691
rect 4814 3655 4852 3657
rect 4814 3621 4816 3655
rect 4850 3621 4852 3655
rect 4814 3563 4852 3621
rect 4848 3529 4852 3563
rect 4814 3513 4852 3529
rect 4886 3629 4950 3663
rect 4886 3595 4916 3629
rect 4886 3587 4950 3595
rect 4886 3553 4903 3587
rect 4937 3553 4950 3587
rect 4614 3467 4780 3477
rect 4886 3471 4950 3553
rect 4648 3433 4780 3467
rect 4614 3417 4780 3433
rect 4331 3337 4348 3371
rect 4382 3337 4398 3371
rect 4437 3337 4459 3371
rect 4493 3337 4572 3371
rect 4636 3365 4710 3381
rect 4247 3281 4297 3323
rect 4636 3331 4658 3365
rect 4692 3331 4710 3365
rect 4746 3371 4780 3417
rect 4857 3455 4950 3471
rect 4891 3421 4950 3455
rect 4857 3405 4950 3421
rect 4984 3529 5018 3697
rect 5054 3707 5056 3741
rect 5090 3707 5117 3741
rect 5054 3691 5117 3707
rect 5163 3749 5231 3757
rect 5163 3715 5179 3749
rect 5213 3715 5231 3749
rect 5163 3678 5231 3715
rect 5163 3645 5179 3678
rect 5052 3644 5179 3645
rect 5213 3644 5231 3678
rect 5052 3629 5231 3644
rect 5086 3607 5231 3629
rect 5086 3595 5179 3607
rect 5052 3573 5179 3595
rect 5213 3573 5231 3607
rect 5265 3719 5299 3791
rect 5445 3749 6147 3791
rect 5265 3639 5299 3685
rect 5265 3589 5299 3605
rect 5333 3743 5399 3748
rect 5333 3709 5349 3743
rect 5383 3709 5399 3743
rect 5333 3675 5399 3709
rect 5333 3641 5349 3675
rect 5383 3641 5399 3675
rect 5333 3607 5399 3641
rect 5052 3570 5231 3573
rect 5193 3529 5231 3570
rect 5333 3573 5349 3607
rect 5383 3579 5399 3607
rect 5445 3715 5463 3749
rect 5497 3715 6095 3749
rect 6129 3715 6147 3749
rect 5445 3647 6147 3715
rect 5445 3613 5463 3647
rect 5497 3613 6095 3647
rect 6129 3613 6147 3647
rect 5383 3573 5411 3579
rect 5445 3573 6147 3613
rect 5333 3563 5411 3573
rect 5368 3553 5411 3563
rect 4984 3513 5159 3529
rect 4984 3479 5125 3513
rect 4984 3463 5159 3479
rect 5193 3513 5343 3529
rect 5193 3479 5309 3513
rect 5193 3463 5343 3479
rect 4984 3371 5018 3463
rect 5193 3429 5233 3463
rect 5377 3437 5411 3553
rect 5366 3429 5411 3437
rect 5167 3426 5233 3429
rect 5167 3392 5183 3426
rect 5217 3392 5233 3426
rect 5335 3428 5411 3429
rect 4746 3337 4777 3371
rect 4811 3337 4827 3371
rect 4861 3337 4880 3371
rect 4914 3337 5018 3371
rect 5073 3371 5115 3387
rect 5073 3337 5078 3371
rect 5112 3337 5115 3371
rect 4636 3281 4710 3331
rect 5073 3281 5115 3337
rect 5167 3358 5233 3392
rect 5167 3324 5183 3358
rect 5217 3324 5233 3358
rect 5267 3387 5301 3403
rect 5267 3281 5301 3353
rect 5335 3394 5351 3428
rect 5385 3412 5411 3428
rect 5445 3505 5523 3539
rect 5557 3505 5622 3539
rect 5656 3505 5721 3539
rect 5755 3505 5775 3539
rect 5445 3435 5775 3505
rect 5809 3503 6147 3573
rect 5809 3469 5829 3503
rect 5863 3469 5932 3503
rect 5966 3469 6035 3503
rect 6069 3469 6147 3503
rect 6273 3741 6329 3757
rect 6273 3707 6295 3741
rect 6273 3673 6329 3707
rect 6273 3639 6295 3673
rect 6273 3605 6329 3639
rect 6363 3749 6505 3791
rect 6363 3715 6381 3749
rect 6415 3715 6455 3749
rect 6489 3715 6505 3749
rect 6363 3681 6505 3715
rect 6363 3647 6381 3681
rect 6415 3647 6455 3681
rect 6489 3647 6505 3681
rect 6363 3636 6505 3647
rect 6539 3749 6605 3757
rect 6539 3715 6555 3749
rect 6589 3715 6605 3749
rect 6723 3749 6789 3791
rect 6539 3681 6605 3715
rect 6539 3647 6555 3681
rect 6589 3647 6605 3681
rect 6273 3571 6295 3605
rect 6539 3613 6605 3647
rect 6539 3602 6555 3613
rect 6273 3470 6329 3571
rect 6375 3579 6555 3602
rect 6589 3579 6605 3613
rect 6375 3559 6605 3579
rect 6644 3723 6687 3742
rect 6644 3689 6653 3723
rect 6375 3513 6432 3559
rect 6409 3479 6432 3513
rect 6469 3519 6563 3525
rect 6644 3519 6687 3689
rect 6723 3715 6739 3749
rect 6773 3715 6789 3749
rect 6723 3681 6789 3715
rect 6723 3647 6739 3681
rect 6773 3647 6789 3681
rect 6825 3749 7159 3791
rect 6825 3715 6843 3749
rect 6877 3715 7107 3749
rect 7141 3715 7159 3749
rect 6825 3647 7159 3715
rect 6825 3613 6843 3647
rect 6877 3613 7107 3647
rect 7141 3613 7159 3647
rect 7211 3741 7245 3757
rect 7211 3673 7245 3707
rect 7279 3725 7345 3791
rect 7279 3691 7295 3725
rect 7329 3691 7345 3725
rect 7379 3741 7416 3757
rect 7413 3707 7416 3741
rect 7379 3673 7416 3707
rect 7464 3749 7517 3791
rect 7464 3715 7483 3749
rect 7464 3699 7517 3715
rect 7551 3741 7601 3757
rect 7551 3707 7567 3741
rect 7898 3749 7932 3791
rect 7245 3655 7344 3657
rect 7245 3639 7302 3655
rect 7211 3623 7302 3639
rect 6745 3519 6791 3587
rect 6825 3573 7159 3613
rect 7298 3621 7302 3623
rect 7336 3621 7344 3655
rect 6503 3513 6563 3519
rect 6503 3485 6513 3513
rect 6469 3479 6513 3485
rect 6547 3479 6563 3513
rect 6597 3513 6687 3519
rect 6597 3479 6613 3513
rect 6647 3483 6687 3513
rect 6725 3513 6745 3519
rect 6647 3479 6663 3483
rect 6725 3479 6741 3513
rect 6779 3485 6791 3519
rect 6775 3479 6791 3485
rect 6825 3505 6845 3539
rect 6879 3505 6975 3539
rect 6273 3451 6341 3470
rect 5385 3394 5401 3412
rect 5335 3383 5401 3394
rect 5335 3360 5365 3383
rect 5335 3326 5351 3360
rect 5399 3349 5401 3383
rect 5385 3326 5401 3349
rect 5335 3325 5401 3326
rect 5445 3376 6147 3435
rect 5445 3342 5463 3376
rect 5497 3342 6095 3376
rect 6129 3342 6147 3376
rect 5445 3281 6147 3342
rect 6273 3417 6285 3451
rect 6319 3428 6341 3451
rect 6273 3394 6291 3417
rect 6325 3394 6341 3428
rect 6375 3445 6432 3479
rect 6375 3429 6517 3445
rect 6375 3407 6479 3429
rect 6273 3360 6341 3394
rect 6457 3395 6479 3407
rect 6513 3395 6517 3429
rect 6457 3379 6517 3395
rect 6555 3429 6791 3445
rect 6555 3425 6739 3429
rect 6555 3391 6571 3425
rect 6605 3407 6739 3425
rect 6605 3391 6621 3407
rect 6723 3395 6739 3407
rect 6773 3395 6791 3429
rect 6457 3377 6520 3379
rect 6457 3375 6522 3377
rect 6457 3374 6524 3375
rect 6273 3326 6291 3360
rect 6325 3326 6341 3360
rect 6273 3315 6341 3326
rect 6375 3357 6409 3373
rect 6375 3281 6409 3323
rect 6457 3372 6525 3374
rect 6457 3371 6526 3372
rect 6457 3369 6527 3371
rect 6457 3368 6528 3369
rect 6457 3361 6529 3368
rect 6457 3327 6479 3361
rect 6513 3327 6529 3361
rect 6457 3315 6529 3327
rect 6655 3357 6689 3373
rect 6655 3281 6689 3323
rect 6723 3361 6791 3395
rect 6723 3327 6739 3361
rect 6773 3327 6791 3361
rect 6723 3315 6791 3327
rect 6825 3435 6975 3505
rect 7009 3503 7159 3573
rect 7009 3469 7105 3503
rect 7139 3469 7159 3503
rect 7194 3587 7264 3589
rect 7194 3553 7205 3587
rect 7239 3553 7264 3587
rect 7194 3513 7264 3553
rect 7194 3479 7208 3513
rect 7242 3479 7264 3513
rect 7194 3459 7264 3479
rect 7298 3528 7344 3621
rect 7298 3494 7310 3528
rect 6825 3383 7159 3435
rect 7298 3425 7344 3494
rect 6825 3349 6843 3383
rect 6877 3349 7107 3383
rect 7141 3349 7159 3383
rect 6825 3281 7159 3349
rect 7211 3391 7344 3425
rect 7413 3639 7416 3673
rect 7551 3672 7601 3707
rect 7643 3702 7659 3736
rect 7693 3702 7864 3736
rect 7379 3587 7416 3639
rect 7540 3646 7601 3672
rect 7690 3655 7796 3668
rect 7379 3553 7381 3587
rect 7415 3553 7416 3587
rect 7211 3383 7245 3391
rect 7379 3383 7416 3553
rect 7450 3581 7506 3597
rect 7450 3547 7472 3581
rect 7450 3519 7506 3547
rect 7450 3485 7472 3519
rect 7450 3407 7506 3485
rect 7540 3425 7574 3646
rect 7690 3621 7722 3655
rect 7756 3629 7796 3655
rect 7608 3587 7656 3608
rect 7608 3553 7619 3587
rect 7653 3553 7656 3587
rect 7608 3551 7656 3553
rect 7608 3517 7615 3551
rect 7649 3517 7656 3551
rect 7608 3489 7656 3517
rect 7690 3455 7724 3621
rect 7758 3595 7796 3629
rect 7830 3579 7864 3702
rect 7898 3681 7932 3715
rect 7898 3631 7932 3647
rect 7966 3741 8016 3757
rect 7966 3707 7982 3741
rect 8274 3741 8337 3791
rect 7966 3691 8016 3707
rect 8061 3697 8077 3731
rect 8111 3697 8238 3731
rect 7830 3563 7932 3579
rect 7830 3561 7898 3563
rect 7540 3399 7585 3425
rect 7619 3421 7635 3455
rect 7669 3421 7724 3455
rect 7619 3411 7724 3421
rect 7758 3529 7898 3561
rect 7758 3527 7932 3529
rect 7211 3333 7245 3349
rect 7279 3323 7295 3357
rect 7329 3323 7345 3357
rect 7413 3349 7416 3383
rect 7379 3333 7416 3349
rect 7467 3357 7517 3373
rect 7279 3281 7345 3323
rect 7467 3323 7483 3357
rect 7551 3371 7585 3399
rect 7758 3371 7792 3527
rect 7898 3513 7932 3527
rect 7834 3477 7874 3483
rect 7966 3477 8000 3691
rect 8034 3655 8072 3657
rect 8034 3621 8036 3655
rect 8070 3621 8072 3655
rect 8034 3563 8072 3621
rect 8068 3529 8072 3563
rect 8034 3513 8072 3529
rect 8106 3629 8170 3663
rect 8106 3595 8136 3629
rect 8106 3587 8170 3595
rect 8106 3553 8123 3587
rect 8157 3553 8170 3587
rect 7834 3467 8000 3477
rect 8106 3471 8170 3553
rect 7868 3433 8000 3467
rect 7834 3417 8000 3433
rect 7551 3337 7568 3371
rect 7602 3337 7618 3371
rect 7657 3337 7679 3371
rect 7713 3337 7792 3371
rect 7856 3365 7930 3381
rect 7467 3281 7517 3323
rect 7856 3331 7878 3365
rect 7912 3331 7930 3365
rect 7966 3371 8000 3417
rect 8077 3455 8170 3471
rect 8111 3421 8170 3455
rect 8077 3405 8170 3421
rect 8204 3529 8238 3697
rect 8274 3707 8276 3741
rect 8310 3707 8337 3741
rect 8274 3691 8337 3707
rect 8383 3749 8451 3757
rect 8383 3715 8399 3749
rect 8433 3715 8451 3749
rect 8383 3678 8451 3715
rect 8383 3645 8399 3678
rect 8272 3644 8399 3645
rect 8433 3644 8451 3678
rect 8272 3629 8451 3644
rect 8306 3607 8451 3629
rect 8306 3595 8399 3607
rect 8272 3573 8399 3595
rect 8433 3573 8451 3607
rect 8485 3719 8519 3791
rect 8485 3639 8519 3685
rect 8485 3589 8519 3605
rect 8553 3743 8619 3748
rect 8553 3709 8569 3743
rect 8603 3723 8619 3743
rect 8553 3689 8585 3709
rect 8553 3675 8619 3689
rect 8553 3641 8569 3675
rect 8603 3641 8619 3675
rect 8553 3607 8619 3641
rect 8272 3570 8451 3573
rect 8413 3529 8451 3570
rect 8553 3573 8569 3607
rect 8603 3579 8619 3607
rect 8849 3720 8907 3791
rect 8849 3686 8861 3720
rect 8895 3686 8907 3720
rect 8849 3627 8907 3686
rect 8849 3593 8861 3627
rect 8895 3593 8907 3627
rect 8603 3573 8631 3579
rect 8553 3563 8631 3573
rect 8588 3553 8631 3563
rect 8849 3558 8907 3593
rect 8941 3749 9643 3791
rect 8941 3715 8959 3749
rect 8993 3715 9591 3749
rect 9625 3715 9643 3749
rect 8941 3647 9643 3715
rect 8941 3613 8959 3647
rect 8993 3613 9591 3647
rect 9625 3613 9643 3647
rect 9787 3741 9821 3757
rect 9787 3673 9821 3707
rect 9855 3725 9921 3791
rect 9855 3691 9871 3725
rect 9905 3691 9921 3725
rect 9955 3741 9992 3757
rect 9989 3707 9992 3741
rect 9955 3673 9992 3707
rect 10040 3749 10093 3791
rect 10040 3715 10059 3749
rect 10040 3699 10093 3715
rect 10127 3741 10177 3757
rect 10127 3707 10143 3741
rect 10474 3749 10508 3791
rect 9821 3655 9920 3657
rect 9821 3639 9878 3655
rect 9787 3623 9878 3639
rect 8941 3573 9643 3613
rect 9874 3621 9878 3623
rect 9912 3621 9920 3655
rect 8204 3513 8379 3529
rect 8204 3479 8345 3513
rect 8204 3463 8379 3479
rect 8413 3513 8563 3529
rect 8413 3479 8529 3513
rect 8413 3463 8563 3479
rect 8204 3371 8238 3463
rect 8413 3429 8453 3463
rect 8597 3437 8631 3553
rect 8586 3429 8631 3437
rect 8387 3426 8453 3429
rect 8387 3392 8403 3426
rect 8437 3392 8453 3426
rect 8555 3428 8631 3429
rect 7966 3337 7997 3371
rect 8031 3337 8047 3371
rect 8081 3337 8100 3371
rect 8134 3337 8238 3371
rect 8293 3371 8335 3387
rect 8293 3337 8298 3371
rect 8332 3337 8335 3371
rect 7856 3281 7930 3331
rect 8293 3281 8335 3337
rect 8387 3358 8453 3392
rect 8387 3324 8403 3358
rect 8437 3324 8453 3358
rect 8487 3387 8521 3403
rect 8487 3281 8521 3353
rect 8555 3394 8571 3428
rect 8605 3412 8631 3428
rect 8941 3505 9019 3539
rect 9053 3505 9118 3539
rect 9152 3505 9217 3539
rect 9251 3505 9271 3539
rect 8941 3435 9271 3505
rect 9305 3503 9643 3573
rect 9305 3469 9325 3503
rect 9359 3469 9428 3503
rect 9462 3469 9531 3503
rect 9565 3469 9643 3503
rect 9770 3587 9840 3589
rect 9770 3553 9781 3587
rect 9815 3553 9840 3587
rect 9770 3513 9840 3553
rect 9770 3479 9784 3513
rect 9818 3479 9840 3513
rect 9770 3459 9840 3479
rect 9874 3528 9920 3621
rect 9874 3494 9886 3528
rect 8605 3394 8621 3412
rect 8555 3360 8621 3394
rect 8555 3326 8571 3360
rect 8605 3326 8621 3360
rect 8555 3325 8621 3326
rect 8849 3409 8907 3426
rect 8849 3375 8861 3409
rect 8895 3375 8907 3409
rect 8849 3281 8907 3375
rect 8941 3376 9643 3435
rect 9874 3425 9920 3494
rect 8941 3342 8959 3376
rect 8993 3342 9591 3376
rect 9625 3342 9643 3376
rect 8941 3281 9643 3342
rect 9787 3391 9920 3425
rect 9989 3639 9992 3673
rect 10127 3672 10177 3707
rect 10219 3702 10235 3736
rect 10269 3702 10440 3736
rect 9955 3587 9992 3639
rect 10116 3646 10177 3672
rect 10266 3655 10372 3668
rect 9955 3553 9957 3587
rect 9991 3553 9992 3587
rect 9787 3383 9821 3391
rect 9955 3383 9992 3553
rect 10026 3581 10082 3597
rect 10026 3547 10048 3581
rect 10026 3519 10082 3547
rect 10026 3485 10048 3519
rect 10026 3407 10082 3485
rect 10116 3425 10150 3646
rect 10266 3621 10298 3655
rect 10332 3629 10372 3655
rect 10184 3587 10232 3608
rect 10184 3553 10195 3587
rect 10229 3553 10232 3587
rect 10184 3551 10232 3553
rect 10184 3517 10191 3551
rect 10225 3517 10232 3551
rect 10184 3489 10232 3517
rect 10266 3455 10300 3621
rect 10334 3595 10372 3629
rect 10406 3579 10440 3702
rect 10474 3681 10508 3715
rect 10474 3631 10508 3647
rect 10542 3741 10592 3757
rect 10542 3707 10558 3741
rect 10850 3741 10913 3791
rect 10542 3691 10592 3707
rect 10637 3697 10653 3731
rect 10687 3697 10814 3731
rect 10406 3563 10508 3579
rect 10406 3561 10474 3563
rect 10116 3399 10161 3425
rect 10195 3421 10211 3455
rect 10245 3421 10300 3455
rect 10195 3411 10300 3421
rect 10334 3529 10474 3561
rect 10334 3527 10508 3529
rect 9787 3333 9821 3349
rect 9855 3323 9871 3357
rect 9905 3323 9921 3357
rect 9989 3349 9992 3383
rect 9955 3333 9992 3349
rect 10043 3357 10093 3373
rect 9855 3281 9921 3323
rect 10043 3323 10059 3357
rect 10127 3371 10161 3399
rect 10334 3371 10368 3527
rect 10474 3513 10508 3527
rect 10410 3477 10450 3483
rect 10542 3477 10576 3691
rect 10610 3655 10648 3657
rect 10610 3621 10612 3655
rect 10646 3621 10648 3655
rect 10610 3563 10648 3621
rect 10644 3529 10648 3563
rect 10610 3513 10648 3529
rect 10682 3629 10746 3663
rect 10682 3595 10712 3629
rect 10682 3587 10746 3595
rect 10682 3553 10699 3587
rect 10733 3553 10746 3587
rect 10410 3467 10576 3477
rect 10682 3471 10746 3553
rect 10444 3433 10576 3467
rect 10410 3417 10576 3433
rect 10127 3337 10144 3371
rect 10178 3337 10194 3371
rect 10233 3337 10255 3371
rect 10289 3337 10368 3371
rect 10432 3365 10506 3381
rect 10043 3281 10093 3323
rect 10432 3331 10454 3365
rect 10488 3331 10506 3365
rect 10542 3371 10576 3417
rect 10653 3455 10746 3471
rect 10687 3421 10746 3455
rect 10653 3405 10746 3421
rect 10780 3529 10814 3697
rect 10850 3707 10852 3741
rect 10886 3707 10913 3741
rect 10850 3691 10913 3707
rect 10959 3749 11027 3757
rect 10959 3715 10975 3749
rect 11009 3715 11027 3749
rect 10959 3678 11027 3715
rect 10959 3645 10975 3678
rect 10848 3644 10975 3645
rect 11009 3644 11027 3678
rect 10848 3629 11027 3644
rect 10882 3607 11027 3629
rect 10882 3595 10975 3607
rect 10848 3573 10975 3595
rect 11009 3573 11027 3607
rect 11061 3719 11095 3791
rect 11241 3749 11759 3791
rect 11061 3639 11095 3685
rect 11061 3589 11095 3605
rect 11129 3743 11195 3748
rect 11129 3709 11145 3743
rect 11179 3723 11195 3743
rect 11129 3689 11161 3709
rect 11129 3675 11195 3689
rect 11129 3641 11145 3675
rect 11179 3641 11195 3675
rect 11129 3607 11195 3641
rect 10848 3570 11027 3573
rect 10989 3529 11027 3570
rect 11129 3573 11145 3607
rect 11179 3579 11195 3607
rect 11241 3715 11259 3749
rect 11293 3715 11707 3749
rect 11741 3715 11759 3749
rect 11241 3647 11759 3715
rect 11241 3613 11259 3647
rect 11293 3613 11707 3647
rect 11741 3613 11759 3647
rect 11811 3741 11845 3757
rect 11811 3673 11845 3707
rect 11879 3725 11945 3791
rect 11879 3691 11895 3725
rect 11929 3691 11945 3725
rect 11979 3741 12016 3757
rect 12013 3707 12016 3741
rect 11979 3673 12016 3707
rect 12064 3749 12117 3791
rect 12064 3715 12083 3749
rect 12064 3699 12117 3715
rect 12151 3741 12201 3757
rect 12151 3707 12167 3741
rect 12498 3749 12532 3791
rect 11845 3655 11944 3657
rect 11845 3639 11902 3655
rect 11811 3623 11902 3639
rect 11179 3573 11207 3579
rect 11241 3573 11759 3613
rect 11898 3621 11902 3623
rect 11936 3621 11944 3655
rect 11129 3563 11207 3573
rect 11164 3553 11207 3563
rect 10780 3513 10955 3529
rect 10780 3479 10921 3513
rect 10780 3463 10955 3479
rect 10989 3513 11139 3529
rect 10989 3479 11105 3513
rect 10989 3463 11139 3479
rect 10780 3371 10814 3463
rect 10989 3429 11029 3463
rect 11173 3437 11207 3553
rect 11162 3429 11207 3437
rect 10963 3426 11029 3429
rect 10963 3392 10979 3426
rect 11013 3392 11029 3426
rect 11131 3428 11207 3429
rect 10542 3337 10573 3371
rect 10607 3337 10623 3371
rect 10657 3337 10676 3371
rect 10710 3337 10814 3371
rect 10869 3371 10911 3387
rect 10869 3337 10874 3371
rect 10908 3337 10911 3371
rect 10432 3281 10506 3331
rect 10869 3281 10911 3337
rect 10963 3358 11029 3392
rect 10963 3324 10979 3358
rect 11013 3324 11029 3358
rect 11063 3387 11097 3403
rect 11063 3281 11097 3353
rect 11131 3394 11147 3428
rect 11181 3412 11207 3428
rect 11241 3505 11319 3539
rect 11353 3505 11429 3539
rect 11463 3505 11483 3539
rect 11241 3435 11483 3505
rect 11517 3503 11759 3573
rect 11517 3469 11537 3503
rect 11571 3469 11647 3503
rect 11681 3469 11759 3503
rect 11794 3587 11864 3589
rect 11794 3553 11805 3587
rect 11839 3553 11864 3587
rect 11794 3513 11864 3553
rect 11794 3479 11808 3513
rect 11842 3479 11864 3513
rect 11794 3459 11864 3479
rect 11898 3528 11944 3621
rect 11898 3494 11910 3528
rect 11181 3394 11197 3412
rect 11131 3360 11197 3394
rect 11131 3326 11147 3360
rect 11181 3326 11197 3360
rect 11131 3325 11197 3326
rect 11241 3376 11759 3435
rect 11898 3425 11944 3494
rect 11241 3342 11259 3376
rect 11293 3342 11707 3376
rect 11741 3342 11759 3376
rect 11241 3281 11759 3342
rect 11811 3391 11944 3425
rect 12013 3639 12016 3673
rect 12151 3672 12201 3707
rect 12243 3702 12259 3736
rect 12293 3702 12464 3736
rect 11979 3587 12016 3639
rect 12140 3646 12201 3672
rect 12290 3655 12396 3668
rect 11979 3553 11981 3587
rect 12015 3553 12016 3587
rect 11811 3383 11845 3391
rect 11979 3383 12016 3553
rect 12050 3581 12106 3597
rect 12050 3547 12072 3581
rect 12050 3519 12106 3547
rect 12050 3485 12072 3519
rect 12050 3407 12106 3485
rect 12140 3425 12174 3646
rect 12290 3621 12322 3655
rect 12356 3629 12396 3655
rect 12208 3587 12256 3608
rect 12208 3553 12219 3587
rect 12253 3553 12256 3587
rect 12208 3551 12256 3553
rect 12208 3517 12215 3551
rect 12249 3517 12256 3551
rect 12208 3489 12256 3517
rect 12290 3455 12324 3621
rect 12358 3595 12396 3629
rect 12430 3579 12464 3702
rect 12498 3681 12532 3715
rect 12498 3631 12532 3647
rect 12566 3741 12616 3757
rect 12566 3707 12582 3741
rect 12874 3741 12937 3791
rect 12566 3691 12616 3707
rect 12661 3697 12677 3731
rect 12711 3697 12838 3731
rect 12430 3563 12532 3579
rect 12430 3561 12498 3563
rect 12140 3399 12185 3425
rect 12219 3421 12235 3455
rect 12269 3421 12324 3455
rect 12219 3411 12324 3421
rect 12358 3529 12498 3561
rect 12358 3527 12532 3529
rect 11811 3333 11845 3349
rect 11879 3323 11895 3357
rect 11929 3323 11945 3357
rect 12013 3349 12016 3383
rect 11979 3333 12016 3349
rect 12067 3357 12117 3373
rect 11879 3281 11945 3323
rect 12067 3323 12083 3357
rect 12151 3371 12185 3399
rect 12358 3371 12392 3527
rect 12498 3513 12532 3527
rect 12434 3477 12474 3483
rect 12566 3477 12600 3691
rect 12634 3655 12672 3657
rect 12634 3621 12636 3655
rect 12670 3621 12672 3655
rect 12634 3563 12672 3621
rect 12668 3529 12672 3563
rect 12634 3513 12672 3529
rect 12706 3629 12770 3663
rect 12706 3595 12736 3629
rect 12706 3587 12770 3595
rect 12706 3553 12723 3587
rect 12757 3553 12770 3587
rect 12434 3467 12600 3477
rect 12706 3471 12770 3553
rect 12468 3433 12600 3467
rect 12434 3417 12600 3433
rect 12151 3337 12168 3371
rect 12202 3337 12218 3371
rect 12257 3337 12279 3371
rect 12313 3337 12392 3371
rect 12456 3365 12530 3381
rect 12067 3281 12117 3323
rect 12456 3331 12478 3365
rect 12512 3331 12530 3365
rect 12566 3371 12600 3417
rect 12677 3455 12770 3471
rect 12711 3421 12770 3455
rect 12677 3405 12770 3421
rect 12804 3529 12838 3697
rect 12874 3707 12876 3741
rect 12910 3707 12937 3741
rect 12874 3691 12937 3707
rect 12983 3749 13051 3757
rect 12983 3715 12999 3749
rect 13033 3715 13051 3749
rect 12983 3678 13051 3715
rect 12983 3645 12999 3678
rect 12872 3644 12999 3645
rect 13033 3644 13051 3678
rect 12872 3629 13051 3644
rect 12906 3607 13051 3629
rect 12906 3595 12999 3607
rect 12872 3573 12999 3595
rect 13033 3573 13051 3607
rect 13085 3719 13119 3791
rect 13265 3749 13967 3791
rect 13085 3639 13119 3685
rect 13085 3589 13119 3605
rect 13153 3743 13219 3748
rect 13153 3709 13169 3743
rect 13203 3723 13219 3743
rect 13153 3689 13185 3709
rect 13153 3675 13219 3689
rect 13153 3641 13169 3675
rect 13203 3641 13219 3675
rect 13153 3607 13219 3641
rect 12872 3570 13051 3573
rect 13013 3529 13051 3570
rect 13153 3573 13169 3607
rect 13203 3579 13219 3607
rect 13265 3715 13283 3749
rect 13317 3715 13915 3749
rect 13949 3715 13967 3749
rect 13265 3647 13967 3715
rect 13265 3613 13283 3647
rect 13317 3613 13915 3647
rect 13949 3613 13967 3647
rect 13203 3573 13231 3579
rect 13265 3573 13967 3613
rect 13153 3563 13231 3573
rect 13188 3553 13231 3563
rect 12804 3513 12979 3529
rect 12804 3479 12945 3513
rect 12804 3463 12979 3479
rect 13013 3513 13163 3529
rect 13013 3479 13129 3513
rect 13013 3463 13163 3479
rect 12804 3371 12838 3463
rect 13013 3429 13053 3463
rect 13197 3437 13231 3553
rect 13186 3429 13231 3437
rect 12987 3426 13053 3429
rect 12987 3392 13003 3426
rect 13037 3392 13053 3426
rect 13155 3428 13231 3429
rect 12566 3337 12597 3371
rect 12631 3337 12647 3371
rect 12681 3337 12700 3371
rect 12734 3337 12838 3371
rect 12893 3371 12935 3387
rect 12893 3337 12898 3371
rect 12932 3337 12935 3371
rect 12456 3281 12530 3331
rect 12893 3281 12935 3337
rect 12987 3358 13053 3392
rect 12987 3324 13003 3358
rect 13037 3324 13053 3358
rect 13087 3387 13121 3403
rect 13087 3281 13121 3353
rect 13155 3394 13171 3428
rect 13205 3412 13231 3428
rect 13265 3505 13343 3539
rect 13377 3505 13442 3539
rect 13476 3505 13541 3539
rect 13575 3505 13595 3539
rect 13265 3435 13595 3505
rect 13629 3503 13967 3573
rect 14001 3720 14059 3791
rect 14001 3686 14013 3720
rect 14047 3686 14059 3720
rect 14093 3749 15162 3791
rect 14093 3715 14111 3749
rect 14145 3715 15111 3749
rect 15145 3715 15162 3749
rect 14093 3704 15162 3715
rect 15197 3749 15715 3791
rect 15197 3715 15215 3749
rect 15249 3715 15663 3749
rect 15697 3715 15715 3749
rect 14001 3627 14059 3686
rect 14001 3593 14013 3627
rect 14047 3593 14059 3627
rect 14001 3558 14059 3593
rect 13629 3469 13649 3503
rect 13683 3469 13752 3503
rect 13786 3469 13855 3503
rect 13889 3469 13967 3503
rect 14410 3539 14478 3556
rect 14410 3505 14427 3539
rect 14461 3505 14478 3539
rect 13205 3394 13221 3412
rect 13155 3360 13221 3394
rect 13155 3326 13171 3360
rect 13205 3326 13221 3360
rect 13155 3325 13221 3326
rect 13265 3376 13967 3435
rect 13265 3342 13283 3376
rect 13317 3342 13915 3376
rect 13949 3342 13967 3376
rect 13265 3281 13967 3342
rect 14001 3409 14059 3426
rect 14001 3375 14013 3409
rect 14047 3375 14059 3409
rect 14410 3390 14478 3505
rect 14774 3503 14844 3704
rect 15197 3647 15715 3715
rect 15197 3613 15215 3647
rect 15249 3613 15663 3647
rect 15697 3613 15715 3647
rect 15197 3573 15715 3613
rect 14774 3469 14791 3503
rect 14825 3469 14844 3503
rect 14774 3454 14844 3469
rect 15197 3505 15275 3539
rect 15309 3505 15385 3539
rect 15419 3505 15439 3539
rect 15197 3435 15439 3505
rect 15473 3503 15715 3573
rect 15473 3469 15493 3503
rect 15527 3469 15603 3503
rect 15637 3469 15715 3503
rect 15749 3741 15803 3757
rect 15749 3707 15767 3741
rect 15801 3707 15803 3741
rect 15749 3660 15803 3707
rect 15749 3626 15767 3660
rect 15801 3626 15803 3660
rect 15837 3741 15903 3791
rect 15837 3707 15853 3741
rect 15887 3707 15903 3741
rect 15837 3673 15903 3707
rect 15837 3639 15853 3673
rect 15887 3639 15903 3673
rect 15939 3741 15973 3757
rect 15939 3673 15973 3707
rect 15749 3576 15803 3626
rect 15939 3605 15973 3639
rect 14001 3281 14059 3375
rect 14093 3376 15162 3390
rect 14093 3342 14111 3376
rect 14145 3342 15111 3376
rect 15145 3342 15162 3376
rect 14093 3281 15162 3342
rect 15197 3376 15715 3435
rect 15197 3342 15215 3376
rect 15249 3342 15663 3376
rect 15697 3342 15715 3376
rect 15197 3281 15715 3342
rect 15749 3416 15783 3576
rect 15840 3571 15973 3605
rect 16025 3749 16359 3791
rect 16025 3715 16043 3749
rect 16077 3715 16307 3749
rect 16341 3715 16359 3749
rect 16025 3647 16359 3715
rect 16025 3613 16043 3647
rect 16077 3613 16307 3647
rect 16341 3613 16359 3647
rect 16025 3573 16359 3613
rect 15840 3542 15874 3571
rect 15817 3526 15874 3542
rect 15851 3492 15874 3526
rect 15817 3476 15874 3492
rect 15840 3425 15874 3476
rect 15921 3519 15987 3535
rect 15921 3513 15945 3519
rect 15921 3479 15937 3513
rect 15979 3485 15987 3519
rect 15971 3479 15987 3485
rect 15921 3461 15987 3479
rect 16025 3505 16045 3539
rect 16079 3505 16175 3539
rect 16025 3435 16175 3505
rect 16209 3503 16359 3573
rect 16209 3469 16305 3503
rect 16339 3469 16359 3503
rect 16393 3749 16485 3757
rect 16393 3715 16435 3749
rect 16469 3715 16485 3749
rect 16393 3681 16485 3715
rect 16393 3647 16435 3681
rect 16469 3647 16485 3681
rect 16523 3749 16589 3791
rect 16523 3715 16539 3749
rect 16573 3715 16589 3749
rect 16523 3681 16589 3715
rect 16523 3647 16539 3681
rect 16573 3647 16589 3681
rect 16629 3707 16689 3723
rect 16629 3673 16647 3707
rect 16681 3673 16689 3707
rect 16393 3519 16443 3647
rect 16629 3613 16689 3673
rect 16723 3707 16779 3791
rect 16723 3673 16731 3707
rect 16765 3673 16779 3707
rect 16723 3657 16779 3673
rect 16853 3749 17187 3791
rect 16853 3715 16871 3749
rect 16905 3715 17135 3749
rect 17169 3715 17187 3749
rect 16501 3579 16689 3613
rect 16853 3647 17187 3715
rect 16853 3613 16871 3647
rect 16905 3613 17135 3647
rect 17169 3613 17187 3647
rect 16501 3529 16535 3579
rect 16763 3529 16816 3601
rect 16853 3573 17187 3613
rect 16393 3485 16405 3519
rect 16439 3485 16443 3519
rect 15749 3387 15801 3416
rect 15840 3391 15973 3425
rect 15749 3383 15767 3387
rect 15749 3349 15761 3383
rect 15939 3370 15973 3391
rect 15795 3349 15801 3353
rect 15749 3315 15801 3349
rect 15837 3323 15853 3357
rect 15887 3323 15903 3357
rect 15837 3281 15903 3323
rect 15939 3315 15973 3336
rect 16025 3383 16359 3435
rect 16025 3349 16043 3383
rect 16077 3349 16307 3383
rect 16341 3349 16359 3383
rect 16025 3281 16359 3349
rect 16393 3373 16443 3485
rect 16477 3513 16535 3529
rect 16477 3479 16479 3513
rect 16513 3479 16535 3513
rect 16569 3519 16637 3529
rect 16569 3513 16589 3519
rect 16569 3479 16587 3513
rect 16623 3485 16637 3519
rect 16621 3479 16637 3485
rect 16681 3519 16816 3529
rect 16715 3513 16816 3519
rect 16715 3485 16728 3513
rect 16681 3479 16728 3485
rect 16762 3479 16816 3513
rect 16853 3505 16873 3539
rect 16907 3505 17003 3539
rect 16477 3463 16535 3479
rect 16501 3445 16535 3463
rect 16501 3407 16779 3445
rect 16713 3385 16779 3407
rect 16393 3357 16505 3373
rect 16393 3323 16455 3357
rect 16489 3323 16505 3357
rect 16393 3315 16505 3323
rect 16539 3357 16589 3373
rect 16573 3323 16589 3357
rect 16713 3351 16731 3385
rect 16765 3351 16779 3385
rect 16713 3335 16779 3351
rect 16853 3435 17003 3505
rect 17037 3503 17187 3573
rect 17037 3469 17133 3503
rect 17167 3469 17187 3503
rect 17221 3749 17313 3757
rect 17221 3715 17263 3749
rect 17297 3715 17313 3749
rect 17221 3681 17313 3715
rect 17221 3647 17263 3681
rect 17297 3647 17313 3681
rect 17351 3749 17417 3791
rect 17351 3715 17367 3749
rect 17401 3715 17417 3749
rect 17351 3681 17417 3715
rect 17351 3647 17367 3681
rect 17401 3647 17417 3681
rect 17457 3707 17517 3723
rect 17457 3673 17475 3707
rect 17509 3673 17517 3707
rect 16853 3383 17187 3435
rect 16853 3349 16871 3383
rect 16905 3349 17135 3383
rect 17169 3349 17187 3383
rect 16539 3281 16589 3323
rect 16853 3281 17187 3349
rect 17221 3383 17271 3647
rect 17457 3613 17517 3673
rect 17551 3707 17607 3791
rect 17551 3673 17559 3707
rect 17593 3673 17607 3707
rect 17551 3657 17607 3673
rect 17681 3749 18383 3791
rect 17681 3715 17699 3749
rect 17733 3715 18331 3749
rect 18365 3715 18383 3749
rect 17329 3579 17517 3613
rect 17681 3647 18383 3715
rect 17681 3613 17699 3647
rect 17733 3613 18331 3647
rect 18365 3613 18383 3647
rect 17591 3587 17644 3601
rect 17329 3529 17363 3579
rect 17591 3553 17601 3587
rect 17635 3553 17644 3587
rect 17681 3573 18383 3613
rect 17591 3529 17644 3553
rect 17305 3513 17363 3529
rect 17305 3479 17307 3513
rect 17341 3479 17363 3513
rect 17397 3519 17465 3529
rect 17397 3513 17417 3519
rect 17397 3479 17415 3513
rect 17451 3485 17465 3519
rect 17449 3479 17465 3485
rect 17509 3513 17644 3529
rect 17509 3479 17556 3513
rect 17590 3479 17644 3513
rect 17681 3505 17759 3539
rect 17793 3505 17858 3539
rect 17892 3505 17957 3539
rect 17991 3505 18011 3539
rect 17305 3463 17363 3479
rect 17329 3445 17363 3463
rect 17329 3407 17607 3445
rect 17221 3349 17233 3383
rect 17267 3373 17271 3383
rect 17541 3385 17607 3407
rect 17267 3357 17333 3373
rect 17267 3349 17283 3357
rect 17221 3323 17283 3349
rect 17317 3323 17333 3357
rect 17221 3315 17333 3323
rect 17367 3357 17417 3373
rect 17401 3323 17417 3357
rect 17541 3351 17559 3385
rect 17593 3351 17607 3385
rect 17541 3335 17607 3351
rect 17681 3435 18011 3505
rect 18045 3503 18383 3573
rect 18045 3469 18065 3503
rect 18099 3469 18168 3503
rect 18202 3469 18271 3503
rect 18305 3469 18383 3503
rect 18601 3749 18843 3791
rect 18601 3715 18619 3749
rect 18653 3715 18791 3749
rect 18825 3715 18843 3749
rect 18601 3654 18843 3715
rect 18601 3620 18619 3654
rect 18653 3620 18791 3654
rect 18825 3620 18843 3654
rect 18601 3573 18843 3620
rect 18601 3499 18705 3573
rect 18601 3465 18651 3499
rect 18685 3465 18705 3499
rect 18739 3505 18759 3539
rect 18793 3505 18843 3539
rect 17681 3376 18383 3435
rect 18739 3431 18843 3505
rect 17681 3342 17699 3376
rect 17733 3342 18331 3376
rect 18365 3342 18383 3376
rect 17367 3281 17417 3323
rect 17681 3281 18383 3342
rect 18601 3378 18843 3431
rect 18601 3344 18619 3378
rect 18653 3344 18791 3378
rect 18825 3344 18843 3378
rect 18601 3281 18843 3344
rect 1104 3247 1133 3281
rect 1167 3247 1225 3281
rect 1259 3247 1317 3281
rect 1351 3247 1409 3281
rect 1443 3247 1501 3281
rect 1535 3247 1593 3281
rect 1627 3247 1685 3281
rect 1719 3247 1777 3281
rect 1811 3247 1869 3281
rect 1903 3247 1961 3281
rect 1995 3247 2053 3281
rect 2087 3247 2145 3281
rect 2179 3247 2237 3281
rect 2271 3247 2329 3281
rect 2363 3247 2421 3281
rect 2455 3247 2513 3281
rect 2547 3247 2605 3281
rect 2639 3247 2697 3281
rect 2731 3247 2789 3281
rect 2823 3247 2881 3281
rect 2915 3247 2973 3281
rect 3007 3247 3065 3281
rect 3099 3247 3157 3281
rect 3191 3247 3249 3281
rect 3283 3247 3341 3281
rect 3375 3247 3433 3281
rect 3467 3247 3525 3281
rect 3559 3247 3617 3281
rect 3651 3247 3709 3281
rect 3743 3247 3801 3281
rect 3835 3247 3893 3281
rect 3927 3247 3985 3281
rect 4019 3247 4077 3281
rect 4111 3247 4169 3281
rect 4203 3247 4261 3281
rect 4295 3247 4353 3281
rect 4387 3247 4445 3281
rect 4479 3247 4537 3281
rect 4571 3247 4629 3281
rect 4663 3247 4721 3281
rect 4755 3247 4813 3281
rect 4847 3247 4905 3281
rect 4939 3247 4997 3281
rect 5031 3247 5089 3281
rect 5123 3247 5181 3281
rect 5215 3247 5273 3281
rect 5307 3247 5365 3281
rect 5399 3247 5457 3281
rect 5491 3247 5549 3281
rect 5583 3247 5641 3281
rect 5675 3247 5733 3281
rect 5767 3247 5825 3281
rect 5859 3247 5917 3281
rect 5951 3247 6009 3281
rect 6043 3247 6101 3281
rect 6135 3247 6193 3281
rect 6227 3247 6285 3281
rect 6319 3247 6377 3281
rect 6411 3247 6469 3281
rect 6503 3247 6561 3281
rect 6595 3247 6653 3281
rect 6687 3247 6745 3281
rect 6779 3247 6837 3281
rect 6871 3247 6929 3281
rect 6963 3247 7021 3281
rect 7055 3247 7113 3281
rect 7147 3247 7205 3281
rect 7239 3247 7297 3281
rect 7331 3247 7389 3281
rect 7423 3247 7481 3281
rect 7515 3247 7573 3281
rect 7607 3247 7665 3281
rect 7699 3247 7757 3281
rect 7791 3247 7849 3281
rect 7883 3247 7941 3281
rect 7975 3247 8033 3281
rect 8067 3247 8125 3281
rect 8159 3247 8217 3281
rect 8251 3247 8309 3281
rect 8343 3247 8401 3281
rect 8435 3247 8493 3281
rect 8527 3247 8585 3281
rect 8619 3247 8677 3281
rect 8711 3247 8769 3281
rect 8803 3247 8861 3281
rect 8895 3247 8953 3281
rect 8987 3247 9045 3281
rect 9079 3247 9137 3281
rect 9171 3247 9229 3281
rect 9263 3247 9321 3281
rect 9355 3247 9413 3281
rect 9447 3247 9505 3281
rect 9539 3247 9597 3281
rect 9631 3247 9689 3281
rect 9723 3247 9781 3281
rect 9815 3247 9873 3281
rect 9907 3247 9965 3281
rect 9999 3247 10057 3281
rect 10091 3247 10149 3281
rect 10183 3247 10241 3281
rect 10275 3247 10333 3281
rect 10367 3247 10425 3281
rect 10459 3247 10517 3281
rect 10551 3247 10609 3281
rect 10643 3247 10701 3281
rect 10735 3247 10793 3281
rect 10827 3247 10885 3281
rect 10919 3247 10977 3281
rect 11011 3247 11069 3281
rect 11103 3247 11161 3281
rect 11195 3247 11253 3281
rect 11287 3247 11345 3281
rect 11379 3247 11437 3281
rect 11471 3247 11529 3281
rect 11563 3247 11621 3281
rect 11655 3247 11713 3281
rect 11747 3247 11805 3281
rect 11839 3247 11897 3281
rect 11931 3247 11989 3281
rect 12023 3247 12081 3281
rect 12115 3247 12173 3281
rect 12207 3247 12265 3281
rect 12299 3247 12357 3281
rect 12391 3247 12449 3281
rect 12483 3247 12541 3281
rect 12575 3247 12633 3281
rect 12667 3247 12725 3281
rect 12759 3247 12817 3281
rect 12851 3247 12909 3281
rect 12943 3247 13001 3281
rect 13035 3247 13093 3281
rect 13127 3247 13185 3281
rect 13219 3247 13277 3281
rect 13311 3247 13369 3281
rect 13403 3247 13461 3281
rect 13495 3247 13553 3281
rect 13587 3247 13645 3281
rect 13679 3247 13737 3281
rect 13771 3247 13829 3281
rect 13863 3247 13921 3281
rect 13955 3247 14013 3281
rect 14047 3247 14105 3281
rect 14139 3247 14197 3281
rect 14231 3247 14289 3281
rect 14323 3247 14381 3281
rect 14415 3247 14473 3281
rect 14507 3247 14565 3281
rect 14599 3247 14657 3281
rect 14691 3247 14749 3281
rect 14783 3247 14841 3281
rect 14875 3247 14933 3281
rect 14967 3247 15025 3281
rect 15059 3247 15117 3281
rect 15151 3247 15209 3281
rect 15243 3247 15301 3281
rect 15335 3247 15393 3281
rect 15427 3247 15485 3281
rect 15519 3247 15577 3281
rect 15611 3247 15669 3281
rect 15703 3247 15761 3281
rect 15795 3247 15853 3281
rect 15887 3247 15945 3281
rect 15979 3247 16037 3281
rect 16071 3247 16129 3281
rect 16163 3247 16221 3281
rect 16255 3247 16313 3281
rect 16347 3247 16405 3281
rect 16439 3247 16497 3281
rect 16531 3247 16589 3281
rect 16623 3247 16681 3281
rect 16715 3247 16773 3281
rect 16807 3247 16865 3281
rect 16899 3247 16957 3281
rect 16991 3247 17049 3281
rect 17083 3247 17141 3281
rect 17175 3247 17233 3281
rect 17267 3247 17325 3281
rect 17359 3247 17417 3281
rect 17451 3247 17509 3281
rect 17543 3247 17601 3281
rect 17635 3247 17693 3281
rect 17727 3247 17785 3281
rect 17819 3247 17877 3281
rect 17911 3247 17969 3281
rect 18003 3247 18061 3281
rect 18095 3247 18153 3281
rect 18187 3247 18245 3281
rect 18279 3247 18337 3281
rect 18371 3247 18429 3281
rect 18463 3247 18521 3281
rect 18555 3247 18613 3281
rect 18647 3247 18705 3281
rect 18739 3247 18797 3281
rect 18831 3247 18860 3281
rect 1121 3184 1363 3247
rect 1121 3150 1139 3184
rect 1173 3150 1311 3184
rect 1345 3150 1363 3184
rect 1121 3097 1363 3150
rect 1397 3179 1731 3247
rect 1397 3145 1415 3179
rect 1449 3145 1679 3179
rect 1713 3145 1731 3179
rect 1121 3023 1225 3097
rect 1397 3093 1731 3145
rect 1857 3197 1909 3213
rect 1857 3163 1875 3197
rect 1857 3147 1909 3163
rect 1951 3201 2006 3247
rect 1951 3167 1961 3201
rect 1995 3167 2006 3201
rect 1951 3151 2006 3167
rect 2048 3197 2089 3213
rect 2048 3163 2055 3197
rect 2123 3201 2190 3247
rect 2123 3167 2139 3201
rect 2173 3167 2190 3201
rect 2225 3179 2559 3247
rect 1121 2989 1171 3023
rect 1205 2989 1225 3023
rect 1259 3029 1279 3063
rect 1313 3029 1363 3063
rect 1259 2955 1363 3029
rect 1397 3023 1547 3093
rect 1397 2989 1417 3023
rect 1451 2989 1547 3023
rect 1581 3025 1677 3059
rect 1711 3025 1731 3059
rect 1581 2955 1731 3025
rect 1121 2908 1363 2955
rect 1121 2874 1139 2908
rect 1173 2874 1311 2908
rect 1345 2874 1363 2908
rect 1121 2813 1363 2874
rect 1121 2779 1139 2813
rect 1173 2779 1311 2813
rect 1345 2779 1363 2813
rect 1121 2737 1363 2779
rect 1397 2915 1731 2955
rect 1397 2881 1415 2915
rect 1449 2881 1679 2915
rect 1713 2881 1731 2915
rect 1397 2813 1731 2881
rect 1397 2779 1415 2813
rect 1449 2779 1679 2813
rect 1713 2779 1731 2813
rect 1397 2737 1731 2779
rect 1857 2965 1891 3147
rect 2048 3133 2089 3163
rect 2225 3145 2243 3179
rect 2277 3145 2507 3179
rect 2541 3145 2559 3179
rect 2611 3201 2671 3247
rect 2611 3167 2628 3201
rect 2662 3167 2671 3201
rect 2611 3151 2671 3167
rect 2705 3192 2757 3208
rect 2705 3158 2714 3192
rect 2748 3158 2757 3192
rect 1925 3049 1997 3115
rect 2048 3111 2185 3133
rect 2048 3099 2145 3111
rect 2117 3077 2145 3099
rect 2179 3077 2185 3111
rect 1925 3015 1929 3049
rect 1963 3043 1997 3049
rect 1925 3009 1961 3015
rect 1995 3009 1997 3043
rect 1925 2999 1997 3009
rect 2033 3049 2083 3065
rect 2067 3015 2083 3049
rect 2033 2965 2083 3015
rect 1857 2932 2083 2965
rect 1857 2898 1875 2932
rect 1909 2931 2083 2932
rect 1909 2898 1911 2931
rect 1857 2827 1911 2898
rect 2117 2893 2185 3077
rect 2225 3093 2559 3145
rect 2705 3117 2757 3158
rect 2791 3201 2843 3247
rect 2791 3167 2800 3201
rect 2834 3167 2843 3201
rect 2791 3151 2843 3167
rect 2879 3192 2931 3208
rect 2879 3158 2886 3192
rect 2920 3158 2931 3192
rect 2879 3117 2931 3158
rect 2965 3201 3015 3247
rect 2965 3167 2972 3201
rect 3006 3167 3015 3201
rect 2965 3151 3015 3167
rect 3051 3192 3103 3208
rect 3051 3158 3058 3192
rect 3092 3179 3103 3192
rect 3051 3145 3065 3158
rect 3099 3145 3103 3179
rect 3137 3201 3187 3247
rect 3137 3167 3144 3201
rect 3178 3167 3187 3201
rect 3137 3151 3187 3167
rect 3223 3192 3275 3208
rect 3223 3158 3230 3192
rect 3264 3158 3275 3192
rect 3051 3117 3103 3145
rect 3223 3117 3275 3158
rect 3309 3201 3358 3247
rect 3309 3167 3315 3201
rect 3349 3167 3358 3201
rect 3309 3151 3358 3167
rect 3392 3192 3447 3208
rect 3392 3158 3401 3192
rect 3435 3158 3447 3192
rect 3392 3117 3447 3158
rect 3481 3201 3530 3247
rect 3481 3167 3487 3201
rect 3521 3167 3530 3201
rect 3481 3151 3530 3167
rect 3564 3192 3616 3208
rect 3564 3158 3573 3192
rect 3607 3158 3616 3192
rect 3564 3117 3616 3158
rect 3650 3201 3702 3247
rect 3650 3167 3659 3201
rect 3693 3167 3702 3201
rect 3650 3151 3702 3167
rect 3736 3192 3788 3208
rect 3736 3158 3745 3192
rect 3779 3158 3788 3192
rect 3736 3117 3788 3158
rect 3822 3201 3874 3247
rect 3822 3167 3831 3201
rect 3865 3167 3874 3201
rect 3822 3151 3874 3167
rect 3908 3192 3960 3208
rect 3908 3158 3917 3192
rect 3951 3158 3960 3192
rect 3908 3117 3960 3158
rect 3994 3192 4046 3247
rect 3994 3158 4003 3192
rect 4037 3158 4046 3192
rect 3994 3135 4046 3158
rect 4080 3192 4130 3211
rect 4080 3158 4089 3192
rect 4123 3158 4130 3192
rect 2225 3023 2375 3093
rect 2611 3083 3960 3117
rect 2225 2989 2245 3023
rect 2279 2989 2375 3023
rect 2409 3025 2505 3059
rect 2539 3025 2559 3059
rect 2409 2955 2559 3025
rect 1857 2793 1875 2827
rect 1909 2793 1911 2827
rect 1857 2777 1911 2793
rect 1945 2859 1961 2893
rect 1995 2859 2011 2893
rect 1945 2825 2011 2859
rect 1945 2791 1961 2825
rect 1995 2791 2011 2825
rect 1945 2737 2011 2791
rect 2052 2858 2185 2893
rect 2225 2915 2559 2955
rect 2611 2965 2844 3083
rect 4080 3049 4130 3158
rect 4166 3192 4218 3247
rect 4166 3158 4175 3192
rect 4209 3158 4218 3192
rect 4166 3142 4218 3158
rect 4252 3192 4302 3211
rect 4252 3158 4261 3192
rect 4295 3158 4302 3192
rect 4252 3049 4302 3158
rect 4338 3205 4399 3247
rect 4338 3171 4347 3205
rect 4381 3171 4399 3205
rect 4338 3145 4399 3171
rect 4433 3186 5502 3247
rect 4433 3152 4451 3186
rect 4485 3152 5451 3186
rect 5485 3152 5502 3186
rect 4433 3138 5502 3152
rect 5537 3186 6239 3247
rect 5537 3152 5555 3186
rect 5589 3152 6187 3186
rect 6221 3152 6239 3186
rect 2878 3015 2898 3049
rect 2932 3015 2966 3049
rect 3000 3015 3034 3049
rect 3068 3015 3102 3049
rect 3136 3015 3170 3049
rect 3204 3015 3238 3049
rect 3272 3015 3306 3049
rect 3340 3015 3374 3049
rect 3408 3015 3442 3049
rect 3476 3015 3510 3049
rect 3544 3015 3578 3049
rect 3612 3015 3646 3049
rect 3680 3015 3714 3049
rect 3748 3015 3782 3049
rect 3816 3015 3850 3049
rect 3884 3015 3918 3049
rect 3952 3015 4302 3049
rect 2878 2999 4302 3015
rect 4336 3077 4353 3111
rect 4387 3077 4399 3111
rect 4336 3049 4399 3077
rect 4336 3015 4345 3049
rect 4379 3015 4399 3049
rect 4336 2999 4399 3015
rect 4750 3023 4818 3138
rect 5537 3093 6239 3152
rect 6273 3153 6331 3247
rect 6273 3119 6285 3153
rect 6319 3119 6331 3153
rect 6273 3102 6331 3119
rect 6365 3186 7067 3247
rect 6365 3152 6383 3186
rect 6417 3152 7015 3186
rect 7049 3152 7067 3186
rect 6365 3093 7067 3152
rect 7193 3207 7343 3213
rect 7193 3173 7211 3207
rect 7245 3173 7286 3207
rect 7320 3173 7343 3207
rect 7193 3139 7343 3173
rect 7193 3105 7211 3139
rect 7245 3105 7286 3139
rect 7320 3105 7343 3139
rect 2611 2943 3960 2965
rect 2611 2920 2714 2943
rect 2225 2881 2243 2915
rect 2277 2881 2507 2915
rect 2541 2881 2559 2915
rect 2699 2909 2714 2920
rect 2748 2920 2886 2943
rect 2748 2909 2757 2920
rect 2052 2827 2089 2858
rect 2052 2793 2055 2827
rect 2052 2777 2089 2793
rect 2123 2788 2139 2822
rect 2173 2788 2190 2822
rect 2123 2737 2190 2788
rect 2225 2813 2559 2881
rect 2225 2779 2243 2813
rect 2277 2779 2507 2813
rect 2541 2779 2559 2813
rect 2225 2737 2559 2779
rect 2611 2837 2665 2886
rect 2611 2803 2628 2837
rect 2662 2803 2665 2837
rect 2611 2737 2665 2803
rect 2699 2857 2757 2909
rect 2879 2909 2886 2920
rect 2920 2917 3058 2943
rect 2920 2909 2931 2917
rect 2699 2823 2714 2857
rect 2748 2823 2757 2857
rect 2699 2772 2757 2823
rect 2791 2837 2842 2883
rect 2791 2803 2800 2837
rect 2834 2803 2842 2837
rect 2791 2738 2842 2803
rect 2879 2857 2931 2909
rect 3051 2909 3058 2917
rect 3092 2917 3230 2943
rect 3092 2909 3103 2917
rect 2879 2823 2886 2857
rect 2920 2823 2931 2857
rect 2879 2772 2931 2823
rect 2965 2837 3014 2883
rect 2965 2803 2972 2837
rect 3006 2803 3014 2837
rect 2965 2738 3014 2803
rect 3051 2857 3103 2909
rect 3223 2909 3230 2917
rect 3264 2917 3401 2943
rect 3264 2909 3275 2917
rect 3051 2823 3058 2857
rect 3092 2823 3103 2857
rect 3051 2772 3103 2823
rect 3137 2837 3186 2883
rect 3137 2803 3144 2837
rect 3178 2803 3186 2837
rect 3137 2738 3186 2803
rect 3223 2857 3275 2909
rect 3392 2909 3401 2917
rect 3435 2917 3573 2943
rect 3435 2909 3444 2917
rect 3223 2823 3230 2857
rect 3264 2823 3275 2857
rect 3223 2772 3275 2823
rect 3309 2837 3358 2883
rect 3309 2803 3315 2837
rect 3349 2803 3358 2837
rect 3309 2738 3358 2803
rect 3392 2857 3444 2909
rect 3564 2909 3573 2917
rect 3607 2917 3745 2943
rect 3607 2909 3616 2917
rect 3392 2823 3401 2857
rect 3435 2823 3444 2857
rect 3392 2772 3444 2823
rect 3478 2837 3530 2883
rect 3478 2803 3487 2837
rect 3521 2803 3530 2837
rect 3478 2738 3530 2803
rect 3564 2857 3616 2909
rect 3736 2909 3745 2917
rect 3779 2917 3917 2943
rect 3779 2909 3788 2917
rect 3564 2823 3573 2857
rect 3607 2823 3616 2857
rect 3564 2772 3616 2823
rect 3650 2837 3702 2883
rect 3650 2803 3659 2837
rect 3693 2803 3702 2837
rect 3650 2738 3702 2803
rect 3736 2857 3788 2909
rect 3908 2909 3917 2917
rect 3951 2909 3960 2943
rect 3736 2823 3745 2857
rect 3779 2823 3788 2857
rect 3736 2772 3788 2823
rect 3822 2837 3874 2883
rect 3822 2803 3831 2837
rect 3865 2803 3874 2837
rect 3822 2738 3874 2803
rect 3908 2857 3960 2909
rect 4080 2897 4130 2999
rect 3908 2823 3917 2857
rect 3951 2823 3960 2857
rect 3908 2772 3960 2823
rect 3994 2881 4046 2897
rect 3994 2847 4003 2881
rect 4037 2847 4046 2881
rect 3994 2813 4046 2847
rect 3994 2779 4003 2813
rect 4037 2779 4046 2813
rect 3994 2738 4046 2779
rect 4080 2863 4089 2897
rect 4123 2863 4130 2897
rect 4080 2829 4130 2863
rect 4080 2795 4089 2829
rect 4123 2795 4130 2829
rect 4080 2772 4130 2795
rect 4166 2881 4218 2899
rect 4166 2847 4175 2881
rect 4209 2847 4218 2881
rect 4166 2813 4218 2847
rect 4166 2779 4175 2813
rect 4209 2779 4218 2813
rect 2791 2737 4046 2738
rect 4166 2737 4218 2779
rect 4253 2889 4302 2999
rect 4750 2989 4767 3023
rect 4801 2989 4818 3023
rect 4750 2972 4818 2989
rect 5114 3059 5184 3074
rect 5114 3025 5131 3059
rect 5165 3025 5184 3059
rect 4253 2855 4261 2889
rect 4295 2855 4302 2889
rect 4253 2821 4302 2855
rect 4253 2787 4261 2821
rect 4295 2787 4302 2821
rect 4253 2771 4302 2787
rect 4338 2881 4397 2899
rect 4338 2847 4347 2881
rect 4381 2847 4397 2881
rect 4338 2813 4397 2847
rect 5114 2824 5184 3025
rect 5537 3023 5867 3093
rect 5537 2989 5615 3023
rect 5649 2989 5714 3023
rect 5748 2989 5813 3023
rect 5847 2989 5867 3023
rect 5901 3025 5921 3059
rect 5955 3025 6024 3059
rect 6058 3025 6127 3059
rect 6161 3025 6239 3059
rect 5901 2955 6239 3025
rect 6365 3023 6695 3093
rect 6365 2989 6443 3023
rect 6477 2989 6542 3023
rect 6576 2989 6641 3023
rect 6675 2989 6695 3023
rect 6729 3025 6749 3059
rect 6783 3025 6852 3059
rect 6886 3025 6955 3059
rect 6989 3025 7067 3059
rect 5537 2915 6239 2955
rect 5537 2881 5555 2915
rect 5589 2881 6187 2915
rect 6221 2881 6239 2915
rect 4338 2779 4347 2813
rect 4381 2779 4397 2813
rect 4338 2737 4397 2779
rect 4433 2813 5502 2824
rect 4433 2779 4451 2813
rect 4485 2779 5451 2813
rect 5485 2779 5502 2813
rect 4433 2737 5502 2779
rect 5537 2813 6239 2881
rect 5537 2779 5555 2813
rect 5589 2779 6187 2813
rect 6221 2779 6239 2813
rect 5537 2737 6239 2779
rect 6273 2935 6331 2970
rect 6729 2955 7067 3025
rect 6273 2901 6285 2935
rect 6319 2901 6331 2935
rect 6273 2842 6331 2901
rect 6273 2808 6285 2842
rect 6319 2808 6331 2842
rect 6273 2737 6331 2808
rect 6365 2915 7067 2955
rect 6365 2881 6383 2915
rect 6417 2881 7015 2915
rect 7049 2881 7067 2915
rect 6365 2813 7067 2881
rect 6365 2779 6383 2813
rect 6417 2779 7015 2813
rect 7049 2779 7067 2813
rect 6365 2737 7067 2779
rect 7193 3043 7343 3105
rect 7193 3009 7297 3043
rect 7331 3009 7343 3043
rect 7193 2771 7343 3009
rect 7377 3179 7711 3247
rect 7377 3145 7395 3179
rect 7429 3145 7659 3179
rect 7693 3145 7711 3179
rect 7745 3205 7806 3247
rect 7745 3171 7763 3205
rect 7797 3171 7806 3205
rect 7745 3145 7806 3171
rect 7842 3192 7892 3211
rect 7842 3158 7849 3192
rect 7883 3158 7892 3192
rect 7377 3093 7711 3145
rect 7377 3023 7527 3093
rect 7377 2989 7397 3023
rect 7431 2989 7527 3023
rect 7561 3025 7657 3059
rect 7691 3025 7711 3059
rect 7561 2955 7711 3025
rect 7745 3049 7808 3111
rect 7745 3043 7765 3049
rect 7745 3009 7757 3043
rect 7799 3015 7808 3049
rect 7791 3009 7808 3015
rect 7745 2999 7808 3009
rect 7842 3049 7892 3158
rect 7926 3192 7978 3247
rect 7926 3158 7935 3192
rect 7969 3158 7978 3192
rect 7926 3142 7978 3158
rect 8014 3192 8064 3211
rect 8014 3158 8021 3192
rect 8055 3158 8064 3192
rect 8014 3049 8064 3158
rect 8098 3192 8150 3247
rect 8098 3158 8107 3192
rect 8141 3158 8150 3192
rect 8098 3135 8150 3158
rect 8184 3192 8236 3208
rect 8184 3158 8193 3192
rect 8227 3158 8236 3192
rect 8184 3117 8236 3158
rect 8270 3201 8322 3247
rect 8270 3167 8279 3201
rect 8313 3167 8322 3201
rect 8270 3151 8322 3167
rect 8356 3192 8408 3208
rect 8356 3158 8365 3192
rect 8399 3158 8408 3192
rect 8356 3117 8408 3158
rect 8442 3201 8494 3247
rect 8442 3167 8451 3201
rect 8485 3167 8494 3201
rect 8442 3151 8494 3167
rect 8528 3192 8580 3208
rect 8528 3158 8537 3192
rect 8571 3158 8580 3192
rect 8528 3117 8580 3158
rect 8614 3201 8663 3247
rect 8614 3167 8623 3201
rect 8657 3167 8663 3201
rect 8614 3151 8663 3167
rect 8697 3192 8752 3208
rect 8697 3158 8709 3192
rect 8743 3158 8752 3192
rect 8697 3117 8752 3158
rect 8786 3201 8835 3247
rect 8786 3167 8795 3201
rect 8829 3167 8835 3201
rect 8786 3151 8835 3167
rect 8869 3192 8921 3208
rect 8869 3158 8880 3192
rect 8914 3158 8921 3192
rect 8869 3117 8921 3158
rect 8957 3201 9007 3247
rect 8957 3167 8966 3201
rect 9000 3167 9007 3201
rect 8957 3151 9007 3167
rect 9041 3192 9093 3208
rect 9041 3179 9052 3192
rect 9041 3145 9045 3179
rect 9086 3158 9093 3192
rect 9079 3145 9093 3158
rect 9129 3201 9179 3247
rect 9129 3167 9138 3201
rect 9172 3167 9179 3201
rect 9129 3151 9179 3167
rect 9213 3192 9265 3208
rect 9213 3158 9224 3192
rect 9258 3158 9265 3192
rect 9041 3117 9093 3145
rect 9213 3117 9265 3158
rect 9301 3201 9353 3247
rect 9301 3167 9310 3201
rect 9344 3167 9353 3201
rect 9301 3151 9353 3167
rect 9387 3192 9439 3208
rect 9387 3158 9396 3192
rect 9430 3158 9439 3192
rect 9387 3117 9439 3158
rect 9473 3201 9533 3247
rect 9473 3167 9482 3201
rect 9516 3167 9533 3201
rect 9473 3151 9533 3167
rect 9585 3186 10654 3247
rect 9585 3152 9603 3186
rect 9637 3152 10603 3186
rect 10637 3152 10654 3186
rect 9585 3138 10654 3152
rect 10689 3186 11391 3247
rect 10689 3152 10707 3186
rect 10741 3152 11339 3186
rect 11373 3152 11391 3186
rect 8184 3083 9533 3117
rect 7842 3015 8192 3049
rect 8226 3015 8260 3049
rect 8294 3015 8328 3049
rect 8362 3015 8396 3049
rect 8430 3015 8464 3049
rect 8498 3015 8532 3049
rect 8566 3015 8600 3049
rect 8634 3015 8668 3049
rect 8702 3015 8736 3049
rect 8770 3015 8804 3049
rect 8838 3015 8872 3049
rect 8906 3015 8940 3049
rect 8974 3015 9008 3049
rect 9042 3015 9076 3049
rect 9110 3015 9144 3049
rect 9178 3015 9212 3049
rect 9246 3015 9266 3049
rect 7842 2999 9266 3015
rect 7377 2915 7711 2955
rect 7377 2881 7395 2915
rect 7429 2881 7659 2915
rect 7693 2881 7711 2915
rect 7377 2813 7711 2881
rect 7377 2779 7395 2813
rect 7429 2779 7659 2813
rect 7693 2779 7711 2813
rect 7377 2737 7711 2779
rect 7747 2881 7806 2899
rect 7747 2847 7763 2881
rect 7797 2847 7806 2881
rect 7747 2813 7806 2847
rect 7747 2779 7763 2813
rect 7797 2779 7806 2813
rect 7747 2737 7806 2779
rect 7842 2889 7891 2999
rect 7842 2855 7849 2889
rect 7883 2855 7891 2889
rect 7842 2821 7891 2855
rect 7842 2787 7849 2821
rect 7883 2787 7891 2821
rect 7842 2771 7891 2787
rect 7926 2881 7978 2899
rect 7926 2847 7935 2881
rect 7969 2847 7978 2881
rect 7926 2813 7978 2847
rect 7926 2779 7935 2813
rect 7969 2779 7978 2813
rect 7926 2737 7978 2779
rect 8014 2897 8064 2999
rect 9300 2965 9533 3083
rect 9902 3023 9970 3138
rect 10689 3093 11391 3152
rect 11425 3153 11483 3247
rect 11787 3205 11853 3247
rect 11425 3119 11437 3153
rect 11471 3119 11483 3153
rect 11425 3102 11483 3119
rect 11719 3179 11753 3195
rect 11787 3171 11803 3205
rect 11837 3171 11853 3205
rect 11975 3205 12025 3247
rect 11887 3179 11924 3195
rect 11719 3137 11753 3145
rect 11921 3145 11924 3179
rect 11975 3171 11991 3205
rect 12364 3197 12438 3247
rect 11975 3155 12025 3171
rect 12059 3157 12076 3191
rect 12110 3157 12126 3191
rect 12165 3157 12187 3191
rect 12221 3157 12300 3191
rect 11719 3103 11852 3137
rect 9902 2989 9919 3023
rect 9953 2989 9970 3023
rect 9902 2972 9970 2989
rect 10266 3059 10336 3074
rect 10266 3025 10283 3059
rect 10317 3025 10336 3059
rect 8184 2943 9533 2965
rect 8184 2909 8193 2943
rect 8227 2917 8365 2943
rect 8227 2909 8236 2917
rect 8014 2863 8021 2897
rect 8055 2863 8064 2897
rect 8014 2829 8064 2863
rect 8014 2795 8021 2829
rect 8055 2795 8064 2829
rect 8014 2772 8064 2795
rect 8098 2881 8150 2897
rect 8098 2847 8107 2881
rect 8141 2847 8150 2881
rect 8098 2813 8150 2847
rect 8098 2779 8107 2813
rect 8141 2779 8150 2813
rect 8098 2738 8150 2779
rect 8184 2857 8236 2909
rect 8356 2909 8365 2917
rect 8399 2917 8537 2943
rect 8399 2909 8408 2917
rect 8184 2823 8193 2857
rect 8227 2823 8236 2857
rect 8184 2772 8236 2823
rect 8270 2837 8322 2883
rect 8270 2803 8279 2837
rect 8313 2803 8322 2837
rect 8270 2738 8322 2803
rect 8356 2857 8408 2909
rect 8528 2909 8537 2917
rect 8571 2917 8709 2943
rect 8571 2909 8580 2917
rect 8356 2823 8365 2857
rect 8399 2823 8408 2857
rect 8356 2772 8408 2823
rect 8442 2837 8494 2883
rect 8442 2803 8451 2837
rect 8485 2803 8494 2837
rect 8442 2738 8494 2803
rect 8528 2857 8580 2909
rect 8700 2909 8709 2917
rect 8743 2917 8880 2943
rect 8743 2909 8752 2917
rect 8528 2823 8537 2857
rect 8571 2823 8580 2857
rect 8528 2772 8580 2823
rect 8614 2837 8666 2883
rect 8614 2803 8623 2837
rect 8657 2803 8666 2837
rect 8614 2738 8666 2803
rect 8700 2857 8752 2909
rect 8869 2909 8880 2917
rect 8914 2917 9052 2943
rect 8914 2909 8921 2917
rect 8700 2823 8709 2857
rect 8743 2823 8752 2857
rect 8700 2772 8752 2823
rect 8786 2837 8835 2883
rect 8786 2803 8795 2837
rect 8829 2803 8835 2837
rect 8786 2738 8835 2803
rect 8869 2857 8921 2909
rect 9041 2909 9052 2917
rect 9086 2917 9224 2943
rect 9086 2909 9093 2917
rect 8869 2823 8880 2857
rect 8914 2823 8921 2857
rect 8869 2772 8921 2823
rect 8958 2837 9007 2883
rect 8958 2803 8966 2837
rect 9000 2803 9007 2837
rect 8958 2738 9007 2803
rect 9041 2857 9093 2909
rect 9213 2909 9224 2917
rect 9258 2920 9396 2943
rect 9258 2909 9265 2920
rect 9041 2823 9052 2857
rect 9086 2823 9093 2857
rect 9041 2772 9093 2823
rect 9130 2837 9179 2883
rect 9130 2803 9138 2837
rect 9172 2803 9179 2837
rect 9130 2738 9179 2803
rect 9213 2857 9265 2909
rect 9387 2909 9396 2920
rect 9430 2920 9533 2943
rect 9430 2909 9445 2920
rect 9213 2823 9224 2857
rect 9258 2823 9265 2857
rect 9213 2772 9265 2823
rect 9302 2837 9353 2883
rect 9302 2803 9310 2837
rect 9344 2803 9353 2837
rect 9302 2738 9353 2803
rect 9387 2857 9445 2909
rect 9387 2823 9396 2857
rect 9430 2823 9445 2857
rect 9387 2772 9445 2823
rect 9479 2837 9533 2886
rect 9479 2803 9482 2837
rect 9516 2803 9533 2837
rect 10266 2824 10336 3025
rect 10689 3023 11019 3093
rect 10689 2989 10767 3023
rect 10801 2989 10866 3023
rect 10900 2989 10965 3023
rect 10999 2989 11019 3023
rect 11053 3025 11073 3059
rect 11107 3025 11176 3059
rect 11210 3025 11279 3059
rect 11313 3025 11391 3059
rect 11053 2955 11391 3025
rect 11702 3049 11772 3069
rect 11702 3043 11716 3049
rect 11702 3009 11713 3043
rect 11750 3015 11772 3049
rect 11747 3009 11772 3015
rect 10689 2915 11391 2955
rect 10689 2881 10707 2915
rect 10741 2881 11339 2915
rect 11373 2881 11391 2915
rect 8098 2737 9353 2738
rect 9479 2737 9533 2803
rect 9585 2813 10654 2824
rect 9585 2779 9603 2813
rect 9637 2779 10603 2813
rect 10637 2779 10654 2813
rect 9585 2737 10654 2779
rect 10689 2813 11391 2881
rect 10689 2779 10707 2813
rect 10741 2779 11339 2813
rect 11373 2779 11391 2813
rect 10689 2737 11391 2779
rect 11425 2935 11483 2970
rect 11702 2939 11772 3009
rect 11806 3034 11852 3103
rect 11806 3000 11818 3034
rect 11425 2901 11437 2935
rect 11471 2901 11483 2935
rect 11806 2907 11852 3000
rect 11806 2905 11810 2907
rect 11425 2842 11483 2901
rect 11425 2808 11437 2842
rect 11471 2808 11483 2842
rect 11425 2737 11483 2808
rect 11719 2889 11810 2905
rect 11753 2873 11810 2889
rect 11844 2873 11852 2907
rect 11753 2871 11852 2873
rect 11887 2975 11924 3145
rect 12059 3129 12093 3157
rect 11887 2941 11889 2975
rect 11923 2941 11924 2975
rect 11887 2889 11924 2941
rect 11958 3111 12014 3121
rect 11992 3077 12014 3111
rect 11958 2981 12014 3077
rect 11958 2947 11980 2981
rect 11958 2931 12014 2947
rect 12048 3103 12093 3129
rect 12127 3107 12232 3117
rect 11719 2821 11753 2855
rect 11921 2855 11924 2889
rect 12048 2882 12082 3103
rect 12127 3073 12143 3107
rect 12177 3073 12232 3107
rect 12116 3011 12164 3039
rect 12116 2977 12123 3011
rect 12157 2977 12164 3011
rect 12116 2975 12164 2977
rect 12116 2941 12127 2975
rect 12161 2941 12164 2975
rect 12116 2920 12164 2941
rect 12198 2907 12232 3073
rect 12266 3001 12300 3157
rect 12364 3163 12386 3197
rect 12420 3163 12438 3197
rect 12801 3191 12843 3247
rect 12364 3147 12438 3163
rect 12474 3157 12505 3191
rect 12539 3157 12555 3191
rect 12589 3157 12608 3191
rect 12642 3157 12746 3191
rect 12474 3111 12508 3157
rect 12342 3095 12508 3111
rect 12376 3061 12508 3095
rect 12342 3051 12508 3061
rect 12585 3107 12678 3123
rect 12619 3073 12678 3107
rect 12585 3057 12678 3073
rect 12342 3045 12382 3051
rect 12406 3001 12440 3015
rect 12266 2999 12440 3001
rect 12266 2967 12406 2999
rect 12338 2965 12406 2967
rect 12338 2949 12440 2965
rect 12048 2856 12109 2882
rect 12198 2873 12230 2907
rect 12266 2899 12304 2933
rect 12264 2873 12304 2899
rect 12198 2860 12304 2873
rect 11719 2771 11753 2787
rect 11787 2803 11803 2837
rect 11837 2803 11853 2837
rect 11787 2737 11853 2803
rect 11887 2821 11924 2855
rect 11921 2787 11924 2821
rect 11887 2771 11924 2787
rect 11972 2813 12025 2829
rect 11972 2779 11991 2813
rect 11972 2737 12025 2779
rect 12059 2821 12109 2856
rect 12338 2826 12372 2949
rect 12059 2787 12075 2821
rect 12151 2792 12167 2826
rect 12201 2792 12372 2826
rect 12406 2881 12440 2897
rect 12406 2813 12440 2847
rect 12059 2771 12109 2787
rect 12406 2737 12440 2779
rect 12474 2837 12508 3051
rect 12542 2999 12580 3015
rect 12576 2965 12580 2999
rect 12542 2907 12580 2965
rect 12542 2873 12544 2907
rect 12578 2873 12580 2907
rect 12542 2871 12580 2873
rect 12614 2975 12678 3057
rect 12614 2941 12631 2975
rect 12665 2941 12678 2975
rect 12614 2933 12678 2941
rect 12614 2899 12644 2933
rect 12614 2865 12678 2899
rect 12712 3065 12746 3157
rect 12801 3157 12806 3191
rect 12840 3157 12843 3191
rect 12801 3141 12843 3157
rect 12895 3170 12911 3204
rect 12945 3170 12961 3204
rect 12895 3136 12961 3170
rect 12895 3102 12911 3136
rect 12945 3102 12961 3136
rect 12995 3175 13029 3247
rect 12995 3125 13029 3141
rect 13063 3202 13129 3203
rect 13063 3168 13079 3202
rect 13113 3179 13129 3202
rect 13063 3145 13093 3168
rect 13127 3145 13129 3179
rect 13063 3134 13129 3145
rect 13173 3186 14242 3247
rect 13173 3152 13191 3186
rect 13225 3152 14191 3186
rect 14225 3152 14242 3186
rect 13173 3138 14242 3152
rect 14277 3186 15346 3247
rect 14277 3152 14295 3186
rect 14329 3152 15295 3186
rect 15329 3152 15346 3186
rect 14277 3138 15346 3152
rect 15381 3186 16450 3247
rect 15381 3152 15399 3186
rect 15433 3152 16399 3186
rect 16433 3152 16450 3186
rect 15381 3138 16450 3152
rect 16577 3153 16635 3247
rect 12895 3099 12961 3102
rect 13063 3100 13079 3134
rect 13113 3116 13129 3134
rect 13113 3100 13139 3116
rect 13063 3099 13139 3100
rect 12921 3065 12961 3099
rect 13094 3091 13139 3099
rect 12712 3049 12887 3065
rect 12712 3015 12853 3049
rect 12712 2999 12887 3015
rect 12921 3049 13071 3065
rect 12921 3015 13037 3049
rect 12921 2999 13071 3015
rect 12474 2821 12524 2837
rect 12712 2831 12746 2999
rect 12921 2958 12959 2999
rect 13105 2975 13139 3091
rect 13096 2965 13139 2975
rect 13490 3023 13558 3138
rect 13490 2989 13507 3023
rect 13541 2989 13558 3023
rect 13490 2972 13558 2989
rect 13854 3059 13924 3074
rect 13854 3025 13871 3059
rect 13905 3025 13924 3059
rect 12780 2955 12959 2958
rect 12780 2933 12907 2955
rect 12814 2921 12907 2933
rect 12941 2921 12959 2955
rect 13061 2955 13139 2965
rect 12814 2899 12959 2921
rect 12780 2884 12959 2899
rect 12780 2883 12907 2884
rect 12891 2850 12907 2883
rect 12941 2850 12959 2884
rect 12474 2787 12490 2821
rect 12569 2797 12585 2831
rect 12619 2797 12746 2831
rect 12782 2821 12845 2837
rect 12474 2771 12524 2787
rect 12782 2787 12784 2821
rect 12818 2787 12845 2821
rect 12782 2737 12845 2787
rect 12891 2813 12959 2850
rect 12891 2779 12907 2813
rect 12941 2779 12959 2813
rect 12891 2771 12959 2779
rect 12993 2923 13027 2939
rect 12993 2843 13027 2889
rect 12993 2737 13027 2809
rect 13061 2921 13077 2955
rect 13111 2949 13139 2955
rect 13111 2921 13127 2949
rect 13061 2887 13127 2921
rect 13061 2853 13077 2887
rect 13111 2853 13127 2887
rect 13061 2819 13127 2853
rect 13854 2824 13924 3025
rect 14594 3023 14662 3138
rect 14594 2989 14611 3023
rect 14645 2989 14662 3023
rect 14594 2972 14662 2989
rect 14958 3059 15028 3074
rect 14958 3025 14975 3059
rect 15009 3025 15028 3059
rect 14958 2824 15028 3025
rect 15698 3023 15766 3138
rect 16577 3119 16589 3153
rect 16623 3119 16635 3153
rect 16577 3102 16635 3119
rect 16853 3175 16905 3213
rect 16853 3141 16871 3175
rect 16941 3205 17007 3247
rect 16941 3171 16957 3205
rect 16991 3171 17007 3205
rect 17043 3192 17077 3213
rect 16853 3112 16905 3141
rect 17043 3137 17077 3158
rect 17129 3186 18198 3247
rect 17129 3152 17147 3186
rect 17181 3152 18147 3186
rect 18181 3152 18198 3186
rect 17129 3138 18198 3152
rect 18233 3179 18567 3247
rect 18233 3145 18251 3179
rect 18285 3145 18515 3179
rect 18549 3145 18567 3179
rect 15698 2989 15715 3023
rect 15749 2989 15766 3023
rect 15698 2972 15766 2989
rect 16062 3059 16132 3074
rect 16062 3025 16079 3059
rect 16113 3025 16132 3059
rect 16062 2824 16132 3025
rect 16577 2935 16635 2970
rect 16577 2901 16589 2935
rect 16623 2901 16635 2935
rect 16577 2842 16635 2901
rect 13061 2785 13077 2819
rect 13111 2785 13127 2819
rect 13061 2780 13127 2785
rect 13173 2813 14242 2824
rect 13173 2779 13191 2813
rect 13225 2779 14191 2813
rect 14225 2779 14242 2813
rect 13173 2737 14242 2779
rect 14277 2813 15346 2824
rect 14277 2779 14295 2813
rect 14329 2779 15295 2813
rect 15329 2779 15346 2813
rect 14277 2737 15346 2779
rect 15381 2813 16450 2824
rect 15381 2779 15399 2813
rect 15433 2779 16399 2813
rect 16433 2779 16450 2813
rect 15381 2737 16450 2779
rect 16577 2808 16589 2842
rect 16623 2808 16635 2842
rect 16577 2737 16635 2808
rect 16853 2952 16887 3112
rect 16944 3103 17077 3137
rect 16944 3052 16978 3103
rect 16921 3036 16978 3052
rect 16955 3002 16978 3036
rect 16921 2986 16978 3002
rect 17025 3049 17091 3067
rect 17025 3015 17041 3049
rect 17075 3043 17091 3049
rect 17025 3009 17049 3015
rect 17083 3009 17091 3043
rect 17025 2993 17091 3009
rect 17446 3023 17514 3138
rect 18233 3093 18567 3145
rect 18601 3184 18843 3247
rect 18601 3150 18619 3184
rect 18653 3150 18791 3184
rect 18825 3150 18843 3184
rect 18601 3097 18843 3150
rect 16944 2957 16978 2986
rect 17446 2989 17463 3023
rect 17497 2989 17514 3023
rect 17446 2972 17514 2989
rect 17810 3059 17880 3074
rect 17810 3025 17827 3059
rect 17861 3025 17880 3059
rect 16853 2902 16907 2952
rect 16944 2923 17077 2957
rect 16853 2868 16871 2902
rect 16905 2868 16907 2902
rect 17043 2889 17077 2923
rect 16853 2839 16907 2868
rect 16853 2805 16865 2839
rect 16899 2821 16907 2839
rect 16853 2787 16871 2805
rect 16905 2787 16907 2821
rect 16853 2771 16907 2787
rect 16941 2855 16957 2889
rect 16991 2855 17007 2889
rect 16941 2821 17007 2855
rect 16941 2787 16957 2821
rect 16991 2787 17007 2821
rect 16941 2737 17007 2787
rect 17043 2821 17077 2855
rect 17810 2824 17880 3025
rect 18233 3023 18383 3093
rect 18233 2989 18253 3023
rect 18287 2989 18383 3023
rect 18417 3025 18513 3059
rect 18547 3025 18567 3059
rect 18417 2955 18567 3025
rect 18233 2915 18567 2955
rect 18233 2881 18251 2915
rect 18285 2881 18515 2915
rect 18549 2881 18567 2915
rect 17043 2771 17077 2787
rect 17129 2813 18198 2824
rect 17129 2779 17147 2813
rect 17181 2779 18147 2813
rect 18181 2779 18198 2813
rect 17129 2737 18198 2779
rect 18233 2813 18567 2881
rect 18233 2779 18251 2813
rect 18285 2779 18515 2813
rect 18549 2779 18567 2813
rect 18233 2737 18567 2779
rect 18601 3029 18651 3063
rect 18685 3029 18705 3063
rect 18601 2955 18705 3029
rect 18739 3023 18843 3097
rect 18739 2989 18759 3023
rect 18793 2989 18843 3023
rect 18601 2908 18843 2955
rect 18601 2874 18619 2908
rect 18653 2874 18791 2908
rect 18825 2874 18843 2908
rect 18601 2813 18843 2874
rect 18601 2779 18619 2813
rect 18653 2779 18791 2813
rect 18825 2779 18843 2813
rect 18601 2737 18843 2779
rect 1104 2703 1133 2737
rect 1167 2703 1225 2737
rect 1259 2703 1317 2737
rect 1351 2703 1409 2737
rect 1443 2703 1501 2737
rect 1535 2703 1593 2737
rect 1627 2703 1685 2737
rect 1719 2703 1777 2737
rect 1811 2703 1869 2737
rect 1903 2703 1961 2737
rect 1995 2703 2053 2737
rect 2087 2703 2145 2737
rect 2179 2703 2237 2737
rect 2271 2703 2329 2737
rect 2363 2703 2421 2737
rect 2455 2703 2513 2737
rect 2547 2703 2605 2737
rect 2639 2703 2697 2737
rect 2731 2703 2789 2737
rect 2823 2703 2881 2737
rect 2915 2703 2973 2737
rect 3007 2703 3065 2737
rect 3099 2703 3157 2737
rect 3191 2703 3249 2737
rect 3283 2703 3341 2737
rect 3375 2703 3433 2737
rect 3467 2703 3525 2737
rect 3559 2703 3617 2737
rect 3651 2703 3709 2737
rect 3743 2703 3801 2737
rect 3835 2703 3893 2737
rect 3927 2703 3985 2737
rect 4019 2703 4077 2737
rect 4111 2703 4169 2737
rect 4203 2703 4261 2737
rect 4295 2703 4353 2737
rect 4387 2703 4445 2737
rect 4479 2703 4537 2737
rect 4571 2703 4629 2737
rect 4663 2703 4721 2737
rect 4755 2703 4813 2737
rect 4847 2703 4905 2737
rect 4939 2703 4997 2737
rect 5031 2703 5089 2737
rect 5123 2703 5181 2737
rect 5215 2703 5273 2737
rect 5307 2703 5365 2737
rect 5399 2703 5457 2737
rect 5491 2703 5549 2737
rect 5583 2703 5641 2737
rect 5675 2703 5733 2737
rect 5767 2703 5825 2737
rect 5859 2703 5917 2737
rect 5951 2703 6009 2737
rect 6043 2703 6101 2737
rect 6135 2703 6193 2737
rect 6227 2703 6285 2737
rect 6319 2703 6377 2737
rect 6411 2703 6469 2737
rect 6503 2703 6561 2737
rect 6595 2703 6653 2737
rect 6687 2703 6745 2737
rect 6779 2703 6837 2737
rect 6871 2703 6929 2737
rect 6963 2703 7021 2737
rect 7055 2703 7113 2737
rect 7147 2703 7205 2737
rect 7239 2703 7297 2737
rect 7331 2703 7389 2737
rect 7423 2703 7481 2737
rect 7515 2703 7573 2737
rect 7607 2703 7665 2737
rect 7699 2703 7757 2737
rect 7791 2703 7849 2737
rect 7883 2703 7941 2737
rect 7975 2703 8033 2737
rect 8067 2703 8125 2737
rect 8159 2703 8217 2737
rect 8251 2703 8309 2737
rect 8343 2703 8401 2737
rect 8435 2703 8493 2737
rect 8527 2703 8585 2737
rect 8619 2703 8677 2737
rect 8711 2703 8769 2737
rect 8803 2703 8861 2737
rect 8895 2703 8953 2737
rect 8987 2703 9045 2737
rect 9079 2703 9137 2737
rect 9171 2703 9229 2737
rect 9263 2703 9321 2737
rect 9355 2703 9413 2737
rect 9447 2703 9505 2737
rect 9539 2703 9597 2737
rect 9631 2703 9689 2737
rect 9723 2703 9781 2737
rect 9815 2703 9873 2737
rect 9907 2703 9965 2737
rect 9999 2703 10057 2737
rect 10091 2703 10149 2737
rect 10183 2703 10241 2737
rect 10275 2703 10333 2737
rect 10367 2703 10425 2737
rect 10459 2703 10517 2737
rect 10551 2703 10609 2737
rect 10643 2703 10701 2737
rect 10735 2703 10793 2737
rect 10827 2703 10885 2737
rect 10919 2703 10977 2737
rect 11011 2703 11069 2737
rect 11103 2703 11161 2737
rect 11195 2703 11253 2737
rect 11287 2703 11345 2737
rect 11379 2703 11437 2737
rect 11471 2703 11529 2737
rect 11563 2703 11621 2737
rect 11655 2703 11713 2737
rect 11747 2703 11805 2737
rect 11839 2703 11897 2737
rect 11931 2703 11989 2737
rect 12023 2703 12081 2737
rect 12115 2703 12173 2737
rect 12207 2703 12265 2737
rect 12299 2703 12357 2737
rect 12391 2703 12449 2737
rect 12483 2703 12541 2737
rect 12575 2703 12633 2737
rect 12667 2703 12725 2737
rect 12759 2703 12817 2737
rect 12851 2703 12909 2737
rect 12943 2703 13001 2737
rect 13035 2703 13093 2737
rect 13127 2703 13185 2737
rect 13219 2703 13277 2737
rect 13311 2703 13369 2737
rect 13403 2703 13461 2737
rect 13495 2703 13553 2737
rect 13587 2703 13645 2737
rect 13679 2703 13737 2737
rect 13771 2703 13829 2737
rect 13863 2703 13921 2737
rect 13955 2703 14013 2737
rect 14047 2703 14105 2737
rect 14139 2703 14197 2737
rect 14231 2703 14289 2737
rect 14323 2703 14381 2737
rect 14415 2703 14473 2737
rect 14507 2703 14565 2737
rect 14599 2703 14657 2737
rect 14691 2703 14749 2737
rect 14783 2703 14841 2737
rect 14875 2703 14933 2737
rect 14967 2703 15025 2737
rect 15059 2703 15117 2737
rect 15151 2703 15209 2737
rect 15243 2703 15301 2737
rect 15335 2703 15393 2737
rect 15427 2703 15485 2737
rect 15519 2703 15577 2737
rect 15611 2703 15669 2737
rect 15703 2703 15761 2737
rect 15795 2703 15853 2737
rect 15887 2703 15945 2737
rect 15979 2703 16037 2737
rect 16071 2703 16129 2737
rect 16163 2703 16221 2737
rect 16255 2703 16313 2737
rect 16347 2703 16405 2737
rect 16439 2703 16497 2737
rect 16531 2703 16589 2737
rect 16623 2703 16681 2737
rect 16715 2703 16773 2737
rect 16807 2703 16865 2737
rect 16899 2703 16957 2737
rect 16991 2703 17049 2737
rect 17083 2703 17141 2737
rect 17175 2703 17233 2737
rect 17267 2703 17325 2737
rect 17359 2703 17417 2737
rect 17451 2703 17509 2737
rect 17543 2703 17601 2737
rect 17635 2703 17693 2737
rect 17727 2703 17785 2737
rect 17819 2703 17877 2737
rect 17911 2703 17969 2737
rect 18003 2703 18061 2737
rect 18095 2703 18153 2737
rect 18187 2703 18245 2737
rect 18279 2703 18337 2737
rect 18371 2703 18429 2737
rect 18463 2703 18521 2737
rect 18555 2703 18613 2737
rect 18647 2703 18705 2737
rect 18739 2703 18797 2737
rect 18831 2703 18860 2737
rect 1121 2661 1363 2703
rect 1121 2627 1139 2661
rect 1173 2627 1311 2661
rect 1345 2627 1363 2661
rect 1121 2566 1363 2627
rect 1121 2532 1139 2566
rect 1173 2532 1311 2566
rect 1345 2532 1363 2566
rect 1121 2485 1363 2532
rect 1397 2661 1915 2703
rect 1397 2627 1415 2661
rect 1449 2627 1863 2661
rect 1897 2627 1915 2661
rect 1397 2559 1915 2627
rect 1397 2525 1415 2559
rect 1449 2525 1863 2559
rect 1897 2525 1915 2559
rect 1397 2485 1915 2525
rect 2053 2655 2119 2660
rect 2053 2635 2069 2655
rect 2103 2621 2119 2655
rect 2087 2601 2119 2621
rect 2053 2587 2119 2601
rect 2053 2553 2069 2587
rect 2103 2553 2119 2587
rect 2053 2519 2119 2553
rect 2053 2491 2069 2519
rect 1121 2417 1171 2451
rect 1205 2417 1225 2451
rect 1121 2343 1225 2417
rect 1259 2411 1363 2485
rect 1259 2377 1279 2411
rect 1313 2377 1363 2411
rect 1397 2417 1475 2451
rect 1509 2417 1585 2451
rect 1619 2417 1639 2451
rect 1397 2347 1639 2417
rect 1673 2415 1915 2485
rect 1673 2381 1693 2415
rect 1727 2381 1803 2415
rect 1837 2381 1915 2415
rect 2041 2485 2069 2491
rect 2103 2485 2119 2519
rect 2153 2631 2187 2703
rect 2153 2551 2187 2597
rect 2153 2501 2187 2517
rect 2221 2661 2289 2669
rect 2221 2627 2239 2661
rect 2273 2627 2289 2661
rect 2221 2590 2289 2627
rect 2335 2653 2398 2703
rect 2335 2619 2362 2653
rect 2396 2619 2398 2653
rect 2656 2653 2706 2669
rect 2335 2603 2398 2619
rect 2434 2609 2561 2643
rect 2595 2609 2611 2643
rect 2690 2619 2706 2653
rect 2221 2556 2239 2590
rect 2273 2557 2289 2590
rect 2273 2556 2400 2557
rect 2221 2541 2400 2556
rect 2221 2519 2366 2541
rect 2041 2475 2119 2485
rect 2221 2485 2239 2519
rect 2273 2507 2366 2519
rect 2273 2485 2400 2507
rect 2221 2482 2400 2485
rect 2041 2465 2084 2475
rect 2041 2349 2075 2465
rect 2221 2441 2259 2482
rect 2434 2441 2468 2609
rect 2656 2603 2706 2619
rect 2109 2425 2259 2441
rect 2143 2391 2259 2425
rect 2109 2375 2259 2391
rect 2293 2425 2468 2441
rect 2327 2391 2468 2425
rect 2293 2375 2468 2391
rect 1121 2290 1363 2343
rect 1121 2256 1139 2290
rect 1173 2256 1311 2290
rect 1345 2256 1363 2290
rect 1121 2193 1363 2256
rect 1397 2288 1915 2347
rect 2041 2341 2086 2349
rect 2219 2341 2259 2375
rect 2041 2340 2117 2341
rect 2041 2324 2067 2340
rect 1397 2254 1415 2288
rect 1449 2254 1863 2288
rect 1897 2254 1915 2288
rect 1397 2193 1915 2254
rect 2051 2306 2067 2324
rect 2101 2306 2117 2340
rect 2219 2338 2285 2341
rect 2051 2272 2117 2306
rect 2051 2238 2067 2272
rect 2101 2238 2117 2272
rect 2051 2237 2117 2238
rect 2151 2299 2185 2315
rect 2151 2193 2185 2265
rect 2219 2304 2235 2338
rect 2269 2304 2285 2338
rect 2219 2270 2285 2304
rect 2219 2236 2235 2270
rect 2269 2236 2285 2270
rect 2337 2283 2379 2299
rect 2337 2249 2340 2283
rect 2374 2249 2379 2283
rect 2434 2283 2468 2375
rect 2502 2541 2566 2575
rect 2536 2507 2566 2541
rect 2502 2499 2566 2507
rect 2502 2465 2515 2499
rect 2549 2465 2566 2499
rect 2502 2383 2566 2465
rect 2600 2567 2638 2569
rect 2600 2533 2602 2567
rect 2636 2533 2638 2567
rect 2600 2475 2638 2533
rect 2600 2441 2604 2475
rect 2600 2425 2638 2441
rect 2672 2389 2706 2603
rect 2740 2661 2774 2703
rect 3071 2653 3121 2669
rect 2740 2593 2774 2627
rect 2740 2543 2774 2559
rect 2808 2614 2979 2648
rect 3013 2614 3029 2648
rect 3105 2619 3121 2653
rect 2808 2491 2842 2614
rect 3071 2584 3121 2619
rect 3155 2661 3208 2703
rect 3189 2627 3208 2661
rect 3155 2611 3208 2627
rect 3256 2653 3293 2669
rect 3256 2619 3259 2653
rect 3256 2585 3293 2619
rect 3327 2637 3393 2703
rect 3327 2603 3343 2637
rect 3377 2603 3393 2637
rect 3427 2653 3461 2669
rect 2876 2567 2982 2580
rect 2876 2541 2916 2567
rect 2876 2507 2914 2541
rect 2950 2533 2982 2567
rect 3071 2558 3132 2584
rect 2740 2475 2842 2491
rect 2774 2473 2842 2475
rect 2774 2441 2914 2473
rect 2740 2439 2914 2441
rect 2740 2425 2774 2439
rect 2798 2389 2838 2395
rect 2502 2367 2595 2383
rect 2502 2333 2561 2367
rect 2502 2317 2595 2333
rect 2672 2379 2838 2389
rect 2672 2345 2804 2379
rect 2672 2329 2838 2345
rect 2672 2283 2706 2329
rect 2434 2249 2538 2283
rect 2572 2249 2591 2283
rect 2625 2249 2641 2283
rect 2675 2249 2706 2283
rect 2742 2277 2816 2293
rect 2337 2193 2379 2249
rect 2742 2243 2760 2277
rect 2794 2243 2816 2277
rect 2880 2283 2914 2439
rect 2948 2367 2982 2533
rect 3016 2499 3064 2520
rect 3016 2465 3019 2499
rect 3053 2465 3064 2499
rect 3016 2463 3064 2465
rect 3016 2429 3023 2463
rect 3057 2429 3064 2463
rect 3016 2401 3064 2429
rect 2948 2333 3003 2367
rect 3037 2333 3053 2367
rect 3098 2337 3132 2558
rect 3256 2551 3259 2585
rect 3427 2585 3461 2619
rect 2948 2323 3053 2333
rect 3087 2311 3132 2337
rect 3166 2493 3222 2509
rect 3200 2459 3222 2493
rect 3166 2431 3222 2459
rect 3166 2397 3177 2431
rect 3211 2397 3222 2431
rect 3166 2319 3222 2397
rect 3256 2499 3293 2551
rect 3256 2465 3257 2499
rect 3291 2465 3293 2499
rect 3087 2283 3121 2311
rect 3256 2295 3293 2465
rect 3328 2567 3427 2569
rect 3328 2533 3336 2567
rect 3370 2551 3427 2567
rect 3370 2535 3461 2551
rect 3697 2632 3755 2703
rect 3697 2598 3709 2632
rect 3743 2598 3755 2632
rect 3697 2539 3755 2598
rect 3370 2533 3374 2535
rect 3328 2440 3374 2533
rect 3697 2505 3709 2539
rect 3743 2505 3755 2539
rect 3362 2406 3374 2440
rect 3328 2337 3374 2406
rect 3408 2499 3478 2501
rect 3408 2465 3433 2499
rect 3467 2465 3478 2499
rect 3697 2470 3755 2505
rect 3408 2425 3478 2465
rect 3408 2391 3430 2425
rect 3464 2391 3478 2425
rect 3408 2371 3478 2391
rect 3328 2303 3461 2337
rect 2880 2249 2959 2283
rect 2993 2249 3015 2283
rect 3054 2249 3070 2283
rect 3104 2249 3121 2283
rect 3155 2269 3205 2285
rect 2742 2193 2816 2243
rect 3189 2235 3205 2269
rect 3256 2261 3259 2295
rect 3427 2295 3461 2303
rect 3256 2245 3293 2261
rect 3155 2193 3205 2235
rect 3327 2235 3343 2269
rect 3377 2235 3393 2269
rect 3427 2245 3461 2261
rect 3697 2321 3755 2338
rect 3697 2287 3709 2321
rect 3743 2287 3755 2321
rect 3327 2193 3393 2235
rect 3697 2193 3755 2287
rect 3973 2335 4123 2669
rect 4157 2661 4491 2703
rect 4157 2627 4175 2661
rect 4209 2627 4439 2661
rect 4473 2627 4491 2661
rect 4157 2559 4491 2627
rect 4157 2525 4175 2559
rect 4209 2525 4439 2559
rect 4473 2525 4491 2559
rect 4635 2653 4669 2669
rect 4635 2585 4669 2619
rect 4703 2637 4769 2703
rect 4703 2603 4719 2637
rect 4753 2603 4769 2637
rect 4803 2653 4840 2669
rect 4837 2619 4840 2653
rect 4803 2585 4840 2619
rect 4888 2661 4941 2703
rect 4888 2627 4907 2661
rect 4888 2611 4941 2627
rect 4975 2653 5025 2669
rect 4975 2619 4991 2653
rect 5322 2661 5356 2703
rect 4669 2567 4768 2569
rect 4669 2551 4726 2567
rect 4635 2535 4726 2551
rect 4157 2485 4491 2525
rect 4722 2533 4726 2535
rect 4760 2533 4768 2567
rect 3973 2301 3991 2335
rect 4025 2301 4066 2335
rect 4100 2301 4123 2335
rect 3973 2295 4123 2301
rect 3973 2261 3985 2295
rect 4019 2267 4123 2295
rect 3973 2233 3991 2261
rect 4025 2233 4066 2267
rect 4100 2233 4123 2267
rect 3973 2227 4123 2233
rect 4157 2417 4177 2451
rect 4211 2417 4307 2451
rect 4157 2347 4307 2417
rect 4341 2415 4491 2485
rect 4341 2381 4437 2415
rect 4471 2381 4491 2415
rect 4618 2499 4688 2501
rect 4618 2465 4629 2499
rect 4663 2465 4688 2499
rect 4618 2425 4688 2465
rect 4618 2391 4632 2425
rect 4666 2391 4688 2425
rect 4618 2371 4688 2391
rect 4722 2440 4768 2533
rect 4722 2406 4734 2440
rect 4157 2295 4491 2347
rect 4722 2337 4768 2406
rect 4157 2261 4175 2295
rect 4209 2261 4439 2295
rect 4473 2261 4491 2295
rect 4157 2193 4491 2261
rect 4635 2303 4768 2337
rect 4837 2551 4840 2585
rect 4975 2584 5025 2619
rect 5067 2614 5083 2648
rect 5117 2614 5288 2648
rect 4803 2499 4840 2551
rect 4964 2558 5025 2584
rect 5114 2567 5220 2580
rect 4803 2465 4805 2499
rect 4839 2465 4840 2499
rect 4635 2295 4669 2303
rect 4803 2295 4840 2465
rect 4874 2493 4930 2509
rect 4874 2459 4896 2493
rect 4874 2363 4930 2459
rect 4908 2329 4930 2363
rect 4874 2319 4930 2329
rect 4964 2337 4998 2558
rect 5114 2533 5146 2567
rect 5180 2541 5220 2567
rect 5032 2499 5080 2520
rect 5032 2465 5043 2499
rect 5077 2465 5080 2499
rect 5032 2463 5080 2465
rect 5032 2429 5039 2463
rect 5073 2429 5080 2463
rect 5032 2401 5080 2429
rect 5114 2367 5148 2533
rect 5182 2507 5220 2541
rect 5254 2491 5288 2614
rect 5322 2593 5356 2627
rect 5322 2543 5356 2559
rect 5390 2653 5440 2669
rect 5390 2619 5406 2653
rect 5698 2653 5761 2703
rect 5390 2603 5440 2619
rect 5485 2609 5501 2643
rect 5535 2609 5662 2643
rect 5254 2475 5356 2491
rect 5254 2473 5322 2475
rect 4964 2311 5009 2337
rect 5043 2333 5059 2367
rect 5093 2333 5148 2367
rect 5043 2323 5148 2333
rect 5182 2441 5322 2473
rect 5182 2439 5356 2441
rect 4635 2245 4669 2261
rect 4703 2235 4719 2269
rect 4753 2235 4769 2269
rect 4837 2261 4840 2295
rect 4803 2245 4840 2261
rect 4891 2269 4941 2285
rect 4703 2193 4769 2235
rect 4891 2235 4907 2269
rect 4975 2283 5009 2311
rect 5182 2283 5216 2439
rect 5322 2425 5356 2439
rect 5258 2389 5298 2395
rect 5390 2389 5424 2603
rect 5458 2567 5496 2569
rect 5458 2533 5460 2567
rect 5494 2533 5496 2567
rect 5458 2475 5496 2533
rect 5492 2441 5496 2475
rect 5458 2425 5496 2441
rect 5530 2541 5594 2575
rect 5530 2507 5560 2541
rect 5530 2499 5594 2507
rect 5530 2465 5547 2499
rect 5581 2465 5594 2499
rect 5258 2379 5424 2389
rect 5530 2383 5594 2465
rect 5292 2345 5424 2379
rect 5258 2329 5424 2345
rect 4975 2249 4992 2283
rect 5026 2249 5042 2283
rect 5081 2249 5103 2283
rect 5137 2249 5216 2283
rect 5280 2277 5354 2293
rect 4891 2193 4941 2235
rect 5280 2243 5302 2277
rect 5336 2243 5354 2277
rect 5390 2283 5424 2329
rect 5501 2367 5594 2383
rect 5535 2333 5594 2367
rect 5501 2317 5594 2333
rect 5628 2441 5662 2609
rect 5698 2619 5700 2653
rect 5734 2619 5761 2653
rect 5698 2603 5761 2619
rect 5807 2661 5875 2669
rect 5807 2627 5823 2661
rect 5857 2627 5875 2661
rect 5807 2590 5875 2627
rect 5807 2557 5823 2590
rect 5696 2556 5823 2557
rect 5857 2556 5875 2590
rect 5696 2541 5875 2556
rect 5730 2519 5875 2541
rect 5730 2507 5823 2519
rect 5696 2485 5823 2507
rect 5857 2485 5875 2519
rect 5909 2631 5943 2703
rect 5909 2551 5943 2597
rect 5909 2501 5943 2517
rect 5977 2655 6043 2660
rect 5977 2621 5993 2655
rect 6027 2635 6043 2655
rect 5977 2601 6009 2621
rect 5977 2587 6043 2601
rect 5977 2553 5993 2587
rect 6027 2553 6043 2587
rect 5977 2519 6043 2553
rect 5696 2482 5875 2485
rect 5837 2441 5875 2482
rect 5977 2485 5993 2519
rect 6027 2491 6043 2519
rect 6273 2632 6331 2703
rect 6273 2598 6285 2632
rect 6319 2598 6331 2632
rect 6273 2539 6331 2598
rect 6273 2505 6285 2539
rect 6319 2505 6331 2539
rect 6027 2485 6055 2491
rect 5977 2475 6055 2485
rect 6012 2465 6055 2475
rect 6273 2470 6331 2505
rect 6365 2661 7067 2703
rect 6365 2627 6383 2661
rect 6417 2627 7015 2661
rect 7049 2627 7067 2661
rect 6365 2559 7067 2627
rect 6365 2525 6383 2559
rect 6417 2525 7015 2559
rect 7049 2525 7067 2559
rect 6365 2485 7067 2525
rect 7205 2655 7271 2660
rect 7205 2621 7221 2655
rect 7255 2621 7271 2655
rect 7205 2587 7271 2621
rect 7205 2553 7221 2587
rect 7255 2553 7271 2587
rect 7205 2519 7271 2553
rect 7205 2491 7221 2519
rect 5628 2425 5803 2441
rect 5628 2391 5769 2425
rect 5628 2375 5803 2391
rect 5837 2425 5987 2441
rect 5837 2391 5953 2425
rect 5837 2375 5987 2391
rect 5628 2283 5662 2375
rect 5837 2341 5877 2375
rect 6021 2349 6055 2465
rect 6010 2341 6055 2349
rect 5811 2338 5877 2341
rect 5811 2304 5827 2338
rect 5861 2304 5877 2338
rect 5979 2340 6055 2341
rect 5390 2249 5421 2283
rect 5455 2249 5471 2283
rect 5505 2249 5524 2283
rect 5558 2249 5662 2283
rect 5717 2283 5759 2299
rect 5717 2249 5722 2283
rect 5756 2249 5759 2283
rect 5280 2193 5354 2243
rect 5717 2193 5759 2249
rect 5811 2270 5877 2304
rect 5811 2236 5827 2270
rect 5861 2236 5877 2270
rect 5911 2299 5945 2315
rect 5911 2193 5945 2265
rect 5979 2306 5995 2340
rect 6029 2324 6055 2340
rect 6365 2417 6443 2451
rect 6477 2417 6542 2451
rect 6576 2417 6641 2451
rect 6675 2417 6695 2451
rect 6365 2347 6695 2417
rect 6729 2415 7067 2485
rect 6729 2381 6749 2415
rect 6783 2381 6852 2415
rect 6886 2381 6955 2415
rect 6989 2381 7067 2415
rect 7193 2485 7221 2491
rect 7255 2485 7271 2519
rect 7305 2631 7339 2703
rect 7305 2551 7339 2597
rect 7305 2501 7339 2517
rect 7373 2661 7441 2669
rect 7373 2627 7391 2661
rect 7425 2627 7441 2661
rect 7373 2590 7441 2627
rect 7487 2653 7550 2703
rect 7487 2619 7514 2653
rect 7548 2619 7550 2653
rect 7808 2653 7858 2669
rect 7487 2603 7550 2619
rect 7586 2609 7713 2643
rect 7747 2609 7763 2643
rect 7842 2619 7858 2653
rect 7373 2556 7391 2590
rect 7425 2557 7441 2590
rect 7425 2556 7552 2557
rect 7373 2541 7552 2556
rect 7373 2519 7518 2541
rect 7193 2475 7271 2485
rect 7373 2485 7391 2519
rect 7425 2507 7518 2519
rect 7425 2485 7552 2507
rect 7373 2482 7552 2485
rect 7193 2465 7236 2475
rect 7193 2349 7227 2465
rect 7373 2441 7411 2482
rect 7586 2441 7620 2609
rect 7808 2603 7858 2619
rect 7261 2425 7411 2441
rect 7295 2391 7411 2425
rect 7261 2375 7411 2391
rect 7445 2425 7620 2441
rect 7479 2391 7620 2425
rect 7445 2375 7620 2391
rect 6029 2306 6045 2324
rect 5979 2272 6045 2306
rect 5979 2238 5995 2272
rect 6029 2238 6045 2272
rect 5979 2237 6045 2238
rect 6273 2321 6331 2338
rect 6273 2287 6285 2321
rect 6319 2287 6331 2321
rect 6273 2193 6331 2287
rect 6365 2288 7067 2347
rect 7193 2341 7238 2349
rect 7371 2341 7411 2375
rect 7193 2340 7269 2341
rect 7193 2324 7219 2340
rect 6365 2254 6383 2288
rect 6417 2254 7015 2288
rect 7049 2254 7067 2288
rect 6365 2193 7067 2254
rect 7203 2306 7219 2324
rect 7253 2306 7269 2340
rect 7371 2338 7437 2341
rect 7203 2295 7269 2306
rect 7203 2261 7205 2295
rect 7239 2272 7269 2295
rect 7203 2238 7219 2261
rect 7253 2238 7269 2272
rect 7203 2237 7269 2238
rect 7303 2299 7337 2315
rect 7303 2193 7337 2265
rect 7371 2304 7387 2338
rect 7421 2304 7437 2338
rect 7371 2270 7437 2304
rect 7371 2236 7387 2270
rect 7421 2236 7437 2270
rect 7489 2283 7531 2299
rect 7489 2249 7492 2283
rect 7526 2249 7531 2283
rect 7586 2283 7620 2375
rect 7654 2541 7718 2575
rect 7688 2507 7718 2541
rect 7654 2499 7718 2507
rect 7654 2465 7667 2499
rect 7701 2465 7718 2499
rect 7654 2383 7718 2465
rect 7752 2567 7790 2569
rect 7752 2533 7754 2567
rect 7788 2533 7790 2567
rect 7752 2475 7790 2533
rect 7752 2441 7756 2475
rect 7752 2425 7790 2441
rect 7824 2389 7858 2603
rect 7892 2661 7926 2703
rect 8223 2653 8273 2669
rect 7892 2593 7926 2627
rect 7892 2543 7926 2559
rect 7960 2614 8131 2648
rect 8165 2614 8181 2648
rect 8257 2619 8273 2653
rect 7960 2491 7994 2614
rect 8223 2584 8273 2619
rect 8307 2661 8360 2703
rect 8341 2627 8360 2661
rect 8307 2611 8360 2627
rect 8408 2653 8445 2669
rect 8408 2619 8411 2653
rect 8408 2585 8445 2619
rect 8479 2637 8545 2703
rect 8479 2603 8495 2637
rect 8529 2603 8545 2637
rect 8579 2653 8613 2669
rect 8028 2567 8134 2580
rect 8028 2541 8068 2567
rect 8028 2507 8066 2541
rect 8102 2533 8134 2567
rect 8223 2558 8284 2584
rect 7892 2475 7994 2491
rect 7926 2473 7994 2475
rect 7926 2441 8066 2473
rect 7892 2439 8066 2441
rect 7892 2425 7926 2439
rect 7950 2389 7990 2395
rect 7654 2367 7747 2383
rect 7654 2333 7713 2367
rect 7654 2317 7747 2333
rect 7824 2379 7990 2389
rect 7824 2345 7956 2379
rect 7824 2329 7990 2345
rect 7824 2283 7858 2329
rect 7586 2249 7690 2283
rect 7724 2249 7743 2283
rect 7777 2249 7793 2283
rect 7827 2249 7858 2283
rect 7894 2277 7968 2293
rect 7489 2193 7531 2249
rect 7894 2243 7912 2277
rect 7946 2243 7968 2277
rect 8032 2283 8066 2439
rect 8100 2367 8134 2533
rect 8168 2499 8216 2520
rect 8168 2465 8171 2499
rect 8205 2465 8216 2499
rect 8168 2463 8216 2465
rect 8168 2429 8175 2463
rect 8209 2429 8216 2463
rect 8168 2401 8216 2429
rect 8100 2333 8155 2367
rect 8189 2333 8205 2367
rect 8250 2337 8284 2558
rect 8408 2551 8411 2585
rect 8579 2585 8613 2619
rect 8100 2323 8205 2333
rect 8239 2311 8284 2337
rect 8318 2493 8374 2509
rect 8352 2459 8374 2493
rect 8318 2363 8374 2459
rect 8318 2329 8340 2363
rect 8318 2319 8374 2329
rect 8408 2499 8445 2551
rect 8408 2465 8409 2499
rect 8443 2465 8445 2499
rect 8239 2283 8273 2311
rect 8408 2295 8445 2465
rect 8480 2567 8579 2569
rect 8480 2533 8488 2567
rect 8522 2551 8579 2567
rect 8522 2535 8613 2551
rect 8849 2632 8907 2703
rect 8849 2598 8861 2632
rect 8895 2598 8907 2632
rect 8849 2539 8907 2598
rect 8522 2533 8526 2535
rect 8480 2440 8526 2533
rect 8849 2505 8861 2539
rect 8895 2505 8907 2539
rect 8514 2406 8526 2440
rect 8480 2337 8526 2406
rect 8560 2431 8630 2501
rect 8849 2470 8907 2505
rect 8941 2661 9643 2703
rect 8941 2627 8959 2661
rect 8993 2627 9591 2661
rect 9625 2627 9643 2661
rect 8941 2559 9643 2627
rect 8941 2525 8959 2559
rect 8993 2525 9591 2559
rect 9625 2525 9643 2559
rect 9787 2653 9821 2669
rect 9787 2585 9821 2619
rect 9855 2637 9921 2703
rect 9855 2603 9871 2637
rect 9905 2603 9921 2637
rect 9955 2653 9992 2669
rect 9989 2619 9992 2653
rect 9955 2585 9992 2619
rect 10040 2661 10093 2703
rect 10040 2627 10059 2661
rect 10040 2611 10093 2627
rect 10127 2653 10177 2669
rect 10127 2619 10143 2653
rect 10474 2661 10508 2703
rect 9821 2567 9920 2569
rect 9821 2551 9878 2567
rect 9787 2535 9878 2551
rect 8941 2485 9643 2525
rect 9874 2533 9878 2535
rect 9912 2533 9920 2567
rect 8560 2425 8585 2431
rect 8560 2391 8582 2425
rect 8619 2397 8630 2431
rect 8616 2391 8630 2397
rect 8560 2371 8630 2391
rect 8941 2417 9019 2451
rect 9053 2417 9118 2451
rect 9152 2417 9217 2451
rect 9251 2417 9271 2451
rect 8941 2347 9271 2417
rect 9305 2415 9643 2485
rect 9305 2381 9325 2415
rect 9359 2381 9428 2415
rect 9462 2381 9531 2415
rect 9565 2381 9643 2415
rect 9770 2431 9840 2501
rect 9770 2397 9781 2431
rect 9815 2425 9840 2431
rect 9770 2391 9784 2397
rect 9818 2391 9840 2425
rect 9770 2371 9840 2391
rect 9874 2440 9920 2533
rect 9874 2406 9886 2440
rect 8480 2303 8613 2337
rect 8032 2249 8111 2283
rect 8145 2249 8167 2283
rect 8206 2249 8222 2283
rect 8256 2249 8273 2283
rect 8307 2269 8357 2285
rect 7894 2193 7968 2243
rect 8341 2235 8357 2269
rect 8408 2261 8411 2295
rect 8579 2295 8613 2303
rect 8408 2245 8445 2261
rect 8307 2193 8357 2235
rect 8479 2235 8495 2269
rect 8529 2235 8545 2269
rect 8579 2245 8613 2261
rect 8849 2321 8907 2338
rect 8849 2287 8861 2321
rect 8895 2287 8907 2321
rect 8479 2193 8545 2235
rect 8849 2193 8907 2287
rect 8941 2288 9643 2347
rect 9874 2337 9920 2406
rect 8941 2254 8959 2288
rect 8993 2254 9591 2288
rect 9625 2254 9643 2288
rect 8941 2193 9643 2254
rect 9787 2303 9920 2337
rect 9989 2551 9992 2585
rect 10127 2584 10177 2619
rect 10219 2614 10235 2648
rect 10269 2614 10440 2648
rect 9955 2499 9992 2551
rect 10116 2558 10177 2584
rect 10266 2567 10372 2580
rect 9955 2465 9957 2499
rect 9991 2465 9992 2499
rect 9787 2295 9821 2303
rect 9955 2295 9992 2465
rect 10026 2493 10082 2509
rect 10026 2459 10048 2493
rect 10026 2363 10082 2459
rect 10026 2329 10048 2363
rect 10026 2319 10082 2329
rect 10116 2337 10150 2558
rect 10266 2533 10298 2567
rect 10332 2541 10372 2567
rect 10184 2499 10232 2520
rect 10184 2465 10195 2499
rect 10229 2465 10232 2499
rect 10184 2463 10232 2465
rect 10184 2429 10191 2463
rect 10225 2429 10232 2463
rect 10184 2401 10232 2429
rect 10266 2367 10300 2533
rect 10334 2507 10372 2541
rect 10406 2491 10440 2614
rect 10474 2593 10508 2627
rect 10474 2543 10508 2559
rect 10542 2653 10592 2669
rect 10542 2619 10558 2653
rect 10850 2653 10913 2703
rect 10542 2603 10592 2619
rect 10637 2609 10653 2643
rect 10687 2609 10814 2643
rect 10406 2475 10508 2491
rect 10406 2473 10474 2475
rect 10116 2311 10161 2337
rect 10195 2333 10211 2367
rect 10245 2333 10300 2367
rect 10195 2323 10300 2333
rect 10334 2441 10474 2473
rect 10334 2439 10508 2441
rect 9787 2245 9821 2261
rect 9855 2235 9871 2269
rect 9905 2235 9921 2269
rect 9989 2261 9992 2295
rect 9955 2245 9992 2261
rect 10043 2269 10093 2285
rect 9855 2193 9921 2235
rect 10043 2235 10059 2269
rect 10127 2283 10161 2311
rect 10334 2283 10368 2439
rect 10474 2425 10508 2439
rect 10410 2389 10450 2395
rect 10542 2389 10576 2603
rect 10610 2567 10648 2569
rect 10610 2533 10612 2567
rect 10646 2533 10648 2567
rect 10610 2475 10648 2533
rect 10644 2441 10648 2475
rect 10610 2425 10648 2441
rect 10682 2541 10746 2575
rect 10682 2507 10712 2541
rect 10682 2499 10746 2507
rect 10682 2465 10699 2499
rect 10733 2465 10746 2499
rect 10410 2379 10576 2389
rect 10682 2383 10746 2465
rect 10444 2345 10576 2379
rect 10410 2329 10576 2345
rect 10127 2249 10144 2283
rect 10178 2249 10194 2283
rect 10233 2249 10255 2283
rect 10289 2249 10368 2283
rect 10432 2277 10506 2293
rect 10043 2193 10093 2235
rect 10432 2243 10454 2277
rect 10488 2243 10506 2277
rect 10542 2283 10576 2329
rect 10653 2367 10746 2383
rect 10687 2333 10746 2367
rect 10653 2317 10746 2333
rect 10780 2441 10814 2609
rect 10850 2619 10852 2653
rect 10886 2619 10913 2653
rect 10850 2603 10913 2619
rect 10959 2661 11027 2669
rect 10959 2627 10975 2661
rect 11009 2627 11027 2661
rect 10959 2590 11027 2627
rect 10959 2557 10975 2590
rect 10848 2556 10975 2557
rect 11009 2556 11027 2590
rect 10848 2541 11027 2556
rect 10882 2519 11027 2541
rect 10882 2507 10975 2519
rect 10848 2485 10975 2507
rect 11009 2485 11027 2519
rect 11061 2631 11095 2703
rect 11061 2551 11095 2597
rect 11061 2501 11095 2517
rect 11129 2655 11195 2660
rect 11129 2621 11145 2655
rect 11179 2621 11195 2655
rect 11129 2587 11195 2621
rect 11129 2553 11145 2587
rect 11179 2567 11195 2587
rect 11129 2533 11161 2553
rect 11129 2519 11195 2533
rect 10848 2482 11027 2485
rect 10989 2441 11027 2482
rect 11129 2485 11145 2519
rect 11179 2491 11195 2519
rect 11425 2632 11483 2703
rect 11425 2598 11437 2632
rect 11471 2598 11483 2632
rect 11425 2539 11483 2598
rect 11425 2505 11437 2539
rect 11471 2505 11483 2539
rect 11179 2485 11207 2491
rect 11129 2475 11207 2485
rect 11164 2465 11207 2475
rect 11425 2470 11483 2505
rect 11517 2661 11851 2703
rect 11517 2627 11535 2661
rect 11569 2627 11799 2661
rect 11833 2627 11851 2661
rect 11517 2559 11851 2627
rect 11517 2525 11535 2559
rect 11569 2525 11799 2559
rect 11833 2525 11851 2559
rect 11517 2485 11851 2525
rect 11897 2655 11963 2660
rect 11897 2635 11913 2655
rect 11947 2621 11963 2655
rect 11931 2601 11963 2621
rect 11897 2587 11963 2601
rect 11897 2553 11913 2587
rect 11947 2553 11963 2587
rect 11897 2519 11963 2553
rect 11897 2491 11913 2519
rect 10780 2425 10955 2441
rect 10780 2391 10921 2425
rect 10780 2375 10955 2391
rect 10989 2425 11139 2441
rect 10989 2391 11105 2425
rect 10989 2375 11139 2391
rect 10780 2283 10814 2375
rect 10989 2341 11029 2375
rect 11173 2349 11207 2465
rect 11162 2341 11207 2349
rect 10963 2338 11029 2341
rect 10963 2304 10979 2338
rect 11013 2304 11029 2338
rect 11131 2340 11207 2341
rect 10542 2249 10573 2283
rect 10607 2249 10623 2283
rect 10657 2249 10676 2283
rect 10710 2249 10814 2283
rect 10869 2283 10911 2299
rect 10869 2249 10874 2283
rect 10908 2249 10911 2283
rect 10432 2193 10506 2243
rect 10869 2193 10911 2249
rect 10963 2270 11029 2304
rect 10963 2236 10979 2270
rect 11013 2236 11029 2270
rect 11063 2299 11097 2315
rect 11063 2193 11097 2265
rect 11131 2306 11147 2340
rect 11181 2324 11207 2340
rect 11517 2417 11537 2451
rect 11571 2417 11667 2451
rect 11517 2347 11667 2417
rect 11701 2415 11851 2485
rect 11701 2381 11797 2415
rect 11831 2381 11851 2415
rect 11885 2485 11913 2491
rect 11947 2485 11963 2519
rect 11997 2631 12031 2703
rect 11997 2551 12031 2597
rect 11997 2501 12031 2517
rect 12065 2661 12133 2669
rect 12065 2627 12083 2661
rect 12117 2627 12133 2661
rect 12065 2590 12133 2627
rect 12179 2653 12242 2703
rect 12179 2619 12206 2653
rect 12240 2619 12242 2653
rect 12500 2653 12550 2669
rect 12179 2603 12242 2619
rect 12278 2609 12405 2643
rect 12439 2609 12455 2643
rect 12534 2619 12550 2653
rect 12065 2556 12083 2590
rect 12117 2557 12133 2590
rect 12117 2556 12244 2557
rect 12065 2541 12244 2556
rect 12065 2519 12210 2541
rect 11885 2475 11963 2485
rect 12065 2485 12083 2519
rect 12117 2507 12210 2519
rect 12117 2485 12244 2507
rect 12065 2482 12244 2485
rect 11885 2465 11928 2475
rect 11885 2349 11919 2465
rect 12065 2441 12103 2482
rect 12278 2441 12312 2609
rect 12500 2603 12550 2619
rect 11953 2425 12103 2441
rect 11987 2391 12103 2425
rect 11953 2375 12103 2391
rect 12137 2425 12312 2441
rect 12171 2391 12312 2425
rect 12137 2375 12312 2391
rect 11181 2306 11197 2324
rect 11131 2272 11197 2306
rect 11131 2238 11147 2272
rect 11181 2238 11197 2272
rect 11131 2237 11197 2238
rect 11425 2321 11483 2338
rect 11425 2287 11437 2321
rect 11471 2287 11483 2321
rect 11425 2193 11483 2287
rect 11517 2295 11851 2347
rect 11885 2341 11930 2349
rect 12063 2341 12103 2375
rect 11885 2340 11961 2341
rect 11885 2324 11911 2340
rect 11517 2261 11535 2295
rect 11569 2261 11799 2295
rect 11833 2261 11851 2295
rect 11517 2193 11851 2261
rect 11895 2306 11911 2324
rect 11945 2306 11961 2340
rect 12063 2338 12129 2341
rect 11895 2272 11961 2306
rect 11895 2238 11911 2272
rect 11945 2238 11961 2272
rect 11895 2237 11961 2238
rect 11995 2299 12029 2315
rect 11995 2193 12029 2265
rect 12063 2304 12079 2338
rect 12113 2304 12129 2338
rect 12063 2270 12129 2304
rect 12063 2236 12079 2270
rect 12113 2236 12129 2270
rect 12181 2283 12223 2299
rect 12181 2249 12184 2283
rect 12218 2249 12223 2283
rect 12278 2283 12312 2375
rect 12346 2541 12410 2575
rect 12380 2507 12410 2541
rect 12346 2499 12410 2507
rect 12346 2465 12359 2499
rect 12393 2465 12410 2499
rect 12346 2383 12410 2465
rect 12444 2567 12482 2569
rect 12444 2533 12446 2567
rect 12480 2533 12482 2567
rect 12444 2475 12482 2533
rect 12444 2441 12448 2475
rect 12444 2425 12482 2441
rect 12516 2389 12550 2603
rect 12584 2661 12618 2703
rect 12915 2653 12965 2669
rect 12584 2593 12618 2627
rect 12584 2543 12618 2559
rect 12652 2614 12823 2648
rect 12857 2614 12873 2648
rect 12949 2619 12965 2653
rect 12652 2491 12686 2614
rect 12915 2584 12965 2619
rect 12999 2661 13052 2703
rect 13033 2627 13052 2661
rect 12999 2611 13052 2627
rect 13100 2653 13137 2669
rect 13100 2619 13103 2653
rect 13100 2585 13137 2619
rect 13171 2637 13237 2703
rect 13171 2603 13187 2637
rect 13221 2603 13237 2637
rect 13271 2653 13305 2669
rect 12720 2567 12826 2580
rect 12720 2541 12760 2567
rect 12720 2507 12758 2541
rect 12794 2533 12826 2567
rect 12915 2558 12976 2584
rect 12584 2475 12686 2491
rect 12618 2473 12686 2475
rect 12618 2441 12758 2473
rect 12584 2439 12758 2441
rect 12584 2425 12618 2439
rect 12642 2389 12682 2395
rect 12346 2367 12439 2383
rect 12346 2333 12405 2367
rect 12346 2317 12439 2333
rect 12516 2379 12682 2389
rect 12516 2345 12648 2379
rect 12516 2329 12682 2345
rect 12516 2283 12550 2329
rect 12278 2249 12382 2283
rect 12416 2249 12435 2283
rect 12469 2249 12485 2283
rect 12519 2249 12550 2283
rect 12586 2277 12660 2293
rect 12181 2193 12223 2249
rect 12586 2243 12604 2277
rect 12638 2243 12660 2277
rect 12724 2283 12758 2439
rect 12792 2367 12826 2533
rect 12860 2499 12908 2520
rect 12860 2465 12863 2499
rect 12897 2465 12908 2499
rect 12860 2463 12908 2465
rect 12860 2429 12867 2463
rect 12901 2429 12908 2463
rect 12860 2401 12908 2429
rect 12792 2333 12847 2367
rect 12881 2333 12897 2367
rect 12942 2337 12976 2558
rect 13100 2551 13103 2585
rect 13271 2585 13305 2619
rect 12792 2323 12897 2333
rect 12931 2311 12976 2337
rect 13010 2493 13066 2509
rect 13044 2459 13066 2493
rect 13010 2363 13066 2459
rect 13010 2329 13032 2363
rect 13010 2319 13066 2329
rect 13100 2499 13137 2551
rect 13100 2465 13101 2499
rect 13135 2465 13137 2499
rect 12931 2283 12965 2311
rect 13100 2295 13137 2465
rect 13172 2567 13271 2569
rect 13172 2533 13180 2567
rect 13214 2551 13271 2567
rect 13214 2535 13305 2551
rect 13357 2661 13875 2703
rect 13357 2627 13375 2661
rect 13409 2627 13823 2661
rect 13857 2627 13875 2661
rect 13357 2559 13875 2627
rect 13214 2533 13218 2535
rect 13172 2440 13218 2533
rect 13357 2525 13375 2559
rect 13409 2525 13823 2559
rect 13857 2525 13875 2559
rect 13206 2406 13218 2440
rect 13172 2337 13218 2406
rect 13252 2431 13322 2501
rect 13357 2485 13875 2525
rect 13252 2425 13277 2431
rect 13252 2391 13274 2425
rect 13311 2397 13322 2431
rect 13308 2391 13322 2397
rect 13252 2371 13322 2391
rect 13357 2417 13435 2451
rect 13469 2417 13545 2451
rect 13579 2417 13599 2451
rect 13357 2347 13599 2417
rect 13633 2415 13875 2485
rect 14001 2632 14059 2703
rect 14001 2598 14013 2632
rect 14047 2598 14059 2632
rect 14001 2539 14059 2598
rect 14001 2505 14013 2539
rect 14047 2505 14059 2539
rect 14001 2470 14059 2505
rect 14277 2660 14381 2669
rect 14277 2635 14331 2660
rect 14277 2601 14289 2635
rect 14323 2626 14331 2635
rect 14365 2626 14381 2660
rect 14323 2601 14381 2626
rect 14277 2592 14381 2601
rect 14277 2558 14331 2592
rect 14365 2558 14381 2592
rect 14415 2660 14481 2703
rect 14415 2626 14431 2660
rect 14465 2626 14481 2660
rect 14415 2592 14481 2626
rect 14553 2661 15622 2703
rect 14553 2627 14571 2661
rect 14605 2627 15571 2661
rect 15605 2627 15622 2661
rect 14553 2616 15622 2627
rect 15657 2661 16359 2703
rect 15657 2627 15675 2661
rect 15709 2627 16307 2661
rect 16341 2627 16359 2661
rect 14415 2558 14431 2592
rect 14465 2558 14481 2592
rect 13633 2381 13653 2415
rect 13687 2381 13763 2415
rect 13797 2381 13875 2415
rect 14277 2359 14381 2558
rect 13172 2303 13305 2337
rect 12724 2249 12803 2283
rect 12837 2249 12859 2283
rect 12898 2249 12914 2283
rect 12948 2249 12965 2283
rect 12999 2269 13049 2285
rect 12586 2193 12660 2243
rect 13033 2235 13049 2269
rect 13100 2261 13103 2295
rect 13271 2295 13305 2303
rect 13100 2245 13137 2261
rect 12999 2193 13049 2235
rect 13171 2235 13187 2269
rect 13221 2235 13237 2269
rect 13271 2245 13305 2261
rect 13357 2288 13875 2347
rect 13357 2254 13375 2288
rect 13409 2254 13823 2288
rect 13857 2254 13875 2288
rect 13171 2193 13237 2235
rect 13357 2193 13875 2254
rect 14001 2321 14059 2338
rect 14415 2329 14519 2524
rect 14001 2287 14013 2321
rect 14047 2287 14059 2321
rect 14001 2193 14059 2287
rect 14313 2291 14331 2325
rect 14365 2291 14381 2325
rect 14313 2257 14381 2291
rect 14313 2223 14331 2257
rect 14365 2223 14381 2257
rect 14415 2295 14431 2329
rect 14465 2295 14519 2329
rect 14870 2451 14938 2468
rect 14870 2417 14887 2451
rect 14921 2417 14938 2451
rect 14870 2302 14938 2417
rect 15234 2415 15304 2616
rect 15657 2559 16359 2627
rect 15657 2525 15675 2559
rect 15709 2525 16307 2559
rect 16341 2525 16359 2559
rect 15657 2485 16359 2525
rect 15234 2381 15251 2415
rect 15285 2381 15304 2415
rect 15234 2366 15304 2381
rect 15657 2417 15735 2451
rect 15769 2417 15834 2451
rect 15868 2417 15933 2451
rect 15967 2417 15987 2451
rect 15657 2347 15987 2417
rect 16021 2415 16359 2485
rect 16577 2632 16635 2703
rect 16577 2598 16589 2632
rect 16623 2598 16635 2632
rect 16577 2539 16635 2598
rect 16577 2505 16589 2539
rect 16623 2505 16635 2539
rect 16577 2470 16635 2505
rect 16853 2653 16907 2669
rect 16853 2635 16871 2653
rect 16853 2601 16865 2635
rect 16905 2619 16907 2653
rect 16899 2601 16907 2619
rect 16853 2572 16907 2601
rect 16853 2538 16871 2572
rect 16905 2538 16907 2572
rect 16941 2653 17007 2703
rect 16941 2619 16957 2653
rect 16991 2619 17007 2653
rect 16941 2585 17007 2619
rect 16941 2551 16957 2585
rect 16991 2551 17007 2585
rect 17043 2653 17077 2669
rect 17043 2585 17077 2619
rect 16853 2488 16907 2538
rect 17043 2517 17077 2551
rect 16021 2381 16041 2415
rect 16075 2381 16144 2415
rect 16178 2381 16247 2415
rect 16281 2381 16359 2415
rect 14415 2261 14519 2295
rect 14415 2227 14431 2261
rect 14465 2227 14519 2261
rect 14553 2288 15622 2302
rect 14553 2254 14571 2288
rect 14605 2254 15571 2288
rect 15605 2254 15622 2288
rect 14313 2193 14381 2223
rect 14553 2193 15622 2254
rect 15657 2288 16359 2347
rect 15657 2254 15675 2288
rect 15709 2254 16307 2288
rect 16341 2254 16359 2288
rect 15657 2193 16359 2254
rect 16577 2321 16635 2338
rect 16577 2287 16589 2321
rect 16623 2287 16635 2321
rect 16577 2193 16635 2287
rect 16853 2328 16887 2488
rect 16944 2483 17077 2517
rect 17129 2661 17463 2703
rect 17129 2627 17147 2661
rect 17181 2627 17411 2661
rect 17445 2627 17463 2661
rect 17129 2559 17463 2627
rect 17129 2525 17147 2559
rect 17181 2525 17411 2559
rect 17445 2525 17463 2559
rect 17129 2485 17463 2525
rect 16944 2454 16978 2483
rect 16921 2438 16978 2454
rect 16955 2404 16978 2438
rect 16921 2388 16978 2404
rect 16944 2337 16978 2388
rect 17025 2431 17091 2447
rect 17025 2425 17049 2431
rect 17025 2391 17041 2425
rect 17083 2397 17091 2431
rect 17075 2391 17091 2397
rect 17025 2373 17091 2391
rect 17129 2417 17149 2451
rect 17183 2417 17279 2451
rect 17129 2347 17279 2417
rect 17313 2415 17463 2485
rect 17515 2653 17549 2669
rect 17515 2585 17549 2619
rect 17592 2653 17658 2703
rect 17592 2619 17608 2653
rect 17642 2619 17658 2653
rect 17592 2585 17658 2619
rect 17592 2551 17608 2585
rect 17642 2551 17658 2585
rect 17692 2637 17743 2669
rect 17692 2603 17694 2637
rect 17728 2603 17743 2637
rect 17692 2556 17743 2603
rect 17515 2517 17549 2551
rect 17692 2522 17694 2556
rect 17728 2522 17743 2556
rect 17515 2483 17658 2517
rect 17692 2488 17743 2522
rect 17313 2381 17409 2415
rect 17443 2381 17463 2415
rect 17497 2431 17568 2447
rect 17497 2397 17509 2431
rect 17543 2425 17568 2431
rect 17497 2391 17517 2397
rect 17551 2391 17568 2425
rect 17497 2373 17568 2391
rect 17624 2441 17658 2483
rect 17624 2425 17675 2441
rect 17624 2391 17641 2425
rect 17624 2375 17675 2391
rect 16853 2299 16905 2328
rect 16944 2303 17077 2337
rect 16853 2265 16871 2299
rect 17043 2282 17077 2303
rect 16853 2227 16905 2265
rect 16941 2235 16957 2269
rect 16991 2235 17007 2269
rect 16941 2193 17007 2235
rect 17043 2227 17077 2248
rect 17129 2295 17463 2347
rect 17624 2337 17658 2375
rect 17709 2342 17743 2488
rect 17778 2661 17830 2703
rect 17812 2627 17830 2661
rect 17778 2593 17830 2627
rect 17812 2559 17830 2593
rect 17778 2525 17830 2559
rect 17812 2491 17830 2525
rect 17778 2473 17830 2491
rect 17865 2661 18567 2703
rect 17865 2627 17883 2661
rect 17917 2627 18515 2661
rect 18549 2627 18567 2661
rect 17865 2559 18567 2627
rect 17865 2525 17883 2559
rect 17917 2525 18515 2559
rect 18549 2525 18567 2559
rect 17865 2485 18567 2525
rect 17865 2417 17943 2451
rect 17977 2417 18042 2451
rect 18076 2417 18141 2451
rect 18175 2417 18195 2451
rect 17129 2261 17147 2295
rect 17181 2261 17411 2295
rect 17445 2261 17463 2295
rect 17129 2193 17463 2261
rect 17515 2303 17658 2337
rect 17515 2282 17549 2303
rect 17692 2299 17743 2342
rect 17692 2295 17694 2299
rect 17515 2227 17549 2248
rect 17592 2235 17608 2269
rect 17642 2235 17658 2269
rect 17592 2193 17658 2235
rect 17692 2261 17693 2295
rect 17728 2265 17743 2299
rect 17727 2261 17743 2265
rect 17692 2227 17743 2261
rect 17778 2341 17830 2361
rect 17812 2307 17830 2341
rect 17778 2273 17830 2307
rect 17812 2239 17830 2273
rect 17778 2193 17830 2239
rect 17865 2347 18195 2417
rect 18229 2415 18567 2485
rect 18229 2381 18249 2415
rect 18283 2381 18352 2415
rect 18386 2381 18455 2415
rect 18489 2381 18567 2415
rect 18601 2661 18843 2703
rect 18601 2627 18619 2661
rect 18653 2627 18791 2661
rect 18825 2627 18843 2661
rect 18601 2566 18843 2627
rect 18601 2532 18619 2566
rect 18653 2532 18791 2566
rect 18825 2532 18843 2566
rect 18601 2485 18843 2532
rect 18601 2411 18705 2485
rect 18601 2377 18651 2411
rect 18685 2377 18705 2411
rect 18739 2417 18759 2451
rect 18793 2417 18843 2451
rect 17865 2288 18567 2347
rect 18739 2343 18843 2417
rect 17865 2254 17883 2288
rect 17917 2254 18515 2288
rect 18549 2254 18567 2288
rect 17865 2193 18567 2254
rect 18601 2290 18843 2343
rect 18601 2256 18619 2290
rect 18653 2256 18791 2290
rect 18825 2256 18843 2290
rect 18601 2193 18843 2256
rect 1104 2159 1133 2193
rect 1167 2159 1225 2193
rect 1259 2159 1317 2193
rect 1351 2159 1409 2193
rect 1443 2159 1501 2193
rect 1535 2159 1593 2193
rect 1627 2159 1685 2193
rect 1719 2159 1777 2193
rect 1811 2159 1869 2193
rect 1903 2159 1961 2193
rect 1995 2159 2053 2193
rect 2087 2159 2145 2193
rect 2179 2159 2237 2193
rect 2271 2159 2329 2193
rect 2363 2159 2421 2193
rect 2455 2159 2513 2193
rect 2547 2159 2605 2193
rect 2639 2159 2697 2193
rect 2731 2159 2789 2193
rect 2823 2159 2881 2193
rect 2915 2159 2973 2193
rect 3007 2159 3065 2193
rect 3099 2159 3157 2193
rect 3191 2159 3249 2193
rect 3283 2159 3341 2193
rect 3375 2159 3433 2193
rect 3467 2159 3525 2193
rect 3559 2159 3617 2193
rect 3651 2159 3709 2193
rect 3743 2159 3801 2193
rect 3835 2159 3893 2193
rect 3927 2159 3985 2193
rect 4019 2159 4077 2193
rect 4111 2159 4169 2193
rect 4203 2159 4261 2193
rect 4295 2159 4353 2193
rect 4387 2159 4445 2193
rect 4479 2159 4537 2193
rect 4571 2159 4629 2193
rect 4663 2159 4721 2193
rect 4755 2159 4813 2193
rect 4847 2159 4905 2193
rect 4939 2159 4997 2193
rect 5031 2159 5089 2193
rect 5123 2159 5181 2193
rect 5215 2159 5273 2193
rect 5307 2159 5365 2193
rect 5399 2159 5457 2193
rect 5491 2159 5549 2193
rect 5583 2159 5641 2193
rect 5675 2159 5733 2193
rect 5767 2159 5825 2193
rect 5859 2159 5917 2193
rect 5951 2159 6009 2193
rect 6043 2159 6101 2193
rect 6135 2159 6193 2193
rect 6227 2159 6285 2193
rect 6319 2159 6377 2193
rect 6411 2159 6469 2193
rect 6503 2159 6561 2193
rect 6595 2159 6653 2193
rect 6687 2159 6745 2193
rect 6779 2159 6837 2193
rect 6871 2159 6929 2193
rect 6963 2159 7021 2193
rect 7055 2159 7113 2193
rect 7147 2159 7205 2193
rect 7239 2159 7297 2193
rect 7331 2159 7389 2193
rect 7423 2159 7481 2193
rect 7515 2159 7573 2193
rect 7607 2159 7665 2193
rect 7699 2159 7757 2193
rect 7791 2159 7849 2193
rect 7883 2159 7941 2193
rect 7975 2159 8033 2193
rect 8067 2159 8125 2193
rect 8159 2159 8217 2193
rect 8251 2159 8309 2193
rect 8343 2159 8401 2193
rect 8435 2159 8493 2193
rect 8527 2159 8585 2193
rect 8619 2159 8677 2193
rect 8711 2159 8769 2193
rect 8803 2159 8861 2193
rect 8895 2159 8953 2193
rect 8987 2159 9045 2193
rect 9079 2159 9137 2193
rect 9171 2159 9229 2193
rect 9263 2159 9321 2193
rect 9355 2159 9413 2193
rect 9447 2159 9505 2193
rect 9539 2159 9597 2193
rect 9631 2159 9689 2193
rect 9723 2159 9781 2193
rect 9815 2159 9873 2193
rect 9907 2159 9965 2193
rect 9999 2159 10057 2193
rect 10091 2159 10149 2193
rect 10183 2159 10241 2193
rect 10275 2159 10333 2193
rect 10367 2159 10425 2193
rect 10459 2159 10517 2193
rect 10551 2159 10609 2193
rect 10643 2159 10701 2193
rect 10735 2159 10793 2193
rect 10827 2159 10885 2193
rect 10919 2159 10977 2193
rect 11011 2159 11069 2193
rect 11103 2159 11161 2193
rect 11195 2159 11253 2193
rect 11287 2159 11345 2193
rect 11379 2159 11437 2193
rect 11471 2159 11529 2193
rect 11563 2159 11621 2193
rect 11655 2159 11713 2193
rect 11747 2159 11805 2193
rect 11839 2159 11897 2193
rect 11931 2159 11989 2193
rect 12023 2159 12081 2193
rect 12115 2159 12173 2193
rect 12207 2159 12265 2193
rect 12299 2159 12357 2193
rect 12391 2159 12449 2193
rect 12483 2159 12541 2193
rect 12575 2159 12633 2193
rect 12667 2159 12725 2193
rect 12759 2159 12817 2193
rect 12851 2159 12909 2193
rect 12943 2159 13001 2193
rect 13035 2159 13093 2193
rect 13127 2159 13185 2193
rect 13219 2159 13277 2193
rect 13311 2159 13369 2193
rect 13403 2159 13461 2193
rect 13495 2159 13553 2193
rect 13587 2159 13645 2193
rect 13679 2159 13737 2193
rect 13771 2159 13829 2193
rect 13863 2159 13921 2193
rect 13955 2159 14013 2193
rect 14047 2159 14105 2193
rect 14139 2159 14197 2193
rect 14231 2159 14289 2193
rect 14323 2159 14381 2193
rect 14415 2159 14473 2193
rect 14507 2159 14565 2193
rect 14599 2159 14657 2193
rect 14691 2159 14749 2193
rect 14783 2159 14841 2193
rect 14875 2159 14933 2193
rect 14967 2159 15025 2193
rect 15059 2159 15117 2193
rect 15151 2159 15209 2193
rect 15243 2159 15301 2193
rect 15335 2159 15393 2193
rect 15427 2159 15485 2193
rect 15519 2159 15577 2193
rect 15611 2159 15669 2193
rect 15703 2159 15761 2193
rect 15795 2159 15853 2193
rect 15887 2159 15945 2193
rect 15979 2159 16037 2193
rect 16071 2159 16129 2193
rect 16163 2159 16221 2193
rect 16255 2159 16313 2193
rect 16347 2159 16405 2193
rect 16439 2159 16497 2193
rect 16531 2159 16589 2193
rect 16623 2159 16681 2193
rect 16715 2159 16773 2193
rect 16807 2159 16865 2193
rect 16899 2159 16957 2193
rect 16991 2159 17049 2193
rect 17083 2159 17141 2193
rect 17175 2159 17233 2193
rect 17267 2159 17325 2193
rect 17359 2159 17417 2193
rect 17451 2159 17509 2193
rect 17543 2159 17601 2193
rect 17635 2159 17693 2193
rect 17727 2159 17785 2193
rect 17819 2159 17877 2193
rect 17911 2159 17969 2193
rect 18003 2159 18061 2193
rect 18095 2159 18153 2193
rect 18187 2159 18245 2193
rect 18279 2159 18337 2193
rect 18371 2159 18429 2193
rect 18463 2159 18521 2193
rect 18555 2159 18613 2193
rect 18647 2159 18705 2193
rect 18739 2159 18797 2193
rect 18831 2159 18860 2193
<< viali >>
rect 1133 7599 1167 7633
rect 1225 7599 1259 7633
rect 1317 7599 1351 7633
rect 1409 7599 1443 7633
rect 1501 7599 1535 7633
rect 1593 7599 1627 7633
rect 1685 7599 1719 7633
rect 1777 7599 1811 7633
rect 1869 7599 1903 7633
rect 1961 7599 1995 7633
rect 2053 7599 2087 7633
rect 2145 7599 2179 7633
rect 2237 7599 2271 7633
rect 2329 7599 2363 7633
rect 2421 7599 2455 7633
rect 2513 7599 2547 7633
rect 2605 7599 2639 7633
rect 2697 7599 2731 7633
rect 2789 7599 2823 7633
rect 2881 7599 2915 7633
rect 2973 7599 3007 7633
rect 3065 7599 3099 7633
rect 3157 7599 3191 7633
rect 3249 7599 3283 7633
rect 3341 7599 3375 7633
rect 3433 7599 3467 7633
rect 3525 7599 3559 7633
rect 3617 7599 3651 7633
rect 3709 7599 3743 7633
rect 3801 7599 3835 7633
rect 3893 7599 3927 7633
rect 3985 7599 4019 7633
rect 4077 7599 4111 7633
rect 4169 7599 4203 7633
rect 4261 7599 4295 7633
rect 4353 7599 4387 7633
rect 4445 7599 4479 7633
rect 4537 7599 4571 7633
rect 4629 7599 4663 7633
rect 4721 7599 4755 7633
rect 4813 7599 4847 7633
rect 4905 7599 4939 7633
rect 4997 7599 5031 7633
rect 5089 7599 5123 7633
rect 5181 7599 5215 7633
rect 5273 7599 5307 7633
rect 5365 7599 5399 7633
rect 5457 7599 5491 7633
rect 5549 7599 5583 7633
rect 5641 7599 5675 7633
rect 5733 7599 5767 7633
rect 5825 7599 5859 7633
rect 5917 7599 5951 7633
rect 6009 7599 6043 7633
rect 6101 7599 6135 7633
rect 6193 7599 6227 7633
rect 6285 7599 6319 7633
rect 6377 7599 6411 7633
rect 6469 7599 6503 7633
rect 6561 7599 6595 7633
rect 6653 7599 6687 7633
rect 6745 7599 6779 7633
rect 6837 7599 6871 7633
rect 6929 7599 6963 7633
rect 7021 7599 7055 7633
rect 7113 7599 7147 7633
rect 7205 7599 7239 7633
rect 7297 7599 7331 7633
rect 7389 7599 7423 7633
rect 7481 7599 7515 7633
rect 7573 7599 7607 7633
rect 7665 7599 7699 7633
rect 7757 7599 7791 7633
rect 7849 7599 7883 7633
rect 7941 7599 7975 7633
rect 8033 7599 8067 7633
rect 8125 7599 8159 7633
rect 8217 7599 8251 7633
rect 8309 7599 8343 7633
rect 8401 7599 8435 7633
rect 8493 7599 8527 7633
rect 8585 7599 8619 7633
rect 8677 7599 8711 7633
rect 8769 7599 8803 7633
rect 8861 7599 8895 7633
rect 8953 7599 8987 7633
rect 9045 7599 9079 7633
rect 9137 7599 9171 7633
rect 9229 7599 9263 7633
rect 9321 7599 9355 7633
rect 9413 7599 9447 7633
rect 9505 7599 9539 7633
rect 9597 7599 9631 7633
rect 9689 7599 9723 7633
rect 9781 7599 9815 7633
rect 9873 7599 9907 7633
rect 9965 7599 9999 7633
rect 10057 7599 10091 7633
rect 10149 7599 10183 7633
rect 10241 7599 10275 7633
rect 10333 7599 10367 7633
rect 10425 7599 10459 7633
rect 10517 7599 10551 7633
rect 10609 7599 10643 7633
rect 10701 7599 10735 7633
rect 10793 7599 10827 7633
rect 10885 7599 10919 7633
rect 10977 7599 11011 7633
rect 11069 7599 11103 7633
rect 11161 7599 11195 7633
rect 11253 7599 11287 7633
rect 11345 7599 11379 7633
rect 11437 7599 11471 7633
rect 11529 7599 11563 7633
rect 11621 7599 11655 7633
rect 11713 7599 11747 7633
rect 11805 7599 11839 7633
rect 11897 7599 11931 7633
rect 11989 7599 12023 7633
rect 12081 7599 12115 7633
rect 12173 7599 12207 7633
rect 12265 7599 12299 7633
rect 12357 7599 12391 7633
rect 12449 7599 12483 7633
rect 12541 7599 12575 7633
rect 12633 7599 12667 7633
rect 12725 7599 12759 7633
rect 12817 7599 12851 7633
rect 12909 7599 12943 7633
rect 13001 7599 13035 7633
rect 13093 7599 13127 7633
rect 13185 7599 13219 7633
rect 13277 7599 13311 7633
rect 13369 7599 13403 7633
rect 13461 7599 13495 7633
rect 13553 7599 13587 7633
rect 13645 7599 13679 7633
rect 13737 7599 13771 7633
rect 13829 7599 13863 7633
rect 13921 7599 13955 7633
rect 14013 7599 14047 7633
rect 14105 7599 14139 7633
rect 14197 7599 14231 7633
rect 14289 7599 14323 7633
rect 14381 7599 14415 7633
rect 14473 7599 14507 7633
rect 14565 7599 14599 7633
rect 14657 7599 14691 7633
rect 14749 7599 14783 7633
rect 14841 7599 14875 7633
rect 14933 7599 14967 7633
rect 15025 7599 15059 7633
rect 15117 7599 15151 7633
rect 15209 7599 15243 7633
rect 15301 7599 15335 7633
rect 15393 7599 15427 7633
rect 15485 7599 15519 7633
rect 15577 7599 15611 7633
rect 15669 7599 15703 7633
rect 15761 7599 15795 7633
rect 15853 7599 15887 7633
rect 15945 7599 15979 7633
rect 16037 7599 16071 7633
rect 16129 7599 16163 7633
rect 16221 7599 16255 7633
rect 16313 7599 16347 7633
rect 16405 7599 16439 7633
rect 16497 7599 16531 7633
rect 16589 7599 16623 7633
rect 16681 7599 16715 7633
rect 16773 7599 16807 7633
rect 16865 7599 16899 7633
rect 16957 7599 16991 7633
rect 17049 7599 17083 7633
rect 17141 7599 17175 7633
rect 17233 7599 17267 7633
rect 17325 7599 17359 7633
rect 17417 7599 17451 7633
rect 17509 7599 17543 7633
rect 17601 7599 17635 7633
rect 17693 7599 17727 7633
rect 17785 7599 17819 7633
rect 17877 7599 17911 7633
rect 17969 7599 18003 7633
rect 18061 7599 18095 7633
rect 18153 7599 18187 7633
rect 18245 7599 18279 7633
rect 18337 7599 18371 7633
rect 18429 7599 18463 7633
rect 18521 7599 18555 7633
rect 18613 7599 18647 7633
rect 18705 7599 18739 7633
rect 18797 7599 18831 7633
rect 1685 7527 1719 7531
rect 1685 7497 1718 7527
rect 1718 7497 1719 7527
rect 1869 7367 1895 7395
rect 1895 7367 1903 7395
rect 1869 7361 1903 7367
rect 4077 7527 4111 7531
rect 4077 7497 4110 7527
rect 4110 7497 4111 7527
rect 4261 7367 4287 7395
rect 4287 7367 4295 7395
rect 4261 7361 4295 7367
rect 5733 7527 5767 7531
rect 5733 7497 5766 7527
rect 5766 7497 5767 7527
rect 5917 7367 5943 7395
rect 5943 7367 5951 7395
rect 5917 7361 5951 7367
rect 8033 7527 8067 7531
rect 8033 7497 8034 7527
rect 8034 7497 8067 7527
rect 7849 7367 7857 7395
rect 7857 7367 7883 7395
rect 7849 7361 7883 7367
rect 9597 7457 9620 7463
rect 9620 7457 9631 7463
rect 9597 7429 9631 7457
rect 10149 7429 10183 7463
rect 12449 7527 12483 7531
rect 12449 7497 12450 7527
rect 12450 7497 12483 7527
rect 10333 7225 10367 7259
rect 12265 7367 12273 7395
rect 12273 7367 12299 7395
rect 12265 7361 12299 7367
rect 14657 7527 14691 7531
rect 14657 7497 14658 7527
rect 14658 7497 14691 7527
rect 14473 7367 14481 7395
rect 14481 7367 14507 7395
rect 14473 7361 14507 7367
rect 17049 7527 17083 7531
rect 17049 7497 17050 7527
rect 17050 7497 17083 7527
rect 16865 7367 16873 7395
rect 16873 7367 16899 7395
rect 16865 7361 16899 7367
rect 18245 7527 18279 7531
rect 18245 7497 18246 7527
rect 18246 7497 18279 7527
rect 18061 7367 18069 7395
rect 18069 7367 18095 7395
rect 18061 7361 18095 7367
rect 1133 7055 1167 7089
rect 1225 7055 1259 7089
rect 1317 7055 1351 7089
rect 1409 7055 1443 7089
rect 1501 7055 1535 7089
rect 1593 7055 1627 7089
rect 1685 7055 1719 7089
rect 1777 7055 1811 7089
rect 1869 7055 1903 7089
rect 1961 7055 1995 7089
rect 2053 7055 2087 7089
rect 2145 7055 2179 7089
rect 2237 7055 2271 7089
rect 2329 7055 2363 7089
rect 2421 7055 2455 7089
rect 2513 7055 2547 7089
rect 2605 7055 2639 7089
rect 2697 7055 2731 7089
rect 2789 7055 2823 7089
rect 2881 7055 2915 7089
rect 2973 7055 3007 7089
rect 3065 7055 3099 7089
rect 3157 7055 3191 7089
rect 3249 7055 3283 7089
rect 3341 7055 3375 7089
rect 3433 7055 3467 7089
rect 3525 7055 3559 7089
rect 3617 7055 3651 7089
rect 3709 7055 3743 7089
rect 3801 7055 3835 7089
rect 3893 7055 3927 7089
rect 3985 7055 4019 7089
rect 4077 7055 4111 7089
rect 4169 7055 4203 7089
rect 4261 7055 4295 7089
rect 4353 7055 4387 7089
rect 4445 7055 4479 7089
rect 4537 7055 4571 7089
rect 4629 7055 4663 7089
rect 4721 7055 4755 7089
rect 4813 7055 4847 7089
rect 4905 7055 4939 7089
rect 4997 7055 5031 7089
rect 5089 7055 5123 7089
rect 5181 7055 5215 7089
rect 5273 7055 5307 7089
rect 5365 7055 5399 7089
rect 5457 7055 5491 7089
rect 5549 7055 5583 7089
rect 5641 7055 5675 7089
rect 5733 7055 5767 7089
rect 5825 7055 5859 7089
rect 5917 7055 5951 7089
rect 6009 7055 6043 7089
rect 6101 7055 6135 7089
rect 6193 7055 6227 7089
rect 6285 7055 6319 7089
rect 6377 7055 6411 7089
rect 6469 7055 6503 7089
rect 6561 7055 6595 7089
rect 6653 7055 6687 7089
rect 6745 7055 6779 7089
rect 6837 7055 6871 7089
rect 6929 7055 6963 7089
rect 7021 7055 7055 7089
rect 7113 7055 7147 7089
rect 7205 7055 7239 7089
rect 7297 7055 7331 7089
rect 7389 7055 7423 7089
rect 7481 7055 7515 7089
rect 7573 7055 7607 7089
rect 7665 7055 7699 7089
rect 7757 7055 7791 7089
rect 7849 7055 7883 7089
rect 7941 7055 7975 7089
rect 8033 7055 8067 7089
rect 8125 7055 8159 7089
rect 8217 7055 8251 7089
rect 8309 7055 8343 7089
rect 8401 7055 8435 7089
rect 8493 7055 8527 7089
rect 8585 7055 8619 7089
rect 8677 7055 8711 7089
rect 8769 7055 8803 7089
rect 8861 7055 8895 7089
rect 8953 7055 8987 7089
rect 9045 7055 9079 7089
rect 9137 7055 9171 7089
rect 9229 7055 9263 7089
rect 9321 7055 9355 7089
rect 9413 7055 9447 7089
rect 9505 7055 9539 7089
rect 9597 7055 9631 7089
rect 9689 7055 9723 7089
rect 9781 7055 9815 7089
rect 9873 7055 9907 7089
rect 9965 7055 9999 7089
rect 10057 7055 10091 7089
rect 10149 7055 10183 7089
rect 10241 7055 10275 7089
rect 10333 7055 10367 7089
rect 10425 7055 10459 7089
rect 10517 7055 10551 7089
rect 10609 7055 10643 7089
rect 10701 7055 10735 7089
rect 10793 7055 10827 7089
rect 10885 7055 10919 7089
rect 10977 7055 11011 7089
rect 11069 7055 11103 7089
rect 11161 7055 11195 7089
rect 11253 7055 11287 7089
rect 11345 7055 11379 7089
rect 11437 7055 11471 7089
rect 11529 7055 11563 7089
rect 11621 7055 11655 7089
rect 11713 7055 11747 7089
rect 11805 7055 11839 7089
rect 11897 7055 11931 7089
rect 11989 7055 12023 7089
rect 12081 7055 12115 7089
rect 12173 7055 12207 7089
rect 12265 7055 12299 7089
rect 12357 7055 12391 7089
rect 12449 7055 12483 7089
rect 12541 7055 12575 7089
rect 12633 7055 12667 7089
rect 12725 7055 12759 7089
rect 12817 7055 12851 7089
rect 12909 7055 12943 7089
rect 13001 7055 13035 7089
rect 13093 7055 13127 7089
rect 13185 7055 13219 7089
rect 13277 7055 13311 7089
rect 13369 7055 13403 7089
rect 13461 7055 13495 7089
rect 13553 7055 13587 7089
rect 13645 7055 13679 7089
rect 13737 7055 13771 7089
rect 13829 7055 13863 7089
rect 13921 7055 13955 7089
rect 14013 7055 14047 7089
rect 14105 7055 14139 7089
rect 14197 7055 14231 7089
rect 14289 7055 14323 7089
rect 14381 7055 14415 7089
rect 14473 7055 14507 7089
rect 14565 7055 14599 7089
rect 14657 7055 14691 7089
rect 14749 7055 14783 7089
rect 14841 7055 14875 7089
rect 14933 7055 14967 7089
rect 15025 7055 15059 7089
rect 15117 7055 15151 7089
rect 15209 7055 15243 7089
rect 15301 7055 15335 7089
rect 15393 7055 15427 7089
rect 15485 7055 15519 7089
rect 15577 7055 15611 7089
rect 15669 7055 15703 7089
rect 15761 7055 15795 7089
rect 15853 7055 15887 7089
rect 15945 7055 15979 7089
rect 16037 7055 16071 7089
rect 16129 7055 16163 7089
rect 16221 7055 16255 7089
rect 16313 7055 16347 7089
rect 16405 7055 16439 7089
rect 16497 7055 16531 7089
rect 16589 7055 16623 7089
rect 16681 7055 16715 7089
rect 16773 7055 16807 7089
rect 16865 7055 16899 7089
rect 16957 7055 16991 7089
rect 17049 7055 17083 7089
rect 17141 7055 17175 7089
rect 17233 7055 17267 7089
rect 17325 7055 17359 7089
rect 17417 7055 17451 7089
rect 17509 7055 17543 7089
rect 17601 7055 17635 7089
rect 17693 7055 17727 7089
rect 17785 7055 17819 7089
rect 17877 7055 17911 7089
rect 17969 7055 18003 7089
rect 18061 7055 18095 7089
rect 18153 7055 18187 7089
rect 18245 7055 18279 7089
rect 18337 7055 18371 7089
rect 18429 7055 18463 7089
rect 18521 7055 18555 7089
rect 18613 7055 18647 7089
rect 18705 7055 18739 7089
rect 18797 7055 18831 7089
rect 1133 6511 1167 6545
rect 1225 6511 1259 6545
rect 1317 6511 1351 6545
rect 1409 6511 1443 6545
rect 1501 6511 1535 6545
rect 1593 6511 1627 6545
rect 1685 6511 1719 6545
rect 1777 6511 1811 6545
rect 1869 6511 1903 6545
rect 1961 6511 1995 6545
rect 2053 6511 2087 6545
rect 2145 6511 2179 6545
rect 2237 6511 2271 6545
rect 2329 6511 2363 6545
rect 2421 6511 2455 6545
rect 2513 6511 2547 6545
rect 2605 6511 2639 6545
rect 2697 6511 2731 6545
rect 2789 6511 2823 6545
rect 2881 6511 2915 6545
rect 2973 6511 3007 6545
rect 3065 6511 3099 6545
rect 3157 6511 3191 6545
rect 3249 6511 3283 6545
rect 3341 6511 3375 6545
rect 3433 6511 3467 6545
rect 3525 6511 3559 6545
rect 3617 6511 3651 6545
rect 3709 6511 3743 6545
rect 3801 6511 3835 6545
rect 3893 6511 3927 6545
rect 3985 6511 4019 6545
rect 4077 6511 4111 6545
rect 4169 6511 4203 6545
rect 4261 6511 4295 6545
rect 4353 6511 4387 6545
rect 4445 6511 4479 6545
rect 4537 6511 4571 6545
rect 4629 6511 4663 6545
rect 4721 6511 4755 6545
rect 4813 6511 4847 6545
rect 4905 6511 4939 6545
rect 4997 6511 5031 6545
rect 5089 6511 5123 6545
rect 5181 6511 5215 6545
rect 5273 6511 5307 6545
rect 5365 6511 5399 6545
rect 5457 6511 5491 6545
rect 5549 6511 5583 6545
rect 5641 6511 5675 6545
rect 5733 6511 5767 6545
rect 5825 6511 5859 6545
rect 5917 6511 5951 6545
rect 6009 6511 6043 6545
rect 6101 6511 6135 6545
rect 6193 6511 6227 6545
rect 6285 6511 6319 6545
rect 6377 6511 6411 6545
rect 6469 6511 6503 6545
rect 6561 6511 6595 6545
rect 6653 6511 6687 6545
rect 6745 6511 6779 6545
rect 6837 6511 6871 6545
rect 6929 6511 6963 6545
rect 7021 6511 7055 6545
rect 7113 6511 7147 6545
rect 7205 6511 7239 6545
rect 7297 6511 7331 6545
rect 7389 6511 7423 6545
rect 7481 6511 7515 6545
rect 7573 6511 7607 6545
rect 7665 6511 7699 6545
rect 7757 6511 7791 6545
rect 7849 6511 7883 6545
rect 7941 6511 7975 6545
rect 8033 6511 8067 6545
rect 8125 6511 8159 6545
rect 8217 6511 8251 6545
rect 8309 6511 8343 6545
rect 8401 6511 8435 6545
rect 8493 6511 8527 6545
rect 8585 6511 8619 6545
rect 8677 6511 8711 6545
rect 8769 6511 8803 6545
rect 8861 6511 8895 6545
rect 8953 6511 8987 6545
rect 9045 6511 9079 6545
rect 9137 6511 9171 6545
rect 9229 6511 9263 6545
rect 9321 6511 9355 6545
rect 9413 6511 9447 6545
rect 9505 6511 9539 6545
rect 9597 6511 9631 6545
rect 9689 6511 9723 6545
rect 9781 6511 9815 6545
rect 9873 6511 9907 6545
rect 9965 6511 9999 6545
rect 10057 6511 10091 6545
rect 10149 6511 10183 6545
rect 10241 6511 10275 6545
rect 10333 6511 10367 6545
rect 10425 6511 10459 6545
rect 10517 6511 10551 6545
rect 10609 6511 10643 6545
rect 10701 6511 10735 6545
rect 10793 6511 10827 6545
rect 10885 6511 10919 6545
rect 10977 6511 11011 6545
rect 11069 6511 11103 6545
rect 11161 6511 11195 6545
rect 11253 6511 11287 6545
rect 11345 6511 11379 6545
rect 11437 6511 11471 6545
rect 11529 6511 11563 6545
rect 11621 6511 11655 6545
rect 11713 6511 11747 6545
rect 11805 6511 11839 6545
rect 11897 6511 11931 6545
rect 11989 6511 12023 6545
rect 12081 6511 12115 6545
rect 12173 6511 12207 6545
rect 12265 6511 12299 6545
rect 12357 6511 12391 6545
rect 12449 6511 12483 6545
rect 12541 6511 12575 6545
rect 12633 6511 12667 6545
rect 12725 6511 12759 6545
rect 12817 6511 12851 6545
rect 12909 6511 12943 6545
rect 13001 6511 13035 6545
rect 13093 6511 13127 6545
rect 13185 6511 13219 6545
rect 13277 6511 13311 6545
rect 13369 6511 13403 6545
rect 13461 6511 13495 6545
rect 13553 6511 13587 6545
rect 13645 6511 13679 6545
rect 13737 6511 13771 6545
rect 13829 6511 13863 6545
rect 13921 6511 13955 6545
rect 14013 6511 14047 6545
rect 14105 6511 14139 6545
rect 14197 6511 14231 6545
rect 14289 6511 14323 6545
rect 14381 6511 14415 6545
rect 14473 6511 14507 6545
rect 14565 6511 14599 6545
rect 14657 6511 14691 6545
rect 14749 6511 14783 6545
rect 14841 6511 14875 6545
rect 14933 6511 14967 6545
rect 15025 6511 15059 6545
rect 15117 6511 15151 6545
rect 15209 6511 15243 6545
rect 15301 6511 15335 6545
rect 15393 6511 15427 6545
rect 15485 6511 15519 6545
rect 15577 6511 15611 6545
rect 15669 6511 15703 6545
rect 15761 6511 15795 6545
rect 15853 6511 15887 6545
rect 15945 6511 15979 6545
rect 16037 6511 16071 6545
rect 16129 6511 16163 6545
rect 16221 6511 16255 6545
rect 16313 6511 16347 6545
rect 16405 6511 16439 6545
rect 16497 6511 16531 6545
rect 16589 6511 16623 6545
rect 16681 6511 16715 6545
rect 16773 6511 16807 6545
rect 16865 6511 16899 6545
rect 16957 6511 16991 6545
rect 17049 6511 17083 6545
rect 17141 6511 17175 6545
rect 17233 6511 17267 6545
rect 17325 6511 17359 6545
rect 17417 6511 17451 6545
rect 17509 6511 17543 6545
rect 17601 6511 17635 6545
rect 17693 6511 17727 6545
rect 17785 6511 17819 6545
rect 17877 6511 17911 6545
rect 17969 6511 18003 6545
rect 18061 6511 18095 6545
rect 18153 6511 18187 6545
rect 18245 6511 18279 6545
rect 18337 6511 18371 6545
rect 18429 6511 18463 6545
rect 18521 6511 18555 6545
rect 18613 6511 18647 6545
rect 18705 6511 18739 6545
rect 18797 6511 18831 6545
rect 1133 5967 1167 6001
rect 1225 5967 1259 6001
rect 1317 5967 1351 6001
rect 1409 5967 1443 6001
rect 1501 5967 1535 6001
rect 1593 5967 1627 6001
rect 1685 5967 1719 6001
rect 1777 5967 1811 6001
rect 1869 5967 1903 6001
rect 1961 5967 1995 6001
rect 2053 5967 2087 6001
rect 2145 5967 2179 6001
rect 2237 5967 2271 6001
rect 2329 5967 2363 6001
rect 2421 5967 2455 6001
rect 2513 5967 2547 6001
rect 2605 5967 2639 6001
rect 2697 5967 2731 6001
rect 2789 5967 2823 6001
rect 2881 5967 2915 6001
rect 2973 5967 3007 6001
rect 3065 5967 3099 6001
rect 3157 5967 3191 6001
rect 3249 5967 3283 6001
rect 3341 5967 3375 6001
rect 3433 5967 3467 6001
rect 3525 5967 3559 6001
rect 3617 5967 3651 6001
rect 3709 5967 3743 6001
rect 3801 5967 3835 6001
rect 3893 5967 3927 6001
rect 3985 5967 4019 6001
rect 4077 5967 4111 6001
rect 4169 5967 4203 6001
rect 4261 5967 4295 6001
rect 4353 5967 4387 6001
rect 4445 5967 4479 6001
rect 4537 5967 4571 6001
rect 4629 5967 4663 6001
rect 4721 5967 4755 6001
rect 4813 5967 4847 6001
rect 4905 5967 4939 6001
rect 4997 5967 5031 6001
rect 5089 5967 5123 6001
rect 5181 5967 5215 6001
rect 5273 5967 5307 6001
rect 5365 5967 5399 6001
rect 5457 5967 5491 6001
rect 5549 5967 5583 6001
rect 5641 5967 5675 6001
rect 5733 5967 5767 6001
rect 5825 5967 5859 6001
rect 5917 5967 5951 6001
rect 6009 5967 6043 6001
rect 6101 5967 6135 6001
rect 6193 5967 6227 6001
rect 6285 5967 6319 6001
rect 6377 5967 6411 6001
rect 6469 5967 6503 6001
rect 6561 5967 6595 6001
rect 6653 5967 6687 6001
rect 6745 5967 6779 6001
rect 6837 5967 6871 6001
rect 6929 5967 6963 6001
rect 7021 5967 7055 6001
rect 7113 5967 7147 6001
rect 7205 5967 7239 6001
rect 7297 5967 7331 6001
rect 7389 5967 7423 6001
rect 7481 5967 7515 6001
rect 7573 5967 7607 6001
rect 7665 5967 7699 6001
rect 7757 5967 7791 6001
rect 7849 5967 7883 6001
rect 7941 5967 7975 6001
rect 8033 5967 8067 6001
rect 8125 5967 8159 6001
rect 8217 5967 8251 6001
rect 8309 5967 8343 6001
rect 8401 5967 8435 6001
rect 8493 5967 8527 6001
rect 8585 5967 8619 6001
rect 8677 5967 8711 6001
rect 8769 5967 8803 6001
rect 8861 5967 8895 6001
rect 8953 5967 8987 6001
rect 9045 5967 9079 6001
rect 9137 5967 9171 6001
rect 9229 5967 9263 6001
rect 9321 5967 9355 6001
rect 9413 5967 9447 6001
rect 9505 5967 9539 6001
rect 9597 5967 9631 6001
rect 9689 5967 9723 6001
rect 9781 5967 9815 6001
rect 9873 5967 9907 6001
rect 9965 5967 9999 6001
rect 10057 5967 10091 6001
rect 10149 5967 10183 6001
rect 10241 5967 10275 6001
rect 10333 5967 10367 6001
rect 10425 5967 10459 6001
rect 10517 5967 10551 6001
rect 10609 5967 10643 6001
rect 10701 5967 10735 6001
rect 10793 5967 10827 6001
rect 10885 5967 10919 6001
rect 10977 5967 11011 6001
rect 11069 5967 11103 6001
rect 11161 5967 11195 6001
rect 11253 5967 11287 6001
rect 11345 5967 11379 6001
rect 11437 5967 11471 6001
rect 11529 5967 11563 6001
rect 11621 5967 11655 6001
rect 11713 5967 11747 6001
rect 11805 5967 11839 6001
rect 11897 5967 11931 6001
rect 11989 5967 12023 6001
rect 12081 5967 12115 6001
rect 12173 5967 12207 6001
rect 12265 5967 12299 6001
rect 12357 5967 12391 6001
rect 12449 5967 12483 6001
rect 12541 5967 12575 6001
rect 12633 5967 12667 6001
rect 12725 5967 12759 6001
rect 12817 5967 12851 6001
rect 12909 5967 12943 6001
rect 13001 5967 13035 6001
rect 13093 5967 13127 6001
rect 13185 5967 13219 6001
rect 13277 5967 13311 6001
rect 13369 5967 13403 6001
rect 13461 5967 13495 6001
rect 13553 5967 13587 6001
rect 13645 5967 13679 6001
rect 13737 5967 13771 6001
rect 13829 5967 13863 6001
rect 13921 5967 13955 6001
rect 14013 5967 14047 6001
rect 14105 5967 14139 6001
rect 14197 5967 14231 6001
rect 14289 5967 14323 6001
rect 14381 5967 14415 6001
rect 14473 5967 14507 6001
rect 14565 5967 14599 6001
rect 14657 5967 14691 6001
rect 14749 5967 14783 6001
rect 14841 5967 14875 6001
rect 14933 5967 14967 6001
rect 15025 5967 15059 6001
rect 15117 5967 15151 6001
rect 15209 5967 15243 6001
rect 15301 5967 15335 6001
rect 15393 5967 15427 6001
rect 15485 5967 15519 6001
rect 15577 5967 15611 6001
rect 15669 5967 15703 6001
rect 15761 5967 15795 6001
rect 15853 5967 15887 6001
rect 15945 5967 15979 6001
rect 16037 5967 16071 6001
rect 16129 5967 16163 6001
rect 16221 5967 16255 6001
rect 16313 5967 16347 6001
rect 16405 5967 16439 6001
rect 16497 5967 16531 6001
rect 16589 5967 16623 6001
rect 16681 5967 16715 6001
rect 16773 5967 16807 6001
rect 16865 5967 16899 6001
rect 16957 5967 16991 6001
rect 17049 5967 17083 6001
rect 17141 5967 17175 6001
rect 17233 5967 17267 6001
rect 17325 5967 17359 6001
rect 17417 5967 17451 6001
rect 17509 5967 17543 6001
rect 17601 5967 17635 6001
rect 17693 5967 17727 6001
rect 17785 5967 17819 6001
rect 17877 5967 17911 6001
rect 17969 5967 18003 6001
rect 18061 5967 18095 6001
rect 18153 5967 18187 6001
rect 18245 5967 18279 6001
rect 18337 5967 18371 6001
rect 18429 5967 18463 6001
rect 18521 5967 18555 6001
rect 18613 5967 18647 6001
rect 18705 5967 18739 6001
rect 18797 5967 18831 6001
rect 2421 5802 2449 5831
rect 2449 5802 2455 5831
rect 2421 5797 2455 5802
rect 2237 5689 2271 5695
rect 2237 5661 2245 5689
rect 2245 5661 2271 5689
rect 3249 5689 3283 5695
rect 3249 5661 3275 5689
rect 3275 5661 3283 5689
rect 3065 5529 3071 5559
rect 3071 5529 3099 5559
rect 3065 5525 3099 5529
rect 6745 5552 6779 5559
rect 6745 5525 6751 5552
rect 6751 5525 6779 5552
rect 7113 5525 7147 5559
rect 7297 5729 7331 5763
rect 7205 5593 7239 5627
rect 10241 5661 10275 5695
rect 9873 5552 9907 5559
rect 9873 5525 9879 5552
rect 9879 5525 9907 5552
rect 10425 5729 10459 5763
rect 10333 5593 10367 5627
rect 11437 5729 11471 5763
rect 11253 5689 11287 5695
rect 11253 5661 11285 5689
rect 11285 5661 11287 5689
rect 11069 5525 11103 5559
rect 12265 5823 12271 5831
rect 12271 5823 12299 5831
rect 12265 5797 12299 5823
rect 12633 5525 12667 5559
rect 12817 5729 12851 5763
rect 12725 5593 12759 5627
rect 14289 5552 14323 5559
rect 14289 5525 14295 5552
rect 14295 5525 14323 5552
rect 14657 5525 14691 5559
rect 14841 5729 14875 5763
rect 14749 5593 14783 5627
rect 1133 5423 1167 5457
rect 1225 5423 1259 5457
rect 1317 5423 1351 5457
rect 1409 5423 1443 5457
rect 1501 5423 1535 5457
rect 1593 5423 1627 5457
rect 1685 5423 1719 5457
rect 1777 5423 1811 5457
rect 1869 5423 1903 5457
rect 1961 5423 1995 5457
rect 2053 5423 2087 5457
rect 2145 5423 2179 5457
rect 2237 5423 2271 5457
rect 2329 5423 2363 5457
rect 2421 5423 2455 5457
rect 2513 5423 2547 5457
rect 2605 5423 2639 5457
rect 2697 5423 2731 5457
rect 2789 5423 2823 5457
rect 2881 5423 2915 5457
rect 2973 5423 3007 5457
rect 3065 5423 3099 5457
rect 3157 5423 3191 5457
rect 3249 5423 3283 5457
rect 3341 5423 3375 5457
rect 3433 5423 3467 5457
rect 3525 5423 3559 5457
rect 3617 5423 3651 5457
rect 3709 5423 3743 5457
rect 3801 5423 3835 5457
rect 3893 5423 3927 5457
rect 3985 5423 4019 5457
rect 4077 5423 4111 5457
rect 4169 5423 4203 5457
rect 4261 5423 4295 5457
rect 4353 5423 4387 5457
rect 4445 5423 4479 5457
rect 4537 5423 4571 5457
rect 4629 5423 4663 5457
rect 4721 5423 4755 5457
rect 4813 5423 4847 5457
rect 4905 5423 4939 5457
rect 4997 5423 5031 5457
rect 5089 5423 5123 5457
rect 5181 5423 5215 5457
rect 5273 5423 5307 5457
rect 5365 5423 5399 5457
rect 5457 5423 5491 5457
rect 5549 5423 5583 5457
rect 5641 5423 5675 5457
rect 5733 5423 5767 5457
rect 5825 5423 5859 5457
rect 5917 5423 5951 5457
rect 6009 5423 6043 5457
rect 6101 5423 6135 5457
rect 6193 5423 6227 5457
rect 6285 5423 6319 5457
rect 6377 5423 6411 5457
rect 6469 5423 6503 5457
rect 6561 5423 6595 5457
rect 6653 5423 6687 5457
rect 6745 5423 6779 5457
rect 6837 5423 6871 5457
rect 6929 5423 6963 5457
rect 7021 5423 7055 5457
rect 7113 5423 7147 5457
rect 7205 5423 7239 5457
rect 7297 5423 7331 5457
rect 7389 5423 7423 5457
rect 7481 5423 7515 5457
rect 7573 5423 7607 5457
rect 7665 5423 7699 5457
rect 7757 5423 7791 5457
rect 7849 5423 7883 5457
rect 7941 5423 7975 5457
rect 8033 5423 8067 5457
rect 8125 5423 8159 5457
rect 8217 5423 8251 5457
rect 8309 5423 8343 5457
rect 8401 5423 8435 5457
rect 8493 5423 8527 5457
rect 8585 5423 8619 5457
rect 8677 5423 8711 5457
rect 8769 5423 8803 5457
rect 8861 5423 8895 5457
rect 8953 5423 8987 5457
rect 9045 5423 9079 5457
rect 9137 5423 9171 5457
rect 9229 5423 9263 5457
rect 9321 5423 9355 5457
rect 9413 5423 9447 5457
rect 9505 5423 9539 5457
rect 9597 5423 9631 5457
rect 9689 5423 9723 5457
rect 9781 5423 9815 5457
rect 9873 5423 9907 5457
rect 9965 5423 9999 5457
rect 10057 5423 10091 5457
rect 10149 5423 10183 5457
rect 10241 5423 10275 5457
rect 10333 5423 10367 5457
rect 10425 5423 10459 5457
rect 10517 5423 10551 5457
rect 10609 5423 10643 5457
rect 10701 5423 10735 5457
rect 10793 5423 10827 5457
rect 10885 5423 10919 5457
rect 10977 5423 11011 5457
rect 11069 5423 11103 5457
rect 11161 5423 11195 5457
rect 11253 5423 11287 5457
rect 11345 5423 11379 5457
rect 11437 5423 11471 5457
rect 11529 5423 11563 5457
rect 11621 5423 11655 5457
rect 11713 5423 11747 5457
rect 11805 5423 11839 5457
rect 11897 5423 11931 5457
rect 11989 5423 12023 5457
rect 12081 5423 12115 5457
rect 12173 5423 12207 5457
rect 12265 5423 12299 5457
rect 12357 5423 12391 5457
rect 12449 5423 12483 5457
rect 12541 5423 12575 5457
rect 12633 5423 12667 5457
rect 12725 5423 12759 5457
rect 12817 5423 12851 5457
rect 12909 5423 12943 5457
rect 13001 5423 13035 5457
rect 13093 5423 13127 5457
rect 13185 5423 13219 5457
rect 13277 5423 13311 5457
rect 13369 5423 13403 5457
rect 13461 5423 13495 5457
rect 13553 5423 13587 5457
rect 13645 5423 13679 5457
rect 13737 5423 13771 5457
rect 13829 5423 13863 5457
rect 13921 5423 13955 5457
rect 14013 5423 14047 5457
rect 14105 5423 14139 5457
rect 14197 5423 14231 5457
rect 14289 5423 14323 5457
rect 14381 5423 14415 5457
rect 14473 5423 14507 5457
rect 14565 5423 14599 5457
rect 14657 5423 14691 5457
rect 14749 5423 14783 5457
rect 14841 5423 14875 5457
rect 14933 5423 14967 5457
rect 15025 5423 15059 5457
rect 15117 5423 15151 5457
rect 15209 5423 15243 5457
rect 15301 5423 15335 5457
rect 15393 5423 15427 5457
rect 15485 5423 15519 5457
rect 15577 5423 15611 5457
rect 15669 5423 15703 5457
rect 15761 5423 15795 5457
rect 15853 5423 15887 5457
rect 15945 5423 15979 5457
rect 16037 5423 16071 5457
rect 16129 5423 16163 5457
rect 16221 5423 16255 5457
rect 16313 5423 16347 5457
rect 16405 5423 16439 5457
rect 16497 5423 16531 5457
rect 16589 5423 16623 5457
rect 16681 5423 16715 5457
rect 16773 5423 16807 5457
rect 16865 5423 16899 5457
rect 16957 5423 16991 5457
rect 17049 5423 17083 5457
rect 17141 5423 17175 5457
rect 17233 5423 17267 5457
rect 17325 5423 17359 5457
rect 17417 5423 17451 5457
rect 17509 5423 17543 5457
rect 17601 5423 17635 5457
rect 17693 5423 17727 5457
rect 17785 5423 17819 5457
rect 17877 5423 17911 5457
rect 17969 5423 18003 5457
rect 18061 5423 18095 5457
rect 18153 5423 18187 5457
rect 18245 5423 18279 5457
rect 18337 5423 18371 5457
rect 18429 5423 18463 5457
rect 18521 5423 18555 5457
rect 18613 5423 18647 5457
rect 18705 5423 18739 5457
rect 18797 5423 18831 5457
rect 2881 5321 2915 5355
rect 2145 5191 2177 5219
rect 2177 5191 2179 5219
rect 2145 5185 2179 5191
rect 2329 5117 2363 5151
rect 1961 4989 1995 5015
rect 1961 4981 1991 4989
rect 1991 4981 1995 4989
rect 3893 5351 3927 5355
rect 3893 5321 3894 5351
rect 3894 5321 3927 5351
rect 3065 5191 3097 5219
rect 3097 5191 3099 5219
rect 3065 5185 3099 5191
rect 3249 5185 3283 5219
rect 3709 5191 3717 5219
rect 3717 5191 3743 5219
rect 3709 5185 3743 5191
rect 4445 5191 4453 5219
rect 4453 5191 4479 5219
rect 4445 5185 4479 5191
rect 4537 4989 4571 5015
rect 4537 4981 4571 4989
rect 7021 5321 7055 5355
rect 6009 5191 6035 5219
rect 6035 5191 6043 5219
rect 6009 5185 6043 5191
rect 5825 4997 5859 5015
rect 5825 4981 5831 4997
rect 5831 4981 5859 4997
rect 6653 4989 6687 5015
rect 6653 4981 6659 4989
rect 6659 4981 6687 4989
rect 7113 5321 7147 5355
rect 7297 5148 7331 5151
rect 7297 5117 7317 5148
rect 7317 5117 7331 5148
rect 7849 4989 7883 5015
rect 7849 4981 7855 4989
rect 7855 4981 7883 4989
rect 8217 5185 8251 5219
rect 8309 5321 8343 5355
rect 8401 5117 8435 5151
rect 9321 5185 9355 5219
rect 9505 5185 9539 5219
rect 9137 4997 9171 5015
rect 9137 4981 9147 4997
rect 9147 4981 9171 4997
rect 9597 5117 9631 5151
rect 10425 4989 10459 5015
rect 10425 4981 10431 4989
rect 10431 4981 10459 4989
rect 10793 5185 10827 5219
rect 10885 5321 10919 5355
rect 10977 5117 11011 5151
rect 13461 5321 13495 5355
rect 13093 4989 13127 5015
rect 13093 4981 13099 4989
rect 13099 4981 13127 4989
rect 13553 5321 13587 5355
rect 13645 5117 13679 5151
rect 1133 4879 1167 4913
rect 1225 4879 1259 4913
rect 1317 4879 1351 4913
rect 1409 4879 1443 4913
rect 1501 4879 1535 4913
rect 1593 4879 1627 4913
rect 1685 4879 1719 4913
rect 1777 4879 1811 4913
rect 1869 4879 1903 4913
rect 1961 4879 1995 4913
rect 2053 4879 2087 4913
rect 2145 4879 2179 4913
rect 2237 4879 2271 4913
rect 2329 4879 2363 4913
rect 2421 4879 2455 4913
rect 2513 4879 2547 4913
rect 2605 4879 2639 4913
rect 2697 4879 2731 4913
rect 2789 4879 2823 4913
rect 2881 4879 2915 4913
rect 2973 4879 3007 4913
rect 3065 4879 3099 4913
rect 3157 4879 3191 4913
rect 3249 4879 3283 4913
rect 3341 4879 3375 4913
rect 3433 4879 3467 4913
rect 3525 4879 3559 4913
rect 3617 4879 3651 4913
rect 3709 4879 3743 4913
rect 3801 4879 3835 4913
rect 3893 4879 3927 4913
rect 3985 4879 4019 4913
rect 4077 4879 4111 4913
rect 4169 4879 4203 4913
rect 4261 4879 4295 4913
rect 4353 4879 4387 4913
rect 4445 4879 4479 4913
rect 4537 4879 4571 4913
rect 4629 4879 4663 4913
rect 4721 4879 4755 4913
rect 4813 4879 4847 4913
rect 4905 4879 4939 4913
rect 4997 4879 5031 4913
rect 5089 4879 5123 4913
rect 5181 4879 5215 4913
rect 5273 4879 5307 4913
rect 5365 4879 5399 4913
rect 5457 4879 5491 4913
rect 5549 4879 5583 4913
rect 5641 4879 5675 4913
rect 5733 4879 5767 4913
rect 5825 4879 5859 4913
rect 5917 4879 5951 4913
rect 6009 4879 6043 4913
rect 6101 4879 6135 4913
rect 6193 4879 6227 4913
rect 6285 4879 6319 4913
rect 6377 4879 6411 4913
rect 6469 4879 6503 4913
rect 6561 4879 6595 4913
rect 6653 4879 6687 4913
rect 6745 4879 6779 4913
rect 6837 4879 6871 4913
rect 6929 4879 6963 4913
rect 7021 4879 7055 4913
rect 7113 4879 7147 4913
rect 7205 4879 7239 4913
rect 7297 4879 7331 4913
rect 7389 4879 7423 4913
rect 7481 4879 7515 4913
rect 7573 4879 7607 4913
rect 7665 4879 7699 4913
rect 7757 4879 7791 4913
rect 7849 4879 7883 4913
rect 7941 4879 7975 4913
rect 8033 4879 8067 4913
rect 8125 4879 8159 4913
rect 8217 4879 8251 4913
rect 8309 4879 8343 4913
rect 8401 4879 8435 4913
rect 8493 4879 8527 4913
rect 8585 4879 8619 4913
rect 8677 4879 8711 4913
rect 8769 4879 8803 4913
rect 8861 4879 8895 4913
rect 8953 4879 8987 4913
rect 9045 4879 9079 4913
rect 9137 4879 9171 4913
rect 9229 4879 9263 4913
rect 9321 4879 9355 4913
rect 9413 4879 9447 4913
rect 9505 4879 9539 4913
rect 9597 4879 9631 4913
rect 9689 4879 9723 4913
rect 9781 4879 9815 4913
rect 9873 4879 9907 4913
rect 9965 4879 9999 4913
rect 10057 4879 10091 4913
rect 10149 4879 10183 4913
rect 10241 4879 10275 4913
rect 10333 4879 10367 4913
rect 10425 4879 10459 4913
rect 10517 4879 10551 4913
rect 10609 4879 10643 4913
rect 10701 4879 10735 4913
rect 10793 4879 10827 4913
rect 10885 4879 10919 4913
rect 10977 4879 11011 4913
rect 11069 4879 11103 4913
rect 11161 4879 11195 4913
rect 11253 4879 11287 4913
rect 11345 4879 11379 4913
rect 11437 4879 11471 4913
rect 11529 4879 11563 4913
rect 11621 4879 11655 4913
rect 11713 4879 11747 4913
rect 11805 4879 11839 4913
rect 11897 4879 11931 4913
rect 11989 4879 12023 4913
rect 12081 4879 12115 4913
rect 12173 4879 12207 4913
rect 12265 4879 12299 4913
rect 12357 4879 12391 4913
rect 12449 4879 12483 4913
rect 12541 4879 12575 4913
rect 12633 4879 12667 4913
rect 12725 4879 12759 4913
rect 12817 4879 12851 4913
rect 12909 4879 12943 4913
rect 13001 4879 13035 4913
rect 13093 4879 13127 4913
rect 13185 4879 13219 4913
rect 13277 4879 13311 4913
rect 13369 4879 13403 4913
rect 13461 4879 13495 4913
rect 13553 4879 13587 4913
rect 13645 4879 13679 4913
rect 13737 4879 13771 4913
rect 13829 4879 13863 4913
rect 13921 4879 13955 4913
rect 14013 4879 14047 4913
rect 14105 4879 14139 4913
rect 14197 4879 14231 4913
rect 14289 4879 14323 4913
rect 14381 4879 14415 4913
rect 14473 4879 14507 4913
rect 14565 4879 14599 4913
rect 14657 4879 14691 4913
rect 14749 4879 14783 4913
rect 14841 4879 14875 4913
rect 14933 4879 14967 4913
rect 15025 4879 15059 4913
rect 15117 4879 15151 4913
rect 15209 4879 15243 4913
rect 15301 4879 15335 4913
rect 15393 4879 15427 4913
rect 15485 4879 15519 4913
rect 15577 4879 15611 4913
rect 15669 4879 15703 4913
rect 15761 4879 15795 4913
rect 15853 4879 15887 4913
rect 15945 4879 15979 4913
rect 16037 4879 16071 4913
rect 16129 4879 16163 4913
rect 16221 4879 16255 4913
rect 16313 4879 16347 4913
rect 16405 4879 16439 4913
rect 16497 4879 16531 4913
rect 16589 4879 16623 4913
rect 16681 4879 16715 4913
rect 16773 4879 16807 4913
rect 16865 4879 16899 4913
rect 16957 4879 16991 4913
rect 17049 4879 17083 4913
rect 17141 4879 17175 4913
rect 17233 4879 17267 4913
rect 17325 4879 17359 4913
rect 17417 4879 17451 4913
rect 17509 4879 17543 4913
rect 17601 4879 17635 4913
rect 17693 4879 17727 4913
rect 17785 4879 17819 4913
rect 17877 4879 17911 4913
rect 17969 4879 18003 4913
rect 18061 4879 18095 4913
rect 18153 4879 18187 4913
rect 18245 4879 18279 4913
rect 18337 4879 18371 4913
rect 18429 4879 18463 4913
rect 18521 4879 18555 4913
rect 18613 4879 18647 4913
rect 18705 4879 18739 4913
rect 18797 4879 18831 4913
rect 2150 4709 2184 4743
rect 2053 4601 2087 4607
rect 2053 4573 2056 4601
rect 2056 4573 2087 4601
rect 2229 4641 2263 4675
rect 2320 4573 2354 4607
rect 2570 4717 2604 4743
rect 2570 4709 2572 4717
rect 2572 4709 2604 4717
rect 2467 4641 2501 4675
rect 2884 4709 2918 4743
rect 2971 4641 3005 4675
rect 3985 4803 4015 4811
rect 4015 4803 4019 4811
rect 3985 4777 4019 4803
rect 3433 4448 3467 4471
rect 3433 4437 3453 4448
rect 3453 4437 3467 4448
rect 4353 4641 4387 4675
rect 4169 4601 4203 4607
rect 4169 4573 4201 4601
rect 4201 4573 4203 4601
rect 5273 4777 5307 4811
rect 5377 4641 5411 4675
rect 5089 4573 5123 4607
rect 4905 4448 4939 4471
rect 4905 4437 4911 4448
rect 4911 4437 4939 4448
rect 6193 4777 6227 4811
rect 6285 4641 6319 4675
rect 6842 4709 6876 4743
rect 6009 4573 6043 4607
rect 5825 4448 5859 4471
rect 5825 4437 5831 4448
rect 5831 4437 5859 4448
rect 6745 4601 6779 4607
rect 6745 4573 6748 4601
rect 6748 4573 6779 4601
rect 6921 4641 6955 4675
rect 7012 4573 7046 4607
rect 7262 4717 7296 4743
rect 7262 4709 7264 4717
rect 7264 4709 7296 4717
rect 7159 4641 7193 4675
rect 7576 4709 7610 4743
rect 7663 4641 7697 4675
rect 9965 4797 9981 4811
rect 9981 4797 9999 4811
rect 9965 4777 9999 4797
rect 8125 4448 8159 4471
rect 8125 4437 8145 4448
rect 8145 4437 8159 4448
rect 10427 4641 10461 4675
rect 10514 4709 10548 4743
rect 10828 4717 10862 4743
rect 10828 4709 10860 4717
rect 10860 4709 10862 4717
rect 10931 4641 10965 4675
rect 11100 4505 11134 4539
rect 11169 4641 11203 4675
rect 11248 4709 11282 4743
rect 11345 4601 11379 4607
rect 11345 4573 11376 4601
rect 11376 4573 11379 4601
rect 12173 4777 12207 4811
rect 12265 4641 12299 4675
rect 11989 4573 12023 4607
rect 11805 4448 11839 4471
rect 11805 4437 11811 4448
rect 11811 4437 11839 4448
rect 13093 4641 13127 4675
rect 12909 4573 12943 4607
rect 13185 4601 13219 4607
rect 13185 4573 13215 4601
rect 13215 4573 13219 4601
rect 12725 4448 12759 4471
rect 12725 4437 12731 4448
rect 12731 4437 12759 4448
rect 14381 4573 14415 4607
rect 14565 4601 14599 4607
rect 14565 4573 14567 4601
rect 14567 4573 14599 4601
rect 14749 4437 14783 4471
rect 1133 4335 1167 4369
rect 1225 4335 1259 4369
rect 1317 4335 1351 4369
rect 1409 4335 1443 4369
rect 1501 4335 1535 4369
rect 1593 4335 1627 4369
rect 1685 4335 1719 4369
rect 1777 4335 1811 4369
rect 1869 4335 1903 4369
rect 1961 4335 1995 4369
rect 2053 4335 2087 4369
rect 2145 4335 2179 4369
rect 2237 4335 2271 4369
rect 2329 4335 2363 4369
rect 2421 4335 2455 4369
rect 2513 4335 2547 4369
rect 2605 4335 2639 4369
rect 2697 4335 2731 4369
rect 2789 4335 2823 4369
rect 2881 4335 2915 4369
rect 2973 4335 3007 4369
rect 3065 4335 3099 4369
rect 3157 4335 3191 4369
rect 3249 4335 3283 4369
rect 3341 4335 3375 4369
rect 3433 4335 3467 4369
rect 3525 4335 3559 4369
rect 3617 4335 3651 4369
rect 3709 4335 3743 4369
rect 3801 4335 3835 4369
rect 3893 4335 3927 4369
rect 3985 4335 4019 4369
rect 4077 4335 4111 4369
rect 4169 4335 4203 4369
rect 4261 4335 4295 4369
rect 4353 4335 4387 4369
rect 4445 4335 4479 4369
rect 4537 4335 4571 4369
rect 4629 4335 4663 4369
rect 4721 4335 4755 4369
rect 4813 4335 4847 4369
rect 4905 4335 4939 4369
rect 4997 4335 5031 4369
rect 5089 4335 5123 4369
rect 5181 4335 5215 4369
rect 5273 4335 5307 4369
rect 5365 4335 5399 4369
rect 5457 4335 5491 4369
rect 5549 4335 5583 4369
rect 5641 4335 5675 4369
rect 5733 4335 5767 4369
rect 5825 4335 5859 4369
rect 5917 4335 5951 4369
rect 6009 4335 6043 4369
rect 6101 4335 6135 4369
rect 6193 4335 6227 4369
rect 6285 4335 6319 4369
rect 6377 4335 6411 4369
rect 6469 4335 6503 4369
rect 6561 4335 6595 4369
rect 6653 4335 6687 4369
rect 6745 4335 6779 4369
rect 6837 4335 6871 4369
rect 6929 4335 6963 4369
rect 7021 4335 7055 4369
rect 7113 4335 7147 4369
rect 7205 4335 7239 4369
rect 7297 4335 7331 4369
rect 7389 4335 7423 4369
rect 7481 4335 7515 4369
rect 7573 4335 7607 4369
rect 7665 4335 7699 4369
rect 7757 4335 7791 4369
rect 7849 4335 7883 4369
rect 7941 4335 7975 4369
rect 8033 4335 8067 4369
rect 8125 4335 8159 4369
rect 8217 4335 8251 4369
rect 8309 4335 8343 4369
rect 8401 4335 8435 4369
rect 8493 4335 8527 4369
rect 8585 4335 8619 4369
rect 8677 4335 8711 4369
rect 8769 4335 8803 4369
rect 8861 4335 8895 4369
rect 8953 4335 8987 4369
rect 9045 4335 9079 4369
rect 9137 4335 9171 4369
rect 9229 4335 9263 4369
rect 9321 4335 9355 4369
rect 9413 4335 9447 4369
rect 9505 4335 9539 4369
rect 9597 4335 9631 4369
rect 9689 4335 9723 4369
rect 9781 4335 9815 4369
rect 9873 4335 9907 4369
rect 9965 4335 9999 4369
rect 10057 4335 10091 4369
rect 10149 4335 10183 4369
rect 10241 4335 10275 4369
rect 10333 4335 10367 4369
rect 10425 4335 10459 4369
rect 10517 4335 10551 4369
rect 10609 4335 10643 4369
rect 10701 4335 10735 4369
rect 10793 4335 10827 4369
rect 10885 4335 10919 4369
rect 10977 4335 11011 4369
rect 11069 4335 11103 4369
rect 11161 4335 11195 4369
rect 11253 4335 11287 4369
rect 11345 4335 11379 4369
rect 11437 4335 11471 4369
rect 11529 4335 11563 4369
rect 11621 4335 11655 4369
rect 11713 4335 11747 4369
rect 11805 4335 11839 4369
rect 11897 4335 11931 4369
rect 11989 4335 12023 4369
rect 12081 4335 12115 4369
rect 12173 4335 12207 4369
rect 12265 4335 12299 4369
rect 12357 4335 12391 4369
rect 12449 4335 12483 4369
rect 12541 4335 12575 4369
rect 12633 4335 12667 4369
rect 12725 4335 12759 4369
rect 12817 4335 12851 4369
rect 12909 4335 12943 4369
rect 13001 4335 13035 4369
rect 13093 4335 13127 4369
rect 13185 4335 13219 4369
rect 13277 4335 13311 4369
rect 13369 4335 13403 4369
rect 13461 4335 13495 4369
rect 13553 4335 13587 4369
rect 13645 4335 13679 4369
rect 13737 4335 13771 4369
rect 13829 4335 13863 4369
rect 13921 4335 13955 4369
rect 14013 4335 14047 4369
rect 14105 4335 14139 4369
rect 14197 4335 14231 4369
rect 14289 4335 14323 4369
rect 14381 4335 14415 4369
rect 14473 4335 14507 4369
rect 14565 4335 14599 4369
rect 14657 4335 14691 4369
rect 14749 4335 14783 4369
rect 14841 4335 14875 4369
rect 14933 4335 14967 4369
rect 15025 4335 15059 4369
rect 15117 4335 15151 4369
rect 15209 4335 15243 4369
rect 15301 4335 15335 4369
rect 15393 4335 15427 4369
rect 15485 4335 15519 4369
rect 15577 4335 15611 4369
rect 15669 4335 15703 4369
rect 15761 4335 15795 4369
rect 15853 4335 15887 4369
rect 15945 4335 15979 4369
rect 16037 4335 16071 4369
rect 16129 4335 16163 4369
rect 16221 4335 16255 4369
rect 16313 4335 16347 4369
rect 16405 4335 16439 4369
rect 16497 4335 16531 4369
rect 16589 4335 16623 4369
rect 16681 4335 16715 4369
rect 16773 4335 16807 4369
rect 16865 4335 16899 4369
rect 16957 4335 16991 4369
rect 17049 4335 17083 4369
rect 17141 4335 17175 4369
rect 17233 4335 17267 4369
rect 17325 4335 17359 4369
rect 17417 4335 17451 4369
rect 17509 4335 17543 4369
rect 17601 4335 17635 4369
rect 17693 4335 17727 4369
rect 17785 4335 17819 4369
rect 17877 4335 17911 4369
rect 17969 4335 18003 4369
rect 18061 4335 18095 4369
rect 18153 4335 18187 4369
rect 18245 4335 18279 4369
rect 18337 4335 18371 4369
rect 18429 4335 18463 4369
rect 18521 4335 18555 4369
rect 18613 4335 18647 4369
rect 18705 4335 18739 4369
rect 18797 4335 18831 4369
rect 1961 4103 1969 4131
rect 1969 4103 1995 4131
rect 1961 4097 1995 4103
rect 2605 4256 2619 4267
rect 2619 4256 2639 4267
rect 2605 4233 2639 4256
rect 2145 3990 2179 3995
rect 2145 3961 2173 3990
rect 2173 3961 2179 3990
rect 3067 4029 3101 4063
rect 3154 3961 3188 3995
rect 3571 4029 3605 4063
rect 3468 3987 3500 3995
rect 3500 3987 3502 3995
rect 3468 3961 3502 3987
rect 3729 4097 3763 4131
rect 3809 4029 3843 4063
rect 4629 4256 4643 4267
rect 4643 4256 4663 4267
rect 4629 4233 4663 4256
rect 3985 4103 4016 4131
rect 4016 4103 4019 4131
rect 3985 4097 4019 4103
rect 3888 3961 3922 3995
rect 5091 4029 5125 4063
rect 5178 3961 5212 3995
rect 5595 4029 5629 4063
rect 5492 3987 5524 3995
rect 5524 3987 5526 3995
rect 5492 3961 5526 3987
rect 5742 4097 5776 4131
rect 5833 4029 5867 4063
rect 6009 4103 6040 4131
rect 6040 4103 6043 4131
rect 6009 4097 6043 4103
rect 5912 3961 5946 3995
rect 7113 4097 7147 4131
rect 7297 4097 7331 4131
rect 6929 3909 6963 3927
rect 6929 3893 6939 3909
rect 6939 3893 6963 3909
rect 7849 4165 7883 4199
rect 7389 4029 7423 4063
rect 9597 4029 9631 4063
rect 10701 4097 10735 4131
rect 10517 3909 10551 3927
rect 10517 3893 10527 3909
rect 10527 3893 10551 3909
rect 10977 4029 11011 4063
rect 11713 4103 11716 4131
rect 11716 4103 11747 4131
rect 11713 4097 11747 4103
rect 10885 3961 10919 3995
rect 11810 3961 11844 3995
rect 11889 4029 11923 4063
rect 11980 4165 12014 4199
rect 12127 4029 12161 4063
rect 12230 3987 12232 3995
rect 12232 3987 12264 3995
rect 12230 3961 12264 3987
rect 12544 3961 12578 3995
rect 12631 4029 12665 4063
rect 13093 4256 13113 4267
rect 13113 4256 13127 4267
rect 13093 4233 13127 4256
rect 15669 4103 15695 4131
rect 15695 4103 15703 4131
rect 15669 4097 15703 4103
rect 17049 4103 17051 4131
rect 17051 4103 17083 4131
rect 17049 4097 17083 4103
rect 15485 3909 15519 3927
rect 15485 3893 15491 3909
rect 15491 3893 15519 3909
rect 16865 4029 16899 4063
rect 17233 3901 17267 3927
rect 17233 3893 17237 3901
rect 17237 3893 17267 3901
rect 1133 3791 1167 3825
rect 1225 3791 1259 3825
rect 1317 3791 1351 3825
rect 1409 3791 1443 3825
rect 1501 3791 1535 3825
rect 1593 3791 1627 3825
rect 1685 3791 1719 3825
rect 1777 3791 1811 3825
rect 1869 3791 1903 3825
rect 1961 3791 1995 3825
rect 2053 3791 2087 3825
rect 2145 3791 2179 3825
rect 2237 3791 2271 3825
rect 2329 3791 2363 3825
rect 2421 3791 2455 3825
rect 2513 3791 2547 3825
rect 2605 3791 2639 3825
rect 2697 3791 2731 3825
rect 2789 3791 2823 3825
rect 2881 3791 2915 3825
rect 2973 3791 3007 3825
rect 3065 3791 3099 3825
rect 3157 3791 3191 3825
rect 3249 3791 3283 3825
rect 3341 3791 3375 3825
rect 3433 3791 3467 3825
rect 3525 3791 3559 3825
rect 3617 3791 3651 3825
rect 3709 3791 3743 3825
rect 3801 3791 3835 3825
rect 3893 3791 3927 3825
rect 3985 3791 4019 3825
rect 4077 3791 4111 3825
rect 4169 3791 4203 3825
rect 4261 3791 4295 3825
rect 4353 3791 4387 3825
rect 4445 3791 4479 3825
rect 4537 3791 4571 3825
rect 4629 3791 4663 3825
rect 4721 3791 4755 3825
rect 4813 3791 4847 3825
rect 4905 3791 4939 3825
rect 4997 3791 5031 3825
rect 5089 3791 5123 3825
rect 5181 3791 5215 3825
rect 5273 3791 5307 3825
rect 5365 3791 5399 3825
rect 5457 3791 5491 3825
rect 5549 3791 5583 3825
rect 5641 3791 5675 3825
rect 5733 3791 5767 3825
rect 5825 3791 5859 3825
rect 5917 3791 5951 3825
rect 6009 3791 6043 3825
rect 6101 3791 6135 3825
rect 6193 3791 6227 3825
rect 6285 3791 6319 3825
rect 6377 3791 6411 3825
rect 6469 3791 6503 3825
rect 6561 3791 6595 3825
rect 6653 3791 6687 3825
rect 6745 3791 6779 3825
rect 6837 3791 6871 3825
rect 6929 3791 6963 3825
rect 7021 3791 7055 3825
rect 7113 3791 7147 3825
rect 7205 3791 7239 3825
rect 7297 3791 7331 3825
rect 7389 3791 7423 3825
rect 7481 3791 7515 3825
rect 7573 3791 7607 3825
rect 7665 3791 7699 3825
rect 7757 3791 7791 3825
rect 7849 3791 7883 3825
rect 7941 3791 7975 3825
rect 8033 3791 8067 3825
rect 8125 3791 8159 3825
rect 8217 3791 8251 3825
rect 8309 3791 8343 3825
rect 8401 3791 8435 3825
rect 8493 3791 8527 3825
rect 8585 3791 8619 3825
rect 8677 3791 8711 3825
rect 8769 3791 8803 3825
rect 8861 3791 8895 3825
rect 8953 3791 8987 3825
rect 9045 3791 9079 3825
rect 9137 3791 9171 3825
rect 9229 3791 9263 3825
rect 9321 3791 9355 3825
rect 9413 3791 9447 3825
rect 9505 3791 9539 3825
rect 9597 3791 9631 3825
rect 9689 3791 9723 3825
rect 9781 3791 9815 3825
rect 9873 3791 9907 3825
rect 9965 3791 9999 3825
rect 10057 3791 10091 3825
rect 10149 3791 10183 3825
rect 10241 3791 10275 3825
rect 10333 3791 10367 3825
rect 10425 3791 10459 3825
rect 10517 3791 10551 3825
rect 10609 3791 10643 3825
rect 10701 3791 10735 3825
rect 10793 3791 10827 3825
rect 10885 3791 10919 3825
rect 10977 3791 11011 3825
rect 11069 3791 11103 3825
rect 11161 3791 11195 3825
rect 11253 3791 11287 3825
rect 11345 3791 11379 3825
rect 11437 3791 11471 3825
rect 11529 3791 11563 3825
rect 11621 3791 11655 3825
rect 11713 3791 11747 3825
rect 11805 3791 11839 3825
rect 11897 3791 11931 3825
rect 11989 3791 12023 3825
rect 12081 3791 12115 3825
rect 12173 3791 12207 3825
rect 12265 3791 12299 3825
rect 12357 3791 12391 3825
rect 12449 3791 12483 3825
rect 12541 3791 12575 3825
rect 12633 3791 12667 3825
rect 12725 3791 12759 3825
rect 12817 3791 12851 3825
rect 12909 3791 12943 3825
rect 13001 3791 13035 3825
rect 13093 3791 13127 3825
rect 13185 3791 13219 3825
rect 13277 3791 13311 3825
rect 13369 3791 13403 3825
rect 13461 3791 13495 3825
rect 13553 3791 13587 3825
rect 13645 3791 13679 3825
rect 13737 3791 13771 3825
rect 13829 3791 13863 3825
rect 13921 3791 13955 3825
rect 14013 3791 14047 3825
rect 14105 3791 14139 3825
rect 14197 3791 14231 3825
rect 14289 3791 14323 3825
rect 14381 3791 14415 3825
rect 14473 3791 14507 3825
rect 14565 3791 14599 3825
rect 14657 3791 14691 3825
rect 14749 3791 14783 3825
rect 14841 3791 14875 3825
rect 14933 3791 14967 3825
rect 15025 3791 15059 3825
rect 15117 3791 15151 3825
rect 15209 3791 15243 3825
rect 15301 3791 15335 3825
rect 15393 3791 15427 3825
rect 15485 3791 15519 3825
rect 15577 3791 15611 3825
rect 15669 3791 15703 3825
rect 15761 3791 15795 3825
rect 15853 3791 15887 3825
rect 15945 3791 15979 3825
rect 16037 3791 16071 3825
rect 16129 3791 16163 3825
rect 16221 3791 16255 3825
rect 16313 3791 16347 3825
rect 16405 3791 16439 3825
rect 16497 3791 16531 3825
rect 16589 3791 16623 3825
rect 16681 3791 16715 3825
rect 16773 3791 16807 3825
rect 16865 3791 16899 3825
rect 16957 3791 16991 3825
rect 17049 3791 17083 3825
rect 17141 3791 17175 3825
rect 17233 3791 17267 3825
rect 17325 3791 17359 3825
rect 17417 3791 17451 3825
rect 17509 3791 17543 3825
rect 17601 3791 17635 3825
rect 17693 3791 17727 3825
rect 17785 3791 17819 3825
rect 17877 3791 17911 3825
rect 17969 3791 18003 3825
rect 18061 3791 18095 3825
rect 18153 3791 18187 3825
rect 18245 3791 18279 3825
rect 18337 3791 18371 3825
rect 18429 3791 18463 3825
rect 18521 3791 18555 3825
rect 18613 3791 18647 3825
rect 18705 3791 18739 3825
rect 18797 3791 18831 3825
rect 2150 3621 2184 3655
rect 2053 3513 2087 3519
rect 2053 3485 2056 3513
rect 2056 3485 2087 3513
rect 2229 3553 2263 3587
rect 2320 3417 2354 3451
rect 2570 3629 2604 3655
rect 2570 3621 2572 3629
rect 2572 3621 2604 3629
rect 2467 3553 2501 3587
rect 2884 3621 2918 3655
rect 2971 3553 3005 3587
rect 3433 3709 3451 3723
rect 3451 3709 3467 3723
rect 3433 3689 3467 3709
rect 4082 3621 4116 3655
rect 3985 3553 4019 3587
rect 4161 3553 4195 3587
rect 4252 3485 4286 3519
rect 4502 3629 4536 3655
rect 4502 3621 4504 3629
rect 4504 3621 4536 3629
rect 4399 3553 4433 3587
rect 4816 3621 4850 3655
rect 4903 3553 4937 3587
rect 6653 3689 6687 3723
rect 7302 3621 7336 3655
rect 6469 3485 6503 3519
rect 6745 3513 6779 3519
rect 6745 3485 6775 3513
rect 6775 3485 6779 3513
rect 5365 3360 5399 3383
rect 5365 3349 5385 3360
rect 5385 3349 5399 3360
rect 6285 3428 6319 3451
rect 6285 3417 6291 3428
rect 6291 3417 6319 3428
rect 7205 3553 7239 3587
rect 7381 3553 7415 3587
rect 7472 3485 7506 3519
rect 7722 3629 7756 3655
rect 7722 3621 7724 3629
rect 7724 3621 7756 3629
rect 7619 3553 7653 3587
rect 8036 3621 8070 3655
rect 8123 3553 8157 3587
rect 8585 3709 8603 3723
rect 8603 3709 8619 3723
rect 8585 3689 8619 3709
rect 9878 3621 9912 3655
rect 9781 3553 9815 3587
rect 9957 3553 9991 3587
rect 10048 3485 10082 3519
rect 10298 3629 10332 3655
rect 10298 3621 10300 3629
rect 10300 3621 10332 3629
rect 10195 3553 10229 3587
rect 10612 3621 10646 3655
rect 10699 3553 10733 3587
rect 11161 3709 11179 3723
rect 11179 3709 11195 3723
rect 11161 3689 11195 3709
rect 11902 3621 11936 3655
rect 11805 3553 11839 3587
rect 11981 3553 12015 3587
rect 12072 3485 12106 3519
rect 12322 3629 12356 3655
rect 12322 3621 12324 3629
rect 12324 3621 12356 3629
rect 12219 3553 12253 3587
rect 12636 3621 12670 3655
rect 12723 3553 12757 3587
rect 13185 3709 13203 3723
rect 13203 3709 13219 3723
rect 13185 3689 13219 3709
rect 15945 3513 15979 3519
rect 15945 3485 15971 3513
rect 15971 3485 15979 3513
rect 16405 3485 16439 3519
rect 15761 3353 15767 3383
rect 15767 3353 15795 3383
rect 15761 3349 15795 3353
rect 16589 3513 16623 3519
rect 16589 3485 16621 3513
rect 16621 3485 16623 3513
rect 16681 3485 16715 3519
rect 17601 3553 17635 3587
rect 17417 3513 17451 3519
rect 17417 3485 17449 3513
rect 17449 3485 17451 3513
rect 17233 3349 17267 3383
rect 1133 3247 1167 3281
rect 1225 3247 1259 3281
rect 1317 3247 1351 3281
rect 1409 3247 1443 3281
rect 1501 3247 1535 3281
rect 1593 3247 1627 3281
rect 1685 3247 1719 3281
rect 1777 3247 1811 3281
rect 1869 3247 1903 3281
rect 1961 3247 1995 3281
rect 2053 3247 2087 3281
rect 2145 3247 2179 3281
rect 2237 3247 2271 3281
rect 2329 3247 2363 3281
rect 2421 3247 2455 3281
rect 2513 3247 2547 3281
rect 2605 3247 2639 3281
rect 2697 3247 2731 3281
rect 2789 3247 2823 3281
rect 2881 3247 2915 3281
rect 2973 3247 3007 3281
rect 3065 3247 3099 3281
rect 3157 3247 3191 3281
rect 3249 3247 3283 3281
rect 3341 3247 3375 3281
rect 3433 3247 3467 3281
rect 3525 3247 3559 3281
rect 3617 3247 3651 3281
rect 3709 3247 3743 3281
rect 3801 3247 3835 3281
rect 3893 3247 3927 3281
rect 3985 3247 4019 3281
rect 4077 3247 4111 3281
rect 4169 3247 4203 3281
rect 4261 3247 4295 3281
rect 4353 3247 4387 3281
rect 4445 3247 4479 3281
rect 4537 3247 4571 3281
rect 4629 3247 4663 3281
rect 4721 3247 4755 3281
rect 4813 3247 4847 3281
rect 4905 3247 4939 3281
rect 4997 3247 5031 3281
rect 5089 3247 5123 3281
rect 5181 3247 5215 3281
rect 5273 3247 5307 3281
rect 5365 3247 5399 3281
rect 5457 3247 5491 3281
rect 5549 3247 5583 3281
rect 5641 3247 5675 3281
rect 5733 3247 5767 3281
rect 5825 3247 5859 3281
rect 5917 3247 5951 3281
rect 6009 3247 6043 3281
rect 6101 3247 6135 3281
rect 6193 3247 6227 3281
rect 6285 3247 6319 3281
rect 6377 3247 6411 3281
rect 6469 3247 6503 3281
rect 6561 3247 6595 3281
rect 6653 3247 6687 3281
rect 6745 3247 6779 3281
rect 6837 3247 6871 3281
rect 6929 3247 6963 3281
rect 7021 3247 7055 3281
rect 7113 3247 7147 3281
rect 7205 3247 7239 3281
rect 7297 3247 7331 3281
rect 7389 3247 7423 3281
rect 7481 3247 7515 3281
rect 7573 3247 7607 3281
rect 7665 3247 7699 3281
rect 7757 3247 7791 3281
rect 7849 3247 7883 3281
rect 7941 3247 7975 3281
rect 8033 3247 8067 3281
rect 8125 3247 8159 3281
rect 8217 3247 8251 3281
rect 8309 3247 8343 3281
rect 8401 3247 8435 3281
rect 8493 3247 8527 3281
rect 8585 3247 8619 3281
rect 8677 3247 8711 3281
rect 8769 3247 8803 3281
rect 8861 3247 8895 3281
rect 8953 3247 8987 3281
rect 9045 3247 9079 3281
rect 9137 3247 9171 3281
rect 9229 3247 9263 3281
rect 9321 3247 9355 3281
rect 9413 3247 9447 3281
rect 9505 3247 9539 3281
rect 9597 3247 9631 3281
rect 9689 3247 9723 3281
rect 9781 3247 9815 3281
rect 9873 3247 9907 3281
rect 9965 3247 9999 3281
rect 10057 3247 10091 3281
rect 10149 3247 10183 3281
rect 10241 3247 10275 3281
rect 10333 3247 10367 3281
rect 10425 3247 10459 3281
rect 10517 3247 10551 3281
rect 10609 3247 10643 3281
rect 10701 3247 10735 3281
rect 10793 3247 10827 3281
rect 10885 3247 10919 3281
rect 10977 3247 11011 3281
rect 11069 3247 11103 3281
rect 11161 3247 11195 3281
rect 11253 3247 11287 3281
rect 11345 3247 11379 3281
rect 11437 3247 11471 3281
rect 11529 3247 11563 3281
rect 11621 3247 11655 3281
rect 11713 3247 11747 3281
rect 11805 3247 11839 3281
rect 11897 3247 11931 3281
rect 11989 3247 12023 3281
rect 12081 3247 12115 3281
rect 12173 3247 12207 3281
rect 12265 3247 12299 3281
rect 12357 3247 12391 3281
rect 12449 3247 12483 3281
rect 12541 3247 12575 3281
rect 12633 3247 12667 3281
rect 12725 3247 12759 3281
rect 12817 3247 12851 3281
rect 12909 3247 12943 3281
rect 13001 3247 13035 3281
rect 13093 3247 13127 3281
rect 13185 3247 13219 3281
rect 13277 3247 13311 3281
rect 13369 3247 13403 3281
rect 13461 3247 13495 3281
rect 13553 3247 13587 3281
rect 13645 3247 13679 3281
rect 13737 3247 13771 3281
rect 13829 3247 13863 3281
rect 13921 3247 13955 3281
rect 14013 3247 14047 3281
rect 14105 3247 14139 3281
rect 14197 3247 14231 3281
rect 14289 3247 14323 3281
rect 14381 3247 14415 3281
rect 14473 3247 14507 3281
rect 14565 3247 14599 3281
rect 14657 3247 14691 3281
rect 14749 3247 14783 3281
rect 14841 3247 14875 3281
rect 14933 3247 14967 3281
rect 15025 3247 15059 3281
rect 15117 3247 15151 3281
rect 15209 3247 15243 3281
rect 15301 3247 15335 3281
rect 15393 3247 15427 3281
rect 15485 3247 15519 3281
rect 15577 3247 15611 3281
rect 15669 3247 15703 3281
rect 15761 3247 15795 3281
rect 15853 3247 15887 3281
rect 15945 3247 15979 3281
rect 16037 3247 16071 3281
rect 16129 3247 16163 3281
rect 16221 3247 16255 3281
rect 16313 3247 16347 3281
rect 16405 3247 16439 3281
rect 16497 3247 16531 3281
rect 16589 3247 16623 3281
rect 16681 3247 16715 3281
rect 16773 3247 16807 3281
rect 16865 3247 16899 3281
rect 16957 3247 16991 3281
rect 17049 3247 17083 3281
rect 17141 3247 17175 3281
rect 17233 3247 17267 3281
rect 17325 3247 17359 3281
rect 17417 3247 17451 3281
rect 17509 3247 17543 3281
rect 17601 3247 17635 3281
rect 17693 3247 17727 3281
rect 17785 3247 17819 3281
rect 17877 3247 17911 3281
rect 17969 3247 18003 3281
rect 18061 3247 18095 3281
rect 18153 3247 18187 3281
rect 18245 3247 18279 3281
rect 18337 3247 18371 3281
rect 18429 3247 18463 3281
rect 18521 3247 18555 3281
rect 18613 3247 18647 3281
rect 18705 3247 18739 3281
rect 18797 3247 18831 3281
rect 2145 3077 2179 3111
rect 1961 3015 1963 3043
rect 1963 3015 1995 3043
rect 1961 3009 1995 3015
rect 3065 3158 3092 3179
rect 3092 3158 3099 3179
rect 3065 3145 3099 3158
rect 4353 3077 4387 3111
rect 7297 3009 7331 3043
rect 7757 3015 7765 3043
rect 7765 3015 7791 3043
rect 7757 3009 7791 3015
rect 9045 3158 9052 3179
rect 9052 3158 9079 3179
rect 9045 3145 9079 3158
rect 11713 3015 11716 3043
rect 11716 3015 11747 3043
rect 11713 3009 11747 3015
rect 11810 2873 11844 2907
rect 11889 2941 11923 2975
rect 11958 3077 11992 3111
rect 12127 2941 12161 2975
rect 12230 2899 12232 2907
rect 12232 2899 12264 2907
rect 12230 2873 12264 2899
rect 12544 2873 12578 2907
rect 12631 2941 12665 2975
rect 13093 3168 13113 3179
rect 13113 3168 13127 3179
rect 13093 3145 13127 3168
rect 17049 3015 17075 3043
rect 17075 3015 17083 3043
rect 17049 3009 17083 3015
rect 16865 2821 16899 2839
rect 16865 2805 16871 2821
rect 16871 2805 16899 2821
rect 1133 2703 1167 2737
rect 1225 2703 1259 2737
rect 1317 2703 1351 2737
rect 1409 2703 1443 2737
rect 1501 2703 1535 2737
rect 1593 2703 1627 2737
rect 1685 2703 1719 2737
rect 1777 2703 1811 2737
rect 1869 2703 1903 2737
rect 1961 2703 1995 2737
rect 2053 2703 2087 2737
rect 2145 2703 2179 2737
rect 2237 2703 2271 2737
rect 2329 2703 2363 2737
rect 2421 2703 2455 2737
rect 2513 2703 2547 2737
rect 2605 2703 2639 2737
rect 2697 2703 2731 2737
rect 2789 2703 2823 2737
rect 2881 2703 2915 2737
rect 2973 2703 3007 2737
rect 3065 2703 3099 2737
rect 3157 2703 3191 2737
rect 3249 2703 3283 2737
rect 3341 2703 3375 2737
rect 3433 2703 3467 2737
rect 3525 2703 3559 2737
rect 3617 2703 3651 2737
rect 3709 2703 3743 2737
rect 3801 2703 3835 2737
rect 3893 2703 3927 2737
rect 3985 2703 4019 2737
rect 4077 2703 4111 2737
rect 4169 2703 4203 2737
rect 4261 2703 4295 2737
rect 4353 2703 4387 2737
rect 4445 2703 4479 2737
rect 4537 2703 4571 2737
rect 4629 2703 4663 2737
rect 4721 2703 4755 2737
rect 4813 2703 4847 2737
rect 4905 2703 4939 2737
rect 4997 2703 5031 2737
rect 5089 2703 5123 2737
rect 5181 2703 5215 2737
rect 5273 2703 5307 2737
rect 5365 2703 5399 2737
rect 5457 2703 5491 2737
rect 5549 2703 5583 2737
rect 5641 2703 5675 2737
rect 5733 2703 5767 2737
rect 5825 2703 5859 2737
rect 5917 2703 5951 2737
rect 6009 2703 6043 2737
rect 6101 2703 6135 2737
rect 6193 2703 6227 2737
rect 6285 2703 6319 2737
rect 6377 2703 6411 2737
rect 6469 2703 6503 2737
rect 6561 2703 6595 2737
rect 6653 2703 6687 2737
rect 6745 2703 6779 2737
rect 6837 2703 6871 2737
rect 6929 2703 6963 2737
rect 7021 2703 7055 2737
rect 7113 2703 7147 2737
rect 7205 2703 7239 2737
rect 7297 2703 7331 2737
rect 7389 2703 7423 2737
rect 7481 2703 7515 2737
rect 7573 2703 7607 2737
rect 7665 2703 7699 2737
rect 7757 2703 7791 2737
rect 7849 2703 7883 2737
rect 7941 2703 7975 2737
rect 8033 2703 8067 2737
rect 8125 2703 8159 2737
rect 8217 2703 8251 2737
rect 8309 2703 8343 2737
rect 8401 2703 8435 2737
rect 8493 2703 8527 2737
rect 8585 2703 8619 2737
rect 8677 2703 8711 2737
rect 8769 2703 8803 2737
rect 8861 2703 8895 2737
rect 8953 2703 8987 2737
rect 9045 2703 9079 2737
rect 9137 2703 9171 2737
rect 9229 2703 9263 2737
rect 9321 2703 9355 2737
rect 9413 2703 9447 2737
rect 9505 2703 9539 2737
rect 9597 2703 9631 2737
rect 9689 2703 9723 2737
rect 9781 2703 9815 2737
rect 9873 2703 9907 2737
rect 9965 2703 9999 2737
rect 10057 2703 10091 2737
rect 10149 2703 10183 2737
rect 10241 2703 10275 2737
rect 10333 2703 10367 2737
rect 10425 2703 10459 2737
rect 10517 2703 10551 2737
rect 10609 2703 10643 2737
rect 10701 2703 10735 2737
rect 10793 2703 10827 2737
rect 10885 2703 10919 2737
rect 10977 2703 11011 2737
rect 11069 2703 11103 2737
rect 11161 2703 11195 2737
rect 11253 2703 11287 2737
rect 11345 2703 11379 2737
rect 11437 2703 11471 2737
rect 11529 2703 11563 2737
rect 11621 2703 11655 2737
rect 11713 2703 11747 2737
rect 11805 2703 11839 2737
rect 11897 2703 11931 2737
rect 11989 2703 12023 2737
rect 12081 2703 12115 2737
rect 12173 2703 12207 2737
rect 12265 2703 12299 2737
rect 12357 2703 12391 2737
rect 12449 2703 12483 2737
rect 12541 2703 12575 2737
rect 12633 2703 12667 2737
rect 12725 2703 12759 2737
rect 12817 2703 12851 2737
rect 12909 2703 12943 2737
rect 13001 2703 13035 2737
rect 13093 2703 13127 2737
rect 13185 2703 13219 2737
rect 13277 2703 13311 2737
rect 13369 2703 13403 2737
rect 13461 2703 13495 2737
rect 13553 2703 13587 2737
rect 13645 2703 13679 2737
rect 13737 2703 13771 2737
rect 13829 2703 13863 2737
rect 13921 2703 13955 2737
rect 14013 2703 14047 2737
rect 14105 2703 14139 2737
rect 14197 2703 14231 2737
rect 14289 2703 14323 2737
rect 14381 2703 14415 2737
rect 14473 2703 14507 2737
rect 14565 2703 14599 2737
rect 14657 2703 14691 2737
rect 14749 2703 14783 2737
rect 14841 2703 14875 2737
rect 14933 2703 14967 2737
rect 15025 2703 15059 2737
rect 15117 2703 15151 2737
rect 15209 2703 15243 2737
rect 15301 2703 15335 2737
rect 15393 2703 15427 2737
rect 15485 2703 15519 2737
rect 15577 2703 15611 2737
rect 15669 2703 15703 2737
rect 15761 2703 15795 2737
rect 15853 2703 15887 2737
rect 15945 2703 15979 2737
rect 16037 2703 16071 2737
rect 16129 2703 16163 2737
rect 16221 2703 16255 2737
rect 16313 2703 16347 2737
rect 16405 2703 16439 2737
rect 16497 2703 16531 2737
rect 16589 2703 16623 2737
rect 16681 2703 16715 2737
rect 16773 2703 16807 2737
rect 16865 2703 16899 2737
rect 16957 2703 16991 2737
rect 17049 2703 17083 2737
rect 17141 2703 17175 2737
rect 17233 2703 17267 2737
rect 17325 2703 17359 2737
rect 17417 2703 17451 2737
rect 17509 2703 17543 2737
rect 17601 2703 17635 2737
rect 17693 2703 17727 2737
rect 17785 2703 17819 2737
rect 17877 2703 17911 2737
rect 17969 2703 18003 2737
rect 18061 2703 18095 2737
rect 18153 2703 18187 2737
rect 18245 2703 18279 2737
rect 18337 2703 18371 2737
rect 18429 2703 18463 2737
rect 18521 2703 18555 2737
rect 18613 2703 18647 2737
rect 18705 2703 18739 2737
rect 18797 2703 18831 2737
rect 2053 2621 2069 2635
rect 2069 2621 2087 2635
rect 2053 2601 2087 2621
rect 2515 2465 2549 2499
rect 2602 2533 2636 2567
rect 2916 2541 2950 2567
rect 2916 2533 2948 2541
rect 2948 2533 2950 2541
rect 3019 2465 3053 2499
rect 3177 2397 3211 2431
rect 3257 2465 3291 2499
rect 3336 2533 3370 2567
rect 3433 2465 3467 2499
rect 4726 2533 4760 2567
rect 3985 2267 4019 2295
rect 3985 2261 3991 2267
rect 3991 2261 4019 2267
rect 4629 2465 4663 2499
rect 4805 2465 4839 2499
rect 4874 2329 4908 2363
rect 5146 2541 5180 2567
rect 5146 2533 5148 2541
rect 5148 2533 5180 2541
rect 5043 2465 5077 2499
rect 5460 2533 5494 2567
rect 5547 2465 5581 2499
rect 6009 2621 6027 2635
rect 6027 2621 6043 2635
rect 6009 2601 6043 2621
rect 7205 2272 7239 2295
rect 7205 2261 7219 2272
rect 7219 2261 7239 2272
rect 7667 2465 7701 2499
rect 7754 2533 7788 2567
rect 8068 2541 8102 2567
rect 8068 2533 8100 2541
rect 8100 2533 8102 2541
rect 8171 2465 8205 2499
rect 8340 2329 8374 2363
rect 8409 2465 8443 2499
rect 8488 2533 8522 2567
rect 9878 2533 9912 2567
rect 8585 2425 8619 2431
rect 8585 2397 8616 2425
rect 8616 2397 8619 2425
rect 9781 2425 9815 2431
rect 9781 2397 9784 2425
rect 9784 2397 9815 2425
rect 9957 2465 9991 2499
rect 10048 2329 10082 2363
rect 10298 2541 10332 2567
rect 10298 2533 10300 2541
rect 10300 2533 10332 2541
rect 10195 2465 10229 2499
rect 10612 2533 10646 2567
rect 10699 2465 10733 2499
rect 11161 2553 11179 2567
rect 11179 2553 11195 2567
rect 11161 2533 11195 2553
rect 11897 2621 11913 2635
rect 11913 2621 11931 2635
rect 11897 2601 11931 2621
rect 12359 2465 12393 2499
rect 12446 2533 12480 2567
rect 12760 2541 12794 2567
rect 12760 2533 12792 2541
rect 12792 2533 12794 2541
rect 12863 2465 12897 2499
rect 13032 2329 13066 2363
rect 13101 2465 13135 2499
rect 13180 2533 13214 2567
rect 13277 2425 13311 2431
rect 13277 2397 13308 2425
rect 13308 2397 13311 2425
rect 14289 2601 14323 2635
rect 16865 2619 16871 2635
rect 16871 2619 16899 2635
rect 16865 2601 16899 2619
rect 17049 2425 17083 2431
rect 17049 2397 17075 2425
rect 17075 2397 17083 2425
rect 17509 2425 17543 2431
rect 17509 2397 17517 2425
rect 17517 2397 17543 2425
rect 17693 2265 17694 2295
rect 17694 2265 17727 2295
rect 17693 2261 17727 2265
rect 1133 2159 1167 2193
rect 1225 2159 1259 2193
rect 1317 2159 1351 2193
rect 1409 2159 1443 2193
rect 1501 2159 1535 2193
rect 1593 2159 1627 2193
rect 1685 2159 1719 2193
rect 1777 2159 1811 2193
rect 1869 2159 1903 2193
rect 1961 2159 1995 2193
rect 2053 2159 2087 2193
rect 2145 2159 2179 2193
rect 2237 2159 2271 2193
rect 2329 2159 2363 2193
rect 2421 2159 2455 2193
rect 2513 2159 2547 2193
rect 2605 2159 2639 2193
rect 2697 2159 2731 2193
rect 2789 2159 2823 2193
rect 2881 2159 2915 2193
rect 2973 2159 3007 2193
rect 3065 2159 3099 2193
rect 3157 2159 3191 2193
rect 3249 2159 3283 2193
rect 3341 2159 3375 2193
rect 3433 2159 3467 2193
rect 3525 2159 3559 2193
rect 3617 2159 3651 2193
rect 3709 2159 3743 2193
rect 3801 2159 3835 2193
rect 3893 2159 3927 2193
rect 3985 2159 4019 2193
rect 4077 2159 4111 2193
rect 4169 2159 4203 2193
rect 4261 2159 4295 2193
rect 4353 2159 4387 2193
rect 4445 2159 4479 2193
rect 4537 2159 4571 2193
rect 4629 2159 4663 2193
rect 4721 2159 4755 2193
rect 4813 2159 4847 2193
rect 4905 2159 4939 2193
rect 4997 2159 5031 2193
rect 5089 2159 5123 2193
rect 5181 2159 5215 2193
rect 5273 2159 5307 2193
rect 5365 2159 5399 2193
rect 5457 2159 5491 2193
rect 5549 2159 5583 2193
rect 5641 2159 5675 2193
rect 5733 2159 5767 2193
rect 5825 2159 5859 2193
rect 5917 2159 5951 2193
rect 6009 2159 6043 2193
rect 6101 2159 6135 2193
rect 6193 2159 6227 2193
rect 6285 2159 6319 2193
rect 6377 2159 6411 2193
rect 6469 2159 6503 2193
rect 6561 2159 6595 2193
rect 6653 2159 6687 2193
rect 6745 2159 6779 2193
rect 6837 2159 6871 2193
rect 6929 2159 6963 2193
rect 7021 2159 7055 2193
rect 7113 2159 7147 2193
rect 7205 2159 7239 2193
rect 7297 2159 7331 2193
rect 7389 2159 7423 2193
rect 7481 2159 7515 2193
rect 7573 2159 7607 2193
rect 7665 2159 7699 2193
rect 7757 2159 7791 2193
rect 7849 2159 7883 2193
rect 7941 2159 7975 2193
rect 8033 2159 8067 2193
rect 8125 2159 8159 2193
rect 8217 2159 8251 2193
rect 8309 2159 8343 2193
rect 8401 2159 8435 2193
rect 8493 2159 8527 2193
rect 8585 2159 8619 2193
rect 8677 2159 8711 2193
rect 8769 2159 8803 2193
rect 8861 2159 8895 2193
rect 8953 2159 8987 2193
rect 9045 2159 9079 2193
rect 9137 2159 9171 2193
rect 9229 2159 9263 2193
rect 9321 2159 9355 2193
rect 9413 2159 9447 2193
rect 9505 2159 9539 2193
rect 9597 2159 9631 2193
rect 9689 2159 9723 2193
rect 9781 2159 9815 2193
rect 9873 2159 9907 2193
rect 9965 2159 9999 2193
rect 10057 2159 10091 2193
rect 10149 2159 10183 2193
rect 10241 2159 10275 2193
rect 10333 2159 10367 2193
rect 10425 2159 10459 2193
rect 10517 2159 10551 2193
rect 10609 2159 10643 2193
rect 10701 2159 10735 2193
rect 10793 2159 10827 2193
rect 10885 2159 10919 2193
rect 10977 2159 11011 2193
rect 11069 2159 11103 2193
rect 11161 2159 11195 2193
rect 11253 2159 11287 2193
rect 11345 2159 11379 2193
rect 11437 2159 11471 2193
rect 11529 2159 11563 2193
rect 11621 2159 11655 2193
rect 11713 2159 11747 2193
rect 11805 2159 11839 2193
rect 11897 2159 11931 2193
rect 11989 2159 12023 2193
rect 12081 2159 12115 2193
rect 12173 2159 12207 2193
rect 12265 2159 12299 2193
rect 12357 2159 12391 2193
rect 12449 2159 12483 2193
rect 12541 2159 12575 2193
rect 12633 2159 12667 2193
rect 12725 2159 12759 2193
rect 12817 2159 12851 2193
rect 12909 2159 12943 2193
rect 13001 2159 13035 2193
rect 13093 2159 13127 2193
rect 13185 2159 13219 2193
rect 13277 2159 13311 2193
rect 13369 2159 13403 2193
rect 13461 2159 13495 2193
rect 13553 2159 13587 2193
rect 13645 2159 13679 2193
rect 13737 2159 13771 2193
rect 13829 2159 13863 2193
rect 13921 2159 13955 2193
rect 14013 2159 14047 2193
rect 14105 2159 14139 2193
rect 14197 2159 14231 2193
rect 14289 2159 14323 2193
rect 14381 2159 14415 2193
rect 14473 2159 14507 2193
rect 14565 2159 14599 2193
rect 14657 2159 14691 2193
rect 14749 2159 14783 2193
rect 14841 2159 14875 2193
rect 14933 2159 14967 2193
rect 15025 2159 15059 2193
rect 15117 2159 15151 2193
rect 15209 2159 15243 2193
rect 15301 2159 15335 2193
rect 15393 2159 15427 2193
rect 15485 2159 15519 2193
rect 15577 2159 15611 2193
rect 15669 2159 15703 2193
rect 15761 2159 15795 2193
rect 15853 2159 15887 2193
rect 15945 2159 15979 2193
rect 16037 2159 16071 2193
rect 16129 2159 16163 2193
rect 16221 2159 16255 2193
rect 16313 2159 16347 2193
rect 16405 2159 16439 2193
rect 16497 2159 16531 2193
rect 16589 2159 16623 2193
rect 16681 2159 16715 2193
rect 16773 2159 16807 2193
rect 16865 2159 16899 2193
rect 16957 2159 16991 2193
rect 17049 2159 17083 2193
rect 17141 2159 17175 2193
rect 17233 2159 17267 2193
rect 17325 2159 17359 2193
rect 17417 2159 17451 2193
rect 17509 2159 17543 2193
rect 17601 2159 17635 2193
rect 17693 2159 17727 2193
rect 17785 2159 17819 2193
rect 17877 2159 17911 2193
rect 17969 2159 18003 2193
rect 18061 2159 18095 2193
rect 18153 2159 18187 2193
rect 18245 2159 18279 2193
rect 18337 2159 18371 2193
rect 18429 2159 18463 2193
rect 18521 2159 18555 2193
rect 18613 2159 18647 2193
rect 18705 2159 18739 2193
rect 18797 2159 18831 2193
<< metal1 >>
rect 1104 7642 19019 7664
rect 1104 7633 5388 7642
rect 1104 7599 1133 7633
rect 1167 7599 1225 7633
rect 1259 7599 1317 7633
rect 1351 7599 1409 7633
rect 1443 7599 1501 7633
rect 1535 7599 1593 7633
rect 1627 7599 1685 7633
rect 1719 7599 1777 7633
rect 1811 7599 1869 7633
rect 1903 7599 1961 7633
rect 1995 7599 2053 7633
rect 2087 7599 2145 7633
rect 2179 7599 2237 7633
rect 2271 7599 2329 7633
rect 2363 7599 2421 7633
rect 2455 7599 2513 7633
rect 2547 7599 2605 7633
rect 2639 7599 2697 7633
rect 2731 7599 2789 7633
rect 2823 7599 2881 7633
rect 2915 7599 2973 7633
rect 3007 7599 3065 7633
rect 3099 7599 3157 7633
rect 3191 7599 3249 7633
rect 3283 7599 3341 7633
rect 3375 7599 3433 7633
rect 3467 7599 3525 7633
rect 3559 7599 3617 7633
rect 3651 7599 3709 7633
rect 3743 7599 3801 7633
rect 3835 7599 3893 7633
rect 3927 7599 3985 7633
rect 4019 7599 4077 7633
rect 4111 7599 4169 7633
rect 4203 7599 4261 7633
rect 4295 7599 4353 7633
rect 4387 7599 4445 7633
rect 4479 7599 4537 7633
rect 4571 7599 4629 7633
rect 4663 7599 4721 7633
rect 4755 7599 4813 7633
rect 4847 7599 4905 7633
rect 4939 7599 4997 7633
rect 5031 7599 5089 7633
rect 5123 7599 5181 7633
rect 5215 7599 5273 7633
rect 5307 7599 5365 7633
rect 1104 7590 5388 7599
rect 5440 7590 5452 7642
rect 5504 7590 5516 7642
rect 5568 7633 5580 7642
rect 5632 7633 5644 7642
rect 5696 7633 9827 7642
rect 9879 7633 9891 7642
rect 5632 7599 5641 7633
rect 5696 7599 5733 7633
rect 5767 7599 5825 7633
rect 5859 7599 5917 7633
rect 5951 7599 6009 7633
rect 6043 7599 6101 7633
rect 6135 7599 6193 7633
rect 6227 7599 6285 7633
rect 6319 7599 6377 7633
rect 6411 7599 6469 7633
rect 6503 7599 6561 7633
rect 6595 7599 6653 7633
rect 6687 7599 6745 7633
rect 6779 7599 6837 7633
rect 6871 7599 6929 7633
rect 6963 7599 7021 7633
rect 7055 7599 7113 7633
rect 7147 7599 7205 7633
rect 7239 7599 7297 7633
rect 7331 7599 7389 7633
rect 7423 7599 7481 7633
rect 7515 7599 7573 7633
rect 7607 7599 7665 7633
rect 7699 7599 7757 7633
rect 7791 7599 7849 7633
rect 7883 7599 7941 7633
rect 7975 7599 8033 7633
rect 8067 7599 8125 7633
rect 8159 7599 8217 7633
rect 8251 7599 8309 7633
rect 8343 7599 8401 7633
rect 8435 7599 8493 7633
rect 8527 7599 8585 7633
rect 8619 7599 8677 7633
rect 8711 7599 8769 7633
rect 8803 7599 8861 7633
rect 8895 7599 8953 7633
rect 8987 7599 9045 7633
rect 9079 7599 9137 7633
rect 9171 7599 9229 7633
rect 9263 7599 9321 7633
rect 9355 7599 9413 7633
rect 9447 7599 9505 7633
rect 9539 7599 9597 7633
rect 9631 7599 9689 7633
rect 9723 7599 9781 7633
rect 9815 7599 9827 7633
rect 5568 7590 5580 7599
rect 5632 7590 5644 7599
rect 5696 7590 9827 7599
rect 9879 7590 9891 7599
rect 9943 7590 9955 7642
rect 10007 7590 10019 7642
rect 10071 7633 10083 7642
rect 10135 7633 14266 7642
rect 14318 7633 14330 7642
rect 14382 7633 14394 7642
rect 10135 7599 10149 7633
rect 10183 7599 10241 7633
rect 10275 7599 10333 7633
rect 10367 7599 10425 7633
rect 10459 7599 10517 7633
rect 10551 7599 10609 7633
rect 10643 7599 10701 7633
rect 10735 7599 10793 7633
rect 10827 7599 10885 7633
rect 10919 7599 10977 7633
rect 11011 7599 11069 7633
rect 11103 7599 11161 7633
rect 11195 7599 11253 7633
rect 11287 7599 11345 7633
rect 11379 7599 11437 7633
rect 11471 7599 11529 7633
rect 11563 7599 11621 7633
rect 11655 7599 11713 7633
rect 11747 7599 11805 7633
rect 11839 7599 11897 7633
rect 11931 7599 11989 7633
rect 12023 7599 12081 7633
rect 12115 7599 12173 7633
rect 12207 7599 12265 7633
rect 12299 7599 12357 7633
rect 12391 7599 12449 7633
rect 12483 7599 12541 7633
rect 12575 7599 12633 7633
rect 12667 7599 12725 7633
rect 12759 7599 12817 7633
rect 12851 7599 12909 7633
rect 12943 7599 13001 7633
rect 13035 7599 13093 7633
rect 13127 7599 13185 7633
rect 13219 7599 13277 7633
rect 13311 7599 13369 7633
rect 13403 7599 13461 7633
rect 13495 7599 13553 7633
rect 13587 7599 13645 7633
rect 13679 7599 13737 7633
rect 13771 7599 13829 7633
rect 13863 7599 13921 7633
rect 13955 7599 14013 7633
rect 14047 7599 14105 7633
rect 14139 7599 14197 7633
rect 14231 7599 14266 7633
rect 14323 7599 14330 7633
rect 10071 7590 10083 7599
rect 10135 7590 14266 7599
rect 14318 7590 14330 7599
rect 14382 7590 14394 7599
rect 14446 7590 14458 7642
rect 14510 7590 14522 7642
rect 14574 7633 18705 7642
rect 14599 7599 14657 7633
rect 14691 7599 14749 7633
rect 14783 7599 14841 7633
rect 14875 7599 14933 7633
rect 14967 7599 15025 7633
rect 15059 7599 15117 7633
rect 15151 7599 15209 7633
rect 15243 7599 15301 7633
rect 15335 7599 15393 7633
rect 15427 7599 15485 7633
rect 15519 7599 15577 7633
rect 15611 7599 15669 7633
rect 15703 7599 15761 7633
rect 15795 7599 15853 7633
rect 15887 7599 15945 7633
rect 15979 7599 16037 7633
rect 16071 7599 16129 7633
rect 16163 7599 16221 7633
rect 16255 7599 16313 7633
rect 16347 7599 16405 7633
rect 16439 7599 16497 7633
rect 16531 7599 16589 7633
rect 16623 7599 16681 7633
rect 16715 7599 16773 7633
rect 16807 7599 16865 7633
rect 16899 7599 16957 7633
rect 16991 7599 17049 7633
rect 17083 7599 17141 7633
rect 17175 7599 17233 7633
rect 17267 7599 17325 7633
rect 17359 7599 17417 7633
rect 17451 7599 17509 7633
rect 17543 7599 17601 7633
rect 17635 7599 17693 7633
rect 17727 7599 17785 7633
rect 17819 7599 17877 7633
rect 17911 7599 17969 7633
rect 18003 7599 18061 7633
rect 18095 7599 18153 7633
rect 18187 7599 18245 7633
rect 18279 7599 18337 7633
rect 18371 7599 18429 7633
rect 18463 7599 18521 7633
rect 18555 7599 18613 7633
rect 18647 7599 18705 7633
rect 14574 7590 18705 7599
rect 18757 7590 18769 7642
rect 18821 7633 18833 7642
rect 18831 7599 18833 7633
rect 18821 7590 18833 7599
rect 18885 7590 18897 7642
rect 18949 7590 18961 7642
rect 19013 7590 19019 7642
rect 1104 7568 19019 7590
rect 1118 7488 1124 7540
rect 1176 7528 1182 7540
rect 1673 7531 1731 7537
rect 1673 7528 1685 7531
rect 1176 7500 1685 7528
rect 1176 7488 1182 7500
rect 1673 7497 1685 7500
rect 1719 7497 1731 7531
rect 1673 7491 1731 7497
rect 3326 7488 3332 7540
rect 3384 7528 3390 7540
rect 4065 7531 4123 7537
rect 4065 7528 4077 7531
rect 3384 7500 4077 7528
rect 3384 7488 3390 7500
rect 4065 7497 4077 7500
rect 4111 7497 4123 7531
rect 5718 7528 5724 7540
rect 5679 7500 5724 7528
rect 4065 7491 4123 7497
rect 5718 7488 5724 7500
rect 5776 7488 5782 7540
rect 7742 7488 7748 7540
rect 7800 7528 7806 7540
rect 8021 7531 8079 7537
rect 8021 7528 8033 7531
rect 7800 7500 8033 7528
rect 7800 7488 7806 7500
rect 8021 7497 8033 7500
rect 8067 7497 8079 7531
rect 12434 7528 12440 7540
rect 12395 7500 12440 7528
rect 8021 7491 8079 7497
rect 12434 7488 12440 7500
rect 12492 7488 12498 7540
rect 14642 7528 14648 7540
rect 14603 7500 14648 7528
rect 14642 7488 14648 7500
rect 14700 7488 14706 7540
rect 16574 7488 16580 7540
rect 16632 7528 16638 7540
rect 17037 7531 17095 7537
rect 17037 7528 17049 7531
rect 16632 7500 17049 7528
rect 16632 7488 16638 7500
rect 17037 7497 17049 7500
rect 17083 7497 17095 7531
rect 17037 7491 17095 7497
rect 18233 7531 18291 7537
rect 18233 7497 18245 7531
rect 18279 7528 18291 7531
rect 18414 7528 18420 7540
rect 18279 7500 18420 7528
rect 18279 7497 18291 7500
rect 18233 7491 18291 7497
rect 18414 7488 18420 7500
rect 18472 7488 18478 7540
rect 9585 7463 9643 7469
rect 9585 7429 9597 7463
rect 9631 7460 9643 7463
rect 10137 7463 10195 7469
rect 10137 7460 10149 7463
rect 9631 7432 10149 7460
rect 9631 7429 9643 7432
rect 9585 7423 9643 7429
rect 10137 7429 10149 7432
rect 10183 7460 10195 7463
rect 10226 7460 10232 7472
rect 10183 7432 10232 7460
rect 10183 7429 10195 7432
rect 10137 7423 10195 7429
rect 10226 7420 10232 7432
rect 10284 7420 10290 7472
rect 1854 7392 1860 7404
rect 1815 7364 1860 7392
rect 1854 7352 1860 7364
rect 1912 7352 1918 7404
rect 4249 7395 4307 7401
rect 4249 7361 4261 7395
rect 4295 7392 4307 7395
rect 4614 7392 4620 7404
rect 4295 7364 4620 7392
rect 4295 7361 4307 7364
rect 4249 7355 4307 7361
rect 4614 7352 4620 7364
rect 4672 7352 4678 7404
rect 5905 7395 5963 7401
rect 5905 7361 5917 7395
rect 5951 7392 5963 7395
rect 6914 7392 6920 7404
rect 5951 7364 6920 7392
rect 5951 7361 5963 7364
rect 5905 7355 5963 7361
rect 6914 7352 6920 7364
rect 6972 7352 6978 7404
rect 7098 7352 7104 7404
rect 7156 7392 7162 7404
rect 7837 7395 7895 7401
rect 7837 7392 7849 7395
rect 7156 7364 7849 7392
rect 7156 7352 7162 7364
rect 7837 7361 7849 7364
rect 7883 7361 7895 7395
rect 7837 7355 7895 7361
rect 10594 7352 10600 7404
rect 10652 7392 10658 7404
rect 12253 7395 12311 7401
rect 12253 7392 12265 7395
rect 10652 7364 12265 7392
rect 10652 7352 10658 7364
rect 12253 7361 12265 7364
rect 12299 7361 12311 7395
rect 12253 7355 12311 7361
rect 12526 7352 12532 7404
rect 12584 7392 12590 7404
rect 14461 7395 14519 7401
rect 14461 7392 14473 7395
rect 12584 7364 14473 7392
rect 12584 7352 12590 7364
rect 14461 7361 14473 7364
rect 14507 7361 14519 7395
rect 14461 7355 14519 7361
rect 14642 7352 14648 7404
rect 14700 7392 14706 7404
rect 16853 7395 16911 7401
rect 16853 7392 16865 7395
rect 14700 7364 16865 7392
rect 14700 7352 14706 7364
rect 16853 7361 16865 7364
rect 16899 7361 16911 7395
rect 16853 7355 16911 7361
rect 18049 7395 18107 7401
rect 18049 7361 18061 7395
rect 18095 7361 18107 7395
rect 18049 7355 18107 7361
rect 13446 7284 13452 7336
rect 13504 7324 13510 7336
rect 18064 7324 18092 7355
rect 13504 7296 18092 7324
rect 13504 7284 13510 7296
rect 10318 7256 10324 7268
rect 10279 7228 10324 7256
rect 10318 7216 10324 7228
rect 10376 7216 10382 7268
rect 1104 7098 18860 7120
rect 1104 7089 3169 7098
rect 1104 7055 1133 7089
rect 1167 7055 1225 7089
rect 1259 7055 1317 7089
rect 1351 7055 1409 7089
rect 1443 7055 1501 7089
rect 1535 7055 1593 7089
rect 1627 7055 1685 7089
rect 1719 7055 1777 7089
rect 1811 7055 1869 7089
rect 1903 7055 1961 7089
rect 1995 7055 2053 7089
rect 2087 7055 2145 7089
rect 2179 7055 2237 7089
rect 2271 7055 2329 7089
rect 2363 7055 2421 7089
rect 2455 7055 2513 7089
rect 2547 7055 2605 7089
rect 2639 7055 2697 7089
rect 2731 7055 2789 7089
rect 2823 7055 2881 7089
rect 2915 7055 2973 7089
rect 3007 7055 3065 7089
rect 3099 7055 3157 7089
rect 1104 7046 3169 7055
rect 3221 7046 3233 7098
rect 3285 7046 3297 7098
rect 3349 7089 3361 7098
rect 3349 7046 3361 7055
rect 3413 7046 3425 7098
rect 3477 7089 7608 7098
rect 3477 7055 3525 7089
rect 3559 7055 3617 7089
rect 3651 7055 3709 7089
rect 3743 7055 3801 7089
rect 3835 7055 3893 7089
rect 3927 7055 3985 7089
rect 4019 7055 4077 7089
rect 4111 7055 4169 7089
rect 4203 7055 4261 7089
rect 4295 7055 4353 7089
rect 4387 7055 4445 7089
rect 4479 7055 4537 7089
rect 4571 7055 4629 7089
rect 4663 7055 4721 7089
rect 4755 7055 4813 7089
rect 4847 7055 4905 7089
rect 4939 7055 4997 7089
rect 5031 7055 5089 7089
rect 5123 7055 5181 7089
rect 5215 7055 5273 7089
rect 5307 7055 5365 7089
rect 5399 7055 5457 7089
rect 5491 7055 5549 7089
rect 5583 7055 5641 7089
rect 5675 7055 5733 7089
rect 5767 7055 5825 7089
rect 5859 7055 5917 7089
rect 5951 7055 6009 7089
rect 6043 7055 6101 7089
rect 6135 7055 6193 7089
rect 6227 7055 6285 7089
rect 6319 7055 6377 7089
rect 6411 7055 6469 7089
rect 6503 7055 6561 7089
rect 6595 7055 6653 7089
rect 6687 7055 6745 7089
rect 6779 7055 6837 7089
rect 6871 7055 6929 7089
rect 6963 7055 7021 7089
rect 7055 7055 7113 7089
rect 7147 7055 7205 7089
rect 7239 7055 7297 7089
rect 7331 7055 7389 7089
rect 7423 7055 7481 7089
rect 7515 7055 7573 7089
rect 7607 7055 7608 7089
rect 3477 7046 7608 7055
rect 7660 7089 7672 7098
rect 7660 7055 7665 7089
rect 7660 7046 7672 7055
rect 7724 7046 7736 7098
rect 7788 7089 7800 7098
rect 7852 7089 7864 7098
rect 7916 7089 12047 7098
rect 12099 7089 12111 7098
rect 12163 7089 12175 7098
rect 7791 7055 7800 7089
rect 7916 7055 7941 7089
rect 7975 7055 8033 7089
rect 8067 7055 8125 7089
rect 8159 7055 8217 7089
rect 8251 7055 8309 7089
rect 8343 7055 8401 7089
rect 8435 7055 8493 7089
rect 8527 7055 8585 7089
rect 8619 7055 8677 7089
rect 8711 7055 8769 7089
rect 8803 7055 8861 7089
rect 8895 7055 8953 7089
rect 8987 7055 9045 7089
rect 9079 7055 9137 7089
rect 9171 7055 9229 7089
rect 9263 7055 9321 7089
rect 9355 7055 9413 7089
rect 9447 7055 9505 7089
rect 9539 7055 9597 7089
rect 9631 7055 9689 7089
rect 9723 7055 9781 7089
rect 9815 7055 9873 7089
rect 9907 7055 9965 7089
rect 9999 7055 10057 7089
rect 10091 7055 10149 7089
rect 10183 7055 10241 7089
rect 10275 7055 10333 7089
rect 10367 7055 10425 7089
rect 10459 7055 10517 7089
rect 10551 7055 10609 7089
rect 10643 7055 10701 7089
rect 10735 7055 10793 7089
rect 10827 7055 10885 7089
rect 10919 7055 10977 7089
rect 11011 7055 11069 7089
rect 11103 7055 11161 7089
rect 11195 7055 11253 7089
rect 11287 7055 11345 7089
rect 11379 7055 11437 7089
rect 11471 7055 11529 7089
rect 11563 7055 11621 7089
rect 11655 7055 11713 7089
rect 11747 7055 11805 7089
rect 11839 7055 11897 7089
rect 11931 7055 11989 7089
rect 12023 7055 12047 7089
rect 12163 7055 12173 7089
rect 7788 7046 7800 7055
rect 7852 7046 7864 7055
rect 7916 7046 12047 7055
rect 12099 7046 12111 7055
rect 12163 7046 12175 7055
rect 12227 7046 12239 7098
rect 12291 7089 12303 7098
rect 12299 7055 12303 7089
rect 12291 7046 12303 7055
rect 12355 7089 16486 7098
rect 12355 7055 12357 7089
rect 12391 7055 12449 7089
rect 12483 7055 12541 7089
rect 12575 7055 12633 7089
rect 12667 7055 12725 7089
rect 12759 7055 12817 7089
rect 12851 7055 12909 7089
rect 12943 7055 13001 7089
rect 13035 7055 13093 7089
rect 13127 7055 13185 7089
rect 13219 7055 13277 7089
rect 13311 7055 13369 7089
rect 13403 7055 13461 7089
rect 13495 7055 13553 7089
rect 13587 7055 13645 7089
rect 13679 7055 13737 7089
rect 13771 7055 13829 7089
rect 13863 7055 13921 7089
rect 13955 7055 14013 7089
rect 14047 7055 14105 7089
rect 14139 7055 14197 7089
rect 14231 7055 14289 7089
rect 14323 7055 14381 7089
rect 14415 7055 14473 7089
rect 14507 7055 14565 7089
rect 14599 7055 14657 7089
rect 14691 7055 14749 7089
rect 14783 7055 14841 7089
rect 14875 7055 14933 7089
rect 14967 7055 15025 7089
rect 15059 7055 15117 7089
rect 15151 7055 15209 7089
rect 15243 7055 15301 7089
rect 15335 7055 15393 7089
rect 15427 7055 15485 7089
rect 15519 7055 15577 7089
rect 15611 7055 15669 7089
rect 15703 7055 15761 7089
rect 15795 7055 15853 7089
rect 15887 7055 15945 7089
rect 15979 7055 16037 7089
rect 16071 7055 16129 7089
rect 16163 7055 16221 7089
rect 16255 7055 16313 7089
rect 16347 7055 16405 7089
rect 16439 7055 16486 7089
rect 12355 7046 16486 7055
rect 16538 7046 16550 7098
rect 16602 7089 16614 7098
rect 16602 7046 16614 7055
rect 16666 7046 16678 7098
rect 16730 7046 16742 7098
rect 16794 7089 18860 7098
rect 16807 7055 16865 7089
rect 16899 7055 16957 7089
rect 16991 7055 17049 7089
rect 17083 7055 17141 7089
rect 17175 7055 17233 7089
rect 17267 7055 17325 7089
rect 17359 7055 17417 7089
rect 17451 7055 17509 7089
rect 17543 7055 17601 7089
rect 17635 7055 17693 7089
rect 17727 7055 17785 7089
rect 17819 7055 17877 7089
rect 17911 7055 17969 7089
rect 18003 7055 18061 7089
rect 18095 7055 18153 7089
rect 18187 7055 18245 7089
rect 18279 7055 18337 7089
rect 18371 7055 18429 7089
rect 18463 7055 18521 7089
rect 18555 7055 18613 7089
rect 18647 7055 18705 7089
rect 18739 7055 18797 7089
rect 18831 7055 18860 7089
rect 16794 7046 18860 7055
rect 1104 7024 18860 7046
rect 1104 6554 19019 6576
rect 1104 6545 5388 6554
rect 1104 6511 1133 6545
rect 1167 6511 1225 6545
rect 1259 6511 1317 6545
rect 1351 6511 1409 6545
rect 1443 6511 1501 6545
rect 1535 6511 1593 6545
rect 1627 6511 1685 6545
rect 1719 6511 1777 6545
rect 1811 6511 1869 6545
rect 1903 6511 1961 6545
rect 1995 6511 2053 6545
rect 2087 6511 2145 6545
rect 2179 6511 2237 6545
rect 2271 6511 2329 6545
rect 2363 6511 2421 6545
rect 2455 6511 2513 6545
rect 2547 6511 2605 6545
rect 2639 6511 2697 6545
rect 2731 6511 2789 6545
rect 2823 6511 2881 6545
rect 2915 6511 2973 6545
rect 3007 6511 3065 6545
rect 3099 6511 3157 6545
rect 3191 6511 3249 6545
rect 3283 6511 3341 6545
rect 3375 6511 3433 6545
rect 3467 6511 3525 6545
rect 3559 6511 3617 6545
rect 3651 6511 3709 6545
rect 3743 6511 3801 6545
rect 3835 6511 3893 6545
rect 3927 6511 3985 6545
rect 4019 6511 4077 6545
rect 4111 6511 4169 6545
rect 4203 6511 4261 6545
rect 4295 6511 4353 6545
rect 4387 6511 4445 6545
rect 4479 6511 4537 6545
rect 4571 6511 4629 6545
rect 4663 6511 4721 6545
rect 4755 6511 4813 6545
rect 4847 6511 4905 6545
rect 4939 6511 4997 6545
rect 5031 6511 5089 6545
rect 5123 6511 5181 6545
rect 5215 6511 5273 6545
rect 5307 6511 5365 6545
rect 1104 6502 5388 6511
rect 5440 6502 5452 6554
rect 5504 6502 5516 6554
rect 5568 6545 5580 6554
rect 5632 6545 5644 6554
rect 5696 6545 9827 6554
rect 9879 6545 9891 6554
rect 5632 6511 5641 6545
rect 5696 6511 5733 6545
rect 5767 6511 5825 6545
rect 5859 6511 5917 6545
rect 5951 6511 6009 6545
rect 6043 6511 6101 6545
rect 6135 6511 6193 6545
rect 6227 6511 6285 6545
rect 6319 6511 6377 6545
rect 6411 6511 6469 6545
rect 6503 6511 6561 6545
rect 6595 6511 6653 6545
rect 6687 6511 6745 6545
rect 6779 6511 6837 6545
rect 6871 6511 6929 6545
rect 6963 6511 7021 6545
rect 7055 6511 7113 6545
rect 7147 6511 7205 6545
rect 7239 6511 7297 6545
rect 7331 6511 7389 6545
rect 7423 6511 7481 6545
rect 7515 6511 7573 6545
rect 7607 6511 7665 6545
rect 7699 6511 7757 6545
rect 7791 6511 7849 6545
rect 7883 6511 7941 6545
rect 7975 6511 8033 6545
rect 8067 6511 8125 6545
rect 8159 6511 8217 6545
rect 8251 6511 8309 6545
rect 8343 6511 8401 6545
rect 8435 6511 8493 6545
rect 8527 6511 8585 6545
rect 8619 6511 8677 6545
rect 8711 6511 8769 6545
rect 8803 6511 8861 6545
rect 8895 6511 8953 6545
rect 8987 6511 9045 6545
rect 9079 6511 9137 6545
rect 9171 6511 9229 6545
rect 9263 6511 9321 6545
rect 9355 6511 9413 6545
rect 9447 6511 9505 6545
rect 9539 6511 9597 6545
rect 9631 6511 9689 6545
rect 9723 6511 9781 6545
rect 9815 6511 9827 6545
rect 5568 6502 5580 6511
rect 5632 6502 5644 6511
rect 5696 6502 9827 6511
rect 9879 6502 9891 6511
rect 9943 6502 9955 6554
rect 10007 6502 10019 6554
rect 10071 6545 10083 6554
rect 10135 6545 14266 6554
rect 14318 6545 14330 6554
rect 14382 6545 14394 6554
rect 10135 6511 10149 6545
rect 10183 6511 10241 6545
rect 10275 6511 10333 6545
rect 10367 6511 10425 6545
rect 10459 6511 10517 6545
rect 10551 6511 10609 6545
rect 10643 6511 10701 6545
rect 10735 6511 10793 6545
rect 10827 6511 10885 6545
rect 10919 6511 10977 6545
rect 11011 6511 11069 6545
rect 11103 6511 11161 6545
rect 11195 6511 11253 6545
rect 11287 6511 11345 6545
rect 11379 6511 11437 6545
rect 11471 6511 11529 6545
rect 11563 6511 11621 6545
rect 11655 6511 11713 6545
rect 11747 6511 11805 6545
rect 11839 6511 11897 6545
rect 11931 6511 11989 6545
rect 12023 6511 12081 6545
rect 12115 6511 12173 6545
rect 12207 6511 12265 6545
rect 12299 6511 12357 6545
rect 12391 6511 12449 6545
rect 12483 6511 12541 6545
rect 12575 6511 12633 6545
rect 12667 6511 12725 6545
rect 12759 6511 12817 6545
rect 12851 6511 12909 6545
rect 12943 6511 13001 6545
rect 13035 6511 13093 6545
rect 13127 6511 13185 6545
rect 13219 6511 13277 6545
rect 13311 6511 13369 6545
rect 13403 6511 13461 6545
rect 13495 6511 13553 6545
rect 13587 6511 13645 6545
rect 13679 6511 13737 6545
rect 13771 6511 13829 6545
rect 13863 6511 13921 6545
rect 13955 6511 14013 6545
rect 14047 6511 14105 6545
rect 14139 6511 14197 6545
rect 14231 6511 14266 6545
rect 14323 6511 14330 6545
rect 10071 6502 10083 6511
rect 10135 6502 14266 6511
rect 14318 6502 14330 6511
rect 14382 6502 14394 6511
rect 14446 6502 14458 6554
rect 14510 6502 14522 6554
rect 14574 6545 18705 6554
rect 14599 6511 14657 6545
rect 14691 6511 14749 6545
rect 14783 6511 14841 6545
rect 14875 6511 14933 6545
rect 14967 6511 15025 6545
rect 15059 6511 15117 6545
rect 15151 6511 15209 6545
rect 15243 6511 15301 6545
rect 15335 6511 15393 6545
rect 15427 6511 15485 6545
rect 15519 6511 15577 6545
rect 15611 6511 15669 6545
rect 15703 6511 15761 6545
rect 15795 6511 15853 6545
rect 15887 6511 15945 6545
rect 15979 6511 16037 6545
rect 16071 6511 16129 6545
rect 16163 6511 16221 6545
rect 16255 6511 16313 6545
rect 16347 6511 16405 6545
rect 16439 6511 16497 6545
rect 16531 6511 16589 6545
rect 16623 6511 16681 6545
rect 16715 6511 16773 6545
rect 16807 6511 16865 6545
rect 16899 6511 16957 6545
rect 16991 6511 17049 6545
rect 17083 6511 17141 6545
rect 17175 6511 17233 6545
rect 17267 6511 17325 6545
rect 17359 6511 17417 6545
rect 17451 6511 17509 6545
rect 17543 6511 17601 6545
rect 17635 6511 17693 6545
rect 17727 6511 17785 6545
rect 17819 6511 17877 6545
rect 17911 6511 17969 6545
rect 18003 6511 18061 6545
rect 18095 6511 18153 6545
rect 18187 6511 18245 6545
rect 18279 6511 18337 6545
rect 18371 6511 18429 6545
rect 18463 6511 18521 6545
rect 18555 6511 18613 6545
rect 18647 6511 18705 6545
rect 14574 6502 18705 6511
rect 18757 6502 18769 6554
rect 18821 6545 18833 6554
rect 18831 6511 18833 6545
rect 18821 6502 18833 6511
rect 18885 6502 18897 6554
rect 18949 6502 18961 6554
rect 19013 6502 19019 6554
rect 1104 6480 19019 6502
rect 1104 6010 18860 6032
rect 1104 6001 3169 6010
rect 1104 5967 1133 6001
rect 1167 5967 1225 6001
rect 1259 5967 1317 6001
rect 1351 5967 1409 6001
rect 1443 5967 1501 6001
rect 1535 5967 1593 6001
rect 1627 5967 1685 6001
rect 1719 5967 1777 6001
rect 1811 5967 1869 6001
rect 1903 5967 1961 6001
rect 1995 5967 2053 6001
rect 2087 5967 2145 6001
rect 2179 5967 2237 6001
rect 2271 5967 2329 6001
rect 2363 5967 2421 6001
rect 2455 5967 2513 6001
rect 2547 5967 2605 6001
rect 2639 5967 2697 6001
rect 2731 5967 2789 6001
rect 2823 5967 2881 6001
rect 2915 5967 2973 6001
rect 3007 5967 3065 6001
rect 3099 5967 3157 6001
rect 1104 5958 3169 5967
rect 3221 5958 3233 6010
rect 3285 5958 3297 6010
rect 3349 6001 3361 6010
rect 3349 5958 3361 5967
rect 3413 5958 3425 6010
rect 3477 6001 7608 6010
rect 3477 5967 3525 6001
rect 3559 5967 3617 6001
rect 3651 5967 3709 6001
rect 3743 5967 3801 6001
rect 3835 5967 3893 6001
rect 3927 5967 3985 6001
rect 4019 5967 4077 6001
rect 4111 5967 4169 6001
rect 4203 5967 4261 6001
rect 4295 5967 4353 6001
rect 4387 5967 4445 6001
rect 4479 5967 4537 6001
rect 4571 5967 4629 6001
rect 4663 5967 4721 6001
rect 4755 5967 4813 6001
rect 4847 5967 4905 6001
rect 4939 5967 4997 6001
rect 5031 5967 5089 6001
rect 5123 5967 5181 6001
rect 5215 5967 5273 6001
rect 5307 5967 5365 6001
rect 5399 5967 5457 6001
rect 5491 5967 5549 6001
rect 5583 5967 5641 6001
rect 5675 5967 5733 6001
rect 5767 5967 5825 6001
rect 5859 5967 5917 6001
rect 5951 5967 6009 6001
rect 6043 5967 6101 6001
rect 6135 5967 6193 6001
rect 6227 5967 6285 6001
rect 6319 5967 6377 6001
rect 6411 5967 6469 6001
rect 6503 5967 6561 6001
rect 6595 5967 6653 6001
rect 6687 5967 6745 6001
rect 6779 5967 6837 6001
rect 6871 5967 6929 6001
rect 6963 5967 7021 6001
rect 7055 5967 7113 6001
rect 7147 5967 7205 6001
rect 7239 5967 7297 6001
rect 7331 5967 7389 6001
rect 7423 5967 7481 6001
rect 7515 5967 7573 6001
rect 7607 5967 7608 6001
rect 3477 5958 7608 5967
rect 7660 6001 7672 6010
rect 7660 5967 7665 6001
rect 7660 5958 7672 5967
rect 7724 5958 7736 6010
rect 7788 6001 7800 6010
rect 7852 6001 7864 6010
rect 7916 6001 12047 6010
rect 12099 6001 12111 6010
rect 12163 6001 12175 6010
rect 7791 5967 7800 6001
rect 7916 5967 7941 6001
rect 7975 5967 8033 6001
rect 8067 5967 8125 6001
rect 8159 5967 8217 6001
rect 8251 5967 8309 6001
rect 8343 5967 8401 6001
rect 8435 5967 8493 6001
rect 8527 5967 8585 6001
rect 8619 5967 8677 6001
rect 8711 5967 8769 6001
rect 8803 5967 8861 6001
rect 8895 5967 8953 6001
rect 8987 5967 9045 6001
rect 9079 5967 9137 6001
rect 9171 5967 9229 6001
rect 9263 5967 9321 6001
rect 9355 5967 9413 6001
rect 9447 5967 9505 6001
rect 9539 5967 9597 6001
rect 9631 5967 9689 6001
rect 9723 5967 9781 6001
rect 9815 5967 9873 6001
rect 9907 5967 9965 6001
rect 9999 5967 10057 6001
rect 10091 5967 10149 6001
rect 10183 5967 10241 6001
rect 10275 5967 10333 6001
rect 10367 5967 10425 6001
rect 10459 5967 10517 6001
rect 10551 5967 10609 6001
rect 10643 5967 10701 6001
rect 10735 5967 10793 6001
rect 10827 5967 10885 6001
rect 10919 5967 10977 6001
rect 11011 5967 11069 6001
rect 11103 5967 11161 6001
rect 11195 5967 11253 6001
rect 11287 5967 11345 6001
rect 11379 5967 11437 6001
rect 11471 5967 11529 6001
rect 11563 5967 11621 6001
rect 11655 5967 11713 6001
rect 11747 5967 11805 6001
rect 11839 5967 11897 6001
rect 11931 5967 11989 6001
rect 12023 5967 12047 6001
rect 12163 5967 12173 6001
rect 7788 5958 7800 5967
rect 7852 5958 7864 5967
rect 7916 5958 12047 5967
rect 12099 5958 12111 5967
rect 12163 5958 12175 5967
rect 12227 5958 12239 6010
rect 12291 6001 12303 6010
rect 12299 5967 12303 6001
rect 12291 5958 12303 5967
rect 12355 6001 16486 6010
rect 12355 5967 12357 6001
rect 12391 5967 12449 6001
rect 12483 5967 12541 6001
rect 12575 5967 12633 6001
rect 12667 5967 12725 6001
rect 12759 5967 12817 6001
rect 12851 5967 12909 6001
rect 12943 5967 13001 6001
rect 13035 5967 13093 6001
rect 13127 5967 13185 6001
rect 13219 5967 13277 6001
rect 13311 5967 13369 6001
rect 13403 5967 13461 6001
rect 13495 5967 13553 6001
rect 13587 5967 13645 6001
rect 13679 5967 13737 6001
rect 13771 5967 13829 6001
rect 13863 5967 13921 6001
rect 13955 5967 14013 6001
rect 14047 5967 14105 6001
rect 14139 5967 14197 6001
rect 14231 5967 14289 6001
rect 14323 5967 14381 6001
rect 14415 5967 14473 6001
rect 14507 5967 14565 6001
rect 14599 5967 14657 6001
rect 14691 5967 14749 6001
rect 14783 5967 14841 6001
rect 14875 5967 14933 6001
rect 14967 5967 15025 6001
rect 15059 5967 15117 6001
rect 15151 5967 15209 6001
rect 15243 5967 15301 6001
rect 15335 5967 15393 6001
rect 15427 5967 15485 6001
rect 15519 5967 15577 6001
rect 15611 5967 15669 6001
rect 15703 5967 15761 6001
rect 15795 5967 15853 6001
rect 15887 5967 15945 6001
rect 15979 5967 16037 6001
rect 16071 5967 16129 6001
rect 16163 5967 16221 6001
rect 16255 5967 16313 6001
rect 16347 5967 16405 6001
rect 16439 5967 16486 6001
rect 12355 5958 16486 5967
rect 16538 5958 16550 6010
rect 16602 6001 16614 6010
rect 16602 5958 16614 5967
rect 16666 5958 16678 6010
rect 16730 5958 16742 6010
rect 16794 6001 18860 6010
rect 16807 5967 16865 6001
rect 16899 5967 16957 6001
rect 16991 5967 17049 6001
rect 17083 5967 17141 6001
rect 17175 5967 17233 6001
rect 17267 5967 17325 6001
rect 17359 5967 17417 6001
rect 17451 5967 17509 6001
rect 17543 5967 17601 6001
rect 17635 5967 17693 6001
rect 17727 5967 17785 6001
rect 17819 5967 17877 6001
rect 17911 5967 17969 6001
rect 18003 5967 18061 6001
rect 18095 5967 18153 6001
rect 18187 5967 18245 6001
rect 18279 5967 18337 6001
rect 18371 5967 18429 6001
rect 18463 5967 18521 6001
rect 18555 5967 18613 6001
rect 18647 5967 18705 6001
rect 18739 5967 18797 6001
rect 18831 5967 18860 6001
rect 16794 5958 18860 5967
rect 1104 5936 18860 5958
rect 2409 5831 2467 5837
rect 2409 5797 2421 5831
rect 2455 5828 2467 5831
rect 7006 5828 7012 5840
rect 2455 5800 7012 5828
rect 2455 5797 2467 5800
rect 2409 5791 2467 5797
rect 7006 5788 7012 5800
rect 7064 5788 7070 5840
rect 10870 5788 10876 5840
rect 10928 5828 10934 5840
rect 12253 5831 12311 5837
rect 12253 5828 12265 5831
rect 10928 5800 12265 5828
rect 10928 5788 10934 5800
rect 12253 5797 12265 5800
rect 12299 5797 12311 5831
rect 12253 5791 12311 5797
rect 5902 5720 5908 5772
rect 5960 5760 5966 5772
rect 6822 5760 6828 5772
rect 5960 5732 6828 5760
rect 5960 5720 5966 5732
rect 6822 5720 6828 5732
rect 6880 5760 6886 5772
rect 7285 5763 7343 5769
rect 7285 5760 7297 5763
rect 6880 5732 7297 5760
rect 6880 5720 6886 5732
rect 7285 5729 7297 5732
rect 7331 5729 7343 5763
rect 10413 5763 10471 5769
rect 10413 5760 10425 5763
rect 7285 5723 7343 5729
rect 9646 5732 10425 5760
rect 2225 5695 2283 5701
rect 2225 5661 2237 5695
rect 2271 5692 2283 5695
rect 2866 5692 2872 5704
rect 2271 5664 2872 5692
rect 2271 5661 2283 5664
rect 2225 5655 2283 5661
rect 2866 5652 2872 5664
rect 2924 5652 2930 5704
rect 3237 5695 3295 5701
rect 3237 5661 3249 5695
rect 3283 5692 3295 5695
rect 3970 5692 3976 5704
rect 3283 5664 3976 5692
rect 3283 5661 3295 5664
rect 3237 5655 3295 5661
rect 3970 5652 3976 5664
rect 4028 5652 4034 5704
rect 5718 5652 5724 5704
rect 5776 5692 5782 5704
rect 9646 5692 9674 5732
rect 10413 5729 10425 5732
rect 10459 5729 10471 5763
rect 10413 5723 10471 5729
rect 10502 5720 10508 5772
rect 10560 5760 10566 5772
rect 11425 5763 11483 5769
rect 11425 5760 11437 5763
rect 10560 5732 11437 5760
rect 10560 5720 10566 5732
rect 11425 5729 11437 5732
rect 11471 5760 11483 5763
rect 12805 5763 12863 5769
rect 12805 5760 12817 5763
rect 11471 5732 12817 5760
rect 11471 5729 11483 5732
rect 11425 5723 11483 5729
rect 12805 5729 12817 5732
rect 12851 5729 12863 5763
rect 14826 5760 14832 5772
rect 14787 5732 14832 5760
rect 12805 5723 12863 5729
rect 14826 5720 14832 5732
rect 14884 5720 14890 5772
rect 10226 5692 10232 5704
rect 5776 5664 9674 5692
rect 10139 5664 10232 5692
rect 5776 5652 5782 5664
rect 10226 5652 10232 5664
rect 10284 5692 10290 5704
rect 10594 5692 10600 5704
rect 10284 5664 10600 5692
rect 10284 5652 10290 5664
rect 10594 5652 10600 5664
rect 10652 5652 10658 5704
rect 11238 5692 11244 5704
rect 11199 5664 11244 5692
rect 11238 5652 11244 5664
rect 11296 5652 11302 5704
rect 7190 5624 7196 5636
rect 7103 5596 7196 5624
rect 7190 5584 7196 5596
rect 7248 5624 7254 5636
rect 8294 5624 8300 5636
rect 7248 5596 8300 5624
rect 7248 5584 7254 5596
rect 8294 5584 8300 5596
rect 8352 5624 8358 5636
rect 10318 5624 10324 5636
rect 8352 5596 10324 5624
rect 8352 5584 8358 5596
rect 10318 5584 10324 5596
rect 10376 5624 10382 5636
rect 10962 5624 10968 5636
rect 10376 5596 10968 5624
rect 10376 5584 10382 5596
rect 10962 5584 10968 5596
rect 11020 5624 11026 5636
rect 12713 5627 12771 5633
rect 12713 5624 12725 5627
rect 11020 5596 12725 5624
rect 11020 5584 11026 5596
rect 12713 5593 12725 5596
rect 12759 5624 12771 5627
rect 13538 5624 13544 5636
rect 12759 5596 13544 5624
rect 12759 5593 12771 5596
rect 12713 5587 12771 5593
rect 13538 5584 13544 5596
rect 13596 5624 13602 5636
rect 14737 5627 14795 5633
rect 14737 5624 14749 5627
rect 13596 5596 14749 5624
rect 13596 5584 13602 5596
rect 14737 5593 14749 5596
rect 14783 5593 14795 5627
rect 14737 5587 14795 5593
rect 3050 5556 3056 5568
rect 3011 5528 3056 5556
rect 3050 5516 3056 5528
rect 3108 5516 3114 5568
rect 5994 5516 6000 5568
rect 6052 5556 6058 5568
rect 6733 5559 6791 5565
rect 6733 5556 6745 5559
rect 6052 5528 6745 5556
rect 6052 5516 6058 5528
rect 6733 5525 6745 5528
rect 6779 5525 6791 5559
rect 7098 5556 7104 5568
rect 7059 5528 7104 5556
rect 6733 5519 6791 5525
rect 7098 5516 7104 5528
rect 7156 5516 7162 5568
rect 9674 5516 9680 5568
rect 9732 5556 9738 5568
rect 9861 5559 9919 5565
rect 9861 5556 9873 5559
rect 9732 5528 9873 5556
rect 9732 5516 9738 5528
rect 9861 5525 9873 5528
rect 9907 5525 9919 5559
rect 11054 5556 11060 5568
rect 11015 5528 11060 5556
rect 9861 5519 9919 5525
rect 11054 5516 11060 5528
rect 11112 5516 11118 5568
rect 12526 5516 12532 5568
rect 12584 5556 12590 5568
rect 12621 5559 12679 5565
rect 12621 5556 12633 5559
rect 12584 5528 12633 5556
rect 12584 5516 12590 5528
rect 12621 5525 12633 5528
rect 12667 5525 12679 5559
rect 12621 5519 12679 5525
rect 13814 5516 13820 5568
rect 13872 5556 13878 5568
rect 14277 5559 14335 5565
rect 14277 5556 14289 5559
rect 13872 5528 14289 5556
rect 13872 5516 13878 5528
rect 14277 5525 14289 5528
rect 14323 5525 14335 5559
rect 14642 5556 14648 5568
rect 14603 5528 14648 5556
rect 14277 5519 14335 5525
rect 14642 5516 14648 5528
rect 14700 5516 14706 5568
rect 1104 5466 19019 5488
rect 1104 5457 5388 5466
rect 1104 5423 1133 5457
rect 1167 5423 1225 5457
rect 1259 5423 1317 5457
rect 1351 5423 1409 5457
rect 1443 5423 1501 5457
rect 1535 5423 1593 5457
rect 1627 5423 1685 5457
rect 1719 5423 1777 5457
rect 1811 5423 1869 5457
rect 1903 5423 1961 5457
rect 1995 5423 2053 5457
rect 2087 5423 2145 5457
rect 2179 5423 2237 5457
rect 2271 5423 2329 5457
rect 2363 5423 2421 5457
rect 2455 5423 2513 5457
rect 2547 5423 2605 5457
rect 2639 5423 2697 5457
rect 2731 5423 2789 5457
rect 2823 5423 2881 5457
rect 2915 5423 2973 5457
rect 3007 5423 3065 5457
rect 3099 5423 3157 5457
rect 3191 5423 3249 5457
rect 3283 5423 3341 5457
rect 3375 5423 3433 5457
rect 3467 5423 3525 5457
rect 3559 5423 3617 5457
rect 3651 5423 3709 5457
rect 3743 5423 3801 5457
rect 3835 5423 3893 5457
rect 3927 5423 3985 5457
rect 4019 5423 4077 5457
rect 4111 5423 4169 5457
rect 4203 5423 4261 5457
rect 4295 5423 4353 5457
rect 4387 5423 4445 5457
rect 4479 5423 4537 5457
rect 4571 5423 4629 5457
rect 4663 5423 4721 5457
rect 4755 5423 4813 5457
rect 4847 5423 4905 5457
rect 4939 5423 4997 5457
rect 5031 5423 5089 5457
rect 5123 5423 5181 5457
rect 5215 5423 5273 5457
rect 5307 5423 5365 5457
rect 1104 5414 5388 5423
rect 5440 5414 5452 5466
rect 5504 5414 5516 5466
rect 5568 5457 5580 5466
rect 5632 5457 5644 5466
rect 5696 5457 9827 5466
rect 9879 5457 9891 5466
rect 5632 5423 5641 5457
rect 5696 5423 5733 5457
rect 5767 5423 5825 5457
rect 5859 5423 5917 5457
rect 5951 5423 6009 5457
rect 6043 5423 6101 5457
rect 6135 5423 6193 5457
rect 6227 5423 6285 5457
rect 6319 5423 6377 5457
rect 6411 5423 6469 5457
rect 6503 5423 6561 5457
rect 6595 5423 6653 5457
rect 6687 5423 6745 5457
rect 6779 5423 6837 5457
rect 6871 5423 6929 5457
rect 6963 5423 7021 5457
rect 7055 5423 7113 5457
rect 7147 5423 7205 5457
rect 7239 5423 7297 5457
rect 7331 5423 7389 5457
rect 7423 5423 7481 5457
rect 7515 5423 7573 5457
rect 7607 5423 7665 5457
rect 7699 5423 7757 5457
rect 7791 5423 7849 5457
rect 7883 5423 7941 5457
rect 7975 5423 8033 5457
rect 8067 5423 8125 5457
rect 8159 5423 8217 5457
rect 8251 5423 8309 5457
rect 8343 5423 8401 5457
rect 8435 5423 8493 5457
rect 8527 5423 8585 5457
rect 8619 5423 8677 5457
rect 8711 5423 8769 5457
rect 8803 5423 8861 5457
rect 8895 5423 8953 5457
rect 8987 5423 9045 5457
rect 9079 5423 9137 5457
rect 9171 5423 9229 5457
rect 9263 5423 9321 5457
rect 9355 5423 9413 5457
rect 9447 5423 9505 5457
rect 9539 5423 9597 5457
rect 9631 5423 9689 5457
rect 9723 5423 9781 5457
rect 9815 5423 9827 5457
rect 5568 5414 5580 5423
rect 5632 5414 5644 5423
rect 5696 5414 9827 5423
rect 9879 5414 9891 5423
rect 9943 5414 9955 5466
rect 10007 5414 10019 5466
rect 10071 5457 10083 5466
rect 10135 5457 14266 5466
rect 14318 5457 14330 5466
rect 14382 5457 14394 5466
rect 10135 5423 10149 5457
rect 10183 5423 10241 5457
rect 10275 5423 10333 5457
rect 10367 5423 10425 5457
rect 10459 5423 10517 5457
rect 10551 5423 10609 5457
rect 10643 5423 10701 5457
rect 10735 5423 10793 5457
rect 10827 5423 10885 5457
rect 10919 5423 10977 5457
rect 11011 5423 11069 5457
rect 11103 5423 11161 5457
rect 11195 5423 11253 5457
rect 11287 5423 11345 5457
rect 11379 5423 11437 5457
rect 11471 5423 11529 5457
rect 11563 5423 11621 5457
rect 11655 5423 11713 5457
rect 11747 5423 11805 5457
rect 11839 5423 11897 5457
rect 11931 5423 11989 5457
rect 12023 5423 12081 5457
rect 12115 5423 12173 5457
rect 12207 5423 12265 5457
rect 12299 5423 12357 5457
rect 12391 5423 12449 5457
rect 12483 5423 12541 5457
rect 12575 5423 12633 5457
rect 12667 5423 12725 5457
rect 12759 5423 12817 5457
rect 12851 5423 12909 5457
rect 12943 5423 13001 5457
rect 13035 5423 13093 5457
rect 13127 5423 13185 5457
rect 13219 5423 13277 5457
rect 13311 5423 13369 5457
rect 13403 5423 13461 5457
rect 13495 5423 13553 5457
rect 13587 5423 13645 5457
rect 13679 5423 13737 5457
rect 13771 5423 13829 5457
rect 13863 5423 13921 5457
rect 13955 5423 14013 5457
rect 14047 5423 14105 5457
rect 14139 5423 14197 5457
rect 14231 5423 14266 5457
rect 14323 5423 14330 5457
rect 10071 5414 10083 5423
rect 10135 5414 14266 5423
rect 14318 5414 14330 5423
rect 14382 5414 14394 5423
rect 14446 5414 14458 5466
rect 14510 5414 14522 5466
rect 14574 5457 18705 5466
rect 14599 5423 14657 5457
rect 14691 5423 14749 5457
rect 14783 5423 14841 5457
rect 14875 5423 14933 5457
rect 14967 5423 15025 5457
rect 15059 5423 15117 5457
rect 15151 5423 15209 5457
rect 15243 5423 15301 5457
rect 15335 5423 15393 5457
rect 15427 5423 15485 5457
rect 15519 5423 15577 5457
rect 15611 5423 15669 5457
rect 15703 5423 15761 5457
rect 15795 5423 15853 5457
rect 15887 5423 15945 5457
rect 15979 5423 16037 5457
rect 16071 5423 16129 5457
rect 16163 5423 16221 5457
rect 16255 5423 16313 5457
rect 16347 5423 16405 5457
rect 16439 5423 16497 5457
rect 16531 5423 16589 5457
rect 16623 5423 16681 5457
rect 16715 5423 16773 5457
rect 16807 5423 16865 5457
rect 16899 5423 16957 5457
rect 16991 5423 17049 5457
rect 17083 5423 17141 5457
rect 17175 5423 17233 5457
rect 17267 5423 17325 5457
rect 17359 5423 17417 5457
rect 17451 5423 17509 5457
rect 17543 5423 17601 5457
rect 17635 5423 17693 5457
rect 17727 5423 17785 5457
rect 17819 5423 17877 5457
rect 17911 5423 17969 5457
rect 18003 5423 18061 5457
rect 18095 5423 18153 5457
rect 18187 5423 18245 5457
rect 18279 5423 18337 5457
rect 18371 5423 18429 5457
rect 18463 5423 18521 5457
rect 18555 5423 18613 5457
rect 18647 5423 18705 5457
rect 14574 5414 18705 5423
rect 18757 5414 18769 5466
rect 18821 5457 18833 5466
rect 18831 5423 18833 5457
rect 18821 5414 18833 5423
rect 18885 5414 18897 5466
rect 18949 5414 18961 5466
rect 19013 5414 19019 5466
rect 1104 5392 19019 5414
rect 2866 5352 2872 5364
rect 2827 5324 2872 5352
rect 2866 5312 2872 5324
rect 2924 5312 2930 5364
rect 3878 5352 3884 5364
rect 3839 5324 3884 5352
rect 3878 5312 3884 5324
rect 3936 5312 3942 5364
rect 7009 5355 7067 5361
rect 7009 5352 7021 5355
rect 6932 5324 7021 5352
rect 6932 5296 6960 5324
rect 7009 5321 7021 5324
rect 7055 5321 7067 5355
rect 7009 5315 7067 5321
rect 7101 5355 7159 5361
rect 7101 5321 7113 5355
rect 7147 5352 7159 5355
rect 7190 5352 7196 5364
rect 7147 5324 7196 5352
rect 7147 5321 7159 5324
rect 7101 5315 7159 5321
rect 7190 5312 7196 5324
rect 7248 5312 7254 5364
rect 8294 5352 8300 5364
rect 8255 5324 8300 5352
rect 8294 5312 8300 5324
rect 8352 5312 8358 5364
rect 10873 5355 10931 5361
rect 10873 5321 10885 5355
rect 10919 5352 10931 5355
rect 10962 5352 10968 5364
rect 10919 5324 10968 5352
rect 10919 5321 10931 5324
rect 10873 5315 10931 5321
rect 10962 5312 10968 5324
rect 11020 5312 11026 5364
rect 13446 5352 13452 5364
rect 13407 5324 13452 5352
rect 13446 5312 13452 5324
rect 13504 5312 13510 5364
rect 13538 5312 13544 5364
rect 13596 5352 13602 5364
rect 13596 5324 13641 5352
rect 13596 5312 13602 5324
rect 5902 5284 5908 5296
rect 3252 5256 5908 5284
rect 2130 5216 2136 5228
rect 2043 5188 2136 5216
rect 2130 5176 2136 5188
rect 2188 5216 2194 5228
rect 3252 5225 3280 5256
rect 5902 5244 5908 5256
rect 5960 5244 5966 5296
rect 6914 5244 6920 5296
rect 6972 5244 6978 5296
rect 11054 5284 11060 5296
rect 7024 5256 11060 5284
rect 3053 5219 3111 5225
rect 3053 5216 3065 5219
rect 2188 5188 3065 5216
rect 2188 5176 2194 5188
rect 3053 5185 3065 5188
rect 3099 5185 3111 5219
rect 3053 5179 3111 5185
rect 3237 5219 3295 5225
rect 3237 5185 3249 5219
rect 3283 5185 3295 5219
rect 3694 5216 3700 5228
rect 3655 5188 3700 5216
rect 3237 5179 3295 5185
rect 2317 5151 2375 5157
rect 2317 5117 2329 5151
rect 2363 5117 2375 5151
rect 3068 5148 3096 5179
rect 3694 5176 3700 5188
rect 3752 5176 3758 5228
rect 3878 5176 3884 5228
rect 3936 5216 3942 5228
rect 4433 5219 4491 5225
rect 4433 5216 4445 5219
rect 3936 5188 4445 5216
rect 3936 5176 3942 5188
rect 4433 5185 4445 5188
rect 4479 5216 4491 5219
rect 5074 5216 5080 5228
rect 4479 5188 5080 5216
rect 4479 5185 4491 5188
rect 4433 5179 4491 5185
rect 5074 5176 5080 5188
rect 5132 5176 5138 5228
rect 5997 5219 6055 5225
rect 5997 5185 6009 5219
rect 6043 5216 6055 5219
rect 6043 5206 6914 5216
rect 7024 5206 7052 5256
rect 11054 5244 11060 5256
rect 11112 5244 11118 5296
rect 8205 5219 8263 5225
rect 8205 5216 8217 5219
rect 6043 5188 7052 5206
rect 6043 5185 6055 5188
rect 5997 5179 6055 5185
rect 6886 5178 7052 5188
rect 7208 5188 8217 5216
rect 3712 5148 3740 5176
rect 3068 5120 3740 5148
rect 2317 5111 2375 5117
rect 2332 5080 2360 5111
rect 4614 5108 4620 5160
rect 4672 5148 4678 5160
rect 4672 5120 7052 5148
rect 4672 5108 4678 5120
rect 2590 5080 2596 5092
rect 2332 5052 2596 5080
rect 2590 5040 2596 5052
rect 2648 5080 2654 5092
rect 5718 5080 5724 5092
rect 2648 5052 5724 5080
rect 2648 5040 2654 5052
rect 5718 5040 5724 5052
rect 5776 5040 5782 5092
rect 7024 5080 7052 5120
rect 7208 5080 7236 5188
rect 8205 5185 8217 5188
rect 8251 5185 8263 5219
rect 9306 5216 9312 5228
rect 9267 5188 9312 5216
rect 8205 5179 8263 5185
rect 9306 5176 9312 5188
rect 9364 5176 9370 5228
rect 9493 5219 9551 5225
rect 9493 5185 9505 5219
rect 9539 5216 9551 5219
rect 9674 5216 9680 5228
rect 9539 5188 9680 5216
rect 9539 5185 9551 5188
rect 9493 5179 9551 5185
rect 9674 5176 9680 5188
rect 9732 5176 9738 5228
rect 9766 5176 9772 5228
rect 9824 5216 9830 5228
rect 10781 5219 10839 5225
rect 10781 5216 10793 5219
rect 9824 5188 10793 5216
rect 9824 5176 9830 5188
rect 10781 5185 10793 5188
rect 10827 5185 10839 5219
rect 10781 5179 10839 5185
rect 7282 5108 7288 5160
rect 7340 5148 7346 5160
rect 8386 5148 8392 5160
rect 7340 5120 7385 5148
rect 8347 5120 8392 5148
rect 7340 5108 7346 5120
rect 8386 5108 8392 5120
rect 8444 5108 8450 5160
rect 9585 5151 9643 5157
rect 9585 5117 9597 5151
rect 9631 5148 9643 5151
rect 9950 5148 9956 5160
rect 9631 5120 9956 5148
rect 9631 5117 9643 5120
rect 9585 5111 9643 5117
rect 9950 5108 9956 5120
rect 10008 5148 10014 5160
rect 10502 5148 10508 5160
rect 10008 5120 10508 5148
rect 10008 5108 10014 5120
rect 10502 5108 10508 5120
rect 10560 5108 10566 5160
rect 10965 5151 11023 5157
rect 10965 5117 10977 5151
rect 11011 5148 11023 5151
rect 11882 5148 11888 5160
rect 11011 5120 11888 5148
rect 11011 5117 11023 5120
rect 10965 5111 11023 5117
rect 11882 5108 11888 5120
rect 11940 5108 11946 5160
rect 12986 5108 12992 5160
rect 13044 5148 13050 5160
rect 13633 5151 13691 5157
rect 13633 5148 13645 5151
rect 13044 5120 13645 5148
rect 13044 5108 13050 5120
rect 13633 5117 13645 5120
rect 13679 5117 13691 5151
rect 13633 5111 13691 5117
rect 7024 5052 7236 5080
rect 11238 5040 11244 5092
rect 11296 5080 11302 5092
rect 14550 5080 14556 5092
rect 11296 5052 14556 5080
rect 11296 5040 11302 5052
rect 14550 5040 14556 5052
rect 14608 5040 14614 5092
rect 1946 5012 1952 5024
rect 1907 4984 1952 5012
rect 1946 4972 1952 4984
rect 2004 4972 2010 5024
rect 4525 5015 4583 5021
rect 4525 4981 4537 5015
rect 4571 5012 4583 5015
rect 4706 5012 4712 5024
rect 4571 4984 4712 5012
rect 4571 4981 4583 4984
rect 4525 4975 4583 4981
rect 4706 4972 4712 4984
rect 4764 4972 4770 5024
rect 4798 4972 4804 5024
rect 4856 5012 4862 5024
rect 5813 5015 5871 5021
rect 5813 5012 5825 5015
rect 4856 4984 5825 5012
rect 4856 4972 4862 4984
rect 5813 4981 5825 4984
rect 5859 4981 5871 5015
rect 6638 5012 6644 5024
rect 6599 4984 6644 5012
rect 5813 4975 5871 4981
rect 6638 4972 6644 4984
rect 6696 4972 6702 5024
rect 6730 4972 6736 5024
rect 6788 5012 6794 5024
rect 7837 5015 7895 5021
rect 7837 5012 7849 5015
rect 6788 4984 7849 5012
rect 6788 4972 6794 4984
rect 7837 4981 7849 4984
rect 7883 4981 7895 5015
rect 9122 5012 9128 5024
rect 9083 4984 9128 5012
rect 7837 4975 7895 4981
rect 9122 4972 9128 4984
rect 9180 4972 9186 5024
rect 9214 4972 9220 5024
rect 9272 5012 9278 5024
rect 10413 5015 10471 5021
rect 10413 5012 10425 5015
rect 9272 4984 10425 5012
rect 9272 4972 9278 4984
rect 10413 4981 10425 4984
rect 10459 4981 10471 5015
rect 13078 5012 13084 5024
rect 13039 4984 13084 5012
rect 10413 4975 10471 4981
rect 13078 4972 13084 4984
rect 13136 4972 13142 5024
rect 1104 4922 18860 4944
rect 1104 4913 3169 4922
rect 1104 4879 1133 4913
rect 1167 4879 1225 4913
rect 1259 4879 1317 4913
rect 1351 4879 1409 4913
rect 1443 4879 1501 4913
rect 1535 4879 1593 4913
rect 1627 4879 1685 4913
rect 1719 4879 1777 4913
rect 1811 4879 1869 4913
rect 1903 4879 1961 4913
rect 1995 4879 2053 4913
rect 2087 4879 2145 4913
rect 2179 4879 2237 4913
rect 2271 4879 2329 4913
rect 2363 4879 2421 4913
rect 2455 4879 2513 4913
rect 2547 4879 2605 4913
rect 2639 4879 2697 4913
rect 2731 4879 2789 4913
rect 2823 4879 2881 4913
rect 2915 4879 2973 4913
rect 3007 4879 3065 4913
rect 3099 4879 3157 4913
rect 1104 4870 3169 4879
rect 3221 4870 3233 4922
rect 3285 4870 3297 4922
rect 3349 4913 3361 4922
rect 3349 4870 3361 4879
rect 3413 4870 3425 4922
rect 3477 4913 7608 4922
rect 3477 4879 3525 4913
rect 3559 4879 3617 4913
rect 3651 4879 3709 4913
rect 3743 4879 3801 4913
rect 3835 4879 3893 4913
rect 3927 4879 3985 4913
rect 4019 4879 4077 4913
rect 4111 4879 4169 4913
rect 4203 4879 4261 4913
rect 4295 4879 4353 4913
rect 4387 4879 4445 4913
rect 4479 4879 4537 4913
rect 4571 4879 4629 4913
rect 4663 4879 4721 4913
rect 4755 4879 4813 4913
rect 4847 4879 4905 4913
rect 4939 4879 4997 4913
rect 5031 4879 5089 4913
rect 5123 4879 5181 4913
rect 5215 4879 5273 4913
rect 5307 4879 5365 4913
rect 5399 4879 5457 4913
rect 5491 4879 5549 4913
rect 5583 4879 5641 4913
rect 5675 4879 5733 4913
rect 5767 4879 5825 4913
rect 5859 4879 5917 4913
rect 5951 4879 6009 4913
rect 6043 4879 6101 4913
rect 6135 4879 6193 4913
rect 6227 4879 6285 4913
rect 6319 4879 6377 4913
rect 6411 4879 6469 4913
rect 6503 4879 6561 4913
rect 6595 4879 6653 4913
rect 6687 4879 6745 4913
rect 6779 4879 6837 4913
rect 6871 4879 6929 4913
rect 6963 4879 7021 4913
rect 7055 4879 7113 4913
rect 7147 4879 7205 4913
rect 7239 4879 7297 4913
rect 7331 4879 7389 4913
rect 7423 4879 7481 4913
rect 7515 4879 7573 4913
rect 7607 4879 7608 4913
rect 3477 4870 7608 4879
rect 7660 4913 7672 4922
rect 7660 4879 7665 4913
rect 7660 4870 7672 4879
rect 7724 4870 7736 4922
rect 7788 4913 7800 4922
rect 7852 4913 7864 4922
rect 7916 4913 12047 4922
rect 12099 4913 12111 4922
rect 12163 4913 12175 4922
rect 7791 4879 7800 4913
rect 7916 4879 7941 4913
rect 7975 4879 8033 4913
rect 8067 4879 8125 4913
rect 8159 4879 8217 4913
rect 8251 4879 8309 4913
rect 8343 4879 8401 4913
rect 8435 4879 8493 4913
rect 8527 4879 8585 4913
rect 8619 4879 8677 4913
rect 8711 4879 8769 4913
rect 8803 4879 8861 4913
rect 8895 4879 8953 4913
rect 8987 4879 9045 4913
rect 9079 4879 9137 4913
rect 9171 4879 9229 4913
rect 9263 4879 9321 4913
rect 9355 4879 9413 4913
rect 9447 4879 9505 4913
rect 9539 4879 9597 4913
rect 9631 4879 9689 4913
rect 9723 4879 9781 4913
rect 9815 4879 9873 4913
rect 9907 4879 9965 4913
rect 9999 4879 10057 4913
rect 10091 4879 10149 4913
rect 10183 4879 10241 4913
rect 10275 4879 10333 4913
rect 10367 4879 10425 4913
rect 10459 4879 10517 4913
rect 10551 4879 10609 4913
rect 10643 4879 10701 4913
rect 10735 4879 10793 4913
rect 10827 4879 10885 4913
rect 10919 4879 10977 4913
rect 11011 4879 11069 4913
rect 11103 4879 11161 4913
rect 11195 4879 11253 4913
rect 11287 4879 11345 4913
rect 11379 4879 11437 4913
rect 11471 4879 11529 4913
rect 11563 4879 11621 4913
rect 11655 4879 11713 4913
rect 11747 4879 11805 4913
rect 11839 4879 11897 4913
rect 11931 4879 11989 4913
rect 12023 4879 12047 4913
rect 12163 4879 12173 4913
rect 7788 4870 7800 4879
rect 7852 4870 7864 4879
rect 7916 4870 12047 4879
rect 12099 4870 12111 4879
rect 12163 4870 12175 4879
rect 12227 4870 12239 4922
rect 12291 4913 12303 4922
rect 12299 4879 12303 4913
rect 12291 4870 12303 4879
rect 12355 4913 16486 4922
rect 12355 4879 12357 4913
rect 12391 4879 12449 4913
rect 12483 4879 12541 4913
rect 12575 4879 12633 4913
rect 12667 4879 12725 4913
rect 12759 4879 12817 4913
rect 12851 4879 12909 4913
rect 12943 4879 13001 4913
rect 13035 4879 13093 4913
rect 13127 4879 13185 4913
rect 13219 4879 13277 4913
rect 13311 4879 13369 4913
rect 13403 4879 13461 4913
rect 13495 4879 13553 4913
rect 13587 4879 13645 4913
rect 13679 4879 13737 4913
rect 13771 4879 13829 4913
rect 13863 4879 13921 4913
rect 13955 4879 14013 4913
rect 14047 4879 14105 4913
rect 14139 4879 14197 4913
rect 14231 4879 14289 4913
rect 14323 4879 14381 4913
rect 14415 4879 14473 4913
rect 14507 4879 14565 4913
rect 14599 4879 14657 4913
rect 14691 4879 14749 4913
rect 14783 4879 14841 4913
rect 14875 4879 14933 4913
rect 14967 4879 15025 4913
rect 15059 4879 15117 4913
rect 15151 4879 15209 4913
rect 15243 4879 15301 4913
rect 15335 4879 15393 4913
rect 15427 4879 15485 4913
rect 15519 4879 15577 4913
rect 15611 4879 15669 4913
rect 15703 4879 15761 4913
rect 15795 4879 15853 4913
rect 15887 4879 15945 4913
rect 15979 4879 16037 4913
rect 16071 4879 16129 4913
rect 16163 4879 16221 4913
rect 16255 4879 16313 4913
rect 16347 4879 16405 4913
rect 16439 4879 16486 4913
rect 12355 4870 16486 4879
rect 16538 4870 16550 4922
rect 16602 4913 16614 4922
rect 16602 4870 16614 4879
rect 16666 4870 16678 4922
rect 16730 4870 16742 4922
rect 16794 4913 18860 4922
rect 16807 4879 16865 4913
rect 16899 4879 16957 4913
rect 16991 4879 17049 4913
rect 17083 4879 17141 4913
rect 17175 4879 17233 4913
rect 17267 4879 17325 4913
rect 17359 4879 17417 4913
rect 17451 4879 17509 4913
rect 17543 4879 17601 4913
rect 17635 4879 17693 4913
rect 17727 4879 17785 4913
rect 17819 4879 17877 4913
rect 17911 4879 17969 4913
rect 18003 4879 18061 4913
rect 18095 4879 18153 4913
rect 18187 4879 18245 4913
rect 18279 4879 18337 4913
rect 18371 4879 18429 4913
rect 18463 4879 18521 4913
rect 18555 4879 18613 4913
rect 18647 4879 18705 4913
rect 18739 4879 18797 4913
rect 18831 4879 18860 4913
rect 16794 4870 18860 4879
rect 1104 4848 18860 4870
rect 3970 4808 3976 4820
rect 3931 4780 3976 4808
rect 3970 4768 3976 4780
rect 4028 4768 4034 4820
rect 5261 4811 5319 4817
rect 5261 4777 5273 4811
rect 5307 4808 5319 4811
rect 5994 4808 6000 4820
rect 5307 4780 6000 4808
rect 5307 4777 5319 4780
rect 5261 4771 5319 4777
rect 5994 4768 6000 4780
rect 6052 4768 6058 4820
rect 6181 4811 6239 4817
rect 6181 4777 6193 4811
rect 6227 4808 6239 4811
rect 6546 4808 6552 4820
rect 6227 4780 6552 4808
rect 6227 4777 6239 4780
rect 6181 4771 6239 4777
rect 6546 4768 6552 4780
rect 6604 4768 6610 4820
rect 9950 4808 9956 4820
rect 6748 4780 7696 4808
rect 9911 4780 9956 4808
rect 2138 4743 2196 4749
rect 2138 4709 2150 4743
rect 2184 4740 2196 4743
rect 2558 4743 2616 4749
rect 2558 4740 2570 4743
rect 2184 4712 2570 4740
rect 2184 4709 2196 4712
rect 2138 4703 2196 4709
rect 2558 4709 2570 4712
rect 2604 4740 2616 4743
rect 2872 4743 2930 4749
rect 2872 4740 2884 4743
rect 2604 4712 2884 4740
rect 2604 4709 2616 4712
rect 2558 4703 2616 4709
rect 2872 4709 2884 4712
rect 2918 4709 2930 4743
rect 2872 4703 2930 4709
rect 3694 4700 3700 4752
rect 3752 4740 3758 4752
rect 6748 4740 6776 4780
rect 3752 4712 6776 4740
rect 6830 4743 6888 4749
rect 3752 4700 3758 4712
rect 2217 4675 2275 4681
rect 2217 4641 2229 4675
rect 2263 4672 2275 4675
rect 2455 4675 2513 4681
rect 2455 4672 2467 4675
rect 2263 4644 2467 4672
rect 2263 4641 2275 4644
rect 2217 4635 2275 4641
rect 2455 4641 2467 4644
rect 2501 4672 2513 4675
rect 2959 4675 3017 4681
rect 2959 4672 2971 4675
rect 2501 4644 2971 4672
rect 2501 4641 2513 4644
rect 2455 4635 2513 4641
rect 2959 4641 2971 4644
rect 3005 4641 3017 4675
rect 2959 4635 3017 4641
rect 2038 4604 2044 4616
rect 1999 4576 2044 4604
rect 2038 4564 2044 4576
rect 2096 4564 2102 4616
rect 2308 4607 2366 4613
rect 2308 4573 2320 4607
rect 2354 4604 2366 4607
rect 3050 4604 3056 4616
rect 2354 4576 3056 4604
rect 2354 4573 2366 4576
rect 2308 4567 2366 4573
rect 3050 4564 3056 4576
rect 3108 4564 3114 4616
rect 4172 4613 4200 4712
rect 6830 4709 6842 4743
rect 6876 4740 6888 4743
rect 7250 4743 7308 4749
rect 7250 4740 7262 4743
rect 6876 4712 7262 4740
rect 6876 4709 6888 4712
rect 6830 4703 6888 4709
rect 7250 4709 7262 4712
rect 7296 4740 7308 4743
rect 7564 4743 7622 4749
rect 7564 4740 7576 4743
rect 7296 4712 7576 4740
rect 7296 4709 7308 4712
rect 7250 4703 7308 4709
rect 7564 4709 7576 4712
rect 7610 4709 7622 4743
rect 7668 4740 7696 4780
rect 9950 4768 9956 4780
rect 10008 4768 10014 4820
rect 11146 4808 11152 4820
rect 10051 4780 11152 4808
rect 10051 4740 10079 4780
rect 11146 4768 11152 4780
rect 11204 4768 11210 4820
rect 12161 4811 12219 4817
rect 12161 4777 12173 4811
rect 12207 4808 12219 4811
rect 13078 4808 13084 4820
rect 12207 4780 13084 4808
rect 12207 4777 12219 4780
rect 12161 4771 12219 4777
rect 13078 4768 13084 4780
rect 13136 4768 13142 4820
rect 7668 4712 10079 4740
rect 10502 4743 10560 4749
rect 7564 4703 7622 4709
rect 10502 4709 10514 4743
rect 10548 4740 10560 4743
rect 10816 4743 10874 4749
rect 10816 4740 10828 4743
rect 10548 4712 10828 4740
rect 10548 4709 10560 4712
rect 10502 4703 10560 4709
rect 10816 4709 10828 4712
rect 10862 4740 10874 4743
rect 11236 4743 11294 4749
rect 11236 4740 11248 4743
rect 10862 4712 11248 4740
rect 10862 4709 10874 4712
rect 10816 4703 10874 4709
rect 11236 4709 11248 4712
rect 11282 4709 11294 4743
rect 12618 4740 12624 4752
rect 11236 4703 11294 4709
rect 12268 4712 12624 4740
rect 4338 4672 4344 4684
rect 4299 4644 4344 4672
rect 4338 4632 4344 4644
rect 4396 4632 4402 4684
rect 5365 4675 5423 4681
rect 5365 4641 5377 4675
rect 5411 4672 5423 4675
rect 5718 4672 5724 4684
rect 5411 4644 5724 4672
rect 5411 4641 5423 4644
rect 5365 4635 5423 4641
rect 5718 4632 5724 4644
rect 5776 4632 5782 4684
rect 6270 4672 6276 4684
rect 6231 4644 6276 4672
rect 6270 4632 6276 4644
rect 6328 4632 6334 4684
rect 12268 4681 12296 4712
rect 12618 4700 12624 4712
rect 12676 4700 12682 4752
rect 17402 4740 17408 4752
rect 13004 4712 17408 4740
rect 6909 4675 6967 4681
rect 6909 4641 6921 4675
rect 6955 4672 6967 4675
rect 7147 4675 7205 4681
rect 7147 4672 7159 4675
rect 6955 4644 7159 4672
rect 6955 4641 6967 4644
rect 6909 4635 6967 4641
rect 7147 4641 7159 4644
rect 7193 4672 7205 4675
rect 7651 4675 7709 4681
rect 7651 4672 7663 4675
rect 7193 4644 7663 4672
rect 7193 4641 7205 4644
rect 7147 4635 7205 4641
rect 7651 4641 7663 4644
rect 7697 4641 7709 4675
rect 7651 4635 7709 4641
rect 10415 4675 10473 4681
rect 10415 4641 10427 4675
rect 10461 4672 10473 4675
rect 10919 4675 10977 4681
rect 10919 4672 10931 4675
rect 10461 4644 10931 4672
rect 10461 4641 10473 4644
rect 10415 4635 10473 4641
rect 10919 4641 10931 4644
rect 10965 4672 10977 4675
rect 11157 4675 11215 4681
rect 11157 4672 11169 4675
rect 10965 4644 11169 4672
rect 10965 4641 10977 4644
rect 10919 4635 10977 4641
rect 11157 4641 11169 4644
rect 11203 4641 11215 4675
rect 11157 4635 11215 4641
rect 12253 4675 12311 4681
rect 12253 4641 12265 4675
rect 12299 4641 12311 4675
rect 13004 4672 13032 4712
rect 17402 4700 17408 4712
rect 17460 4700 17466 4752
rect 12253 4635 12311 4641
rect 12912 4644 13032 4672
rect 13081 4675 13139 4681
rect 4157 4607 4215 4613
rect 4157 4573 4169 4607
rect 4203 4573 4215 4607
rect 5074 4604 5080 4616
rect 5035 4576 5080 4604
rect 4157 4567 4215 4573
rect 5074 4564 5080 4576
rect 5132 4564 5138 4616
rect 5997 4607 6055 4613
rect 5997 4573 6009 4607
rect 6043 4604 6055 4607
rect 6086 4604 6092 4616
rect 6043 4576 6092 4604
rect 6043 4573 6055 4576
rect 5997 4567 6055 4573
rect 6086 4564 6092 4576
rect 6144 4564 6150 4616
rect 6730 4604 6736 4616
rect 6691 4576 6736 4604
rect 6730 4564 6736 4576
rect 6788 4564 6794 4616
rect 7006 4613 7012 4616
rect 7000 4567 7012 4613
rect 7064 4604 7070 4616
rect 11330 4604 11336 4616
rect 7064 4576 7100 4604
rect 11291 4576 11336 4604
rect 7006 4564 7012 4567
rect 7064 4564 7070 4576
rect 11330 4564 11336 4576
rect 11388 4564 11394 4616
rect 11422 4564 11428 4616
rect 11480 4604 11486 4616
rect 12912 4613 12940 4644
rect 13081 4641 13093 4675
rect 13127 4672 13139 4675
rect 13814 4672 13820 4684
rect 13127 4644 13820 4672
rect 13127 4641 13139 4644
rect 13081 4635 13139 4641
rect 13814 4632 13820 4644
rect 13872 4632 13878 4684
rect 11977 4607 12035 4613
rect 11977 4604 11989 4607
rect 11480 4576 11989 4604
rect 11480 4564 11486 4576
rect 11977 4573 11989 4576
rect 12023 4573 12035 4607
rect 12897 4607 12955 4613
rect 12897 4604 12909 4607
rect 11977 4567 12035 4573
rect 12544 4576 12909 4604
rect 6546 4536 6552 4548
rect 3436 4508 6552 4536
rect 3436 4477 3464 4508
rect 6546 4496 6552 4508
rect 6604 4496 6610 4548
rect 11088 4539 11146 4545
rect 11088 4505 11100 4539
rect 11134 4536 11146 4539
rect 11698 4536 11704 4548
rect 11134 4508 11704 4536
rect 11134 4505 11146 4508
rect 11088 4499 11146 4505
rect 11698 4496 11704 4508
rect 11756 4496 11762 4548
rect 11992 4536 12020 4567
rect 12544 4536 12572 4576
rect 12897 4573 12909 4576
rect 12943 4573 12955 4607
rect 12897 4567 12955 4573
rect 12986 4564 12992 4616
rect 13044 4604 13050 4616
rect 13173 4607 13231 4613
rect 13173 4604 13185 4607
rect 13044 4576 13185 4604
rect 13044 4564 13050 4576
rect 13173 4573 13185 4576
rect 13219 4573 13231 4607
rect 13173 4567 13231 4573
rect 13262 4564 13268 4616
rect 13320 4604 13326 4616
rect 14369 4607 14427 4613
rect 14369 4604 14381 4607
rect 13320 4576 14381 4604
rect 13320 4564 13326 4576
rect 14369 4573 14381 4576
rect 14415 4573 14427 4607
rect 14550 4604 14556 4616
rect 14511 4576 14556 4604
rect 14369 4567 14427 4573
rect 14550 4564 14556 4576
rect 14608 4604 14614 4616
rect 14734 4604 14740 4616
rect 14608 4576 14740 4604
rect 14608 4564 14614 4576
rect 14734 4564 14740 4576
rect 14792 4564 14798 4616
rect 11992 4508 12572 4536
rect 12618 4496 12624 4548
rect 12676 4536 12682 4548
rect 13280 4536 13308 4564
rect 12676 4508 13308 4536
rect 12676 4496 12682 4508
rect 3421 4471 3479 4477
rect 3421 4437 3433 4471
rect 3467 4437 3479 4471
rect 3421 4431 3479 4437
rect 4246 4428 4252 4480
rect 4304 4468 4310 4480
rect 4893 4471 4951 4477
rect 4893 4468 4905 4471
rect 4304 4440 4905 4468
rect 4304 4428 4310 4440
rect 4893 4437 4905 4440
rect 4939 4437 4951 4471
rect 4893 4431 4951 4437
rect 5718 4428 5724 4480
rect 5776 4468 5782 4480
rect 5813 4471 5871 4477
rect 5813 4468 5825 4471
rect 5776 4440 5825 4468
rect 5776 4428 5782 4440
rect 5813 4437 5825 4440
rect 5859 4437 5871 4471
rect 5813 4431 5871 4437
rect 7282 4428 7288 4480
rect 7340 4468 7346 4480
rect 8113 4471 8171 4477
rect 8113 4468 8125 4471
rect 7340 4440 8125 4468
rect 7340 4428 7346 4440
rect 8113 4437 8125 4440
rect 8159 4437 8171 4471
rect 8113 4431 8171 4437
rect 11793 4471 11851 4477
rect 11793 4437 11805 4471
rect 11839 4468 11851 4471
rect 11974 4468 11980 4480
rect 11839 4440 11980 4468
rect 11839 4437 11851 4440
rect 11793 4431 11851 4437
rect 11974 4428 11980 4440
rect 12032 4428 12038 4480
rect 12434 4428 12440 4480
rect 12492 4468 12498 4480
rect 12713 4471 12771 4477
rect 12713 4468 12725 4471
rect 12492 4440 12725 4468
rect 12492 4428 12498 4440
rect 12713 4437 12725 4440
rect 12759 4437 12771 4471
rect 12713 4431 12771 4437
rect 14737 4471 14795 4477
rect 14737 4437 14749 4471
rect 14783 4468 14795 4471
rect 15654 4468 15660 4480
rect 14783 4440 15660 4468
rect 14783 4437 14795 4440
rect 14737 4431 14795 4437
rect 15654 4428 15660 4440
rect 15712 4428 15718 4480
rect 1104 4378 19019 4400
rect 1104 4369 5388 4378
rect 1104 4335 1133 4369
rect 1167 4335 1225 4369
rect 1259 4335 1317 4369
rect 1351 4335 1409 4369
rect 1443 4335 1501 4369
rect 1535 4335 1593 4369
rect 1627 4335 1685 4369
rect 1719 4335 1777 4369
rect 1811 4335 1869 4369
rect 1903 4335 1961 4369
rect 1995 4335 2053 4369
rect 2087 4335 2145 4369
rect 2179 4335 2237 4369
rect 2271 4335 2329 4369
rect 2363 4335 2421 4369
rect 2455 4335 2513 4369
rect 2547 4335 2605 4369
rect 2639 4335 2697 4369
rect 2731 4335 2789 4369
rect 2823 4335 2881 4369
rect 2915 4335 2973 4369
rect 3007 4335 3065 4369
rect 3099 4335 3157 4369
rect 3191 4335 3249 4369
rect 3283 4335 3341 4369
rect 3375 4335 3433 4369
rect 3467 4335 3525 4369
rect 3559 4335 3617 4369
rect 3651 4335 3709 4369
rect 3743 4335 3801 4369
rect 3835 4335 3893 4369
rect 3927 4335 3985 4369
rect 4019 4335 4077 4369
rect 4111 4335 4169 4369
rect 4203 4335 4261 4369
rect 4295 4335 4353 4369
rect 4387 4335 4445 4369
rect 4479 4335 4537 4369
rect 4571 4335 4629 4369
rect 4663 4335 4721 4369
rect 4755 4335 4813 4369
rect 4847 4335 4905 4369
rect 4939 4335 4997 4369
rect 5031 4335 5089 4369
rect 5123 4335 5181 4369
rect 5215 4335 5273 4369
rect 5307 4335 5365 4369
rect 1104 4326 5388 4335
rect 5440 4326 5452 4378
rect 5504 4326 5516 4378
rect 5568 4369 5580 4378
rect 5632 4369 5644 4378
rect 5696 4369 9827 4378
rect 9879 4369 9891 4378
rect 5632 4335 5641 4369
rect 5696 4335 5733 4369
rect 5767 4335 5825 4369
rect 5859 4335 5917 4369
rect 5951 4335 6009 4369
rect 6043 4335 6101 4369
rect 6135 4335 6193 4369
rect 6227 4335 6285 4369
rect 6319 4335 6377 4369
rect 6411 4335 6469 4369
rect 6503 4335 6561 4369
rect 6595 4335 6653 4369
rect 6687 4335 6745 4369
rect 6779 4335 6837 4369
rect 6871 4335 6929 4369
rect 6963 4335 7021 4369
rect 7055 4335 7113 4369
rect 7147 4335 7205 4369
rect 7239 4335 7297 4369
rect 7331 4335 7389 4369
rect 7423 4335 7481 4369
rect 7515 4335 7573 4369
rect 7607 4335 7665 4369
rect 7699 4335 7757 4369
rect 7791 4335 7849 4369
rect 7883 4335 7941 4369
rect 7975 4335 8033 4369
rect 8067 4335 8125 4369
rect 8159 4335 8217 4369
rect 8251 4335 8309 4369
rect 8343 4335 8401 4369
rect 8435 4335 8493 4369
rect 8527 4335 8585 4369
rect 8619 4335 8677 4369
rect 8711 4335 8769 4369
rect 8803 4335 8861 4369
rect 8895 4335 8953 4369
rect 8987 4335 9045 4369
rect 9079 4335 9137 4369
rect 9171 4335 9229 4369
rect 9263 4335 9321 4369
rect 9355 4335 9413 4369
rect 9447 4335 9505 4369
rect 9539 4335 9597 4369
rect 9631 4335 9689 4369
rect 9723 4335 9781 4369
rect 9815 4335 9827 4369
rect 5568 4326 5580 4335
rect 5632 4326 5644 4335
rect 5696 4326 9827 4335
rect 9879 4326 9891 4335
rect 9943 4326 9955 4378
rect 10007 4326 10019 4378
rect 10071 4369 10083 4378
rect 10135 4369 14266 4378
rect 14318 4369 14330 4378
rect 14382 4369 14394 4378
rect 10135 4335 10149 4369
rect 10183 4335 10241 4369
rect 10275 4335 10333 4369
rect 10367 4335 10425 4369
rect 10459 4335 10517 4369
rect 10551 4335 10609 4369
rect 10643 4335 10701 4369
rect 10735 4335 10793 4369
rect 10827 4335 10885 4369
rect 10919 4335 10977 4369
rect 11011 4335 11069 4369
rect 11103 4335 11161 4369
rect 11195 4335 11253 4369
rect 11287 4335 11345 4369
rect 11379 4335 11437 4369
rect 11471 4335 11529 4369
rect 11563 4335 11621 4369
rect 11655 4335 11713 4369
rect 11747 4335 11805 4369
rect 11839 4335 11897 4369
rect 11931 4335 11989 4369
rect 12023 4335 12081 4369
rect 12115 4335 12173 4369
rect 12207 4335 12265 4369
rect 12299 4335 12357 4369
rect 12391 4335 12449 4369
rect 12483 4335 12541 4369
rect 12575 4335 12633 4369
rect 12667 4335 12725 4369
rect 12759 4335 12817 4369
rect 12851 4335 12909 4369
rect 12943 4335 13001 4369
rect 13035 4335 13093 4369
rect 13127 4335 13185 4369
rect 13219 4335 13277 4369
rect 13311 4335 13369 4369
rect 13403 4335 13461 4369
rect 13495 4335 13553 4369
rect 13587 4335 13645 4369
rect 13679 4335 13737 4369
rect 13771 4335 13829 4369
rect 13863 4335 13921 4369
rect 13955 4335 14013 4369
rect 14047 4335 14105 4369
rect 14139 4335 14197 4369
rect 14231 4335 14266 4369
rect 14323 4335 14330 4369
rect 10071 4326 10083 4335
rect 10135 4326 14266 4335
rect 14318 4326 14330 4335
rect 14382 4326 14394 4335
rect 14446 4326 14458 4378
rect 14510 4326 14522 4378
rect 14574 4369 18705 4378
rect 14599 4335 14657 4369
rect 14691 4335 14749 4369
rect 14783 4335 14841 4369
rect 14875 4335 14933 4369
rect 14967 4335 15025 4369
rect 15059 4335 15117 4369
rect 15151 4335 15209 4369
rect 15243 4335 15301 4369
rect 15335 4335 15393 4369
rect 15427 4335 15485 4369
rect 15519 4335 15577 4369
rect 15611 4335 15669 4369
rect 15703 4335 15761 4369
rect 15795 4335 15853 4369
rect 15887 4335 15945 4369
rect 15979 4335 16037 4369
rect 16071 4335 16129 4369
rect 16163 4335 16221 4369
rect 16255 4335 16313 4369
rect 16347 4335 16405 4369
rect 16439 4335 16497 4369
rect 16531 4335 16589 4369
rect 16623 4335 16681 4369
rect 16715 4335 16773 4369
rect 16807 4335 16865 4369
rect 16899 4335 16957 4369
rect 16991 4335 17049 4369
rect 17083 4335 17141 4369
rect 17175 4335 17233 4369
rect 17267 4335 17325 4369
rect 17359 4335 17417 4369
rect 17451 4335 17509 4369
rect 17543 4335 17601 4369
rect 17635 4335 17693 4369
rect 17727 4335 17785 4369
rect 17819 4335 17877 4369
rect 17911 4335 17969 4369
rect 18003 4335 18061 4369
rect 18095 4335 18153 4369
rect 18187 4335 18245 4369
rect 18279 4335 18337 4369
rect 18371 4335 18429 4369
rect 18463 4335 18521 4369
rect 18555 4335 18613 4369
rect 18647 4335 18705 4369
rect 14574 4326 18705 4335
rect 18757 4326 18769 4378
rect 18821 4369 18833 4378
rect 18831 4335 18833 4369
rect 18821 4326 18833 4335
rect 18885 4326 18897 4378
rect 18949 4326 18961 4378
rect 19013 4326 19019 4378
rect 1104 4304 19019 4326
rect 2590 4264 2596 4276
rect 2551 4236 2596 4264
rect 2590 4224 2596 4236
rect 2648 4224 2654 4276
rect 4614 4264 4620 4276
rect 4575 4236 4620 4264
rect 4614 4224 4620 4236
rect 4672 4224 4678 4276
rect 4706 4224 4712 4276
rect 4764 4264 4770 4276
rect 11514 4264 11520 4276
rect 4764 4236 11520 4264
rect 4764 4224 4770 4236
rect 11514 4224 11520 4236
rect 11572 4224 11578 4276
rect 13081 4267 13139 4273
rect 13081 4233 13093 4267
rect 13127 4264 13139 4267
rect 13446 4264 13452 4276
rect 13127 4236 13452 4264
rect 13127 4233 13139 4236
rect 13081 4227 13139 4233
rect 13446 4224 13452 4236
rect 13504 4224 13510 4276
rect 4798 4196 4804 4208
rect 3804 4168 4804 4196
rect 1946 4128 1952 4140
rect 1907 4100 1952 4128
rect 1946 4088 1952 4100
rect 2004 4088 2010 4140
rect 3717 4131 3775 4137
rect 3717 4097 3729 4131
rect 3763 4128 3775 4131
rect 3804 4128 3832 4168
rect 4798 4156 4804 4168
rect 4856 4156 4862 4208
rect 5552 4168 6040 4196
rect 3970 4128 3976 4140
rect 3763 4100 3832 4128
rect 3883 4100 3976 4128
rect 3763 4097 3775 4100
rect 3717 4091 3775 4097
rect 3970 4088 3976 4100
rect 4028 4128 4034 4140
rect 5552 4128 5580 4168
rect 4028 4100 5580 4128
rect 4028 4088 4034 4100
rect 5718 4088 5724 4140
rect 5776 4137 5782 4140
rect 6012 4137 6040 4168
rect 6086 4156 6092 4208
rect 6144 4196 6150 4208
rect 6144 4168 7144 4196
rect 6144 4156 6150 4168
rect 5776 4128 5788 4137
rect 5997 4131 6055 4137
rect 5776 4100 5821 4128
rect 5776 4091 5788 4100
rect 5997 4097 6009 4131
rect 6043 4128 6055 4131
rect 6730 4128 6736 4140
rect 6043 4100 6736 4128
rect 6043 4097 6055 4100
rect 5997 4091 6055 4097
rect 5776 4088 5782 4091
rect 6730 4088 6736 4100
rect 6788 4088 6794 4140
rect 7116 4137 7144 4168
rect 7374 4156 7380 4208
rect 7432 4196 7438 4208
rect 7837 4199 7895 4205
rect 7837 4196 7849 4199
rect 7432 4168 7849 4196
rect 7432 4156 7438 4168
rect 7837 4165 7849 4168
rect 7883 4165 7895 4199
rect 7837 4159 7895 4165
rect 9306 4156 9312 4208
rect 9364 4196 9370 4208
rect 11422 4196 11428 4208
rect 9364 4168 11428 4196
rect 9364 4156 9370 4168
rect 7101 4131 7159 4137
rect 7101 4097 7113 4131
rect 7147 4128 7159 4131
rect 7190 4128 7196 4140
rect 7147 4100 7196 4128
rect 7147 4097 7159 4100
rect 7101 4091 7159 4097
rect 7190 4088 7196 4100
rect 7248 4088 7254 4140
rect 7285 4131 7343 4137
rect 7285 4097 7297 4131
rect 7331 4128 7343 4131
rect 9214 4128 9220 4140
rect 7331 4100 9220 4128
rect 7331 4097 7343 4100
rect 7285 4091 7343 4097
rect 9214 4088 9220 4100
rect 9272 4088 9278 4140
rect 10704 4137 10732 4168
rect 11422 4156 11428 4168
rect 11480 4156 11486 4208
rect 11974 4205 11980 4208
rect 11968 4196 11980 4205
rect 11935 4168 11980 4196
rect 11968 4159 11980 4168
rect 11974 4156 11980 4159
rect 12032 4156 12038 4208
rect 15488 4168 15792 4196
rect 10689 4131 10747 4137
rect 10689 4097 10701 4131
rect 10735 4097 10747 4131
rect 11330 4128 11336 4140
rect 10689 4091 10747 4097
rect 10888 4100 11336 4128
rect 3055 4063 3113 4069
rect 3055 4029 3067 4063
rect 3101 4060 3113 4063
rect 3559 4063 3617 4069
rect 3559 4060 3571 4063
rect 3101 4032 3571 4060
rect 3101 4029 3113 4032
rect 3055 4023 3113 4029
rect 3559 4029 3571 4032
rect 3605 4060 3617 4063
rect 3797 4063 3855 4069
rect 3797 4060 3809 4063
rect 3605 4032 3809 4060
rect 3605 4029 3617 4032
rect 3559 4023 3617 4029
rect 3797 4029 3809 4032
rect 3843 4029 3855 4063
rect 3797 4023 3855 4029
rect 5079 4063 5137 4069
rect 5079 4029 5091 4063
rect 5125 4060 5137 4063
rect 5583 4063 5641 4069
rect 5583 4060 5595 4063
rect 5125 4032 5595 4060
rect 5125 4029 5137 4032
rect 5079 4023 5137 4029
rect 5583 4029 5595 4032
rect 5629 4060 5641 4063
rect 5821 4063 5879 4069
rect 5821 4060 5833 4063
rect 5629 4032 5833 4060
rect 5629 4029 5641 4032
rect 5583 4023 5641 4029
rect 5821 4029 5833 4032
rect 5867 4029 5879 4063
rect 5821 4023 5879 4029
rect 6454 4020 6460 4072
rect 6512 4060 6518 4072
rect 6914 4060 6920 4072
rect 6512 4032 6920 4060
rect 6512 4020 6518 4032
rect 6914 4020 6920 4032
rect 6972 4020 6978 4072
rect 7377 4063 7435 4069
rect 7377 4060 7389 4063
rect 7208 4032 7389 4060
rect 2133 3995 2191 4001
rect 2133 3961 2145 3995
rect 2179 3992 2191 3995
rect 3142 3995 3200 4001
rect 2179 3964 2774 3992
rect 2179 3961 2191 3964
rect 2133 3955 2191 3961
rect 2746 3924 2774 3964
rect 3142 3961 3154 3995
rect 3188 3992 3200 3995
rect 3456 3995 3514 4001
rect 3456 3992 3468 3995
rect 3188 3964 3468 3992
rect 3188 3961 3200 3964
rect 3142 3955 3200 3961
rect 3456 3961 3468 3964
rect 3502 3992 3514 3995
rect 3876 3995 3934 4001
rect 3876 3992 3888 3995
rect 3502 3964 3888 3992
rect 3502 3961 3514 3964
rect 3456 3955 3514 3961
rect 3876 3961 3888 3964
rect 3922 3961 3934 3995
rect 3876 3955 3934 3961
rect 5166 3995 5224 4001
rect 5166 3961 5178 3995
rect 5212 3992 5224 3995
rect 5480 3995 5538 4001
rect 5480 3992 5492 3995
rect 5212 3964 5492 3992
rect 5212 3961 5224 3964
rect 5166 3955 5224 3961
rect 5480 3961 5492 3964
rect 5526 3992 5538 3995
rect 5900 3995 5958 4001
rect 5900 3992 5912 3995
rect 5526 3964 5912 3992
rect 5526 3961 5538 3964
rect 5480 3955 5538 3961
rect 5900 3961 5912 3964
rect 5946 3961 5958 3995
rect 5900 3955 5958 3961
rect 6546 3952 6552 4004
rect 6604 3992 6610 4004
rect 7208 3992 7236 4032
rect 7377 4029 7389 4032
rect 7423 4060 7435 4063
rect 8386 4060 8392 4072
rect 7423 4032 8392 4060
rect 7423 4029 7435 4032
rect 7377 4023 7435 4029
rect 8386 4020 8392 4032
rect 8444 4020 8450 4072
rect 9582 4060 9588 4072
rect 9543 4032 9588 4060
rect 9582 4020 9588 4032
rect 9640 4060 9646 4072
rect 10888 4060 10916 4100
rect 11330 4088 11336 4100
rect 11388 4128 11394 4140
rect 11701 4131 11759 4137
rect 11701 4128 11713 4131
rect 11388 4100 11713 4128
rect 11388 4088 11394 4100
rect 11701 4097 11713 4100
rect 11747 4128 11759 4131
rect 11790 4128 11796 4140
rect 11747 4100 11796 4128
rect 11747 4097 11759 4100
rect 11701 4091 11759 4097
rect 11790 4088 11796 4100
rect 11848 4088 11854 4140
rect 14826 4088 14832 4140
rect 14884 4128 14890 4140
rect 15488 4128 15516 4168
rect 15654 4128 15660 4140
rect 14884 4100 15516 4128
rect 15615 4100 15660 4128
rect 14884 4088 14890 4100
rect 15654 4088 15660 4100
rect 15712 4088 15718 4140
rect 9640 4032 10916 4060
rect 9640 4020 9646 4032
rect 10962 4020 10968 4072
rect 11020 4060 11026 4072
rect 11877 4063 11935 4069
rect 11020 4032 11065 4060
rect 11020 4020 11026 4032
rect 11877 4029 11889 4063
rect 11923 4060 11935 4063
rect 12115 4063 12173 4069
rect 12115 4060 12127 4063
rect 11923 4032 12127 4060
rect 11923 4029 11935 4032
rect 11877 4023 11935 4029
rect 12115 4029 12127 4032
rect 12161 4060 12173 4063
rect 12619 4063 12677 4069
rect 12619 4060 12631 4063
rect 12161 4032 12631 4060
rect 12161 4029 12173 4032
rect 12115 4023 12173 4029
rect 12619 4029 12631 4032
rect 12665 4029 12677 4063
rect 12619 4023 12677 4029
rect 14734 4020 14740 4072
rect 14792 4060 14798 4072
rect 15764 4060 15792 4168
rect 17037 4131 17095 4137
rect 17037 4097 17049 4131
rect 17083 4097 17095 4131
rect 17037 4091 17095 4097
rect 16853 4063 16911 4069
rect 16853 4060 16865 4063
rect 14792 4032 15700 4060
rect 15764 4032 16865 4060
rect 14792 4020 14798 4032
rect 10870 3992 10876 4004
rect 6604 3964 7236 3992
rect 10831 3964 10876 3992
rect 6604 3952 6610 3964
rect 10870 3952 10876 3964
rect 10928 3952 10934 4004
rect 11798 3995 11856 4001
rect 11798 3961 11810 3995
rect 11844 3992 11856 3995
rect 12218 3995 12276 4001
rect 12218 3992 12230 3995
rect 11844 3964 12230 3992
rect 11844 3961 11856 3964
rect 11798 3955 11856 3961
rect 12218 3961 12230 3964
rect 12264 3992 12276 3995
rect 12532 3995 12590 4001
rect 12532 3992 12544 3995
rect 12264 3964 12544 3992
rect 12264 3961 12276 3964
rect 12218 3955 12276 3961
rect 12532 3961 12544 3964
rect 12578 3961 12590 3995
rect 15672 3992 15700 4032
rect 16853 4029 16865 4032
rect 16899 4029 16911 4063
rect 16853 4023 16911 4029
rect 16390 3992 16396 4004
rect 15672 3964 16396 3992
rect 12532 3955 12590 3961
rect 16390 3952 16396 3964
rect 16448 3992 16454 4004
rect 17052 3992 17080 4091
rect 16448 3964 17080 3992
rect 16448 3952 16454 3964
rect 4522 3924 4528 3936
rect 2746 3896 4528 3924
rect 4522 3884 4528 3896
rect 4580 3884 4586 3936
rect 6914 3924 6920 3936
rect 6875 3896 6920 3924
rect 6914 3884 6920 3896
rect 6972 3884 6978 3936
rect 10502 3924 10508 3936
rect 10463 3896 10508 3924
rect 10502 3884 10508 3896
rect 10560 3884 10566 3936
rect 11606 3884 11612 3936
rect 11664 3924 11670 3936
rect 15473 3927 15531 3933
rect 15473 3924 15485 3927
rect 11664 3896 15485 3924
rect 11664 3884 11670 3896
rect 15473 3893 15485 3896
rect 15519 3893 15531 3927
rect 17218 3924 17224 3936
rect 17179 3896 17224 3924
rect 15473 3887 15531 3893
rect 17218 3884 17224 3896
rect 17276 3884 17282 3936
rect 1104 3834 18860 3856
rect 1104 3825 3169 3834
rect 1104 3791 1133 3825
rect 1167 3791 1225 3825
rect 1259 3791 1317 3825
rect 1351 3791 1409 3825
rect 1443 3791 1501 3825
rect 1535 3791 1593 3825
rect 1627 3791 1685 3825
rect 1719 3791 1777 3825
rect 1811 3791 1869 3825
rect 1903 3791 1961 3825
rect 1995 3791 2053 3825
rect 2087 3791 2145 3825
rect 2179 3791 2237 3825
rect 2271 3791 2329 3825
rect 2363 3791 2421 3825
rect 2455 3791 2513 3825
rect 2547 3791 2605 3825
rect 2639 3791 2697 3825
rect 2731 3791 2789 3825
rect 2823 3791 2881 3825
rect 2915 3791 2973 3825
rect 3007 3791 3065 3825
rect 3099 3791 3157 3825
rect 1104 3782 3169 3791
rect 3221 3782 3233 3834
rect 3285 3782 3297 3834
rect 3349 3825 3361 3834
rect 3349 3782 3361 3791
rect 3413 3782 3425 3834
rect 3477 3825 7608 3834
rect 3477 3791 3525 3825
rect 3559 3791 3617 3825
rect 3651 3791 3709 3825
rect 3743 3791 3801 3825
rect 3835 3791 3893 3825
rect 3927 3791 3985 3825
rect 4019 3791 4077 3825
rect 4111 3791 4169 3825
rect 4203 3791 4261 3825
rect 4295 3791 4353 3825
rect 4387 3791 4445 3825
rect 4479 3791 4537 3825
rect 4571 3791 4629 3825
rect 4663 3791 4721 3825
rect 4755 3791 4813 3825
rect 4847 3791 4905 3825
rect 4939 3791 4997 3825
rect 5031 3791 5089 3825
rect 5123 3791 5181 3825
rect 5215 3791 5273 3825
rect 5307 3791 5365 3825
rect 5399 3791 5457 3825
rect 5491 3791 5549 3825
rect 5583 3791 5641 3825
rect 5675 3791 5733 3825
rect 5767 3791 5825 3825
rect 5859 3791 5917 3825
rect 5951 3791 6009 3825
rect 6043 3791 6101 3825
rect 6135 3791 6193 3825
rect 6227 3791 6285 3825
rect 6319 3791 6377 3825
rect 6411 3791 6469 3825
rect 6503 3791 6561 3825
rect 6595 3791 6653 3825
rect 6687 3791 6745 3825
rect 6779 3791 6837 3825
rect 6871 3791 6929 3825
rect 6963 3791 7021 3825
rect 7055 3791 7113 3825
rect 7147 3791 7205 3825
rect 7239 3791 7297 3825
rect 7331 3791 7389 3825
rect 7423 3791 7481 3825
rect 7515 3791 7573 3825
rect 7607 3791 7608 3825
rect 3477 3782 7608 3791
rect 7660 3825 7672 3834
rect 7660 3791 7665 3825
rect 7660 3782 7672 3791
rect 7724 3782 7736 3834
rect 7788 3825 7800 3834
rect 7852 3825 7864 3834
rect 7916 3825 12047 3834
rect 12099 3825 12111 3834
rect 12163 3825 12175 3834
rect 7791 3791 7800 3825
rect 7916 3791 7941 3825
rect 7975 3791 8033 3825
rect 8067 3791 8125 3825
rect 8159 3791 8217 3825
rect 8251 3791 8309 3825
rect 8343 3791 8401 3825
rect 8435 3791 8493 3825
rect 8527 3791 8585 3825
rect 8619 3791 8677 3825
rect 8711 3791 8769 3825
rect 8803 3791 8861 3825
rect 8895 3791 8953 3825
rect 8987 3791 9045 3825
rect 9079 3791 9137 3825
rect 9171 3791 9229 3825
rect 9263 3791 9321 3825
rect 9355 3791 9413 3825
rect 9447 3791 9505 3825
rect 9539 3791 9597 3825
rect 9631 3791 9689 3825
rect 9723 3791 9781 3825
rect 9815 3791 9873 3825
rect 9907 3791 9965 3825
rect 9999 3791 10057 3825
rect 10091 3791 10149 3825
rect 10183 3791 10241 3825
rect 10275 3791 10333 3825
rect 10367 3791 10425 3825
rect 10459 3791 10517 3825
rect 10551 3791 10609 3825
rect 10643 3791 10701 3825
rect 10735 3791 10793 3825
rect 10827 3791 10885 3825
rect 10919 3791 10977 3825
rect 11011 3791 11069 3825
rect 11103 3791 11161 3825
rect 11195 3791 11253 3825
rect 11287 3791 11345 3825
rect 11379 3791 11437 3825
rect 11471 3791 11529 3825
rect 11563 3791 11621 3825
rect 11655 3791 11713 3825
rect 11747 3791 11805 3825
rect 11839 3791 11897 3825
rect 11931 3791 11989 3825
rect 12023 3791 12047 3825
rect 12163 3791 12173 3825
rect 7788 3782 7800 3791
rect 7852 3782 7864 3791
rect 7916 3782 12047 3791
rect 12099 3782 12111 3791
rect 12163 3782 12175 3791
rect 12227 3782 12239 3834
rect 12291 3825 12303 3834
rect 12299 3791 12303 3825
rect 12291 3782 12303 3791
rect 12355 3825 16486 3834
rect 12355 3791 12357 3825
rect 12391 3791 12449 3825
rect 12483 3791 12541 3825
rect 12575 3791 12633 3825
rect 12667 3791 12725 3825
rect 12759 3791 12817 3825
rect 12851 3791 12909 3825
rect 12943 3791 13001 3825
rect 13035 3791 13093 3825
rect 13127 3791 13185 3825
rect 13219 3791 13277 3825
rect 13311 3791 13369 3825
rect 13403 3791 13461 3825
rect 13495 3791 13553 3825
rect 13587 3791 13645 3825
rect 13679 3791 13737 3825
rect 13771 3791 13829 3825
rect 13863 3791 13921 3825
rect 13955 3791 14013 3825
rect 14047 3791 14105 3825
rect 14139 3791 14197 3825
rect 14231 3791 14289 3825
rect 14323 3791 14381 3825
rect 14415 3791 14473 3825
rect 14507 3791 14565 3825
rect 14599 3791 14657 3825
rect 14691 3791 14749 3825
rect 14783 3791 14841 3825
rect 14875 3791 14933 3825
rect 14967 3791 15025 3825
rect 15059 3791 15117 3825
rect 15151 3791 15209 3825
rect 15243 3791 15301 3825
rect 15335 3791 15393 3825
rect 15427 3791 15485 3825
rect 15519 3791 15577 3825
rect 15611 3791 15669 3825
rect 15703 3791 15761 3825
rect 15795 3791 15853 3825
rect 15887 3791 15945 3825
rect 15979 3791 16037 3825
rect 16071 3791 16129 3825
rect 16163 3791 16221 3825
rect 16255 3791 16313 3825
rect 16347 3791 16405 3825
rect 16439 3791 16486 3825
rect 12355 3782 16486 3791
rect 16538 3782 16550 3834
rect 16602 3825 16614 3834
rect 16602 3782 16614 3791
rect 16666 3782 16678 3834
rect 16730 3782 16742 3834
rect 16794 3825 18860 3834
rect 16807 3791 16865 3825
rect 16899 3791 16957 3825
rect 16991 3791 17049 3825
rect 17083 3791 17141 3825
rect 17175 3791 17233 3825
rect 17267 3791 17325 3825
rect 17359 3791 17417 3825
rect 17451 3791 17509 3825
rect 17543 3791 17601 3825
rect 17635 3791 17693 3825
rect 17727 3791 17785 3825
rect 17819 3791 17877 3825
rect 17911 3791 17969 3825
rect 18003 3791 18061 3825
rect 18095 3791 18153 3825
rect 18187 3791 18245 3825
rect 18279 3791 18337 3825
rect 18371 3791 18429 3825
rect 18463 3791 18521 3825
rect 18555 3791 18613 3825
rect 18647 3791 18705 3825
rect 18739 3791 18797 3825
rect 18831 3791 18860 3825
rect 16794 3782 18860 3791
rect 1104 3760 18860 3782
rect 3421 3723 3479 3729
rect 3421 3689 3433 3723
rect 3467 3720 3479 3723
rect 6454 3720 6460 3732
rect 3467 3692 6460 3720
rect 3467 3689 3479 3692
rect 3421 3683 3479 3689
rect 6454 3680 6460 3692
rect 6512 3680 6518 3732
rect 6638 3720 6644 3732
rect 6599 3692 6644 3720
rect 6638 3680 6644 3692
rect 6696 3680 6702 3732
rect 8573 3723 8631 3729
rect 8573 3689 8585 3723
rect 8619 3720 8631 3723
rect 10134 3720 10140 3732
rect 8619 3692 10140 3720
rect 8619 3689 8631 3692
rect 8573 3683 8631 3689
rect 10134 3680 10140 3692
rect 10192 3680 10198 3732
rect 11149 3723 11207 3729
rect 11149 3689 11161 3723
rect 11195 3720 11207 3723
rect 12526 3720 12532 3732
rect 11195 3692 12532 3720
rect 11195 3689 11207 3692
rect 11149 3683 11207 3689
rect 12526 3680 12532 3692
rect 12584 3680 12590 3732
rect 13173 3723 13231 3729
rect 13173 3689 13185 3723
rect 13219 3720 13231 3723
rect 14642 3720 14648 3732
rect 13219 3692 14648 3720
rect 13219 3689 13231 3692
rect 13173 3683 13231 3689
rect 14642 3680 14648 3692
rect 14700 3680 14706 3732
rect 2138 3655 2196 3661
rect 2138 3621 2150 3655
rect 2184 3652 2196 3655
rect 2558 3655 2616 3661
rect 2558 3652 2570 3655
rect 2184 3624 2570 3652
rect 2184 3621 2196 3624
rect 2138 3615 2196 3621
rect 2558 3621 2570 3624
rect 2604 3652 2616 3655
rect 2872 3655 2930 3661
rect 2872 3652 2884 3655
rect 2604 3624 2884 3652
rect 2604 3621 2616 3624
rect 2558 3615 2616 3621
rect 2872 3621 2884 3624
rect 2918 3621 2930 3655
rect 2872 3615 2930 3621
rect 4070 3655 4128 3661
rect 4070 3621 4082 3655
rect 4116 3652 4128 3655
rect 4490 3655 4548 3661
rect 4490 3652 4502 3655
rect 4116 3624 4502 3652
rect 4116 3621 4128 3624
rect 4070 3615 4128 3621
rect 4490 3621 4502 3624
rect 4536 3652 4548 3655
rect 4804 3655 4862 3661
rect 4804 3652 4816 3655
rect 4536 3624 4816 3652
rect 4536 3621 4548 3624
rect 4490 3615 4548 3621
rect 4804 3621 4816 3624
rect 4850 3621 4862 3655
rect 4804 3615 4862 3621
rect 6730 3612 6736 3664
rect 6788 3612 6794 3664
rect 7290 3655 7348 3661
rect 7290 3621 7302 3655
rect 7336 3652 7348 3655
rect 7710 3655 7768 3661
rect 7710 3652 7722 3655
rect 7336 3624 7722 3652
rect 7336 3621 7348 3624
rect 7290 3615 7348 3621
rect 7710 3621 7722 3624
rect 7756 3652 7768 3655
rect 8024 3655 8082 3661
rect 8024 3652 8036 3655
rect 7756 3624 8036 3652
rect 7756 3621 7768 3624
rect 7710 3615 7768 3621
rect 8024 3621 8036 3624
rect 8070 3621 8082 3655
rect 8024 3615 8082 3621
rect 9866 3655 9924 3661
rect 9866 3621 9878 3655
rect 9912 3652 9924 3655
rect 10286 3655 10344 3661
rect 10286 3652 10298 3655
rect 9912 3624 10298 3652
rect 9912 3621 9924 3624
rect 9866 3615 9924 3621
rect 10286 3621 10298 3624
rect 10332 3652 10344 3655
rect 10600 3655 10658 3661
rect 10600 3652 10612 3655
rect 10332 3624 10612 3652
rect 10332 3621 10344 3624
rect 10286 3615 10344 3621
rect 10600 3621 10612 3624
rect 10646 3621 10658 3655
rect 10600 3615 10658 3621
rect 11890 3655 11948 3661
rect 11890 3621 11902 3655
rect 11936 3652 11948 3655
rect 12310 3655 12368 3661
rect 12310 3652 12322 3655
rect 11936 3624 12322 3652
rect 11936 3621 11948 3624
rect 11890 3615 11948 3621
rect 12310 3621 12322 3624
rect 12356 3652 12368 3655
rect 12624 3655 12682 3661
rect 12624 3652 12636 3655
rect 12356 3624 12636 3652
rect 12356 3621 12368 3624
rect 12310 3615 12368 3621
rect 12624 3621 12636 3624
rect 12670 3621 12682 3655
rect 12624 3615 12682 3621
rect 2217 3587 2275 3593
rect 2217 3553 2229 3587
rect 2263 3584 2275 3587
rect 2455 3587 2513 3593
rect 2455 3584 2467 3587
rect 2263 3556 2467 3584
rect 2263 3553 2275 3556
rect 2217 3547 2275 3553
rect 2455 3553 2467 3556
rect 2501 3584 2513 3587
rect 2959 3587 3017 3593
rect 2959 3584 2971 3587
rect 2501 3556 2971 3584
rect 2501 3553 2513 3556
rect 2455 3547 2513 3553
rect 2959 3553 2971 3556
rect 3005 3553 3017 3587
rect 3970 3584 3976 3596
rect 3931 3556 3976 3584
rect 2959 3547 3017 3553
rect 3970 3544 3976 3556
rect 4028 3544 4034 3596
rect 4149 3587 4207 3593
rect 4149 3553 4161 3587
rect 4195 3584 4207 3587
rect 4387 3587 4445 3593
rect 4387 3584 4399 3587
rect 4195 3556 4399 3584
rect 4195 3553 4207 3556
rect 4149 3547 4207 3553
rect 4387 3553 4399 3556
rect 4433 3584 4445 3587
rect 4891 3587 4949 3593
rect 4891 3584 4903 3587
rect 4433 3556 4903 3584
rect 4433 3553 4445 3556
rect 4387 3547 4445 3553
rect 4891 3553 4903 3556
rect 4937 3553 4949 3587
rect 6748 3584 6776 3612
rect 7193 3587 7251 3593
rect 7193 3584 7205 3587
rect 6748 3556 7205 3584
rect 4891 3547 4949 3553
rect 7193 3553 7205 3556
rect 7239 3553 7251 3587
rect 7193 3547 7251 3553
rect 7369 3587 7427 3593
rect 7369 3553 7381 3587
rect 7415 3584 7427 3587
rect 7607 3587 7665 3593
rect 7607 3584 7619 3587
rect 7415 3556 7619 3584
rect 7415 3553 7427 3556
rect 7369 3547 7427 3553
rect 7607 3553 7619 3556
rect 7653 3584 7665 3587
rect 8111 3587 8169 3593
rect 8111 3584 8123 3587
rect 7653 3556 8123 3584
rect 7653 3553 7665 3556
rect 7607 3547 7665 3553
rect 8111 3553 8123 3556
rect 8157 3553 8169 3587
rect 8111 3547 8169 3553
rect 9582 3544 9588 3596
rect 9640 3584 9646 3596
rect 9769 3587 9827 3593
rect 9769 3584 9781 3587
rect 9640 3556 9781 3584
rect 9640 3544 9646 3556
rect 9769 3553 9781 3556
rect 9815 3553 9827 3587
rect 9769 3547 9827 3553
rect 9945 3587 10003 3593
rect 9945 3553 9957 3587
rect 9991 3584 10003 3587
rect 10183 3587 10241 3593
rect 10183 3584 10195 3587
rect 9991 3556 10195 3584
rect 9991 3553 10003 3556
rect 9945 3547 10003 3553
rect 10183 3553 10195 3556
rect 10229 3584 10241 3587
rect 10687 3587 10745 3593
rect 10687 3584 10699 3587
rect 10229 3556 10699 3584
rect 10229 3553 10241 3556
rect 10183 3547 10241 3553
rect 10687 3553 10699 3556
rect 10733 3553 10745 3587
rect 11790 3584 11796 3596
rect 11751 3556 11796 3584
rect 10687 3547 10745 3553
rect 11790 3544 11796 3556
rect 11848 3544 11854 3596
rect 11969 3587 12027 3593
rect 11969 3553 11981 3587
rect 12015 3584 12027 3587
rect 12207 3587 12265 3593
rect 12207 3584 12219 3587
rect 12015 3556 12219 3584
rect 12015 3553 12027 3556
rect 11969 3547 12027 3553
rect 12207 3553 12219 3556
rect 12253 3584 12265 3587
rect 12711 3587 12769 3593
rect 12711 3584 12723 3587
rect 12253 3556 12723 3584
rect 12253 3553 12265 3556
rect 12207 3547 12265 3553
rect 12711 3553 12723 3556
rect 12757 3553 12769 3587
rect 17494 3584 17500 3596
rect 12711 3547 12769 3553
rect 12820 3556 17500 3584
rect 2038 3516 2044 3528
rect 1999 3488 2044 3516
rect 2038 3476 2044 3488
rect 2096 3476 2102 3528
rect 4246 3525 4252 3528
rect 4240 3516 4252 3525
rect 4207 3488 4252 3516
rect 4240 3479 4252 3488
rect 4246 3476 4252 3479
rect 4304 3476 4310 3528
rect 6086 3476 6092 3528
rect 6144 3516 6150 3528
rect 6457 3519 6515 3525
rect 6457 3516 6469 3519
rect 6144 3488 6469 3516
rect 6144 3476 6150 3488
rect 6457 3485 6469 3488
rect 6503 3485 6515 3519
rect 6457 3479 6515 3485
rect 6546 3476 6552 3528
rect 6604 3516 6610 3528
rect 6733 3519 6791 3525
rect 6733 3516 6745 3519
rect 6604 3488 6745 3516
rect 6604 3476 6610 3488
rect 6733 3485 6745 3488
rect 6779 3516 6791 3519
rect 6822 3516 6828 3528
rect 6779 3488 6828 3516
rect 6779 3485 6791 3488
rect 6733 3479 6791 3485
rect 6822 3476 6828 3488
rect 6880 3476 6886 3528
rect 7460 3519 7518 3525
rect 7460 3485 7472 3519
rect 7506 3516 7518 3519
rect 9122 3516 9128 3528
rect 7506 3488 9128 3516
rect 7506 3485 7518 3488
rect 7460 3479 7518 3485
rect 9122 3476 9128 3488
rect 9180 3476 9186 3528
rect 10036 3519 10094 3525
rect 10036 3485 10048 3519
rect 10082 3516 10094 3519
rect 10502 3516 10508 3528
rect 10082 3488 10508 3516
rect 10082 3485 10094 3488
rect 10036 3479 10094 3485
rect 10502 3476 10508 3488
rect 10560 3476 10566 3528
rect 12060 3519 12118 3525
rect 12060 3485 12072 3519
rect 12106 3516 12118 3519
rect 12434 3516 12440 3528
rect 12106 3488 12440 3516
rect 12106 3485 12118 3488
rect 12060 3479 12118 3485
rect 12434 3476 12440 3488
rect 12492 3476 12498 3528
rect 2308 3451 2366 3457
rect 2308 3417 2320 3451
rect 2354 3448 2366 3451
rect 6273 3451 6331 3457
rect 6273 3448 6285 3451
rect 2354 3420 6285 3448
rect 2354 3417 2366 3420
rect 2308 3411 2366 3417
rect 6273 3417 6285 3420
rect 6319 3417 6331 3451
rect 6273 3411 6331 3417
rect 5353 3383 5411 3389
rect 5353 3349 5365 3383
rect 5399 3380 5411 3383
rect 7098 3380 7104 3392
rect 5399 3352 7104 3380
rect 5399 3349 5411 3352
rect 5353 3343 5411 3349
rect 7098 3340 7104 3352
rect 7156 3340 7162 3392
rect 8386 3340 8392 3392
rect 8444 3380 8450 3392
rect 12820 3380 12848 3556
rect 17494 3544 17500 3556
rect 17552 3584 17558 3596
rect 17589 3587 17647 3593
rect 17589 3584 17601 3587
rect 17552 3556 17601 3584
rect 17552 3544 17558 3556
rect 17589 3553 17601 3556
rect 17635 3553 17647 3587
rect 17589 3547 17647 3553
rect 15933 3519 15991 3525
rect 15933 3485 15945 3519
rect 15979 3516 15991 3519
rect 16393 3519 16451 3525
rect 16393 3516 16405 3519
rect 15979 3488 16405 3516
rect 15979 3485 15991 3488
rect 15933 3479 15991 3485
rect 16393 3485 16405 3488
rect 16439 3485 16451 3519
rect 16393 3479 16451 3485
rect 16482 3476 16488 3528
rect 16540 3516 16546 3528
rect 16577 3519 16635 3525
rect 16577 3516 16589 3519
rect 16540 3488 16589 3516
rect 16540 3476 16546 3488
rect 16577 3485 16589 3488
rect 16623 3485 16635 3519
rect 16577 3479 16635 3485
rect 16669 3519 16727 3525
rect 16669 3485 16681 3519
rect 16715 3485 16727 3519
rect 17402 3516 17408 3528
rect 17363 3488 17408 3516
rect 16669 3479 16727 3485
rect 12986 3408 12992 3460
rect 13044 3448 13050 3460
rect 16684 3448 16712 3479
rect 17402 3476 17408 3488
rect 17460 3476 17466 3528
rect 13044 3420 16712 3448
rect 13044 3408 13050 3420
rect 15746 3380 15752 3392
rect 8444 3352 12848 3380
rect 15707 3352 15752 3380
rect 8444 3340 8450 3352
rect 15746 3340 15752 3352
rect 15804 3340 15810 3392
rect 17034 3340 17040 3392
rect 17092 3380 17098 3392
rect 17221 3383 17279 3389
rect 17221 3380 17233 3383
rect 17092 3352 17233 3380
rect 17092 3340 17098 3352
rect 17221 3349 17233 3352
rect 17267 3349 17279 3383
rect 17221 3343 17279 3349
rect 1104 3290 19019 3312
rect 1104 3281 5388 3290
rect 1104 3247 1133 3281
rect 1167 3247 1225 3281
rect 1259 3247 1317 3281
rect 1351 3247 1409 3281
rect 1443 3247 1501 3281
rect 1535 3247 1593 3281
rect 1627 3247 1685 3281
rect 1719 3247 1777 3281
rect 1811 3247 1869 3281
rect 1903 3247 1961 3281
rect 1995 3247 2053 3281
rect 2087 3247 2145 3281
rect 2179 3247 2237 3281
rect 2271 3247 2329 3281
rect 2363 3247 2421 3281
rect 2455 3247 2513 3281
rect 2547 3247 2605 3281
rect 2639 3247 2697 3281
rect 2731 3247 2789 3281
rect 2823 3247 2881 3281
rect 2915 3247 2973 3281
rect 3007 3247 3065 3281
rect 3099 3247 3157 3281
rect 3191 3247 3249 3281
rect 3283 3247 3341 3281
rect 3375 3247 3433 3281
rect 3467 3247 3525 3281
rect 3559 3247 3617 3281
rect 3651 3247 3709 3281
rect 3743 3247 3801 3281
rect 3835 3247 3893 3281
rect 3927 3247 3985 3281
rect 4019 3247 4077 3281
rect 4111 3247 4169 3281
rect 4203 3247 4261 3281
rect 4295 3247 4353 3281
rect 4387 3247 4445 3281
rect 4479 3247 4537 3281
rect 4571 3247 4629 3281
rect 4663 3247 4721 3281
rect 4755 3247 4813 3281
rect 4847 3247 4905 3281
rect 4939 3247 4997 3281
rect 5031 3247 5089 3281
rect 5123 3247 5181 3281
rect 5215 3247 5273 3281
rect 5307 3247 5365 3281
rect 1104 3238 5388 3247
rect 5440 3238 5452 3290
rect 5504 3238 5516 3290
rect 5568 3281 5580 3290
rect 5632 3281 5644 3290
rect 5696 3281 9827 3290
rect 9879 3281 9891 3290
rect 5632 3247 5641 3281
rect 5696 3247 5733 3281
rect 5767 3247 5825 3281
rect 5859 3247 5917 3281
rect 5951 3247 6009 3281
rect 6043 3247 6101 3281
rect 6135 3247 6193 3281
rect 6227 3247 6285 3281
rect 6319 3247 6377 3281
rect 6411 3247 6469 3281
rect 6503 3247 6561 3281
rect 6595 3247 6653 3281
rect 6687 3247 6745 3281
rect 6779 3247 6837 3281
rect 6871 3247 6929 3281
rect 6963 3247 7021 3281
rect 7055 3247 7113 3281
rect 7147 3247 7205 3281
rect 7239 3247 7297 3281
rect 7331 3247 7389 3281
rect 7423 3247 7481 3281
rect 7515 3247 7573 3281
rect 7607 3247 7665 3281
rect 7699 3247 7757 3281
rect 7791 3247 7849 3281
rect 7883 3247 7941 3281
rect 7975 3247 8033 3281
rect 8067 3247 8125 3281
rect 8159 3247 8217 3281
rect 8251 3247 8309 3281
rect 8343 3247 8401 3281
rect 8435 3247 8493 3281
rect 8527 3247 8585 3281
rect 8619 3247 8677 3281
rect 8711 3247 8769 3281
rect 8803 3247 8861 3281
rect 8895 3247 8953 3281
rect 8987 3247 9045 3281
rect 9079 3247 9137 3281
rect 9171 3247 9229 3281
rect 9263 3247 9321 3281
rect 9355 3247 9413 3281
rect 9447 3247 9505 3281
rect 9539 3247 9597 3281
rect 9631 3247 9689 3281
rect 9723 3247 9781 3281
rect 9815 3247 9827 3281
rect 5568 3238 5580 3247
rect 5632 3238 5644 3247
rect 5696 3238 9827 3247
rect 9879 3238 9891 3247
rect 9943 3238 9955 3290
rect 10007 3238 10019 3290
rect 10071 3281 10083 3290
rect 10135 3281 14266 3290
rect 14318 3281 14330 3290
rect 14382 3281 14394 3290
rect 10135 3247 10149 3281
rect 10183 3247 10241 3281
rect 10275 3247 10333 3281
rect 10367 3247 10425 3281
rect 10459 3247 10517 3281
rect 10551 3247 10609 3281
rect 10643 3247 10701 3281
rect 10735 3247 10793 3281
rect 10827 3247 10885 3281
rect 10919 3247 10977 3281
rect 11011 3247 11069 3281
rect 11103 3247 11161 3281
rect 11195 3247 11253 3281
rect 11287 3247 11345 3281
rect 11379 3247 11437 3281
rect 11471 3247 11529 3281
rect 11563 3247 11621 3281
rect 11655 3247 11713 3281
rect 11747 3247 11805 3281
rect 11839 3247 11897 3281
rect 11931 3247 11989 3281
rect 12023 3247 12081 3281
rect 12115 3247 12173 3281
rect 12207 3247 12265 3281
rect 12299 3247 12357 3281
rect 12391 3247 12449 3281
rect 12483 3247 12541 3281
rect 12575 3247 12633 3281
rect 12667 3247 12725 3281
rect 12759 3247 12817 3281
rect 12851 3247 12909 3281
rect 12943 3247 13001 3281
rect 13035 3247 13093 3281
rect 13127 3247 13185 3281
rect 13219 3247 13277 3281
rect 13311 3247 13369 3281
rect 13403 3247 13461 3281
rect 13495 3247 13553 3281
rect 13587 3247 13645 3281
rect 13679 3247 13737 3281
rect 13771 3247 13829 3281
rect 13863 3247 13921 3281
rect 13955 3247 14013 3281
rect 14047 3247 14105 3281
rect 14139 3247 14197 3281
rect 14231 3247 14266 3281
rect 14323 3247 14330 3281
rect 10071 3238 10083 3247
rect 10135 3238 14266 3247
rect 14318 3238 14330 3247
rect 14382 3238 14394 3247
rect 14446 3238 14458 3290
rect 14510 3238 14522 3290
rect 14574 3281 18705 3290
rect 14599 3247 14657 3281
rect 14691 3247 14749 3281
rect 14783 3247 14841 3281
rect 14875 3247 14933 3281
rect 14967 3247 15025 3281
rect 15059 3247 15117 3281
rect 15151 3247 15209 3281
rect 15243 3247 15301 3281
rect 15335 3247 15393 3281
rect 15427 3247 15485 3281
rect 15519 3247 15577 3281
rect 15611 3247 15669 3281
rect 15703 3247 15761 3281
rect 15795 3247 15853 3281
rect 15887 3247 15945 3281
rect 15979 3247 16037 3281
rect 16071 3247 16129 3281
rect 16163 3247 16221 3281
rect 16255 3247 16313 3281
rect 16347 3247 16405 3281
rect 16439 3247 16497 3281
rect 16531 3247 16589 3281
rect 16623 3247 16681 3281
rect 16715 3247 16773 3281
rect 16807 3247 16865 3281
rect 16899 3247 16957 3281
rect 16991 3247 17049 3281
rect 17083 3247 17141 3281
rect 17175 3247 17233 3281
rect 17267 3247 17325 3281
rect 17359 3247 17417 3281
rect 17451 3247 17509 3281
rect 17543 3247 17601 3281
rect 17635 3247 17693 3281
rect 17727 3247 17785 3281
rect 17819 3247 17877 3281
rect 17911 3247 17969 3281
rect 18003 3247 18061 3281
rect 18095 3247 18153 3281
rect 18187 3247 18245 3281
rect 18279 3247 18337 3281
rect 18371 3247 18429 3281
rect 18463 3247 18521 3281
rect 18555 3247 18613 3281
rect 18647 3247 18705 3281
rect 14574 3238 18705 3247
rect 18757 3238 18769 3290
rect 18821 3281 18833 3290
rect 18831 3247 18833 3281
rect 18821 3238 18833 3247
rect 18885 3238 18897 3290
rect 18949 3238 18961 3290
rect 19013 3238 19019 3290
rect 1104 3216 19019 3238
rect 2038 3136 2044 3188
rect 2096 3176 2102 3188
rect 3053 3179 3111 3185
rect 3053 3176 3065 3179
rect 2096 3148 3065 3176
rect 2096 3136 2102 3148
rect 3053 3145 3065 3148
rect 3099 3176 3111 3179
rect 3970 3176 3976 3188
rect 3099 3148 3976 3176
rect 3099 3145 3111 3148
rect 3053 3139 3111 3145
rect 3970 3136 3976 3148
rect 4028 3136 4034 3188
rect 9033 3179 9091 3185
rect 9033 3145 9045 3179
rect 9079 3145 9091 3179
rect 9033 3139 9091 3145
rect 2130 3108 2136 3120
rect 2091 3080 2136 3108
rect 2130 3068 2136 3080
rect 2188 3068 2194 3120
rect 4341 3111 4399 3117
rect 4341 3077 4353 3111
rect 4387 3108 4399 3111
rect 7374 3108 7380 3120
rect 4387 3080 7380 3108
rect 4387 3077 4399 3080
rect 4341 3071 4399 3077
rect 7374 3068 7380 3080
rect 7432 3108 7438 3120
rect 9048 3108 9076 3139
rect 9858 3136 9864 3188
rect 9916 3176 9922 3188
rect 10962 3176 10968 3188
rect 9916 3148 10968 3176
rect 9916 3136 9922 3148
rect 10962 3136 10968 3148
rect 11020 3176 11026 3188
rect 13081 3179 13139 3185
rect 11020 3148 12940 3176
rect 11020 3136 11026 3148
rect 7432 3080 9076 3108
rect 7432 3068 7438 3080
rect 11514 3068 11520 3120
rect 11572 3108 11578 3120
rect 11946 3111 12004 3117
rect 11946 3108 11958 3111
rect 11572 3080 11958 3108
rect 11572 3068 11578 3080
rect 11946 3077 11958 3080
rect 11992 3077 12004 3111
rect 12912 3108 12940 3148
rect 13081 3145 13093 3179
rect 13127 3176 13139 3179
rect 13262 3176 13268 3188
rect 13127 3148 13268 3176
rect 13127 3145 13139 3148
rect 13081 3139 13139 3145
rect 13262 3136 13268 3148
rect 13320 3136 13326 3188
rect 14826 3108 14832 3120
rect 12912 3080 14832 3108
rect 11946 3071 12004 3077
rect 14826 3068 14832 3080
rect 14884 3068 14890 3120
rect 1949 3043 2007 3049
rect 1949 3009 1961 3043
rect 1995 3040 2007 3043
rect 2498 3040 2504 3052
rect 1995 3012 2504 3040
rect 1995 3009 2007 3012
rect 1949 3003 2007 3009
rect 2498 3000 2504 3012
rect 2556 3000 2562 3052
rect 7285 3043 7343 3049
rect 7285 3009 7297 3043
rect 7331 3040 7343 3043
rect 7466 3040 7472 3052
rect 7331 3012 7472 3040
rect 7331 3009 7343 3012
rect 7285 3003 7343 3009
rect 7466 3000 7472 3012
rect 7524 3040 7530 3052
rect 7745 3043 7803 3049
rect 7745 3040 7757 3043
rect 7524 3012 7757 3040
rect 7524 3000 7530 3012
rect 7745 3009 7757 3012
rect 7791 3009 7803 3043
rect 7745 3003 7803 3009
rect 11701 3043 11759 3049
rect 11701 3009 11713 3043
rect 11747 3040 11759 3043
rect 11790 3040 11796 3052
rect 11747 3012 11796 3040
rect 11747 3009 11759 3012
rect 11701 3003 11759 3009
rect 11790 3000 11796 3012
rect 11848 3000 11854 3052
rect 17034 3040 17040 3052
rect 16995 3012 17040 3040
rect 17034 3000 17040 3012
rect 17092 3000 17098 3052
rect 11877 2975 11935 2981
rect 11877 2941 11889 2975
rect 11923 2972 11935 2975
rect 12115 2975 12173 2981
rect 12115 2972 12127 2975
rect 11923 2944 12127 2972
rect 11923 2941 11935 2944
rect 11877 2935 11935 2941
rect 12115 2941 12127 2944
rect 12161 2972 12173 2975
rect 12619 2975 12677 2981
rect 12619 2972 12631 2975
rect 12161 2944 12631 2972
rect 12161 2941 12173 2944
rect 12115 2935 12173 2941
rect 12619 2941 12631 2944
rect 12665 2941 12677 2975
rect 12619 2935 12677 2941
rect 11798 2907 11856 2913
rect 11798 2873 11810 2907
rect 11844 2904 11856 2907
rect 12218 2907 12276 2913
rect 12218 2904 12230 2907
rect 11844 2876 12230 2904
rect 11844 2873 11856 2876
rect 11798 2867 11856 2873
rect 12218 2873 12230 2876
rect 12264 2904 12276 2907
rect 12532 2907 12590 2913
rect 12532 2904 12544 2907
rect 12264 2876 12544 2904
rect 12264 2873 12276 2876
rect 12218 2867 12276 2873
rect 12532 2873 12544 2876
rect 12578 2873 12590 2907
rect 14274 2904 14280 2916
rect 12532 2867 12590 2873
rect 12636 2876 14280 2904
rect 12434 2796 12440 2848
rect 12492 2836 12498 2848
rect 12636 2836 12664 2876
rect 14274 2864 14280 2876
rect 14332 2864 14338 2916
rect 12492 2808 12664 2836
rect 12492 2796 12498 2808
rect 14734 2796 14740 2848
rect 14792 2836 14798 2848
rect 16853 2839 16911 2845
rect 16853 2836 16865 2839
rect 14792 2808 16865 2836
rect 14792 2796 14798 2808
rect 16853 2805 16865 2808
rect 16899 2805 16911 2839
rect 16853 2799 16911 2805
rect 1104 2746 18860 2768
rect 1104 2737 3169 2746
rect 1104 2703 1133 2737
rect 1167 2703 1225 2737
rect 1259 2703 1317 2737
rect 1351 2703 1409 2737
rect 1443 2703 1501 2737
rect 1535 2703 1593 2737
rect 1627 2703 1685 2737
rect 1719 2703 1777 2737
rect 1811 2703 1869 2737
rect 1903 2703 1961 2737
rect 1995 2703 2053 2737
rect 2087 2703 2145 2737
rect 2179 2703 2237 2737
rect 2271 2703 2329 2737
rect 2363 2703 2421 2737
rect 2455 2703 2513 2737
rect 2547 2703 2605 2737
rect 2639 2703 2697 2737
rect 2731 2703 2789 2737
rect 2823 2703 2881 2737
rect 2915 2703 2973 2737
rect 3007 2703 3065 2737
rect 3099 2703 3157 2737
rect 1104 2694 3169 2703
rect 3221 2694 3233 2746
rect 3285 2694 3297 2746
rect 3349 2737 3361 2746
rect 3349 2694 3361 2703
rect 3413 2694 3425 2746
rect 3477 2737 7608 2746
rect 3477 2703 3525 2737
rect 3559 2703 3617 2737
rect 3651 2703 3709 2737
rect 3743 2703 3801 2737
rect 3835 2703 3893 2737
rect 3927 2703 3985 2737
rect 4019 2703 4077 2737
rect 4111 2703 4169 2737
rect 4203 2703 4261 2737
rect 4295 2703 4353 2737
rect 4387 2703 4445 2737
rect 4479 2703 4537 2737
rect 4571 2703 4629 2737
rect 4663 2703 4721 2737
rect 4755 2703 4813 2737
rect 4847 2703 4905 2737
rect 4939 2703 4997 2737
rect 5031 2703 5089 2737
rect 5123 2703 5181 2737
rect 5215 2703 5273 2737
rect 5307 2703 5365 2737
rect 5399 2703 5457 2737
rect 5491 2703 5549 2737
rect 5583 2703 5641 2737
rect 5675 2703 5733 2737
rect 5767 2703 5825 2737
rect 5859 2703 5917 2737
rect 5951 2703 6009 2737
rect 6043 2703 6101 2737
rect 6135 2703 6193 2737
rect 6227 2703 6285 2737
rect 6319 2703 6377 2737
rect 6411 2703 6469 2737
rect 6503 2703 6561 2737
rect 6595 2703 6653 2737
rect 6687 2703 6745 2737
rect 6779 2703 6837 2737
rect 6871 2703 6929 2737
rect 6963 2703 7021 2737
rect 7055 2703 7113 2737
rect 7147 2703 7205 2737
rect 7239 2703 7297 2737
rect 7331 2703 7389 2737
rect 7423 2703 7481 2737
rect 7515 2703 7573 2737
rect 7607 2703 7608 2737
rect 3477 2694 7608 2703
rect 7660 2737 7672 2746
rect 7660 2703 7665 2737
rect 7660 2694 7672 2703
rect 7724 2694 7736 2746
rect 7788 2737 7800 2746
rect 7852 2737 7864 2746
rect 7916 2737 12047 2746
rect 12099 2737 12111 2746
rect 12163 2737 12175 2746
rect 7791 2703 7800 2737
rect 7916 2703 7941 2737
rect 7975 2703 8033 2737
rect 8067 2703 8125 2737
rect 8159 2703 8217 2737
rect 8251 2703 8309 2737
rect 8343 2703 8401 2737
rect 8435 2703 8493 2737
rect 8527 2703 8585 2737
rect 8619 2703 8677 2737
rect 8711 2703 8769 2737
rect 8803 2703 8861 2737
rect 8895 2703 8953 2737
rect 8987 2703 9045 2737
rect 9079 2703 9137 2737
rect 9171 2703 9229 2737
rect 9263 2703 9321 2737
rect 9355 2703 9413 2737
rect 9447 2703 9505 2737
rect 9539 2703 9597 2737
rect 9631 2703 9689 2737
rect 9723 2703 9781 2737
rect 9815 2703 9873 2737
rect 9907 2703 9965 2737
rect 9999 2703 10057 2737
rect 10091 2703 10149 2737
rect 10183 2703 10241 2737
rect 10275 2703 10333 2737
rect 10367 2703 10425 2737
rect 10459 2703 10517 2737
rect 10551 2703 10609 2737
rect 10643 2703 10701 2737
rect 10735 2703 10793 2737
rect 10827 2703 10885 2737
rect 10919 2703 10977 2737
rect 11011 2703 11069 2737
rect 11103 2703 11161 2737
rect 11195 2703 11253 2737
rect 11287 2703 11345 2737
rect 11379 2703 11437 2737
rect 11471 2703 11529 2737
rect 11563 2703 11621 2737
rect 11655 2703 11713 2737
rect 11747 2703 11805 2737
rect 11839 2703 11897 2737
rect 11931 2703 11989 2737
rect 12023 2703 12047 2737
rect 12163 2703 12173 2737
rect 7788 2694 7800 2703
rect 7852 2694 7864 2703
rect 7916 2694 12047 2703
rect 12099 2694 12111 2703
rect 12163 2694 12175 2703
rect 12227 2694 12239 2746
rect 12291 2737 12303 2746
rect 12299 2703 12303 2737
rect 12291 2694 12303 2703
rect 12355 2737 16486 2746
rect 12355 2703 12357 2737
rect 12391 2703 12449 2737
rect 12483 2703 12541 2737
rect 12575 2703 12633 2737
rect 12667 2703 12725 2737
rect 12759 2703 12817 2737
rect 12851 2703 12909 2737
rect 12943 2703 13001 2737
rect 13035 2703 13093 2737
rect 13127 2703 13185 2737
rect 13219 2703 13277 2737
rect 13311 2703 13369 2737
rect 13403 2703 13461 2737
rect 13495 2703 13553 2737
rect 13587 2703 13645 2737
rect 13679 2703 13737 2737
rect 13771 2703 13829 2737
rect 13863 2703 13921 2737
rect 13955 2703 14013 2737
rect 14047 2703 14105 2737
rect 14139 2703 14197 2737
rect 14231 2703 14289 2737
rect 14323 2703 14381 2737
rect 14415 2703 14473 2737
rect 14507 2703 14565 2737
rect 14599 2703 14657 2737
rect 14691 2703 14749 2737
rect 14783 2703 14841 2737
rect 14875 2703 14933 2737
rect 14967 2703 15025 2737
rect 15059 2703 15117 2737
rect 15151 2703 15209 2737
rect 15243 2703 15301 2737
rect 15335 2703 15393 2737
rect 15427 2703 15485 2737
rect 15519 2703 15577 2737
rect 15611 2703 15669 2737
rect 15703 2703 15761 2737
rect 15795 2703 15853 2737
rect 15887 2703 15945 2737
rect 15979 2703 16037 2737
rect 16071 2703 16129 2737
rect 16163 2703 16221 2737
rect 16255 2703 16313 2737
rect 16347 2703 16405 2737
rect 16439 2703 16486 2737
rect 12355 2694 16486 2703
rect 16538 2694 16550 2746
rect 16602 2737 16614 2746
rect 16602 2694 16614 2703
rect 16666 2694 16678 2746
rect 16730 2694 16742 2746
rect 16794 2737 18860 2746
rect 16807 2703 16865 2737
rect 16899 2703 16957 2737
rect 16991 2703 17049 2737
rect 17083 2703 17141 2737
rect 17175 2703 17233 2737
rect 17267 2703 17325 2737
rect 17359 2703 17417 2737
rect 17451 2703 17509 2737
rect 17543 2703 17601 2737
rect 17635 2703 17693 2737
rect 17727 2703 17785 2737
rect 17819 2703 17877 2737
rect 17911 2703 17969 2737
rect 18003 2703 18061 2737
rect 18095 2703 18153 2737
rect 18187 2703 18245 2737
rect 18279 2703 18337 2737
rect 18371 2703 18429 2737
rect 18463 2703 18521 2737
rect 18555 2703 18613 2737
rect 18647 2703 18705 2737
rect 18739 2703 18797 2737
rect 18831 2703 18860 2737
rect 16794 2694 18860 2703
rect 1104 2672 18860 2694
rect 1854 2592 1860 2644
rect 1912 2632 1918 2644
rect 2041 2635 2099 2641
rect 2041 2632 2053 2635
rect 1912 2604 2053 2632
rect 1912 2592 1918 2604
rect 2041 2601 2053 2604
rect 2087 2632 2099 2635
rect 5997 2635 6055 2641
rect 2087 2604 5948 2632
rect 2087 2601 2099 2604
rect 2041 2595 2099 2601
rect 2590 2567 2648 2573
rect 2590 2533 2602 2567
rect 2636 2564 2648 2567
rect 2904 2567 2962 2573
rect 2904 2564 2916 2567
rect 2636 2536 2916 2564
rect 2636 2533 2648 2536
rect 2590 2527 2648 2533
rect 2904 2533 2916 2536
rect 2950 2564 2962 2567
rect 3324 2567 3382 2573
rect 3324 2564 3336 2567
rect 2950 2536 3336 2564
rect 2950 2533 2962 2536
rect 2904 2527 2962 2533
rect 3324 2533 3336 2536
rect 3370 2533 3382 2567
rect 3324 2527 3382 2533
rect 4714 2567 4772 2573
rect 4714 2533 4726 2567
rect 4760 2564 4772 2567
rect 5134 2567 5192 2573
rect 5134 2564 5146 2567
rect 4760 2536 5146 2564
rect 4760 2533 4772 2536
rect 4714 2527 4772 2533
rect 5134 2533 5146 2536
rect 5180 2564 5192 2567
rect 5448 2567 5506 2573
rect 5448 2564 5460 2567
rect 5180 2536 5460 2564
rect 5180 2533 5192 2536
rect 5134 2527 5192 2533
rect 5448 2533 5460 2536
rect 5494 2533 5506 2567
rect 5920 2564 5948 2604
rect 5997 2601 6009 2635
rect 6043 2632 6055 2635
rect 6546 2632 6552 2644
rect 6043 2604 6552 2632
rect 6043 2601 6055 2604
rect 5997 2595 6055 2601
rect 6546 2592 6552 2604
rect 6604 2592 6610 2644
rect 9674 2632 9680 2644
rect 6886 2604 9680 2632
rect 6886 2564 6914 2604
rect 9674 2592 9680 2604
rect 9732 2592 9738 2644
rect 10042 2592 10048 2644
rect 10100 2632 10106 2644
rect 11606 2632 11612 2644
rect 10100 2604 11612 2632
rect 10100 2592 10106 2604
rect 11606 2592 11612 2604
rect 11664 2592 11670 2644
rect 11882 2632 11888 2644
rect 11843 2604 11888 2632
rect 11882 2592 11888 2604
rect 11940 2592 11946 2644
rect 12986 2632 12992 2644
rect 12360 2604 12992 2632
rect 5920 2536 6914 2564
rect 7742 2567 7800 2573
rect 5448 2527 5506 2533
rect 7742 2533 7754 2567
rect 7788 2564 7800 2567
rect 8056 2567 8114 2573
rect 8056 2564 8068 2567
rect 7788 2536 8068 2564
rect 7788 2533 7800 2536
rect 7742 2527 7800 2533
rect 8056 2533 8068 2536
rect 8102 2564 8114 2567
rect 8476 2567 8534 2573
rect 8476 2564 8488 2567
rect 8102 2536 8488 2564
rect 8102 2533 8114 2536
rect 8056 2527 8114 2533
rect 8476 2533 8488 2536
rect 8522 2533 8534 2567
rect 8476 2527 8534 2533
rect 9866 2567 9924 2573
rect 9866 2533 9878 2567
rect 9912 2564 9924 2567
rect 10286 2567 10344 2573
rect 10286 2564 10298 2567
rect 9912 2536 10298 2564
rect 9912 2533 9924 2536
rect 9866 2527 9924 2533
rect 10286 2533 10298 2536
rect 10332 2564 10344 2567
rect 10600 2567 10658 2573
rect 10600 2564 10612 2567
rect 10332 2536 10612 2564
rect 10332 2533 10344 2536
rect 10286 2527 10344 2533
rect 10600 2533 10612 2536
rect 10646 2533 10658 2567
rect 10600 2527 10658 2533
rect 11149 2567 11207 2573
rect 11149 2533 11161 2567
rect 11195 2564 11207 2567
rect 12360 2564 12388 2604
rect 12986 2592 12992 2604
rect 13044 2592 13050 2644
rect 14274 2632 14280 2644
rect 14235 2604 14280 2632
rect 14274 2592 14280 2604
rect 14332 2592 14338 2644
rect 16850 2632 16856 2644
rect 16811 2604 16856 2632
rect 16850 2592 16856 2604
rect 16908 2592 16914 2644
rect 11195 2536 12388 2564
rect 12434 2567 12492 2573
rect 11195 2533 11207 2536
rect 11149 2527 11207 2533
rect 12434 2533 12446 2567
rect 12480 2564 12492 2567
rect 12748 2567 12806 2573
rect 12748 2564 12760 2567
rect 12480 2536 12760 2564
rect 12480 2533 12492 2536
rect 12434 2527 12492 2533
rect 12748 2533 12760 2536
rect 12794 2564 12806 2567
rect 13168 2567 13226 2573
rect 13168 2564 13180 2567
rect 12794 2536 13180 2564
rect 12794 2533 12806 2536
rect 12748 2527 12806 2533
rect 13168 2533 13180 2536
rect 13214 2533 13226 2567
rect 13168 2527 13226 2533
rect 2503 2499 2561 2505
rect 2503 2465 2515 2499
rect 2549 2496 2561 2499
rect 3007 2499 3065 2505
rect 3007 2496 3019 2499
rect 2549 2468 3019 2496
rect 2549 2465 2561 2468
rect 2503 2459 2561 2465
rect 3007 2465 3019 2468
rect 3053 2496 3065 2499
rect 3245 2499 3303 2505
rect 3245 2496 3257 2499
rect 3053 2468 3257 2496
rect 3053 2465 3065 2468
rect 3007 2459 3065 2465
rect 3245 2465 3257 2468
rect 3291 2465 3303 2499
rect 3245 2459 3303 2465
rect 3421 2499 3479 2505
rect 3421 2465 3433 2499
rect 3467 2496 3479 2499
rect 3970 2496 3976 2508
rect 3467 2468 3976 2496
rect 3467 2465 3479 2468
rect 3421 2459 3479 2465
rect 3970 2456 3976 2468
rect 4028 2496 4034 2508
rect 4617 2499 4675 2505
rect 4617 2496 4629 2499
rect 4028 2468 4629 2496
rect 4028 2456 4034 2468
rect 4617 2465 4629 2468
rect 4663 2465 4675 2499
rect 4617 2459 4675 2465
rect 4793 2499 4851 2505
rect 4793 2465 4805 2499
rect 4839 2496 4851 2499
rect 5031 2499 5089 2505
rect 5031 2496 5043 2499
rect 4839 2468 5043 2496
rect 4839 2465 4851 2468
rect 4793 2459 4851 2465
rect 5031 2465 5043 2468
rect 5077 2496 5089 2499
rect 5535 2499 5593 2505
rect 5535 2496 5547 2499
rect 5077 2468 5547 2496
rect 5077 2465 5089 2468
rect 5031 2459 5089 2465
rect 5535 2465 5547 2468
rect 5581 2465 5593 2499
rect 5535 2459 5593 2465
rect 7655 2499 7713 2505
rect 7655 2465 7667 2499
rect 7701 2496 7713 2499
rect 8159 2499 8217 2505
rect 8159 2496 8171 2499
rect 7701 2468 8171 2496
rect 7701 2465 7713 2468
rect 7655 2459 7713 2465
rect 8159 2465 8171 2468
rect 8205 2496 8217 2499
rect 8397 2499 8455 2505
rect 8397 2496 8409 2499
rect 8205 2468 8409 2496
rect 8205 2465 8217 2468
rect 8159 2459 8217 2465
rect 8397 2465 8409 2468
rect 8443 2465 8455 2499
rect 8397 2459 8455 2465
rect 9945 2499 10003 2505
rect 9945 2465 9957 2499
rect 9991 2496 10003 2499
rect 10183 2499 10241 2505
rect 10183 2496 10195 2499
rect 9991 2468 10195 2496
rect 9991 2465 10003 2468
rect 9945 2459 10003 2465
rect 10183 2465 10195 2468
rect 10229 2496 10241 2499
rect 10687 2499 10745 2505
rect 10687 2496 10699 2499
rect 10229 2468 10699 2496
rect 10229 2465 10241 2468
rect 10183 2459 10241 2465
rect 10687 2465 10699 2468
rect 10733 2465 10745 2499
rect 10687 2459 10745 2465
rect 12347 2499 12405 2505
rect 12347 2465 12359 2499
rect 12393 2496 12405 2499
rect 12851 2499 12909 2505
rect 12851 2496 12863 2499
rect 12393 2468 12863 2496
rect 12393 2465 12405 2468
rect 12347 2459 12405 2465
rect 12851 2465 12863 2468
rect 12897 2496 12909 2499
rect 13089 2499 13147 2505
rect 13089 2496 13101 2499
rect 12897 2468 13101 2496
rect 12897 2465 12909 2468
rect 12851 2459 12909 2465
rect 13089 2465 13101 2468
rect 13135 2465 13147 2499
rect 13089 2459 13147 2465
rect 3165 2431 3223 2437
rect 3165 2397 3177 2431
rect 3211 2428 3223 2431
rect 6914 2428 6920 2440
rect 3211 2400 6920 2428
rect 3211 2397 3223 2400
rect 3165 2391 3223 2397
rect 6914 2388 6920 2400
rect 6972 2388 6978 2440
rect 8573 2431 8631 2437
rect 8573 2397 8585 2431
rect 8619 2428 8631 2431
rect 9769 2431 9827 2437
rect 9769 2428 9781 2431
rect 8619 2400 9781 2428
rect 8619 2397 8631 2400
rect 8573 2391 8631 2397
rect 9769 2397 9781 2400
rect 9815 2428 9827 2431
rect 11698 2428 11704 2440
rect 9815 2400 11704 2428
rect 9815 2397 9827 2400
rect 9769 2391 9827 2397
rect 11698 2388 11704 2400
rect 11756 2428 11762 2440
rect 13265 2431 13323 2437
rect 13265 2428 13277 2431
rect 11756 2400 13277 2428
rect 11756 2388 11762 2400
rect 13265 2397 13277 2400
rect 13311 2397 13323 2431
rect 13265 2391 13323 2397
rect 17037 2431 17095 2437
rect 17037 2397 17049 2431
rect 17083 2428 17095 2431
rect 17218 2428 17224 2440
rect 17083 2400 17224 2428
rect 17083 2397 17095 2400
rect 17037 2391 17095 2397
rect 17218 2388 17224 2400
rect 17276 2388 17282 2440
rect 17494 2428 17500 2440
rect 17455 2400 17500 2428
rect 17494 2388 17500 2400
rect 17552 2388 17558 2440
rect 4522 2320 4528 2372
rect 4580 2360 4586 2372
rect 10042 2369 10048 2372
rect 4862 2363 4920 2369
rect 4862 2360 4874 2363
rect 4580 2332 4874 2360
rect 4580 2320 4586 2332
rect 4862 2329 4874 2332
rect 4908 2329 4920 2363
rect 4862 2323 4920 2329
rect 8328 2363 8386 2369
rect 8328 2329 8340 2363
rect 8374 2360 8386 2363
rect 8374 2332 9996 2360
rect 8374 2329 8386 2332
rect 8328 2323 8386 2329
rect 2498 2252 2504 2304
rect 2556 2292 2562 2304
rect 3973 2295 4031 2301
rect 3973 2292 3985 2295
rect 2556 2264 3985 2292
rect 2556 2252 2562 2264
rect 3973 2261 3985 2264
rect 4019 2261 4031 2295
rect 3973 2255 4031 2261
rect 7193 2295 7251 2301
rect 7193 2261 7205 2295
rect 7239 2292 7251 2295
rect 9858 2292 9864 2304
rect 7239 2264 9864 2292
rect 7239 2261 7251 2264
rect 7193 2255 7251 2261
rect 9858 2252 9864 2264
rect 9916 2252 9922 2304
rect 9968 2292 9996 2332
rect 10036 2323 10048 2369
rect 10100 2360 10106 2372
rect 13020 2363 13078 2369
rect 10100 2332 10136 2360
rect 10042 2320 10048 2323
rect 10100 2320 10106 2332
rect 13020 2329 13032 2363
rect 13066 2360 13078 2363
rect 14734 2360 14740 2372
rect 13066 2332 14740 2360
rect 13066 2329 13078 2332
rect 13020 2323 13078 2329
rect 14734 2320 14740 2332
rect 14792 2320 14798 2372
rect 15746 2292 15752 2304
rect 9968 2264 15752 2292
rect 15746 2252 15752 2264
rect 15804 2252 15810 2304
rect 17402 2252 17408 2304
rect 17460 2292 17466 2304
rect 17681 2295 17739 2301
rect 17681 2292 17693 2295
rect 17460 2264 17693 2292
rect 17460 2252 17466 2264
rect 17681 2261 17693 2264
rect 17727 2261 17739 2295
rect 17681 2255 17739 2261
rect 1104 2202 19019 2224
rect 1104 2193 5388 2202
rect 1104 2159 1133 2193
rect 1167 2159 1225 2193
rect 1259 2159 1317 2193
rect 1351 2159 1409 2193
rect 1443 2159 1501 2193
rect 1535 2159 1593 2193
rect 1627 2159 1685 2193
rect 1719 2159 1777 2193
rect 1811 2159 1869 2193
rect 1903 2159 1961 2193
rect 1995 2159 2053 2193
rect 2087 2159 2145 2193
rect 2179 2159 2237 2193
rect 2271 2159 2329 2193
rect 2363 2159 2421 2193
rect 2455 2159 2513 2193
rect 2547 2159 2605 2193
rect 2639 2159 2697 2193
rect 2731 2159 2789 2193
rect 2823 2159 2881 2193
rect 2915 2159 2973 2193
rect 3007 2159 3065 2193
rect 3099 2159 3157 2193
rect 3191 2159 3249 2193
rect 3283 2159 3341 2193
rect 3375 2159 3433 2193
rect 3467 2159 3525 2193
rect 3559 2159 3617 2193
rect 3651 2159 3709 2193
rect 3743 2159 3801 2193
rect 3835 2159 3893 2193
rect 3927 2159 3985 2193
rect 4019 2159 4077 2193
rect 4111 2159 4169 2193
rect 4203 2159 4261 2193
rect 4295 2159 4353 2193
rect 4387 2159 4445 2193
rect 4479 2159 4537 2193
rect 4571 2159 4629 2193
rect 4663 2159 4721 2193
rect 4755 2159 4813 2193
rect 4847 2159 4905 2193
rect 4939 2159 4997 2193
rect 5031 2159 5089 2193
rect 5123 2159 5181 2193
rect 5215 2159 5273 2193
rect 5307 2159 5365 2193
rect 1104 2150 5388 2159
rect 5440 2150 5452 2202
rect 5504 2150 5516 2202
rect 5568 2193 5580 2202
rect 5632 2193 5644 2202
rect 5696 2193 9827 2202
rect 9879 2193 9891 2202
rect 5632 2159 5641 2193
rect 5696 2159 5733 2193
rect 5767 2159 5825 2193
rect 5859 2159 5917 2193
rect 5951 2159 6009 2193
rect 6043 2159 6101 2193
rect 6135 2159 6193 2193
rect 6227 2159 6285 2193
rect 6319 2159 6377 2193
rect 6411 2159 6469 2193
rect 6503 2159 6561 2193
rect 6595 2159 6653 2193
rect 6687 2159 6745 2193
rect 6779 2159 6837 2193
rect 6871 2159 6929 2193
rect 6963 2159 7021 2193
rect 7055 2159 7113 2193
rect 7147 2159 7205 2193
rect 7239 2159 7297 2193
rect 7331 2159 7389 2193
rect 7423 2159 7481 2193
rect 7515 2159 7573 2193
rect 7607 2159 7665 2193
rect 7699 2159 7757 2193
rect 7791 2159 7849 2193
rect 7883 2159 7941 2193
rect 7975 2159 8033 2193
rect 8067 2159 8125 2193
rect 8159 2159 8217 2193
rect 8251 2159 8309 2193
rect 8343 2159 8401 2193
rect 8435 2159 8493 2193
rect 8527 2159 8585 2193
rect 8619 2159 8677 2193
rect 8711 2159 8769 2193
rect 8803 2159 8861 2193
rect 8895 2159 8953 2193
rect 8987 2159 9045 2193
rect 9079 2159 9137 2193
rect 9171 2159 9229 2193
rect 9263 2159 9321 2193
rect 9355 2159 9413 2193
rect 9447 2159 9505 2193
rect 9539 2159 9597 2193
rect 9631 2159 9689 2193
rect 9723 2159 9781 2193
rect 9815 2159 9827 2193
rect 5568 2150 5580 2159
rect 5632 2150 5644 2159
rect 5696 2150 9827 2159
rect 9879 2150 9891 2159
rect 9943 2150 9955 2202
rect 10007 2150 10019 2202
rect 10071 2193 10083 2202
rect 10135 2193 14266 2202
rect 14318 2193 14330 2202
rect 14382 2193 14394 2202
rect 10135 2159 10149 2193
rect 10183 2159 10241 2193
rect 10275 2159 10333 2193
rect 10367 2159 10425 2193
rect 10459 2159 10517 2193
rect 10551 2159 10609 2193
rect 10643 2159 10701 2193
rect 10735 2159 10793 2193
rect 10827 2159 10885 2193
rect 10919 2159 10977 2193
rect 11011 2159 11069 2193
rect 11103 2159 11161 2193
rect 11195 2159 11253 2193
rect 11287 2159 11345 2193
rect 11379 2159 11437 2193
rect 11471 2159 11529 2193
rect 11563 2159 11621 2193
rect 11655 2159 11713 2193
rect 11747 2159 11805 2193
rect 11839 2159 11897 2193
rect 11931 2159 11989 2193
rect 12023 2159 12081 2193
rect 12115 2159 12173 2193
rect 12207 2159 12265 2193
rect 12299 2159 12357 2193
rect 12391 2159 12449 2193
rect 12483 2159 12541 2193
rect 12575 2159 12633 2193
rect 12667 2159 12725 2193
rect 12759 2159 12817 2193
rect 12851 2159 12909 2193
rect 12943 2159 13001 2193
rect 13035 2159 13093 2193
rect 13127 2159 13185 2193
rect 13219 2159 13277 2193
rect 13311 2159 13369 2193
rect 13403 2159 13461 2193
rect 13495 2159 13553 2193
rect 13587 2159 13645 2193
rect 13679 2159 13737 2193
rect 13771 2159 13829 2193
rect 13863 2159 13921 2193
rect 13955 2159 14013 2193
rect 14047 2159 14105 2193
rect 14139 2159 14197 2193
rect 14231 2159 14266 2193
rect 14323 2159 14330 2193
rect 10071 2150 10083 2159
rect 10135 2150 14266 2159
rect 14318 2150 14330 2159
rect 14382 2150 14394 2159
rect 14446 2150 14458 2202
rect 14510 2150 14522 2202
rect 14574 2193 18705 2202
rect 14599 2159 14657 2193
rect 14691 2159 14749 2193
rect 14783 2159 14841 2193
rect 14875 2159 14933 2193
rect 14967 2159 15025 2193
rect 15059 2159 15117 2193
rect 15151 2159 15209 2193
rect 15243 2159 15301 2193
rect 15335 2159 15393 2193
rect 15427 2159 15485 2193
rect 15519 2159 15577 2193
rect 15611 2159 15669 2193
rect 15703 2159 15761 2193
rect 15795 2159 15853 2193
rect 15887 2159 15945 2193
rect 15979 2159 16037 2193
rect 16071 2159 16129 2193
rect 16163 2159 16221 2193
rect 16255 2159 16313 2193
rect 16347 2159 16405 2193
rect 16439 2159 16497 2193
rect 16531 2159 16589 2193
rect 16623 2159 16681 2193
rect 16715 2159 16773 2193
rect 16807 2159 16865 2193
rect 16899 2159 16957 2193
rect 16991 2159 17049 2193
rect 17083 2159 17141 2193
rect 17175 2159 17233 2193
rect 17267 2159 17325 2193
rect 17359 2159 17417 2193
rect 17451 2159 17509 2193
rect 17543 2159 17601 2193
rect 17635 2159 17693 2193
rect 17727 2159 17785 2193
rect 17819 2159 17877 2193
rect 17911 2159 17969 2193
rect 18003 2159 18061 2193
rect 18095 2159 18153 2193
rect 18187 2159 18245 2193
rect 18279 2159 18337 2193
rect 18371 2159 18429 2193
rect 18463 2159 18521 2193
rect 18555 2159 18613 2193
rect 18647 2159 18705 2193
rect 14574 2150 18705 2159
rect 18757 2150 18769 2202
rect 18821 2193 18833 2202
rect 18831 2159 18833 2193
rect 18821 2150 18833 2159
rect 18885 2150 18897 2202
rect 18949 2150 18961 2202
rect 19013 2150 19019 2202
rect 1104 2128 19019 2150
<< via1 >>
rect 5388 7633 5440 7642
rect 5388 7599 5399 7633
rect 5399 7599 5440 7633
rect 5388 7590 5440 7599
rect 5452 7633 5504 7642
rect 5452 7599 5457 7633
rect 5457 7599 5491 7633
rect 5491 7599 5504 7633
rect 5452 7590 5504 7599
rect 5516 7633 5568 7642
rect 5580 7633 5632 7642
rect 5644 7633 5696 7642
rect 9827 7633 9879 7642
rect 9891 7633 9943 7642
rect 5516 7599 5549 7633
rect 5549 7599 5568 7633
rect 5580 7599 5583 7633
rect 5583 7599 5632 7633
rect 5644 7599 5675 7633
rect 5675 7599 5696 7633
rect 9827 7599 9873 7633
rect 9873 7599 9879 7633
rect 9891 7599 9907 7633
rect 9907 7599 9943 7633
rect 5516 7590 5568 7599
rect 5580 7590 5632 7599
rect 5644 7590 5696 7599
rect 9827 7590 9879 7599
rect 9891 7590 9943 7599
rect 9955 7633 10007 7642
rect 9955 7599 9965 7633
rect 9965 7599 9999 7633
rect 9999 7599 10007 7633
rect 9955 7590 10007 7599
rect 10019 7633 10071 7642
rect 10083 7633 10135 7642
rect 14266 7633 14318 7642
rect 14330 7633 14382 7642
rect 14394 7633 14446 7642
rect 10019 7599 10057 7633
rect 10057 7599 10071 7633
rect 10083 7599 10091 7633
rect 10091 7599 10135 7633
rect 14266 7599 14289 7633
rect 14289 7599 14318 7633
rect 14330 7599 14381 7633
rect 14381 7599 14382 7633
rect 14394 7599 14415 7633
rect 14415 7599 14446 7633
rect 10019 7590 10071 7599
rect 10083 7590 10135 7599
rect 14266 7590 14318 7599
rect 14330 7590 14382 7599
rect 14394 7590 14446 7599
rect 14458 7633 14510 7642
rect 14458 7599 14473 7633
rect 14473 7599 14507 7633
rect 14507 7599 14510 7633
rect 14458 7590 14510 7599
rect 14522 7633 14574 7642
rect 18705 7633 18757 7642
rect 14522 7599 14565 7633
rect 14565 7599 14574 7633
rect 18705 7599 18739 7633
rect 18739 7599 18757 7633
rect 14522 7590 14574 7599
rect 18705 7590 18757 7599
rect 18769 7633 18821 7642
rect 18769 7599 18797 7633
rect 18797 7599 18821 7633
rect 18769 7590 18821 7599
rect 18833 7590 18885 7642
rect 18897 7590 18949 7642
rect 18961 7590 19013 7642
rect 1124 7488 1176 7540
rect 3332 7488 3384 7540
rect 5724 7531 5776 7540
rect 5724 7497 5733 7531
rect 5733 7497 5767 7531
rect 5767 7497 5776 7531
rect 5724 7488 5776 7497
rect 7748 7488 7800 7540
rect 12440 7531 12492 7540
rect 12440 7497 12449 7531
rect 12449 7497 12483 7531
rect 12483 7497 12492 7531
rect 12440 7488 12492 7497
rect 14648 7531 14700 7540
rect 14648 7497 14657 7531
rect 14657 7497 14691 7531
rect 14691 7497 14700 7531
rect 14648 7488 14700 7497
rect 16580 7488 16632 7540
rect 18420 7488 18472 7540
rect 10232 7420 10284 7472
rect 1860 7395 1912 7404
rect 1860 7361 1869 7395
rect 1869 7361 1903 7395
rect 1903 7361 1912 7395
rect 1860 7352 1912 7361
rect 4620 7352 4672 7404
rect 6920 7352 6972 7404
rect 7104 7352 7156 7404
rect 10600 7352 10652 7404
rect 12532 7352 12584 7404
rect 14648 7352 14700 7404
rect 13452 7284 13504 7336
rect 10324 7259 10376 7268
rect 10324 7225 10333 7259
rect 10333 7225 10367 7259
rect 10367 7225 10376 7259
rect 10324 7216 10376 7225
rect 3169 7089 3221 7098
rect 3169 7055 3191 7089
rect 3191 7055 3221 7089
rect 3169 7046 3221 7055
rect 3233 7089 3285 7098
rect 3233 7055 3249 7089
rect 3249 7055 3283 7089
rect 3283 7055 3285 7089
rect 3233 7046 3285 7055
rect 3297 7089 3349 7098
rect 3361 7089 3413 7098
rect 3297 7055 3341 7089
rect 3341 7055 3349 7089
rect 3361 7055 3375 7089
rect 3375 7055 3413 7089
rect 3297 7046 3349 7055
rect 3361 7046 3413 7055
rect 3425 7089 3477 7098
rect 3425 7055 3433 7089
rect 3433 7055 3467 7089
rect 3467 7055 3477 7089
rect 3425 7046 3477 7055
rect 7608 7046 7660 7098
rect 7672 7089 7724 7098
rect 7672 7055 7699 7089
rect 7699 7055 7724 7089
rect 7672 7046 7724 7055
rect 7736 7089 7788 7098
rect 7800 7089 7852 7098
rect 7864 7089 7916 7098
rect 12047 7089 12099 7098
rect 12111 7089 12163 7098
rect 12175 7089 12227 7098
rect 7736 7055 7757 7089
rect 7757 7055 7788 7089
rect 7800 7055 7849 7089
rect 7849 7055 7852 7089
rect 7864 7055 7883 7089
rect 7883 7055 7916 7089
rect 12047 7055 12081 7089
rect 12081 7055 12099 7089
rect 12111 7055 12115 7089
rect 12115 7055 12163 7089
rect 12175 7055 12207 7089
rect 12207 7055 12227 7089
rect 7736 7046 7788 7055
rect 7800 7046 7852 7055
rect 7864 7046 7916 7055
rect 12047 7046 12099 7055
rect 12111 7046 12163 7055
rect 12175 7046 12227 7055
rect 12239 7089 12291 7098
rect 12239 7055 12265 7089
rect 12265 7055 12291 7089
rect 12239 7046 12291 7055
rect 12303 7046 12355 7098
rect 16486 7089 16538 7098
rect 16486 7055 16497 7089
rect 16497 7055 16531 7089
rect 16531 7055 16538 7089
rect 16486 7046 16538 7055
rect 16550 7089 16602 7098
rect 16614 7089 16666 7098
rect 16550 7055 16589 7089
rect 16589 7055 16602 7089
rect 16614 7055 16623 7089
rect 16623 7055 16666 7089
rect 16550 7046 16602 7055
rect 16614 7046 16666 7055
rect 16678 7089 16730 7098
rect 16678 7055 16681 7089
rect 16681 7055 16715 7089
rect 16715 7055 16730 7089
rect 16678 7046 16730 7055
rect 16742 7089 16794 7098
rect 16742 7055 16773 7089
rect 16773 7055 16794 7089
rect 16742 7046 16794 7055
rect 5388 6545 5440 6554
rect 5388 6511 5399 6545
rect 5399 6511 5440 6545
rect 5388 6502 5440 6511
rect 5452 6545 5504 6554
rect 5452 6511 5457 6545
rect 5457 6511 5491 6545
rect 5491 6511 5504 6545
rect 5452 6502 5504 6511
rect 5516 6545 5568 6554
rect 5580 6545 5632 6554
rect 5644 6545 5696 6554
rect 9827 6545 9879 6554
rect 9891 6545 9943 6554
rect 5516 6511 5549 6545
rect 5549 6511 5568 6545
rect 5580 6511 5583 6545
rect 5583 6511 5632 6545
rect 5644 6511 5675 6545
rect 5675 6511 5696 6545
rect 9827 6511 9873 6545
rect 9873 6511 9879 6545
rect 9891 6511 9907 6545
rect 9907 6511 9943 6545
rect 5516 6502 5568 6511
rect 5580 6502 5632 6511
rect 5644 6502 5696 6511
rect 9827 6502 9879 6511
rect 9891 6502 9943 6511
rect 9955 6545 10007 6554
rect 9955 6511 9965 6545
rect 9965 6511 9999 6545
rect 9999 6511 10007 6545
rect 9955 6502 10007 6511
rect 10019 6545 10071 6554
rect 10083 6545 10135 6554
rect 14266 6545 14318 6554
rect 14330 6545 14382 6554
rect 14394 6545 14446 6554
rect 10019 6511 10057 6545
rect 10057 6511 10071 6545
rect 10083 6511 10091 6545
rect 10091 6511 10135 6545
rect 14266 6511 14289 6545
rect 14289 6511 14318 6545
rect 14330 6511 14381 6545
rect 14381 6511 14382 6545
rect 14394 6511 14415 6545
rect 14415 6511 14446 6545
rect 10019 6502 10071 6511
rect 10083 6502 10135 6511
rect 14266 6502 14318 6511
rect 14330 6502 14382 6511
rect 14394 6502 14446 6511
rect 14458 6545 14510 6554
rect 14458 6511 14473 6545
rect 14473 6511 14507 6545
rect 14507 6511 14510 6545
rect 14458 6502 14510 6511
rect 14522 6545 14574 6554
rect 18705 6545 18757 6554
rect 14522 6511 14565 6545
rect 14565 6511 14574 6545
rect 18705 6511 18739 6545
rect 18739 6511 18757 6545
rect 14522 6502 14574 6511
rect 18705 6502 18757 6511
rect 18769 6545 18821 6554
rect 18769 6511 18797 6545
rect 18797 6511 18821 6545
rect 18769 6502 18821 6511
rect 18833 6502 18885 6554
rect 18897 6502 18949 6554
rect 18961 6502 19013 6554
rect 3169 6001 3221 6010
rect 3169 5967 3191 6001
rect 3191 5967 3221 6001
rect 3169 5958 3221 5967
rect 3233 6001 3285 6010
rect 3233 5967 3249 6001
rect 3249 5967 3283 6001
rect 3283 5967 3285 6001
rect 3233 5958 3285 5967
rect 3297 6001 3349 6010
rect 3361 6001 3413 6010
rect 3297 5967 3341 6001
rect 3341 5967 3349 6001
rect 3361 5967 3375 6001
rect 3375 5967 3413 6001
rect 3297 5958 3349 5967
rect 3361 5958 3413 5967
rect 3425 6001 3477 6010
rect 3425 5967 3433 6001
rect 3433 5967 3467 6001
rect 3467 5967 3477 6001
rect 3425 5958 3477 5967
rect 7608 5958 7660 6010
rect 7672 6001 7724 6010
rect 7672 5967 7699 6001
rect 7699 5967 7724 6001
rect 7672 5958 7724 5967
rect 7736 6001 7788 6010
rect 7800 6001 7852 6010
rect 7864 6001 7916 6010
rect 12047 6001 12099 6010
rect 12111 6001 12163 6010
rect 12175 6001 12227 6010
rect 7736 5967 7757 6001
rect 7757 5967 7788 6001
rect 7800 5967 7849 6001
rect 7849 5967 7852 6001
rect 7864 5967 7883 6001
rect 7883 5967 7916 6001
rect 12047 5967 12081 6001
rect 12081 5967 12099 6001
rect 12111 5967 12115 6001
rect 12115 5967 12163 6001
rect 12175 5967 12207 6001
rect 12207 5967 12227 6001
rect 7736 5958 7788 5967
rect 7800 5958 7852 5967
rect 7864 5958 7916 5967
rect 12047 5958 12099 5967
rect 12111 5958 12163 5967
rect 12175 5958 12227 5967
rect 12239 6001 12291 6010
rect 12239 5967 12265 6001
rect 12265 5967 12291 6001
rect 12239 5958 12291 5967
rect 12303 5958 12355 6010
rect 16486 6001 16538 6010
rect 16486 5967 16497 6001
rect 16497 5967 16531 6001
rect 16531 5967 16538 6001
rect 16486 5958 16538 5967
rect 16550 6001 16602 6010
rect 16614 6001 16666 6010
rect 16550 5967 16589 6001
rect 16589 5967 16602 6001
rect 16614 5967 16623 6001
rect 16623 5967 16666 6001
rect 16550 5958 16602 5967
rect 16614 5958 16666 5967
rect 16678 6001 16730 6010
rect 16678 5967 16681 6001
rect 16681 5967 16715 6001
rect 16715 5967 16730 6001
rect 16678 5958 16730 5967
rect 16742 6001 16794 6010
rect 16742 5967 16773 6001
rect 16773 5967 16794 6001
rect 16742 5958 16794 5967
rect 7012 5788 7064 5840
rect 10876 5788 10928 5840
rect 5908 5720 5960 5772
rect 6828 5720 6880 5772
rect 2872 5652 2924 5704
rect 3976 5652 4028 5704
rect 5724 5652 5776 5704
rect 10508 5720 10560 5772
rect 14832 5763 14884 5772
rect 14832 5729 14841 5763
rect 14841 5729 14875 5763
rect 14875 5729 14884 5763
rect 14832 5720 14884 5729
rect 10232 5695 10284 5704
rect 10232 5661 10241 5695
rect 10241 5661 10275 5695
rect 10275 5661 10284 5695
rect 10232 5652 10284 5661
rect 10600 5652 10652 5704
rect 11244 5695 11296 5704
rect 11244 5661 11253 5695
rect 11253 5661 11287 5695
rect 11287 5661 11296 5695
rect 11244 5652 11296 5661
rect 7196 5627 7248 5636
rect 7196 5593 7205 5627
rect 7205 5593 7239 5627
rect 7239 5593 7248 5627
rect 7196 5584 7248 5593
rect 8300 5584 8352 5636
rect 10324 5627 10376 5636
rect 10324 5593 10333 5627
rect 10333 5593 10367 5627
rect 10367 5593 10376 5627
rect 10324 5584 10376 5593
rect 10968 5584 11020 5636
rect 13544 5584 13596 5636
rect 3056 5559 3108 5568
rect 3056 5525 3065 5559
rect 3065 5525 3099 5559
rect 3099 5525 3108 5559
rect 3056 5516 3108 5525
rect 6000 5516 6052 5568
rect 7104 5559 7156 5568
rect 7104 5525 7113 5559
rect 7113 5525 7147 5559
rect 7147 5525 7156 5559
rect 7104 5516 7156 5525
rect 9680 5516 9732 5568
rect 11060 5559 11112 5568
rect 11060 5525 11069 5559
rect 11069 5525 11103 5559
rect 11103 5525 11112 5559
rect 11060 5516 11112 5525
rect 12532 5516 12584 5568
rect 13820 5516 13872 5568
rect 14648 5559 14700 5568
rect 14648 5525 14657 5559
rect 14657 5525 14691 5559
rect 14691 5525 14700 5559
rect 14648 5516 14700 5525
rect 5388 5457 5440 5466
rect 5388 5423 5399 5457
rect 5399 5423 5440 5457
rect 5388 5414 5440 5423
rect 5452 5457 5504 5466
rect 5452 5423 5457 5457
rect 5457 5423 5491 5457
rect 5491 5423 5504 5457
rect 5452 5414 5504 5423
rect 5516 5457 5568 5466
rect 5580 5457 5632 5466
rect 5644 5457 5696 5466
rect 9827 5457 9879 5466
rect 9891 5457 9943 5466
rect 5516 5423 5549 5457
rect 5549 5423 5568 5457
rect 5580 5423 5583 5457
rect 5583 5423 5632 5457
rect 5644 5423 5675 5457
rect 5675 5423 5696 5457
rect 9827 5423 9873 5457
rect 9873 5423 9879 5457
rect 9891 5423 9907 5457
rect 9907 5423 9943 5457
rect 5516 5414 5568 5423
rect 5580 5414 5632 5423
rect 5644 5414 5696 5423
rect 9827 5414 9879 5423
rect 9891 5414 9943 5423
rect 9955 5457 10007 5466
rect 9955 5423 9965 5457
rect 9965 5423 9999 5457
rect 9999 5423 10007 5457
rect 9955 5414 10007 5423
rect 10019 5457 10071 5466
rect 10083 5457 10135 5466
rect 14266 5457 14318 5466
rect 14330 5457 14382 5466
rect 14394 5457 14446 5466
rect 10019 5423 10057 5457
rect 10057 5423 10071 5457
rect 10083 5423 10091 5457
rect 10091 5423 10135 5457
rect 14266 5423 14289 5457
rect 14289 5423 14318 5457
rect 14330 5423 14381 5457
rect 14381 5423 14382 5457
rect 14394 5423 14415 5457
rect 14415 5423 14446 5457
rect 10019 5414 10071 5423
rect 10083 5414 10135 5423
rect 14266 5414 14318 5423
rect 14330 5414 14382 5423
rect 14394 5414 14446 5423
rect 14458 5457 14510 5466
rect 14458 5423 14473 5457
rect 14473 5423 14507 5457
rect 14507 5423 14510 5457
rect 14458 5414 14510 5423
rect 14522 5457 14574 5466
rect 18705 5457 18757 5466
rect 14522 5423 14565 5457
rect 14565 5423 14574 5457
rect 18705 5423 18739 5457
rect 18739 5423 18757 5457
rect 14522 5414 14574 5423
rect 18705 5414 18757 5423
rect 18769 5457 18821 5466
rect 18769 5423 18797 5457
rect 18797 5423 18821 5457
rect 18769 5414 18821 5423
rect 18833 5414 18885 5466
rect 18897 5414 18949 5466
rect 18961 5414 19013 5466
rect 2872 5355 2924 5364
rect 2872 5321 2881 5355
rect 2881 5321 2915 5355
rect 2915 5321 2924 5355
rect 2872 5312 2924 5321
rect 3884 5355 3936 5364
rect 3884 5321 3893 5355
rect 3893 5321 3927 5355
rect 3927 5321 3936 5355
rect 3884 5312 3936 5321
rect 7196 5312 7248 5364
rect 8300 5355 8352 5364
rect 8300 5321 8309 5355
rect 8309 5321 8343 5355
rect 8343 5321 8352 5355
rect 8300 5312 8352 5321
rect 10968 5312 11020 5364
rect 13452 5355 13504 5364
rect 13452 5321 13461 5355
rect 13461 5321 13495 5355
rect 13495 5321 13504 5355
rect 13452 5312 13504 5321
rect 13544 5355 13596 5364
rect 13544 5321 13553 5355
rect 13553 5321 13587 5355
rect 13587 5321 13596 5355
rect 13544 5312 13596 5321
rect 2136 5219 2188 5228
rect 2136 5185 2145 5219
rect 2145 5185 2179 5219
rect 2179 5185 2188 5219
rect 5908 5244 5960 5296
rect 6920 5244 6972 5296
rect 2136 5176 2188 5185
rect 3700 5219 3752 5228
rect 3700 5185 3709 5219
rect 3709 5185 3743 5219
rect 3743 5185 3752 5219
rect 3700 5176 3752 5185
rect 3884 5176 3936 5228
rect 5080 5176 5132 5228
rect 11060 5244 11112 5296
rect 4620 5108 4672 5160
rect 2596 5040 2648 5092
rect 5724 5040 5776 5092
rect 9312 5219 9364 5228
rect 9312 5185 9321 5219
rect 9321 5185 9355 5219
rect 9355 5185 9364 5219
rect 9312 5176 9364 5185
rect 9680 5176 9732 5228
rect 9772 5176 9824 5228
rect 7288 5151 7340 5160
rect 7288 5117 7297 5151
rect 7297 5117 7331 5151
rect 7331 5117 7340 5151
rect 8392 5151 8444 5160
rect 7288 5108 7340 5117
rect 8392 5117 8401 5151
rect 8401 5117 8435 5151
rect 8435 5117 8444 5151
rect 8392 5108 8444 5117
rect 9956 5108 10008 5160
rect 10508 5108 10560 5160
rect 11888 5108 11940 5160
rect 12992 5108 13044 5160
rect 11244 5040 11296 5092
rect 14556 5040 14608 5092
rect 1952 5015 2004 5024
rect 1952 4981 1961 5015
rect 1961 4981 1995 5015
rect 1995 4981 2004 5015
rect 1952 4972 2004 4981
rect 4712 4972 4764 5024
rect 4804 4972 4856 5024
rect 6644 5015 6696 5024
rect 6644 4981 6653 5015
rect 6653 4981 6687 5015
rect 6687 4981 6696 5015
rect 6644 4972 6696 4981
rect 6736 4972 6788 5024
rect 9128 5015 9180 5024
rect 9128 4981 9137 5015
rect 9137 4981 9171 5015
rect 9171 4981 9180 5015
rect 9128 4972 9180 4981
rect 9220 4972 9272 5024
rect 13084 5015 13136 5024
rect 13084 4981 13093 5015
rect 13093 4981 13127 5015
rect 13127 4981 13136 5015
rect 13084 4972 13136 4981
rect 3169 4913 3221 4922
rect 3169 4879 3191 4913
rect 3191 4879 3221 4913
rect 3169 4870 3221 4879
rect 3233 4913 3285 4922
rect 3233 4879 3249 4913
rect 3249 4879 3283 4913
rect 3283 4879 3285 4913
rect 3233 4870 3285 4879
rect 3297 4913 3349 4922
rect 3361 4913 3413 4922
rect 3297 4879 3341 4913
rect 3341 4879 3349 4913
rect 3361 4879 3375 4913
rect 3375 4879 3413 4913
rect 3297 4870 3349 4879
rect 3361 4870 3413 4879
rect 3425 4913 3477 4922
rect 3425 4879 3433 4913
rect 3433 4879 3467 4913
rect 3467 4879 3477 4913
rect 3425 4870 3477 4879
rect 7608 4870 7660 4922
rect 7672 4913 7724 4922
rect 7672 4879 7699 4913
rect 7699 4879 7724 4913
rect 7672 4870 7724 4879
rect 7736 4913 7788 4922
rect 7800 4913 7852 4922
rect 7864 4913 7916 4922
rect 12047 4913 12099 4922
rect 12111 4913 12163 4922
rect 12175 4913 12227 4922
rect 7736 4879 7757 4913
rect 7757 4879 7788 4913
rect 7800 4879 7849 4913
rect 7849 4879 7852 4913
rect 7864 4879 7883 4913
rect 7883 4879 7916 4913
rect 12047 4879 12081 4913
rect 12081 4879 12099 4913
rect 12111 4879 12115 4913
rect 12115 4879 12163 4913
rect 12175 4879 12207 4913
rect 12207 4879 12227 4913
rect 7736 4870 7788 4879
rect 7800 4870 7852 4879
rect 7864 4870 7916 4879
rect 12047 4870 12099 4879
rect 12111 4870 12163 4879
rect 12175 4870 12227 4879
rect 12239 4913 12291 4922
rect 12239 4879 12265 4913
rect 12265 4879 12291 4913
rect 12239 4870 12291 4879
rect 12303 4870 12355 4922
rect 16486 4913 16538 4922
rect 16486 4879 16497 4913
rect 16497 4879 16531 4913
rect 16531 4879 16538 4913
rect 16486 4870 16538 4879
rect 16550 4913 16602 4922
rect 16614 4913 16666 4922
rect 16550 4879 16589 4913
rect 16589 4879 16602 4913
rect 16614 4879 16623 4913
rect 16623 4879 16666 4913
rect 16550 4870 16602 4879
rect 16614 4870 16666 4879
rect 16678 4913 16730 4922
rect 16678 4879 16681 4913
rect 16681 4879 16715 4913
rect 16715 4879 16730 4913
rect 16678 4870 16730 4879
rect 16742 4913 16794 4922
rect 16742 4879 16773 4913
rect 16773 4879 16794 4913
rect 16742 4870 16794 4879
rect 3976 4811 4028 4820
rect 3976 4777 3985 4811
rect 3985 4777 4019 4811
rect 4019 4777 4028 4811
rect 3976 4768 4028 4777
rect 6000 4768 6052 4820
rect 6552 4768 6604 4820
rect 9956 4811 10008 4820
rect 3700 4700 3752 4752
rect 2044 4607 2096 4616
rect 2044 4573 2053 4607
rect 2053 4573 2087 4607
rect 2087 4573 2096 4607
rect 2044 4564 2096 4573
rect 3056 4564 3108 4616
rect 9956 4777 9965 4811
rect 9965 4777 9999 4811
rect 9999 4777 10008 4811
rect 9956 4768 10008 4777
rect 11152 4768 11204 4820
rect 13084 4768 13136 4820
rect 4344 4675 4396 4684
rect 4344 4641 4353 4675
rect 4353 4641 4387 4675
rect 4387 4641 4396 4675
rect 4344 4632 4396 4641
rect 5724 4632 5776 4684
rect 6276 4675 6328 4684
rect 6276 4641 6285 4675
rect 6285 4641 6319 4675
rect 6319 4641 6328 4675
rect 6276 4632 6328 4641
rect 12624 4700 12676 4752
rect 17408 4700 17460 4752
rect 5080 4607 5132 4616
rect 5080 4573 5089 4607
rect 5089 4573 5123 4607
rect 5123 4573 5132 4607
rect 5080 4564 5132 4573
rect 6092 4564 6144 4616
rect 6736 4607 6788 4616
rect 6736 4573 6745 4607
rect 6745 4573 6779 4607
rect 6779 4573 6788 4607
rect 6736 4564 6788 4573
rect 7012 4607 7064 4616
rect 7012 4573 7046 4607
rect 7046 4573 7064 4607
rect 11336 4607 11388 4616
rect 7012 4564 7064 4573
rect 11336 4573 11345 4607
rect 11345 4573 11379 4607
rect 11379 4573 11388 4607
rect 11336 4564 11388 4573
rect 11428 4564 11480 4616
rect 13820 4632 13872 4684
rect 6552 4496 6604 4548
rect 11704 4496 11756 4548
rect 12992 4564 13044 4616
rect 13268 4564 13320 4616
rect 14556 4607 14608 4616
rect 14556 4573 14565 4607
rect 14565 4573 14599 4607
rect 14599 4573 14608 4607
rect 14556 4564 14608 4573
rect 14740 4564 14792 4616
rect 12624 4496 12676 4548
rect 4252 4428 4304 4480
rect 5724 4428 5776 4480
rect 7288 4428 7340 4480
rect 11980 4428 12032 4480
rect 12440 4428 12492 4480
rect 15660 4428 15712 4480
rect 5388 4369 5440 4378
rect 5388 4335 5399 4369
rect 5399 4335 5440 4369
rect 5388 4326 5440 4335
rect 5452 4369 5504 4378
rect 5452 4335 5457 4369
rect 5457 4335 5491 4369
rect 5491 4335 5504 4369
rect 5452 4326 5504 4335
rect 5516 4369 5568 4378
rect 5580 4369 5632 4378
rect 5644 4369 5696 4378
rect 9827 4369 9879 4378
rect 9891 4369 9943 4378
rect 5516 4335 5549 4369
rect 5549 4335 5568 4369
rect 5580 4335 5583 4369
rect 5583 4335 5632 4369
rect 5644 4335 5675 4369
rect 5675 4335 5696 4369
rect 9827 4335 9873 4369
rect 9873 4335 9879 4369
rect 9891 4335 9907 4369
rect 9907 4335 9943 4369
rect 5516 4326 5568 4335
rect 5580 4326 5632 4335
rect 5644 4326 5696 4335
rect 9827 4326 9879 4335
rect 9891 4326 9943 4335
rect 9955 4369 10007 4378
rect 9955 4335 9965 4369
rect 9965 4335 9999 4369
rect 9999 4335 10007 4369
rect 9955 4326 10007 4335
rect 10019 4369 10071 4378
rect 10083 4369 10135 4378
rect 14266 4369 14318 4378
rect 14330 4369 14382 4378
rect 14394 4369 14446 4378
rect 10019 4335 10057 4369
rect 10057 4335 10071 4369
rect 10083 4335 10091 4369
rect 10091 4335 10135 4369
rect 14266 4335 14289 4369
rect 14289 4335 14318 4369
rect 14330 4335 14381 4369
rect 14381 4335 14382 4369
rect 14394 4335 14415 4369
rect 14415 4335 14446 4369
rect 10019 4326 10071 4335
rect 10083 4326 10135 4335
rect 14266 4326 14318 4335
rect 14330 4326 14382 4335
rect 14394 4326 14446 4335
rect 14458 4369 14510 4378
rect 14458 4335 14473 4369
rect 14473 4335 14507 4369
rect 14507 4335 14510 4369
rect 14458 4326 14510 4335
rect 14522 4369 14574 4378
rect 18705 4369 18757 4378
rect 14522 4335 14565 4369
rect 14565 4335 14574 4369
rect 18705 4335 18739 4369
rect 18739 4335 18757 4369
rect 14522 4326 14574 4335
rect 18705 4326 18757 4335
rect 18769 4369 18821 4378
rect 18769 4335 18797 4369
rect 18797 4335 18821 4369
rect 18769 4326 18821 4335
rect 18833 4326 18885 4378
rect 18897 4326 18949 4378
rect 18961 4326 19013 4378
rect 2596 4267 2648 4276
rect 2596 4233 2605 4267
rect 2605 4233 2639 4267
rect 2639 4233 2648 4267
rect 2596 4224 2648 4233
rect 4620 4267 4672 4276
rect 4620 4233 4629 4267
rect 4629 4233 4663 4267
rect 4663 4233 4672 4267
rect 4620 4224 4672 4233
rect 4712 4224 4764 4276
rect 11520 4224 11572 4276
rect 13452 4224 13504 4276
rect 1952 4131 2004 4140
rect 1952 4097 1961 4131
rect 1961 4097 1995 4131
rect 1995 4097 2004 4131
rect 1952 4088 2004 4097
rect 4804 4156 4856 4208
rect 3976 4131 4028 4140
rect 3976 4097 3985 4131
rect 3985 4097 4019 4131
rect 4019 4097 4028 4131
rect 3976 4088 4028 4097
rect 5724 4131 5776 4140
rect 6092 4156 6144 4208
rect 5724 4097 5742 4131
rect 5742 4097 5776 4131
rect 5724 4088 5776 4097
rect 6736 4088 6788 4140
rect 7380 4156 7432 4208
rect 9312 4156 9364 4208
rect 7196 4088 7248 4140
rect 9220 4088 9272 4140
rect 11428 4156 11480 4208
rect 11980 4199 12032 4208
rect 11980 4165 12014 4199
rect 12014 4165 12032 4199
rect 11980 4156 12032 4165
rect 6460 4020 6512 4072
rect 6920 4020 6972 4072
rect 6552 3952 6604 4004
rect 8392 4020 8444 4072
rect 9588 4063 9640 4072
rect 9588 4029 9597 4063
rect 9597 4029 9631 4063
rect 9631 4029 9640 4063
rect 11336 4088 11388 4140
rect 11796 4088 11848 4140
rect 14832 4088 14884 4140
rect 15660 4131 15712 4140
rect 15660 4097 15669 4131
rect 15669 4097 15703 4131
rect 15703 4097 15712 4131
rect 15660 4088 15712 4097
rect 9588 4020 9640 4029
rect 10968 4063 11020 4072
rect 10968 4029 10977 4063
rect 10977 4029 11011 4063
rect 11011 4029 11020 4063
rect 10968 4020 11020 4029
rect 14740 4020 14792 4072
rect 10876 3995 10928 4004
rect 10876 3961 10885 3995
rect 10885 3961 10919 3995
rect 10919 3961 10928 3995
rect 10876 3952 10928 3961
rect 16396 3952 16448 4004
rect 4528 3884 4580 3936
rect 6920 3927 6972 3936
rect 6920 3893 6929 3927
rect 6929 3893 6963 3927
rect 6963 3893 6972 3927
rect 6920 3884 6972 3893
rect 10508 3927 10560 3936
rect 10508 3893 10517 3927
rect 10517 3893 10551 3927
rect 10551 3893 10560 3927
rect 10508 3884 10560 3893
rect 11612 3884 11664 3936
rect 17224 3927 17276 3936
rect 17224 3893 17233 3927
rect 17233 3893 17267 3927
rect 17267 3893 17276 3927
rect 17224 3884 17276 3893
rect 3169 3825 3221 3834
rect 3169 3791 3191 3825
rect 3191 3791 3221 3825
rect 3169 3782 3221 3791
rect 3233 3825 3285 3834
rect 3233 3791 3249 3825
rect 3249 3791 3283 3825
rect 3283 3791 3285 3825
rect 3233 3782 3285 3791
rect 3297 3825 3349 3834
rect 3361 3825 3413 3834
rect 3297 3791 3341 3825
rect 3341 3791 3349 3825
rect 3361 3791 3375 3825
rect 3375 3791 3413 3825
rect 3297 3782 3349 3791
rect 3361 3782 3413 3791
rect 3425 3825 3477 3834
rect 3425 3791 3433 3825
rect 3433 3791 3467 3825
rect 3467 3791 3477 3825
rect 3425 3782 3477 3791
rect 7608 3782 7660 3834
rect 7672 3825 7724 3834
rect 7672 3791 7699 3825
rect 7699 3791 7724 3825
rect 7672 3782 7724 3791
rect 7736 3825 7788 3834
rect 7800 3825 7852 3834
rect 7864 3825 7916 3834
rect 12047 3825 12099 3834
rect 12111 3825 12163 3834
rect 12175 3825 12227 3834
rect 7736 3791 7757 3825
rect 7757 3791 7788 3825
rect 7800 3791 7849 3825
rect 7849 3791 7852 3825
rect 7864 3791 7883 3825
rect 7883 3791 7916 3825
rect 12047 3791 12081 3825
rect 12081 3791 12099 3825
rect 12111 3791 12115 3825
rect 12115 3791 12163 3825
rect 12175 3791 12207 3825
rect 12207 3791 12227 3825
rect 7736 3782 7788 3791
rect 7800 3782 7852 3791
rect 7864 3782 7916 3791
rect 12047 3782 12099 3791
rect 12111 3782 12163 3791
rect 12175 3782 12227 3791
rect 12239 3825 12291 3834
rect 12239 3791 12265 3825
rect 12265 3791 12291 3825
rect 12239 3782 12291 3791
rect 12303 3782 12355 3834
rect 16486 3825 16538 3834
rect 16486 3791 16497 3825
rect 16497 3791 16531 3825
rect 16531 3791 16538 3825
rect 16486 3782 16538 3791
rect 16550 3825 16602 3834
rect 16614 3825 16666 3834
rect 16550 3791 16589 3825
rect 16589 3791 16602 3825
rect 16614 3791 16623 3825
rect 16623 3791 16666 3825
rect 16550 3782 16602 3791
rect 16614 3782 16666 3791
rect 16678 3825 16730 3834
rect 16678 3791 16681 3825
rect 16681 3791 16715 3825
rect 16715 3791 16730 3825
rect 16678 3782 16730 3791
rect 16742 3825 16794 3834
rect 16742 3791 16773 3825
rect 16773 3791 16794 3825
rect 16742 3782 16794 3791
rect 6460 3680 6512 3732
rect 6644 3723 6696 3732
rect 6644 3689 6653 3723
rect 6653 3689 6687 3723
rect 6687 3689 6696 3723
rect 6644 3680 6696 3689
rect 10140 3680 10192 3732
rect 12532 3680 12584 3732
rect 14648 3680 14700 3732
rect 6736 3612 6788 3664
rect 3976 3587 4028 3596
rect 3976 3553 3985 3587
rect 3985 3553 4019 3587
rect 4019 3553 4028 3587
rect 3976 3544 4028 3553
rect 9588 3544 9640 3596
rect 11796 3587 11848 3596
rect 11796 3553 11805 3587
rect 11805 3553 11839 3587
rect 11839 3553 11848 3587
rect 11796 3544 11848 3553
rect 2044 3519 2096 3528
rect 2044 3485 2053 3519
rect 2053 3485 2087 3519
rect 2087 3485 2096 3519
rect 2044 3476 2096 3485
rect 4252 3519 4304 3528
rect 4252 3485 4286 3519
rect 4286 3485 4304 3519
rect 4252 3476 4304 3485
rect 6092 3476 6144 3528
rect 6552 3476 6604 3528
rect 6828 3476 6880 3528
rect 9128 3476 9180 3528
rect 10508 3476 10560 3528
rect 12440 3476 12492 3528
rect 7104 3340 7156 3392
rect 8392 3340 8444 3392
rect 17500 3544 17552 3596
rect 16488 3476 16540 3528
rect 17408 3519 17460 3528
rect 12992 3408 13044 3460
rect 17408 3485 17417 3519
rect 17417 3485 17451 3519
rect 17451 3485 17460 3519
rect 17408 3476 17460 3485
rect 15752 3383 15804 3392
rect 15752 3349 15761 3383
rect 15761 3349 15795 3383
rect 15795 3349 15804 3383
rect 15752 3340 15804 3349
rect 17040 3340 17092 3392
rect 5388 3281 5440 3290
rect 5388 3247 5399 3281
rect 5399 3247 5440 3281
rect 5388 3238 5440 3247
rect 5452 3281 5504 3290
rect 5452 3247 5457 3281
rect 5457 3247 5491 3281
rect 5491 3247 5504 3281
rect 5452 3238 5504 3247
rect 5516 3281 5568 3290
rect 5580 3281 5632 3290
rect 5644 3281 5696 3290
rect 9827 3281 9879 3290
rect 9891 3281 9943 3290
rect 5516 3247 5549 3281
rect 5549 3247 5568 3281
rect 5580 3247 5583 3281
rect 5583 3247 5632 3281
rect 5644 3247 5675 3281
rect 5675 3247 5696 3281
rect 9827 3247 9873 3281
rect 9873 3247 9879 3281
rect 9891 3247 9907 3281
rect 9907 3247 9943 3281
rect 5516 3238 5568 3247
rect 5580 3238 5632 3247
rect 5644 3238 5696 3247
rect 9827 3238 9879 3247
rect 9891 3238 9943 3247
rect 9955 3281 10007 3290
rect 9955 3247 9965 3281
rect 9965 3247 9999 3281
rect 9999 3247 10007 3281
rect 9955 3238 10007 3247
rect 10019 3281 10071 3290
rect 10083 3281 10135 3290
rect 14266 3281 14318 3290
rect 14330 3281 14382 3290
rect 14394 3281 14446 3290
rect 10019 3247 10057 3281
rect 10057 3247 10071 3281
rect 10083 3247 10091 3281
rect 10091 3247 10135 3281
rect 14266 3247 14289 3281
rect 14289 3247 14318 3281
rect 14330 3247 14381 3281
rect 14381 3247 14382 3281
rect 14394 3247 14415 3281
rect 14415 3247 14446 3281
rect 10019 3238 10071 3247
rect 10083 3238 10135 3247
rect 14266 3238 14318 3247
rect 14330 3238 14382 3247
rect 14394 3238 14446 3247
rect 14458 3281 14510 3290
rect 14458 3247 14473 3281
rect 14473 3247 14507 3281
rect 14507 3247 14510 3281
rect 14458 3238 14510 3247
rect 14522 3281 14574 3290
rect 18705 3281 18757 3290
rect 14522 3247 14565 3281
rect 14565 3247 14574 3281
rect 18705 3247 18739 3281
rect 18739 3247 18757 3281
rect 14522 3238 14574 3247
rect 18705 3238 18757 3247
rect 18769 3281 18821 3290
rect 18769 3247 18797 3281
rect 18797 3247 18821 3281
rect 18769 3238 18821 3247
rect 18833 3238 18885 3290
rect 18897 3238 18949 3290
rect 18961 3238 19013 3290
rect 2044 3136 2096 3188
rect 3976 3136 4028 3188
rect 2136 3111 2188 3120
rect 2136 3077 2145 3111
rect 2145 3077 2179 3111
rect 2179 3077 2188 3111
rect 2136 3068 2188 3077
rect 7380 3068 7432 3120
rect 9864 3136 9916 3188
rect 10968 3136 11020 3188
rect 11520 3068 11572 3120
rect 13268 3136 13320 3188
rect 14832 3068 14884 3120
rect 2504 3000 2556 3052
rect 7472 3000 7524 3052
rect 11796 3000 11848 3052
rect 17040 3043 17092 3052
rect 17040 3009 17049 3043
rect 17049 3009 17083 3043
rect 17083 3009 17092 3043
rect 17040 3000 17092 3009
rect 12440 2796 12492 2848
rect 14280 2864 14332 2916
rect 14740 2796 14792 2848
rect 3169 2737 3221 2746
rect 3169 2703 3191 2737
rect 3191 2703 3221 2737
rect 3169 2694 3221 2703
rect 3233 2737 3285 2746
rect 3233 2703 3249 2737
rect 3249 2703 3283 2737
rect 3283 2703 3285 2737
rect 3233 2694 3285 2703
rect 3297 2737 3349 2746
rect 3361 2737 3413 2746
rect 3297 2703 3341 2737
rect 3341 2703 3349 2737
rect 3361 2703 3375 2737
rect 3375 2703 3413 2737
rect 3297 2694 3349 2703
rect 3361 2694 3413 2703
rect 3425 2737 3477 2746
rect 3425 2703 3433 2737
rect 3433 2703 3467 2737
rect 3467 2703 3477 2737
rect 3425 2694 3477 2703
rect 7608 2694 7660 2746
rect 7672 2737 7724 2746
rect 7672 2703 7699 2737
rect 7699 2703 7724 2737
rect 7672 2694 7724 2703
rect 7736 2737 7788 2746
rect 7800 2737 7852 2746
rect 7864 2737 7916 2746
rect 12047 2737 12099 2746
rect 12111 2737 12163 2746
rect 12175 2737 12227 2746
rect 7736 2703 7757 2737
rect 7757 2703 7788 2737
rect 7800 2703 7849 2737
rect 7849 2703 7852 2737
rect 7864 2703 7883 2737
rect 7883 2703 7916 2737
rect 12047 2703 12081 2737
rect 12081 2703 12099 2737
rect 12111 2703 12115 2737
rect 12115 2703 12163 2737
rect 12175 2703 12207 2737
rect 12207 2703 12227 2737
rect 7736 2694 7788 2703
rect 7800 2694 7852 2703
rect 7864 2694 7916 2703
rect 12047 2694 12099 2703
rect 12111 2694 12163 2703
rect 12175 2694 12227 2703
rect 12239 2737 12291 2746
rect 12239 2703 12265 2737
rect 12265 2703 12291 2737
rect 12239 2694 12291 2703
rect 12303 2694 12355 2746
rect 16486 2737 16538 2746
rect 16486 2703 16497 2737
rect 16497 2703 16531 2737
rect 16531 2703 16538 2737
rect 16486 2694 16538 2703
rect 16550 2737 16602 2746
rect 16614 2737 16666 2746
rect 16550 2703 16589 2737
rect 16589 2703 16602 2737
rect 16614 2703 16623 2737
rect 16623 2703 16666 2737
rect 16550 2694 16602 2703
rect 16614 2694 16666 2703
rect 16678 2737 16730 2746
rect 16678 2703 16681 2737
rect 16681 2703 16715 2737
rect 16715 2703 16730 2737
rect 16678 2694 16730 2703
rect 16742 2737 16794 2746
rect 16742 2703 16773 2737
rect 16773 2703 16794 2737
rect 16742 2694 16794 2703
rect 1860 2592 1912 2644
rect 6552 2592 6604 2644
rect 9680 2592 9732 2644
rect 10048 2592 10100 2644
rect 11612 2592 11664 2644
rect 11888 2635 11940 2644
rect 11888 2601 11897 2635
rect 11897 2601 11931 2635
rect 11931 2601 11940 2635
rect 11888 2592 11940 2601
rect 12992 2592 13044 2644
rect 14280 2635 14332 2644
rect 14280 2601 14289 2635
rect 14289 2601 14323 2635
rect 14323 2601 14332 2635
rect 14280 2592 14332 2601
rect 16856 2635 16908 2644
rect 16856 2601 16865 2635
rect 16865 2601 16899 2635
rect 16899 2601 16908 2635
rect 16856 2592 16908 2601
rect 3976 2456 4028 2508
rect 6920 2388 6972 2440
rect 11704 2388 11756 2440
rect 17224 2388 17276 2440
rect 17500 2431 17552 2440
rect 17500 2397 17509 2431
rect 17509 2397 17543 2431
rect 17543 2397 17552 2431
rect 17500 2388 17552 2397
rect 4528 2320 4580 2372
rect 2504 2252 2556 2304
rect 9864 2252 9916 2304
rect 10048 2363 10100 2372
rect 10048 2329 10082 2363
rect 10082 2329 10100 2363
rect 10048 2320 10100 2329
rect 14740 2320 14792 2372
rect 15752 2252 15804 2304
rect 17408 2252 17460 2304
rect 5388 2193 5440 2202
rect 5388 2159 5399 2193
rect 5399 2159 5440 2193
rect 5388 2150 5440 2159
rect 5452 2193 5504 2202
rect 5452 2159 5457 2193
rect 5457 2159 5491 2193
rect 5491 2159 5504 2193
rect 5452 2150 5504 2159
rect 5516 2193 5568 2202
rect 5580 2193 5632 2202
rect 5644 2193 5696 2202
rect 9827 2193 9879 2202
rect 9891 2193 9943 2202
rect 5516 2159 5549 2193
rect 5549 2159 5568 2193
rect 5580 2159 5583 2193
rect 5583 2159 5632 2193
rect 5644 2159 5675 2193
rect 5675 2159 5696 2193
rect 9827 2159 9873 2193
rect 9873 2159 9879 2193
rect 9891 2159 9907 2193
rect 9907 2159 9943 2193
rect 5516 2150 5568 2159
rect 5580 2150 5632 2159
rect 5644 2150 5696 2159
rect 9827 2150 9879 2159
rect 9891 2150 9943 2159
rect 9955 2193 10007 2202
rect 9955 2159 9965 2193
rect 9965 2159 9999 2193
rect 9999 2159 10007 2193
rect 9955 2150 10007 2159
rect 10019 2193 10071 2202
rect 10083 2193 10135 2202
rect 14266 2193 14318 2202
rect 14330 2193 14382 2202
rect 14394 2193 14446 2202
rect 10019 2159 10057 2193
rect 10057 2159 10071 2193
rect 10083 2159 10091 2193
rect 10091 2159 10135 2193
rect 14266 2159 14289 2193
rect 14289 2159 14318 2193
rect 14330 2159 14381 2193
rect 14381 2159 14382 2193
rect 14394 2159 14415 2193
rect 14415 2159 14446 2193
rect 10019 2150 10071 2159
rect 10083 2150 10135 2159
rect 14266 2150 14318 2159
rect 14330 2150 14382 2159
rect 14394 2150 14446 2159
rect 14458 2193 14510 2202
rect 14458 2159 14473 2193
rect 14473 2159 14507 2193
rect 14507 2159 14510 2193
rect 14458 2150 14510 2159
rect 14522 2193 14574 2202
rect 18705 2193 18757 2202
rect 14522 2159 14565 2193
rect 14565 2159 14574 2193
rect 18705 2159 18739 2193
rect 18739 2159 18757 2193
rect 14522 2150 14574 2159
rect 18705 2150 18757 2159
rect 18769 2193 18821 2202
rect 18769 2159 18797 2193
rect 18797 2159 18821 2193
rect 18769 2150 18821 2159
rect 18833 2150 18885 2202
rect 18897 2150 18949 2202
rect 18961 2150 19013 2202
<< metal2 >>
rect 1122 9200 1178 10000
rect 3330 9200 3386 10000
rect 5538 9330 5594 10000
rect 5538 9302 5764 9330
rect 5538 9200 5594 9302
rect 1136 7546 1164 9200
rect 3344 7546 3372 9200
rect 5388 7644 5696 7653
rect 5388 7642 5394 7644
rect 5450 7642 5474 7644
rect 5530 7642 5554 7644
rect 5610 7642 5634 7644
rect 5690 7642 5696 7644
rect 5450 7590 5452 7642
rect 5632 7590 5634 7642
rect 5388 7588 5394 7590
rect 5450 7588 5474 7590
rect 5530 7588 5554 7590
rect 5610 7588 5634 7590
rect 5690 7588 5696 7590
rect 5388 7579 5696 7588
rect 5736 7546 5764 9302
rect 7746 9200 7802 10000
rect 9954 9330 10010 10000
rect 12162 9330 12218 10000
rect 14370 9330 14426 10000
rect 9954 9302 10272 9330
rect 9954 9200 10010 9302
rect 7760 7546 7788 9200
rect 9827 7644 10135 7653
rect 9827 7642 9833 7644
rect 9889 7642 9913 7644
rect 9969 7642 9993 7644
rect 10049 7642 10073 7644
rect 10129 7642 10135 7644
rect 9889 7590 9891 7642
rect 10071 7590 10073 7642
rect 9827 7588 9833 7590
rect 9889 7588 9913 7590
rect 9969 7588 9993 7590
rect 10049 7588 10073 7590
rect 10129 7588 10135 7590
rect 9827 7579 10135 7588
rect 1124 7540 1176 7546
rect 1124 7482 1176 7488
rect 3332 7540 3384 7546
rect 3332 7482 3384 7488
rect 5724 7540 5776 7546
rect 5724 7482 5776 7488
rect 7748 7540 7800 7546
rect 7748 7482 7800 7488
rect 10244 7478 10272 9302
rect 12162 9302 12388 9330
rect 12162 9200 12218 9302
rect 12360 7528 12388 9302
rect 14370 9302 14688 9330
rect 14370 9200 14426 9302
rect 14266 7644 14574 7653
rect 14266 7642 14272 7644
rect 14328 7642 14352 7644
rect 14408 7642 14432 7644
rect 14488 7642 14512 7644
rect 14568 7642 14574 7644
rect 14328 7590 14330 7642
rect 14510 7590 14512 7642
rect 14266 7588 14272 7590
rect 14328 7588 14352 7590
rect 14408 7588 14432 7590
rect 14488 7588 14512 7590
rect 14568 7588 14574 7590
rect 14266 7579 14574 7588
rect 14660 7546 14688 9302
rect 16578 9200 16634 10000
rect 18786 9330 18842 10000
rect 18432 9302 18842 9330
rect 16592 7546 16620 9200
rect 18432 7546 18460 9302
rect 18786 9200 18842 9302
rect 18705 7644 19013 7653
rect 18705 7642 18711 7644
rect 18767 7642 18791 7644
rect 18847 7642 18871 7644
rect 18927 7642 18951 7644
rect 19007 7642 19013 7644
rect 18767 7590 18769 7642
rect 18949 7590 18951 7642
rect 18705 7588 18711 7590
rect 18767 7588 18791 7590
rect 18847 7588 18871 7590
rect 18927 7588 18951 7590
rect 19007 7588 19013 7590
rect 18705 7579 19013 7588
rect 12440 7540 12492 7546
rect 12360 7500 12440 7528
rect 12440 7482 12492 7488
rect 14648 7540 14700 7546
rect 14648 7482 14700 7488
rect 16580 7540 16632 7546
rect 16580 7482 16632 7488
rect 18420 7540 18472 7546
rect 18420 7482 18472 7488
rect 10232 7472 10284 7478
rect 10232 7414 10284 7420
rect 1860 7404 1912 7410
rect 1860 7346 1912 7352
rect 4620 7404 4672 7410
rect 4620 7346 4672 7352
rect 6920 7404 6972 7410
rect 6920 7346 6972 7352
rect 7104 7404 7156 7410
rect 7104 7346 7156 7352
rect 10600 7404 10652 7410
rect 10600 7346 10652 7352
rect 12532 7404 12584 7410
rect 12532 7346 12584 7352
rect 14648 7404 14700 7410
rect 14648 7346 14700 7352
rect 1872 2650 1900 7346
rect 3169 7100 3477 7109
rect 3169 7098 3175 7100
rect 3231 7098 3255 7100
rect 3311 7098 3335 7100
rect 3391 7098 3415 7100
rect 3471 7098 3477 7100
rect 3231 7046 3233 7098
rect 3413 7046 3415 7098
rect 3169 7044 3175 7046
rect 3231 7044 3255 7046
rect 3311 7044 3335 7046
rect 3391 7044 3415 7046
rect 3471 7044 3477 7046
rect 3169 7035 3477 7044
rect 3169 6012 3477 6021
rect 3169 6010 3175 6012
rect 3231 6010 3255 6012
rect 3311 6010 3335 6012
rect 3391 6010 3415 6012
rect 3471 6010 3477 6012
rect 3231 5958 3233 6010
rect 3413 5958 3415 6010
rect 3169 5956 3175 5958
rect 3231 5956 3255 5958
rect 3311 5956 3335 5958
rect 3391 5956 3415 5958
rect 3471 5956 3477 5958
rect 3169 5947 3477 5956
rect 2872 5704 2924 5710
rect 2872 5646 2924 5652
rect 3976 5704 4028 5710
rect 3976 5646 4028 5652
rect 2884 5370 2912 5646
rect 3056 5568 3108 5574
rect 3056 5510 3108 5516
rect 2872 5364 2924 5370
rect 2872 5306 2924 5312
rect 2136 5228 2188 5234
rect 2136 5170 2188 5176
rect 1952 5024 2004 5030
rect 1952 4966 2004 4972
rect 1964 4146 1992 4966
rect 2044 4616 2096 4622
rect 2044 4558 2096 4564
rect 1952 4140 2004 4146
rect 1952 4082 2004 4088
rect 2056 3534 2084 4558
rect 2044 3528 2096 3534
rect 2044 3470 2096 3476
rect 2056 3194 2084 3470
rect 2044 3188 2096 3194
rect 2044 3130 2096 3136
rect 2148 3126 2176 5170
rect 2596 5092 2648 5098
rect 2596 5034 2648 5040
rect 2608 4282 2636 5034
rect 3068 4622 3096 5510
rect 3884 5364 3936 5370
rect 3884 5306 3936 5312
rect 3896 5234 3924 5306
rect 3700 5228 3752 5234
rect 3700 5170 3752 5176
rect 3884 5228 3936 5234
rect 3884 5170 3936 5176
rect 3169 4924 3477 4933
rect 3169 4922 3175 4924
rect 3231 4922 3255 4924
rect 3311 4922 3335 4924
rect 3391 4922 3415 4924
rect 3471 4922 3477 4924
rect 3231 4870 3233 4922
rect 3413 4870 3415 4922
rect 3169 4868 3175 4870
rect 3231 4868 3255 4870
rect 3311 4868 3335 4870
rect 3391 4868 3415 4870
rect 3471 4868 3477 4870
rect 3169 4859 3477 4868
rect 3712 4758 3740 5170
rect 3988 4826 4016 5646
rect 4632 5166 4660 7346
rect 5388 6556 5696 6565
rect 5388 6554 5394 6556
rect 5450 6554 5474 6556
rect 5530 6554 5554 6556
rect 5610 6554 5634 6556
rect 5690 6554 5696 6556
rect 5450 6502 5452 6554
rect 5632 6502 5634 6554
rect 5388 6500 5394 6502
rect 5450 6500 5474 6502
rect 5530 6500 5554 6502
rect 5610 6500 5634 6502
rect 5690 6500 5696 6502
rect 5388 6491 5696 6500
rect 5908 5772 5960 5778
rect 5908 5714 5960 5720
rect 6828 5772 6880 5778
rect 6828 5714 6880 5720
rect 5724 5704 5776 5710
rect 5724 5646 5776 5652
rect 5388 5468 5696 5477
rect 5388 5466 5394 5468
rect 5450 5466 5474 5468
rect 5530 5466 5554 5468
rect 5610 5466 5634 5468
rect 5690 5466 5696 5468
rect 5450 5414 5452 5466
rect 5632 5414 5634 5466
rect 5388 5412 5394 5414
rect 5450 5412 5474 5414
rect 5530 5412 5554 5414
rect 5610 5412 5634 5414
rect 5690 5412 5696 5414
rect 5388 5403 5696 5412
rect 5080 5228 5132 5234
rect 5080 5170 5132 5176
rect 4620 5160 4672 5166
rect 4620 5102 4672 5108
rect 3976 4820 4028 4826
rect 3976 4762 4028 4768
rect 3700 4752 3752 4758
rect 3700 4694 3752 4700
rect 4342 4720 4398 4729
rect 4342 4655 4344 4664
rect 4396 4655 4398 4664
rect 4344 4626 4396 4632
rect 3056 4616 3108 4622
rect 3056 4558 3108 4564
rect 4252 4480 4304 4486
rect 4252 4422 4304 4428
rect 2596 4276 2648 4282
rect 2596 4218 2648 4224
rect 3976 4140 4028 4146
rect 3976 4082 4028 4088
rect 3169 3836 3477 3845
rect 3169 3834 3175 3836
rect 3231 3834 3255 3836
rect 3311 3834 3335 3836
rect 3391 3834 3415 3836
rect 3471 3834 3477 3836
rect 3231 3782 3233 3834
rect 3413 3782 3415 3834
rect 3169 3780 3175 3782
rect 3231 3780 3255 3782
rect 3311 3780 3335 3782
rect 3391 3780 3415 3782
rect 3471 3780 3477 3782
rect 3169 3771 3477 3780
rect 3988 3602 4016 4082
rect 3976 3596 4028 3602
rect 3976 3538 4028 3544
rect 3988 3194 4016 3538
rect 4264 3534 4292 4422
rect 4632 4282 4660 5102
rect 4712 5024 4764 5030
rect 4712 4966 4764 4972
rect 4804 5024 4856 5030
rect 4804 4966 4856 4972
rect 4724 4282 4752 4966
rect 4620 4276 4672 4282
rect 4620 4218 4672 4224
rect 4712 4276 4764 4282
rect 4712 4218 4764 4224
rect 4816 4214 4844 4966
rect 5092 4622 5120 5170
rect 5736 5098 5764 5646
rect 5920 5302 5948 5714
rect 6000 5568 6052 5574
rect 6000 5510 6052 5516
rect 5908 5296 5960 5302
rect 5908 5238 5960 5244
rect 5724 5092 5776 5098
rect 5724 5034 5776 5040
rect 5736 4690 5764 5034
rect 6012 4826 6040 5510
rect 6564 5086 6776 5114
rect 6564 4826 6592 5086
rect 6748 5030 6776 5086
rect 6644 5024 6696 5030
rect 6644 4966 6696 4972
rect 6736 5024 6788 5030
rect 6736 4966 6788 4972
rect 6000 4820 6052 4826
rect 6000 4762 6052 4768
rect 6552 4820 6604 4826
rect 6552 4762 6604 4768
rect 6274 4720 6330 4729
rect 5724 4684 5776 4690
rect 6274 4655 6276 4664
rect 5724 4626 5776 4632
rect 6328 4655 6330 4664
rect 6276 4626 6328 4632
rect 5080 4616 5132 4622
rect 5078 4584 5080 4593
rect 6092 4616 6144 4622
rect 5132 4584 5134 4593
rect 5078 4519 5134 4528
rect 6090 4584 6092 4593
rect 6144 4584 6146 4593
rect 6090 4519 6146 4528
rect 6552 4548 6604 4554
rect 5724 4480 5776 4486
rect 5724 4422 5776 4428
rect 5388 4380 5696 4389
rect 5388 4378 5394 4380
rect 5450 4378 5474 4380
rect 5530 4378 5554 4380
rect 5610 4378 5634 4380
rect 5690 4378 5696 4380
rect 5450 4326 5452 4378
rect 5632 4326 5634 4378
rect 5388 4324 5394 4326
rect 5450 4324 5474 4326
rect 5530 4324 5554 4326
rect 5610 4324 5634 4326
rect 5690 4324 5696 4326
rect 5388 4315 5696 4324
rect 4804 4208 4856 4214
rect 4804 4150 4856 4156
rect 5736 4146 5764 4422
rect 6104 4214 6132 4519
rect 6552 4490 6604 4496
rect 6092 4208 6144 4214
rect 6092 4150 6144 4156
rect 5724 4140 5776 4146
rect 5724 4082 5776 4088
rect 4528 3936 4580 3942
rect 4528 3878 4580 3884
rect 4252 3528 4304 3534
rect 4252 3470 4304 3476
rect 3976 3188 4028 3194
rect 3976 3130 4028 3136
rect 2136 3120 2188 3126
rect 2136 3062 2188 3068
rect 2504 3052 2556 3058
rect 2504 2994 2556 3000
rect 1860 2644 1912 2650
rect 1860 2586 1912 2592
rect 2516 2310 2544 2994
rect 3169 2748 3477 2757
rect 3169 2746 3175 2748
rect 3231 2746 3255 2748
rect 3311 2746 3335 2748
rect 3391 2746 3415 2748
rect 3471 2746 3477 2748
rect 3231 2694 3233 2746
rect 3413 2694 3415 2746
rect 3169 2692 3175 2694
rect 3231 2692 3255 2694
rect 3311 2692 3335 2694
rect 3391 2692 3415 2694
rect 3471 2692 3477 2694
rect 3169 2683 3477 2692
rect 3988 2514 4016 3130
rect 3976 2508 4028 2514
rect 3976 2450 4028 2456
rect 4540 2378 4568 3878
rect 6104 3534 6132 4150
rect 6460 4072 6512 4078
rect 6460 4014 6512 4020
rect 6472 3738 6500 4014
rect 6564 4010 6592 4490
rect 6552 4004 6604 4010
rect 6552 3946 6604 3952
rect 6656 3738 6684 4966
rect 6736 4616 6788 4622
rect 6736 4558 6788 4564
rect 6748 4146 6776 4558
rect 6736 4140 6788 4146
rect 6736 4082 6788 4088
rect 6460 3732 6512 3738
rect 6460 3674 6512 3680
rect 6644 3732 6696 3738
rect 6644 3674 6696 3680
rect 6748 3670 6776 4082
rect 6736 3664 6788 3670
rect 6736 3606 6788 3612
rect 6840 3534 6868 5714
rect 6932 5302 6960 7346
rect 7012 5840 7064 5846
rect 7012 5782 7064 5788
rect 6920 5296 6972 5302
rect 6920 5238 6972 5244
rect 6932 4078 6960 5238
rect 7024 4622 7052 5782
rect 7116 5574 7144 7346
rect 10324 7268 10376 7274
rect 10324 7210 10376 7216
rect 7608 7100 7916 7109
rect 7608 7098 7614 7100
rect 7670 7098 7694 7100
rect 7750 7098 7774 7100
rect 7830 7098 7854 7100
rect 7910 7098 7916 7100
rect 7670 7046 7672 7098
rect 7852 7046 7854 7098
rect 7608 7044 7614 7046
rect 7670 7044 7694 7046
rect 7750 7044 7774 7046
rect 7830 7044 7854 7046
rect 7910 7044 7916 7046
rect 7608 7035 7916 7044
rect 9827 6556 10135 6565
rect 9827 6554 9833 6556
rect 9889 6554 9913 6556
rect 9969 6554 9993 6556
rect 10049 6554 10073 6556
rect 10129 6554 10135 6556
rect 9889 6502 9891 6554
rect 10071 6502 10073 6554
rect 9827 6500 9833 6502
rect 9889 6500 9913 6502
rect 9969 6500 9993 6502
rect 10049 6500 10073 6502
rect 10129 6500 10135 6502
rect 9827 6491 10135 6500
rect 7608 6012 7916 6021
rect 7608 6010 7614 6012
rect 7670 6010 7694 6012
rect 7750 6010 7774 6012
rect 7830 6010 7854 6012
rect 7910 6010 7916 6012
rect 7670 5958 7672 6010
rect 7852 5958 7854 6010
rect 7608 5956 7614 5958
rect 7670 5956 7694 5958
rect 7750 5956 7774 5958
rect 7830 5956 7854 5958
rect 7910 5956 7916 5958
rect 7608 5947 7916 5956
rect 10232 5704 10284 5710
rect 10232 5646 10284 5652
rect 7196 5636 7248 5642
rect 7196 5578 7248 5584
rect 8300 5636 8352 5642
rect 8300 5578 8352 5584
rect 7104 5568 7156 5574
rect 7104 5510 7156 5516
rect 7012 4616 7064 4622
rect 7012 4558 7064 4564
rect 6920 4072 6972 4078
rect 6920 4014 6972 4020
rect 6920 3936 6972 3942
rect 6920 3878 6972 3884
rect 6092 3528 6144 3534
rect 6092 3470 6144 3476
rect 6552 3528 6604 3534
rect 6552 3470 6604 3476
rect 6828 3528 6880 3534
rect 6828 3470 6880 3476
rect 5388 3292 5696 3301
rect 5388 3290 5394 3292
rect 5450 3290 5474 3292
rect 5530 3290 5554 3292
rect 5610 3290 5634 3292
rect 5690 3290 5696 3292
rect 5450 3238 5452 3290
rect 5632 3238 5634 3290
rect 5388 3236 5394 3238
rect 5450 3236 5474 3238
rect 5530 3236 5554 3238
rect 5610 3236 5634 3238
rect 5690 3236 5696 3238
rect 5388 3227 5696 3236
rect 6564 2650 6592 3470
rect 6552 2644 6604 2650
rect 6552 2586 6604 2592
rect 6932 2446 6960 3878
rect 7116 3398 7144 5510
rect 7208 5370 7236 5578
rect 8312 5370 8340 5578
rect 9680 5568 9732 5574
rect 9680 5510 9732 5516
rect 7196 5364 7248 5370
rect 7196 5306 7248 5312
rect 8300 5364 8352 5370
rect 8300 5306 8352 5312
rect 9692 5234 9720 5510
rect 9827 5468 10135 5477
rect 9827 5466 9833 5468
rect 9889 5466 9913 5468
rect 9969 5466 9993 5468
rect 10049 5466 10073 5468
rect 10129 5466 10135 5468
rect 9889 5414 9891 5466
rect 10071 5414 10073 5466
rect 9827 5412 9833 5414
rect 9889 5412 9913 5414
rect 9969 5412 9993 5414
rect 10049 5412 10073 5414
rect 10129 5412 10135 5414
rect 9827 5403 10135 5412
rect 9312 5228 9364 5234
rect 9312 5170 9364 5176
rect 9680 5228 9732 5234
rect 9680 5170 9732 5176
rect 9772 5228 9824 5234
rect 9772 5170 9824 5176
rect 7288 5160 7340 5166
rect 7288 5102 7340 5108
rect 8392 5160 8444 5166
rect 8392 5102 8444 5108
rect 7300 4729 7328 5102
rect 7608 4924 7916 4933
rect 7608 4922 7614 4924
rect 7670 4922 7694 4924
rect 7750 4922 7774 4924
rect 7830 4922 7854 4924
rect 7910 4922 7916 4924
rect 7670 4870 7672 4922
rect 7852 4870 7854 4922
rect 7608 4868 7614 4870
rect 7670 4868 7694 4870
rect 7750 4868 7774 4870
rect 7830 4868 7854 4870
rect 7910 4868 7916 4870
rect 7608 4859 7916 4868
rect 7286 4720 7342 4729
rect 7286 4655 7342 4664
rect 7300 4486 7328 4655
rect 7288 4480 7340 4486
rect 7288 4422 7340 4428
rect 7380 4208 7432 4214
rect 7194 4176 7250 4185
rect 7380 4150 7432 4156
rect 7194 4111 7196 4120
rect 7248 4111 7250 4120
rect 7196 4082 7248 4088
rect 7104 3392 7156 3398
rect 7104 3334 7156 3340
rect 7392 3126 7420 4150
rect 8404 4078 8432 5102
rect 9128 5024 9180 5030
rect 9128 4966 9180 4972
rect 9220 5024 9272 5030
rect 9220 4966 9272 4972
rect 8392 4072 8444 4078
rect 8392 4014 8444 4020
rect 7608 3836 7916 3845
rect 7608 3834 7614 3836
rect 7670 3834 7694 3836
rect 7750 3834 7774 3836
rect 7830 3834 7854 3836
rect 7910 3834 7916 3836
rect 7670 3782 7672 3834
rect 7852 3782 7854 3834
rect 7608 3780 7614 3782
rect 7670 3780 7694 3782
rect 7750 3780 7774 3782
rect 7830 3780 7854 3782
rect 7910 3780 7916 3782
rect 7608 3771 7916 3780
rect 8404 3398 8432 4014
rect 9140 3534 9168 4966
rect 9232 4146 9260 4966
rect 9324 4214 9352 5170
rect 9784 4468 9812 5170
rect 9956 5160 10008 5166
rect 9956 5102 10008 5108
rect 9968 4826 9996 5102
rect 9956 4820 10008 4826
rect 9956 4762 10008 4768
rect 9692 4440 9812 4468
rect 9312 4208 9364 4214
rect 9310 4176 9312 4185
rect 9364 4176 9366 4185
rect 9220 4140 9272 4146
rect 9310 4111 9366 4120
rect 9220 4082 9272 4088
rect 9588 4072 9640 4078
rect 9588 4014 9640 4020
rect 9600 3602 9628 4014
rect 9588 3596 9640 3602
rect 9588 3538 9640 3544
rect 9128 3528 9180 3534
rect 9128 3470 9180 3476
rect 8392 3392 8444 3398
rect 8392 3334 8444 3340
rect 7380 3120 7432 3126
rect 7380 3062 7432 3068
rect 7472 3052 7524 3058
rect 7472 2994 7524 3000
rect 6920 2440 6972 2446
rect 6920 2382 6972 2388
rect 4528 2372 4580 2378
rect 4528 2314 4580 2320
rect 2504 2304 2556 2310
rect 2504 2246 2556 2252
rect 2516 800 2544 2246
rect 5388 2204 5696 2213
rect 5388 2202 5394 2204
rect 5450 2202 5474 2204
rect 5530 2202 5554 2204
rect 5610 2202 5634 2204
rect 5690 2202 5696 2204
rect 5450 2150 5452 2202
rect 5632 2150 5634 2202
rect 5388 2148 5394 2150
rect 5450 2148 5474 2150
rect 5530 2148 5554 2150
rect 5610 2148 5634 2150
rect 5690 2148 5696 2150
rect 5388 2139 5696 2148
rect 7484 800 7512 2994
rect 7608 2748 7916 2757
rect 7608 2746 7614 2748
rect 7670 2746 7694 2748
rect 7750 2746 7774 2748
rect 7830 2746 7854 2748
rect 7910 2746 7916 2748
rect 7670 2694 7672 2746
rect 7852 2694 7854 2746
rect 7608 2692 7614 2694
rect 7670 2692 7694 2694
rect 7750 2692 7774 2694
rect 7830 2692 7854 2694
rect 7910 2692 7916 2694
rect 7608 2683 7916 2692
rect 9692 2650 9720 4440
rect 9827 4380 10135 4389
rect 9827 4378 9833 4380
rect 9889 4378 9913 4380
rect 9969 4378 9993 4380
rect 10049 4378 10073 4380
rect 10129 4378 10135 4380
rect 9889 4326 9891 4378
rect 10071 4326 10073 4378
rect 9827 4324 9833 4326
rect 9889 4324 9913 4326
rect 9969 4324 9993 4326
rect 10049 4324 10073 4326
rect 10129 4324 10135 4326
rect 9827 4315 10135 4324
rect 10140 3732 10192 3738
rect 10244 3720 10272 5646
rect 10336 5642 10364 7210
rect 10508 5772 10560 5778
rect 10508 5714 10560 5720
rect 10324 5636 10376 5642
rect 10324 5578 10376 5584
rect 10520 5166 10548 5714
rect 10612 5710 10640 7346
rect 12047 7100 12355 7109
rect 12047 7098 12053 7100
rect 12109 7098 12133 7100
rect 12189 7098 12213 7100
rect 12269 7098 12293 7100
rect 12349 7098 12355 7100
rect 12109 7046 12111 7098
rect 12291 7046 12293 7098
rect 12047 7044 12053 7046
rect 12109 7044 12133 7046
rect 12189 7044 12213 7046
rect 12269 7044 12293 7046
rect 12349 7044 12355 7046
rect 12047 7035 12355 7044
rect 12047 6012 12355 6021
rect 12047 6010 12053 6012
rect 12109 6010 12133 6012
rect 12189 6010 12213 6012
rect 12269 6010 12293 6012
rect 12349 6010 12355 6012
rect 12109 5958 12111 6010
rect 12291 5958 12293 6010
rect 12047 5956 12053 5958
rect 12109 5956 12133 5958
rect 12189 5956 12213 5958
rect 12269 5956 12293 5958
rect 12349 5956 12355 5958
rect 12047 5947 12355 5956
rect 10876 5840 10928 5846
rect 10876 5782 10928 5788
rect 10600 5704 10652 5710
rect 10600 5646 10652 5652
rect 10508 5160 10560 5166
rect 10508 5102 10560 5108
rect 10888 4010 10916 5782
rect 11244 5704 11296 5710
rect 11244 5646 11296 5652
rect 10968 5636 11020 5642
rect 10968 5578 11020 5584
rect 10980 5370 11008 5578
rect 11060 5568 11112 5574
rect 11060 5510 11112 5516
rect 10968 5364 11020 5370
rect 10968 5306 11020 5312
rect 11072 5302 11100 5510
rect 11060 5296 11112 5302
rect 11060 5238 11112 5244
rect 11256 5098 11284 5646
rect 12544 5574 12572 7346
rect 13452 7336 13504 7342
rect 13452 7278 13504 7284
rect 12532 5568 12584 5574
rect 12532 5510 12584 5516
rect 11888 5160 11940 5166
rect 11888 5102 11940 5108
rect 11244 5092 11296 5098
rect 11164 5052 11244 5080
rect 11164 4826 11192 5052
rect 11244 5034 11296 5040
rect 11152 4820 11204 4826
rect 11152 4762 11204 4768
rect 11336 4616 11388 4622
rect 11336 4558 11388 4564
rect 11428 4616 11480 4622
rect 11428 4558 11480 4564
rect 11348 4146 11376 4558
rect 11440 4214 11468 4558
rect 11704 4548 11756 4554
rect 11704 4490 11756 4496
rect 11520 4276 11572 4282
rect 11520 4218 11572 4224
rect 11428 4208 11480 4214
rect 11428 4150 11480 4156
rect 11336 4140 11388 4146
rect 11336 4082 11388 4088
rect 10968 4072 11020 4078
rect 10968 4014 11020 4020
rect 10876 4004 10928 4010
rect 10876 3946 10928 3952
rect 10508 3936 10560 3942
rect 10508 3878 10560 3884
rect 10192 3692 10272 3720
rect 10140 3674 10192 3680
rect 10520 3534 10548 3878
rect 10508 3528 10560 3534
rect 10508 3470 10560 3476
rect 9827 3292 10135 3301
rect 9827 3290 9833 3292
rect 9889 3290 9913 3292
rect 9969 3290 9993 3292
rect 10049 3290 10073 3292
rect 10129 3290 10135 3292
rect 9889 3238 9891 3290
rect 10071 3238 10073 3290
rect 9827 3236 9833 3238
rect 9889 3236 9913 3238
rect 9969 3236 9993 3238
rect 10049 3236 10073 3238
rect 10129 3236 10135 3238
rect 9827 3227 10135 3236
rect 10980 3194 11008 4014
rect 9864 3188 9916 3194
rect 9864 3130 9916 3136
rect 10968 3188 11020 3194
rect 10968 3130 11020 3136
rect 9680 2644 9732 2650
rect 9680 2586 9732 2592
rect 9876 2310 9904 3130
rect 11532 3126 11560 4218
rect 11612 3936 11664 3942
rect 11612 3878 11664 3884
rect 11520 3120 11572 3126
rect 11520 3062 11572 3068
rect 11624 2650 11652 3878
rect 11716 2961 11744 4490
rect 11796 4140 11848 4146
rect 11796 4082 11848 4088
rect 11808 3602 11836 4082
rect 11796 3596 11848 3602
rect 11796 3538 11848 3544
rect 11808 3058 11836 3538
rect 11796 3052 11848 3058
rect 11796 2994 11848 3000
rect 11702 2952 11758 2961
rect 11702 2887 11758 2896
rect 11808 2774 11836 2994
rect 11716 2746 11836 2774
rect 10048 2644 10100 2650
rect 10048 2586 10100 2592
rect 11612 2644 11664 2650
rect 11612 2586 11664 2592
rect 10060 2378 10088 2586
rect 11716 2446 11744 2746
rect 11900 2650 11928 5102
rect 12047 4924 12355 4933
rect 12047 4922 12053 4924
rect 12109 4922 12133 4924
rect 12189 4922 12213 4924
rect 12269 4922 12293 4924
rect 12349 4922 12355 4924
rect 12109 4870 12111 4922
rect 12291 4870 12293 4922
rect 12047 4868 12053 4870
rect 12109 4868 12133 4870
rect 12189 4868 12213 4870
rect 12269 4868 12293 4870
rect 12349 4868 12355 4870
rect 12047 4859 12355 4868
rect 11980 4480 12032 4486
rect 11980 4422 12032 4428
rect 12440 4480 12492 4486
rect 12440 4422 12492 4428
rect 11992 4214 12020 4422
rect 11980 4208 12032 4214
rect 11980 4150 12032 4156
rect 12047 3836 12355 3845
rect 12047 3834 12053 3836
rect 12109 3834 12133 3836
rect 12189 3834 12213 3836
rect 12269 3834 12293 3836
rect 12349 3834 12355 3836
rect 12109 3782 12111 3834
rect 12291 3782 12293 3834
rect 12047 3780 12053 3782
rect 12109 3780 12133 3782
rect 12189 3780 12213 3782
rect 12269 3780 12293 3782
rect 12349 3780 12355 3782
rect 12047 3771 12355 3780
rect 12452 3534 12480 4422
rect 12544 3738 12572 5510
rect 13464 5370 13492 7278
rect 14266 6556 14574 6565
rect 14266 6554 14272 6556
rect 14328 6554 14352 6556
rect 14408 6554 14432 6556
rect 14488 6554 14512 6556
rect 14568 6554 14574 6556
rect 14328 6502 14330 6554
rect 14510 6502 14512 6554
rect 14266 6500 14272 6502
rect 14328 6500 14352 6502
rect 14408 6500 14432 6502
rect 14488 6500 14512 6502
rect 14568 6500 14574 6502
rect 14266 6491 14574 6500
rect 13544 5636 13596 5642
rect 13544 5578 13596 5584
rect 13556 5370 13584 5578
rect 14660 5574 14688 7346
rect 16486 7100 16794 7109
rect 16486 7098 16492 7100
rect 16548 7098 16572 7100
rect 16628 7098 16652 7100
rect 16708 7098 16732 7100
rect 16788 7098 16794 7100
rect 16548 7046 16550 7098
rect 16730 7046 16732 7098
rect 16486 7044 16492 7046
rect 16548 7044 16572 7046
rect 16628 7044 16652 7046
rect 16708 7044 16732 7046
rect 16788 7044 16794 7046
rect 16486 7035 16794 7044
rect 18705 6556 19013 6565
rect 18705 6554 18711 6556
rect 18767 6554 18791 6556
rect 18847 6554 18871 6556
rect 18927 6554 18951 6556
rect 19007 6554 19013 6556
rect 18767 6502 18769 6554
rect 18949 6502 18951 6554
rect 18705 6500 18711 6502
rect 18767 6500 18791 6502
rect 18847 6500 18871 6502
rect 18927 6500 18951 6502
rect 19007 6500 19013 6502
rect 18705 6491 19013 6500
rect 16486 6012 16794 6021
rect 16486 6010 16492 6012
rect 16548 6010 16572 6012
rect 16628 6010 16652 6012
rect 16708 6010 16732 6012
rect 16788 6010 16794 6012
rect 16548 5958 16550 6010
rect 16730 5958 16732 6010
rect 16486 5956 16492 5958
rect 16548 5956 16572 5958
rect 16628 5956 16652 5958
rect 16708 5956 16732 5958
rect 16788 5956 16794 5958
rect 16486 5947 16794 5956
rect 14832 5772 14884 5778
rect 14832 5714 14884 5720
rect 13820 5568 13872 5574
rect 13820 5510 13872 5516
rect 14648 5568 14700 5574
rect 14648 5510 14700 5516
rect 13452 5364 13504 5370
rect 13452 5306 13504 5312
rect 13544 5364 13596 5370
rect 13544 5306 13596 5312
rect 12992 5160 13044 5166
rect 12992 5102 13044 5108
rect 12624 4752 12676 4758
rect 12624 4694 12676 4700
rect 12636 4554 12664 4694
rect 13004 4622 13032 5102
rect 13084 5024 13136 5030
rect 13084 4966 13136 4972
rect 13096 4826 13124 4966
rect 13084 4820 13136 4826
rect 13084 4762 13136 4768
rect 12992 4616 13044 4622
rect 12992 4558 13044 4564
rect 13268 4616 13320 4622
rect 13268 4558 13320 4564
rect 12624 4548 12676 4554
rect 12624 4490 12676 4496
rect 12532 3732 12584 3738
rect 12532 3674 12584 3680
rect 12440 3528 12492 3534
rect 12440 3470 12492 3476
rect 13004 3466 13032 4558
rect 12992 3460 13044 3466
rect 12992 3402 13044 3408
rect 12440 2848 12492 2854
rect 12440 2790 12492 2796
rect 12047 2748 12355 2757
rect 12047 2746 12053 2748
rect 12109 2746 12133 2748
rect 12189 2746 12213 2748
rect 12269 2746 12293 2748
rect 12349 2746 12355 2748
rect 12109 2694 12111 2746
rect 12291 2694 12293 2746
rect 12047 2692 12053 2694
rect 12109 2692 12133 2694
rect 12189 2692 12213 2694
rect 12269 2692 12293 2694
rect 12349 2692 12355 2694
rect 12047 2683 12355 2692
rect 11888 2644 11940 2650
rect 11888 2586 11940 2592
rect 11704 2440 11756 2446
rect 11704 2382 11756 2388
rect 10048 2372 10100 2378
rect 10048 2314 10100 2320
rect 9864 2304 9916 2310
rect 9864 2246 9916 2252
rect 9827 2204 10135 2213
rect 9827 2202 9833 2204
rect 9889 2202 9913 2204
rect 9969 2202 9993 2204
rect 10049 2202 10073 2204
rect 10129 2202 10135 2204
rect 9889 2150 9891 2202
rect 10071 2150 10073 2202
rect 9827 2148 9833 2150
rect 9889 2148 9913 2150
rect 9969 2148 9993 2150
rect 10049 2148 10073 2150
rect 10129 2148 10135 2150
rect 9827 2139 10135 2148
rect 12452 800 12480 2790
rect 13004 2650 13032 3402
rect 13280 3194 13308 4558
rect 13464 4282 13492 5306
rect 13832 4690 13860 5510
rect 14266 5468 14574 5477
rect 14266 5466 14272 5468
rect 14328 5466 14352 5468
rect 14408 5466 14432 5468
rect 14488 5466 14512 5468
rect 14568 5466 14574 5468
rect 14328 5414 14330 5466
rect 14510 5414 14512 5466
rect 14266 5412 14272 5414
rect 14328 5412 14352 5414
rect 14408 5412 14432 5414
rect 14488 5412 14512 5414
rect 14568 5412 14574 5414
rect 14266 5403 14574 5412
rect 14556 5092 14608 5098
rect 14556 5034 14608 5040
rect 13820 4684 13872 4690
rect 13820 4626 13872 4632
rect 14568 4622 14596 5034
rect 14556 4616 14608 4622
rect 14556 4558 14608 4564
rect 14266 4380 14574 4389
rect 14266 4378 14272 4380
rect 14328 4378 14352 4380
rect 14408 4378 14432 4380
rect 14488 4378 14512 4380
rect 14568 4378 14574 4380
rect 14328 4326 14330 4378
rect 14510 4326 14512 4378
rect 14266 4324 14272 4326
rect 14328 4324 14352 4326
rect 14408 4324 14432 4326
rect 14488 4324 14512 4326
rect 14568 4324 14574 4326
rect 14266 4315 14574 4324
rect 13452 4276 13504 4282
rect 13452 4218 13504 4224
rect 14660 3738 14688 5510
rect 14740 4616 14792 4622
rect 14740 4558 14792 4564
rect 14752 4078 14780 4558
rect 14844 4146 14872 5714
rect 18705 5468 19013 5477
rect 18705 5466 18711 5468
rect 18767 5466 18791 5468
rect 18847 5466 18871 5468
rect 18927 5466 18951 5468
rect 19007 5466 19013 5468
rect 18767 5414 18769 5466
rect 18949 5414 18951 5466
rect 18705 5412 18711 5414
rect 18767 5412 18791 5414
rect 18847 5412 18871 5414
rect 18927 5412 18951 5414
rect 19007 5412 19013 5414
rect 18705 5403 19013 5412
rect 16486 4924 16794 4933
rect 16486 4922 16492 4924
rect 16548 4922 16572 4924
rect 16628 4922 16652 4924
rect 16708 4922 16732 4924
rect 16788 4922 16794 4924
rect 16548 4870 16550 4922
rect 16730 4870 16732 4922
rect 16486 4868 16492 4870
rect 16548 4868 16572 4870
rect 16628 4868 16652 4870
rect 16708 4868 16732 4870
rect 16788 4868 16794 4870
rect 16486 4859 16794 4868
rect 17408 4752 17460 4758
rect 17408 4694 17460 4700
rect 15660 4480 15712 4486
rect 15660 4422 15712 4428
rect 15672 4146 15700 4422
rect 14832 4140 14884 4146
rect 14832 4082 14884 4088
rect 15660 4140 15712 4146
rect 15660 4082 15712 4088
rect 14740 4072 14792 4078
rect 14740 4014 14792 4020
rect 14648 3732 14700 3738
rect 14648 3674 14700 3680
rect 14266 3292 14574 3301
rect 14266 3290 14272 3292
rect 14328 3290 14352 3292
rect 14408 3290 14432 3292
rect 14488 3290 14512 3292
rect 14568 3290 14574 3292
rect 14328 3238 14330 3290
rect 14510 3238 14512 3290
rect 14266 3236 14272 3238
rect 14328 3236 14352 3238
rect 14408 3236 14432 3238
rect 14488 3236 14512 3238
rect 14568 3236 14574 3238
rect 14266 3227 14574 3236
rect 13268 3188 13320 3194
rect 13268 3130 13320 3136
rect 14844 3126 14872 4082
rect 16396 4004 16448 4010
rect 16396 3946 16448 3952
rect 16408 3516 16436 3946
rect 17224 3936 17276 3942
rect 17224 3878 17276 3884
rect 16486 3836 16794 3845
rect 16486 3834 16492 3836
rect 16548 3834 16572 3836
rect 16628 3834 16652 3836
rect 16708 3834 16732 3836
rect 16788 3834 16794 3836
rect 16548 3782 16550 3834
rect 16730 3782 16732 3834
rect 16486 3780 16492 3782
rect 16548 3780 16572 3782
rect 16628 3780 16652 3782
rect 16708 3780 16732 3782
rect 16788 3780 16794 3782
rect 16486 3771 16794 3780
rect 16488 3528 16540 3534
rect 16408 3488 16488 3516
rect 16488 3470 16540 3476
rect 15752 3392 15804 3398
rect 15752 3334 15804 3340
rect 17040 3392 17092 3398
rect 17040 3334 17092 3340
rect 14832 3120 14884 3126
rect 14832 3062 14884 3068
rect 14280 2916 14332 2922
rect 14280 2858 14332 2864
rect 14292 2650 14320 2858
rect 14740 2848 14792 2854
rect 14740 2790 14792 2796
rect 12992 2644 13044 2650
rect 12992 2586 13044 2592
rect 14280 2644 14332 2650
rect 14280 2586 14332 2592
rect 14752 2378 14780 2790
rect 14740 2372 14792 2378
rect 14740 2314 14792 2320
rect 15764 2310 15792 3334
rect 17052 3058 17080 3334
rect 17040 3052 17092 3058
rect 17040 2994 17092 3000
rect 16854 2952 16910 2961
rect 16854 2887 16910 2896
rect 16486 2748 16794 2757
rect 16486 2746 16492 2748
rect 16548 2746 16572 2748
rect 16628 2746 16652 2748
rect 16708 2746 16732 2748
rect 16788 2746 16794 2748
rect 16548 2694 16550 2746
rect 16730 2694 16732 2746
rect 16486 2692 16492 2694
rect 16548 2692 16572 2694
rect 16628 2692 16652 2694
rect 16708 2692 16732 2694
rect 16788 2692 16794 2694
rect 16486 2683 16794 2692
rect 16868 2650 16896 2887
rect 16856 2644 16908 2650
rect 16856 2586 16908 2592
rect 17236 2446 17264 3878
rect 17420 3534 17448 4694
rect 18705 4380 19013 4389
rect 18705 4378 18711 4380
rect 18767 4378 18791 4380
rect 18847 4378 18871 4380
rect 18927 4378 18951 4380
rect 19007 4378 19013 4380
rect 18767 4326 18769 4378
rect 18949 4326 18951 4378
rect 18705 4324 18711 4326
rect 18767 4324 18791 4326
rect 18847 4324 18871 4326
rect 18927 4324 18951 4326
rect 19007 4324 19013 4326
rect 18705 4315 19013 4324
rect 17500 3596 17552 3602
rect 17500 3538 17552 3544
rect 17408 3528 17460 3534
rect 17408 3470 17460 3476
rect 17512 2446 17540 3538
rect 18705 3292 19013 3301
rect 18705 3290 18711 3292
rect 18767 3290 18791 3292
rect 18847 3290 18871 3292
rect 18927 3290 18951 3292
rect 19007 3290 19013 3292
rect 18767 3238 18769 3290
rect 18949 3238 18951 3290
rect 18705 3236 18711 3238
rect 18767 3236 18791 3238
rect 18847 3236 18871 3238
rect 18927 3236 18951 3238
rect 19007 3236 19013 3238
rect 18705 3227 19013 3236
rect 17224 2440 17276 2446
rect 17224 2382 17276 2388
rect 17500 2440 17552 2446
rect 17500 2382 17552 2388
rect 15752 2304 15804 2310
rect 15752 2246 15804 2252
rect 17408 2304 17460 2310
rect 17408 2246 17460 2252
rect 14266 2204 14574 2213
rect 14266 2202 14272 2204
rect 14328 2202 14352 2204
rect 14408 2202 14432 2204
rect 14488 2202 14512 2204
rect 14568 2202 14574 2204
rect 14328 2150 14330 2202
rect 14510 2150 14512 2202
rect 14266 2148 14272 2150
rect 14328 2148 14352 2150
rect 14408 2148 14432 2150
rect 14488 2148 14512 2150
rect 14568 2148 14574 2150
rect 14266 2139 14574 2148
rect 17420 800 17448 2246
rect 18705 2204 19013 2213
rect 18705 2202 18711 2204
rect 18767 2202 18791 2204
rect 18847 2202 18871 2204
rect 18927 2202 18951 2204
rect 19007 2202 19013 2204
rect 18767 2150 18769 2202
rect 18949 2150 18951 2202
rect 18705 2148 18711 2150
rect 18767 2148 18791 2150
rect 18847 2148 18871 2150
rect 18927 2148 18951 2150
rect 19007 2148 19013 2150
rect 18705 2139 19013 2148
rect 2502 0 2558 800
rect 7470 0 7526 800
rect 12438 0 12494 800
rect 17406 0 17462 800
<< via2 >>
rect 5394 7642 5450 7644
rect 5474 7642 5530 7644
rect 5554 7642 5610 7644
rect 5634 7642 5690 7644
rect 5394 7590 5440 7642
rect 5440 7590 5450 7642
rect 5474 7590 5504 7642
rect 5504 7590 5516 7642
rect 5516 7590 5530 7642
rect 5554 7590 5568 7642
rect 5568 7590 5580 7642
rect 5580 7590 5610 7642
rect 5634 7590 5644 7642
rect 5644 7590 5690 7642
rect 5394 7588 5450 7590
rect 5474 7588 5530 7590
rect 5554 7588 5610 7590
rect 5634 7588 5690 7590
rect 9833 7642 9889 7644
rect 9913 7642 9969 7644
rect 9993 7642 10049 7644
rect 10073 7642 10129 7644
rect 9833 7590 9879 7642
rect 9879 7590 9889 7642
rect 9913 7590 9943 7642
rect 9943 7590 9955 7642
rect 9955 7590 9969 7642
rect 9993 7590 10007 7642
rect 10007 7590 10019 7642
rect 10019 7590 10049 7642
rect 10073 7590 10083 7642
rect 10083 7590 10129 7642
rect 9833 7588 9889 7590
rect 9913 7588 9969 7590
rect 9993 7588 10049 7590
rect 10073 7588 10129 7590
rect 14272 7642 14328 7644
rect 14352 7642 14408 7644
rect 14432 7642 14488 7644
rect 14512 7642 14568 7644
rect 14272 7590 14318 7642
rect 14318 7590 14328 7642
rect 14352 7590 14382 7642
rect 14382 7590 14394 7642
rect 14394 7590 14408 7642
rect 14432 7590 14446 7642
rect 14446 7590 14458 7642
rect 14458 7590 14488 7642
rect 14512 7590 14522 7642
rect 14522 7590 14568 7642
rect 14272 7588 14328 7590
rect 14352 7588 14408 7590
rect 14432 7588 14488 7590
rect 14512 7588 14568 7590
rect 18711 7642 18767 7644
rect 18791 7642 18847 7644
rect 18871 7642 18927 7644
rect 18951 7642 19007 7644
rect 18711 7590 18757 7642
rect 18757 7590 18767 7642
rect 18791 7590 18821 7642
rect 18821 7590 18833 7642
rect 18833 7590 18847 7642
rect 18871 7590 18885 7642
rect 18885 7590 18897 7642
rect 18897 7590 18927 7642
rect 18951 7590 18961 7642
rect 18961 7590 19007 7642
rect 18711 7588 18767 7590
rect 18791 7588 18847 7590
rect 18871 7588 18927 7590
rect 18951 7588 19007 7590
rect 3175 7098 3231 7100
rect 3255 7098 3311 7100
rect 3335 7098 3391 7100
rect 3415 7098 3471 7100
rect 3175 7046 3221 7098
rect 3221 7046 3231 7098
rect 3255 7046 3285 7098
rect 3285 7046 3297 7098
rect 3297 7046 3311 7098
rect 3335 7046 3349 7098
rect 3349 7046 3361 7098
rect 3361 7046 3391 7098
rect 3415 7046 3425 7098
rect 3425 7046 3471 7098
rect 3175 7044 3231 7046
rect 3255 7044 3311 7046
rect 3335 7044 3391 7046
rect 3415 7044 3471 7046
rect 3175 6010 3231 6012
rect 3255 6010 3311 6012
rect 3335 6010 3391 6012
rect 3415 6010 3471 6012
rect 3175 5958 3221 6010
rect 3221 5958 3231 6010
rect 3255 5958 3285 6010
rect 3285 5958 3297 6010
rect 3297 5958 3311 6010
rect 3335 5958 3349 6010
rect 3349 5958 3361 6010
rect 3361 5958 3391 6010
rect 3415 5958 3425 6010
rect 3425 5958 3471 6010
rect 3175 5956 3231 5958
rect 3255 5956 3311 5958
rect 3335 5956 3391 5958
rect 3415 5956 3471 5958
rect 3175 4922 3231 4924
rect 3255 4922 3311 4924
rect 3335 4922 3391 4924
rect 3415 4922 3471 4924
rect 3175 4870 3221 4922
rect 3221 4870 3231 4922
rect 3255 4870 3285 4922
rect 3285 4870 3297 4922
rect 3297 4870 3311 4922
rect 3335 4870 3349 4922
rect 3349 4870 3361 4922
rect 3361 4870 3391 4922
rect 3415 4870 3425 4922
rect 3425 4870 3471 4922
rect 3175 4868 3231 4870
rect 3255 4868 3311 4870
rect 3335 4868 3391 4870
rect 3415 4868 3471 4870
rect 5394 6554 5450 6556
rect 5474 6554 5530 6556
rect 5554 6554 5610 6556
rect 5634 6554 5690 6556
rect 5394 6502 5440 6554
rect 5440 6502 5450 6554
rect 5474 6502 5504 6554
rect 5504 6502 5516 6554
rect 5516 6502 5530 6554
rect 5554 6502 5568 6554
rect 5568 6502 5580 6554
rect 5580 6502 5610 6554
rect 5634 6502 5644 6554
rect 5644 6502 5690 6554
rect 5394 6500 5450 6502
rect 5474 6500 5530 6502
rect 5554 6500 5610 6502
rect 5634 6500 5690 6502
rect 5394 5466 5450 5468
rect 5474 5466 5530 5468
rect 5554 5466 5610 5468
rect 5634 5466 5690 5468
rect 5394 5414 5440 5466
rect 5440 5414 5450 5466
rect 5474 5414 5504 5466
rect 5504 5414 5516 5466
rect 5516 5414 5530 5466
rect 5554 5414 5568 5466
rect 5568 5414 5580 5466
rect 5580 5414 5610 5466
rect 5634 5414 5644 5466
rect 5644 5414 5690 5466
rect 5394 5412 5450 5414
rect 5474 5412 5530 5414
rect 5554 5412 5610 5414
rect 5634 5412 5690 5414
rect 4342 4684 4398 4720
rect 4342 4664 4344 4684
rect 4344 4664 4396 4684
rect 4396 4664 4398 4684
rect 3175 3834 3231 3836
rect 3255 3834 3311 3836
rect 3335 3834 3391 3836
rect 3415 3834 3471 3836
rect 3175 3782 3221 3834
rect 3221 3782 3231 3834
rect 3255 3782 3285 3834
rect 3285 3782 3297 3834
rect 3297 3782 3311 3834
rect 3335 3782 3349 3834
rect 3349 3782 3361 3834
rect 3361 3782 3391 3834
rect 3415 3782 3425 3834
rect 3425 3782 3471 3834
rect 3175 3780 3231 3782
rect 3255 3780 3311 3782
rect 3335 3780 3391 3782
rect 3415 3780 3471 3782
rect 6274 4684 6330 4720
rect 6274 4664 6276 4684
rect 6276 4664 6328 4684
rect 6328 4664 6330 4684
rect 5078 4564 5080 4584
rect 5080 4564 5132 4584
rect 5132 4564 5134 4584
rect 5078 4528 5134 4564
rect 6090 4564 6092 4584
rect 6092 4564 6144 4584
rect 6144 4564 6146 4584
rect 6090 4528 6146 4564
rect 5394 4378 5450 4380
rect 5474 4378 5530 4380
rect 5554 4378 5610 4380
rect 5634 4378 5690 4380
rect 5394 4326 5440 4378
rect 5440 4326 5450 4378
rect 5474 4326 5504 4378
rect 5504 4326 5516 4378
rect 5516 4326 5530 4378
rect 5554 4326 5568 4378
rect 5568 4326 5580 4378
rect 5580 4326 5610 4378
rect 5634 4326 5644 4378
rect 5644 4326 5690 4378
rect 5394 4324 5450 4326
rect 5474 4324 5530 4326
rect 5554 4324 5610 4326
rect 5634 4324 5690 4326
rect 3175 2746 3231 2748
rect 3255 2746 3311 2748
rect 3335 2746 3391 2748
rect 3415 2746 3471 2748
rect 3175 2694 3221 2746
rect 3221 2694 3231 2746
rect 3255 2694 3285 2746
rect 3285 2694 3297 2746
rect 3297 2694 3311 2746
rect 3335 2694 3349 2746
rect 3349 2694 3361 2746
rect 3361 2694 3391 2746
rect 3415 2694 3425 2746
rect 3425 2694 3471 2746
rect 3175 2692 3231 2694
rect 3255 2692 3311 2694
rect 3335 2692 3391 2694
rect 3415 2692 3471 2694
rect 7614 7098 7670 7100
rect 7694 7098 7750 7100
rect 7774 7098 7830 7100
rect 7854 7098 7910 7100
rect 7614 7046 7660 7098
rect 7660 7046 7670 7098
rect 7694 7046 7724 7098
rect 7724 7046 7736 7098
rect 7736 7046 7750 7098
rect 7774 7046 7788 7098
rect 7788 7046 7800 7098
rect 7800 7046 7830 7098
rect 7854 7046 7864 7098
rect 7864 7046 7910 7098
rect 7614 7044 7670 7046
rect 7694 7044 7750 7046
rect 7774 7044 7830 7046
rect 7854 7044 7910 7046
rect 9833 6554 9889 6556
rect 9913 6554 9969 6556
rect 9993 6554 10049 6556
rect 10073 6554 10129 6556
rect 9833 6502 9879 6554
rect 9879 6502 9889 6554
rect 9913 6502 9943 6554
rect 9943 6502 9955 6554
rect 9955 6502 9969 6554
rect 9993 6502 10007 6554
rect 10007 6502 10019 6554
rect 10019 6502 10049 6554
rect 10073 6502 10083 6554
rect 10083 6502 10129 6554
rect 9833 6500 9889 6502
rect 9913 6500 9969 6502
rect 9993 6500 10049 6502
rect 10073 6500 10129 6502
rect 7614 6010 7670 6012
rect 7694 6010 7750 6012
rect 7774 6010 7830 6012
rect 7854 6010 7910 6012
rect 7614 5958 7660 6010
rect 7660 5958 7670 6010
rect 7694 5958 7724 6010
rect 7724 5958 7736 6010
rect 7736 5958 7750 6010
rect 7774 5958 7788 6010
rect 7788 5958 7800 6010
rect 7800 5958 7830 6010
rect 7854 5958 7864 6010
rect 7864 5958 7910 6010
rect 7614 5956 7670 5958
rect 7694 5956 7750 5958
rect 7774 5956 7830 5958
rect 7854 5956 7910 5958
rect 5394 3290 5450 3292
rect 5474 3290 5530 3292
rect 5554 3290 5610 3292
rect 5634 3290 5690 3292
rect 5394 3238 5440 3290
rect 5440 3238 5450 3290
rect 5474 3238 5504 3290
rect 5504 3238 5516 3290
rect 5516 3238 5530 3290
rect 5554 3238 5568 3290
rect 5568 3238 5580 3290
rect 5580 3238 5610 3290
rect 5634 3238 5644 3290
rect 5644 3238 5690 3290
rect 5394 3236 5450 3238
rect 5474 3236 5530 3238
rect 5554 3236 5610 3238
rect 5634 3236 5690 3238
rect 9833 5466 9889 5468
rect 9913 5466 9969 5468
rect 9993 5466 10049 5468
rect 10073 5466 10129 5468
rect 9833 5414 9879 5466
rect 9879 5414 9889 5466
rect 9913 5414 9943 5466
rect 9943 5414 9955 5466
rect 9955 5414 9969 5466
rect 9993 5414 10007 5466
rect 10007 5414 10019 5466
rect 10019 5414 10049 5466
rect 10073 5414 10083 5466
rect 10083 5414 10129 5466
rect 9833 5412 9889 5414
rect 9913 5412 9969 5414
rect 9993 5412 10049 5414
rect 10073 5412 10129 5414
rect 7614 4922 7670 4924
rect 7694 4922 7750 4924
rect 7774 4922 7830 4924
rect 7854 4922 7910 4924
rect 7614 4870 7660 4922
rect 7660 4870 7670 4922
rect 7694 4870 7724 4922
rect 7724 4870 7736 4922
rect 7736 4870 7750 4922
rect 7774 4870 7788 4922
rect 7788 4870 7800 4922
rect 7800 4870 7830 4922
rect 7854 4870 7864 4922
rect 7864 4870 7910 4922
rect 7614 4868 7670 4870
rect 7694 4868 7750 4870
rect 7774 4868 7830 4870
rect 7854 4868 7910 4870
rect 7286 4664 7342 4720
rect 7194 4140 7250 4176
rect 7194 4120 7196 4140
rect 7196 4120 7248 4140
rect 7248 4120 7250 4140
rect 7614 3834 7670 3836
rect 7694 3834 7750 3836
rect 7774 3834 7830 3836
rect 7854 3834 7910 3836
rect 7614 3782 7660 3834
rect 7660 3782 7670 3834
rect 7694 3782 7724 3834
rect 7724 3782 7736 3834
rect 7736 3782 7750 3834
rect 7774 3782 7788 3834
rect 7788 3782 7800 3834
rect 7800 3782 7830 3834
rect 7854 3782 7864 3834
rect 7864 3782 7910 3834
rect 7614 3780 7670 3782
rect 7694 3780 7750 3782
rect 7774 3780 7830 3782
rect 7854 3780 7910 3782
rect 9310 4156 9312 4176
rect 9312 4156 9364 4176
rect 9364 4156 9366 4176
rect 9310 4120 9366 4156
rect 5394 2202 5450 2204
rect 5474 2202 5530 2204
rect 5554 2202 5610 2204
rect 5634 2202 5690 2204
rect 5394 2150 5440 2202
rect 5440 2150 5450 2202
rect 5474 2150 5504 2202
rect 5504 2150 5516 2202
rect 5516 2150 5530 2202
rect 5554 2150 5568 2202
rect 5568 2150 5580 2202
rect 5580 2150 5610 2202
rect 5634 2150 5644 2202
rect 5644 2150 5690 2202
rect 5394 2148 5450 2150
rect 5474 2148 5530 2150
rect 5554 2148 5610 2150
rect 5634 2148 5690 2150
rect 7614 2746 7670 2748
rect 7694 2746 7750 2748
rect 7774 2746 7830 2748
rect 7854 2746 7910 2748
rect 7614 2694 7660 2746
rect 7660 2694 7670 2746
rect 7694 2694 7724 2746
rect 7724 2694 7736 2746
rect 7736 2694 7750 2746
rect 7774 2694 7788 2746
rect 7788 2694 7800 2746
rect 7800 2694 7830 2746
rect 7854 2694 7864 2746
rect 7864 2694 7910 2746
rect 7614 2692 7670 2694
rect 7694 2692 7750 2694
rect 7774 2692 7830 2694
rect 7854 2692 7910 2694
rect 9833 4378 9889 4380
rect 9913 4378 9969 4380
rect 9993 4378 10049 4380
rect 10073 4378 10129 4380
rect 9833 4326 9879 4378
rect 9879 4326 9889 4378
rect 9913 4326 9943 4378
rect 9943 4326 9955 4378
rect 9955 4326 9969 4378
rect 9993 4326 10007 4378
rect 10007 4326 10019 4378
rect 10019 4326 10049 4378
rect 10073 4326 10083 4378
rect 10083 4326 10129 4378
rect 9833 4324 9889 4326
rect 9913 4324 9969 4326
rect 9993 4324 10049 4326
rect 10073 4324 10129 4326
rect 12053 7098 12109 7100
rect 12133 7098 12189 7100
rect 12213 7098 12269 7100
rect 12293 7098 12349 7100
rect 12053 7046 12099 7098
rect 12099 7046 12109 7098
rect 12133 7046 12163 7098
rect 12163 7046 12175 7098
rect 12175 7046 12189 7098
rect 12213 7046 12227 7098
rect 12227 7046 12239 7098
rect 12239 7046 12269 7098
rect 12293 7046 12303 7098
rect 12303 7046 12349 7098
rect 12053 7044 12109 7046
rect 12133 7044 12189 7046
rect 12213 7044 12269 7046
rect 12293 7044 12349 7046
rect 12053 6010 12109 6012
rect 12133 6010 12189 6012
rect 12213 6010 12269 6012
rect 12293 6010 12349 6012
rect 12053 5958 12099 6010
rect 12099 5958 12109 6010
rect 12133 5958 12163 6010
rect 12163 5958 12175 6010
rect 12175 5958 12189 6010
rect 12213 5958 12227 6010
rect 12227 5958 12239 6010
rect 12239 5958 12269 6010
rect 12293 5958 12303 6010
rect 12303 5958 12349 6010
rect 12053 5956 12109 5958
rect 12133 5956 12189 5958
rect 12213 5956 12269 5958
rect 12293 5956 12349 5958
rect 9833 3290 9889 3292
rect 9913 3290 9969 3292
rect 9993 3290 10049 3292
rect 10073 3290 10129 3292
rect 9833 3238 9879 3290
rect 9879 3238 9889 3290
rect 9913 3238 9943 3290
rect 9943 3238 9955 3290
rect 9955 3238 9969 3290
rect 9993 3238 10007 3290
rect 10007 3238 10019 3290
rect 10019 3238 10049 3290
rect 10073 3238 10083 3290
rect 10083 3238 10129 3290
rect 9833 3236 9889 3238
rect 9913 3236 9969 3238
rect 9993 3236 10049 3238
rect 10073 3236 10129 3238
rect 11702 2896 11758 2952
rect 12053 4922 12109 4924
rect 12133 4922 12189 4924
rect 12213 4922 12269 4924
rect 12293 4922 12349 4924
rect 12053 4870 12099 4922
rect 12099 4870 12109 4922
rect 12133 4870 12163 4922
rect 12163 4870 12175 4922
rect 12175 4870 12189 4922
rect 12213 4870 12227 4922
rect 12227 4870 12239 4922
rect 12239 4870 12269 4922
rect 12293 4870 12303 4922
rect 12303 4870 12349 4922
rect 12053 4868 12109 4870
rect 12133 4868 12189 4870
rect 12213 4868 12269 4870
rect 12293 4868 12349 4870
rect 12053 3834 12109 3836
rect 12133 3834 12189 3836
rect 12213 3834 12269 3836
rect 12293 3834 12349 3836
rect 12053 3782 12099 3834
rect 12099 3782 12109 3834
rect 12133 3782 12163 3834
rect 12163 3782 12175 3834
rect 12175 3782 12189 3834
rect 12213 3782 12227 3834
rect 12227 3782 12239 3834
rect 12239 3782 12269 3834
rect 12293 3782 12303 3834
rect 12303 3782 12349 3834
rect 12053 3780 12109 3782
rect 12133 3780 12189 3782
rect 12213 3780 12269 3782
rect 12293 3780 12349 3782
rect 14272 6554 14328 6556
rect 14352 6554 14408 6556
rect 14432 6554 14488 6556
rect 14512 6554 14568 6556
rect 14272 6502 14318 6554
rect 14318 6502 14328 6554
rect 14352 6502 14382 6554
rect 14382 6502 14394 6554
rect 14394 6502 14408 6554
rect 14432 6502 14446 6554
rect 14446 6502 14458 6554
rect 14458 6502 14488 6554
rect 14512 6502 14522 6554
rect 14522 6502 14568 6554
rect 14272 6500 14328 6502
rect 14352 6500 14408 6502
rect 14432 6500 14488 6502
rect 14512 6500 14568 6502
rect 16492 7098 16548 7100
rect 16572 7098 16628 7100
rect 16652 7098 16708 7100
rect 16732 7098 16788 7100
rect 16492 7046 16538 7098
rect 16538 7046 16548 7098
rect 16572 7046 16602 7098
rect 16602 7046 16614 7098
rect 16614 7046 16628 7098
rect 16652 7046 16666 7098
rect 16666 7046 16678 7098
rect 16678 7046 16708 7098
rect 16732 7046 16742 7098
rect 16742 7046 16788 7098
rect 16492 7044 16548 7046
rect 16572 7044 16628 7046
rect 16652 7044 16708 7046
rect 16732 7044 16788 7046
rect 18711 6554 18767 6556
rect 18791 6554 18847 6556
rect 18871 6554 18927 6556
rect 18951 6554 19007 6556
rect 18711 6502 18757 6554
rect 18757 6502 18767 6554
rect 18791 6502 18821 6554
rect 18821 6502 18833 6554
rect 18833 6502 18847 6554
rect 18871 6502 18885 6554
rect 18885 6502 18897 6554
rect 18897 6502 18927 6554
rect 18951 6502 18961 6554
rect 18961 6502 19007 6554
rect 18711 6500 18767 6502
rect 18791 6500 18847 6502
rect 18871 6500 18927 6502
rect 18951 6500 19007 6502
rect 16492 6010 16548 6012
rect 16572 6010 16628 6012
rect 16652 6010 16708 6012
rect 16732 6010 16788 6012
rect 16492 5958 16538 6010
rect 16538 5958 16548 6010
rect 16572 5958 16602 6010
rect 16602 5958 16614 6010
rect 16614 5958 16628 6010
rect 16652 5958 16666 6010
rect 16666 5958 16678 6010
rect 16678 5958 16708 6010
rect 16732 5958 16742 6010
rect 16742 5958 16788 6010
rect 16492 5956 16548 5958
rect 16572 5956 16628 5958
rect 16652 5956 16708 5958
rect 16732 5956 16788 5958
rect 12053 2746 12109 2748
rect 12133 2746 12189 2748
rect 12213 2746 12269 2748
rect 12293 2746 12349 2748
rect 12053 2694 12099 2746
rect 12099 2694 12109 2746
rect 12133 2694 12163 2746
rect 12163 2694 12175 2746
rect 12175 2694 12189 2746
rect 12213 2694 12227 2746
rect 12227 2694 12239 2746
rect 12239 2694 12269 2746
rect 12293 2694 12303 2746
rect 12303 2694 12349 2746
rect 12053 2692 12109 2694
rect 12133 2692 12189 2694
rect 12213 2692 12269 2694
rect 12293 2692 12349 2694
rect 9833 2202 9889 2204
rect 9913 2202 9969 2204
rect 9993 2202 10049 2204
rect 10073 2202 10129 2204
rect 9833 2150 9879 2202
rect 9879 2150 9889 2202
rect 9913 2150 9943 2202
rect 9943 2150 9955 2202
rect 9955 2150 9969 2202
rect 9993 2150 10007 2202
rect 10007 2150 10019 2202
rect 10019 2150 10049 2202
rect 10073 2150 10083 2202
rect 10083 2150 10129 2202
rect 9833 2148 9889 2150
rect 9913 2148 9969 2150
rect 9993 2148 10049 2150
rect 10073 2148 10129 2150
rect 14272 5466 14328 5468
rect 14352 5466 14408 5468
rect 14432 5466 14488 5468
rect 14512 5466 14568 5468
rect 14272 5414 14318 5466
rect 14318 5414 14328 5466
rect 14352 5414 14382 5466
rect 14382 5414 14394 5466
rect 14394 5414 14408 5466
rect 14432 5414 14446 5466
rect 14446 5414 14458 5466
rect 14458 5414 14488 5466
rect 14512 5414 14522 5466
rect 14522 5414 14568 5466
rect 14272 5412 14328 5414
rect 14352 5412 14408 5414
rect 14432 5412 14488 5414
rect 14512 5412 14568 5414
rect 14272 4378 14328 4380
rect 14352 4378 14408 4380
rect 14432 4378 14488 4380
rect 14512 4378 14568 4380
rect 14272 4326 14318 4378
rect 14318 4326 14328 4378
rect 14352 4326 14382 4378
rect 14382 4326 14394 4378
rect 14394 4326 14408 4378
rect 14432 4326 14446 4378
rect 14446 4326 14458 4378
rect 14458 4326 14488 4378
rect 14512 4326 14522 4378
rect 14522 4326 14568 4378
rect 14272 4324 14328 4326
rect 14352 4324 14408 4326
rect 14432 4324 14488 4326
rect 14512 4324 14568 4326
rect 18711 5466 18767 5468
rect 18791 5466 18847 5468
rect 18871 5466 18927 5468
rect 18951 5466 19007 5468
rect 18711 5414 18757 5466
rect 18757 5414 18767 5466
rect 18791 5414 18821 5466
rect 18821 5414 18833 5466
rect 18833 5414 18847 5466
rect 18871 5414 18885 5466
rect 18885 5414 18897 5466
rect 18897 5414 18927 5466
rect 18951 5414 18961 5466
rect 18961 5414 19007 5466
rect 18711 5412 18767 5414
rect 18791 5412 18847 5414
rect 18871 5412 18927 5414
rect 18951 5412 19007 5414
rect 16492 4922 16548 4924
rect 16572 4922 16628 4924
rect 16652 4922 16708 4924
rect 16732 4922 16788 4924
rect 16492 4870 16538 4922
rect 16538 4870 16548 4922
rect 16572 4870 16602 4922
rect 16602 4870 16614 4922
rect 16614 4870 16628 4922
rect 16652 4870 16666 4922
rect 16666 4870 16678 4922
rect 16678 4870 16708 4922
rect 16732 4870 16742 4922
rect 16742 4870 16788 4922
rect 16492 4868 16548 4870
rect 16572 4868 16628 4870
rect 16652 4868 16708 4870
rect 16732 4868 16788 4870
rect 14272 3290 14328 3292
rect 14352 3290 14408 3292
rect 14432 3290 14488 3292
rect 14512 3290 14568 3292
rect 14272 3238 14318 3290
rect 14318 3238 14328 3290
rect 14352 3238 14382 3290
rect 14382 3238 14394 3290
rect 14394 3238 14408 3290
rect 14432 3238 14446 3290
rect 14446 3238 14458 3290
rect 14458 3238 14488 3290
rect 14512 3238 14522 3290
rect 14522 3238 14568 3290
rect 14272 3236 14328 3238
rect 14352 3236 14408 3238
rect 14432 3236 14488 3238
rect 14512 3236 14568 3238
rect 16492 3834 16548 3836
rect 16572 3834 16628 3836
rect 16652 3834 16708 3836
rect 16732 3834 16788 3836
rect 16492 3782 16538 3834
rect 16538 3782 16548 3834
rect 16572 3782 16602 3834
rect 16602 3782 16614 3834
rect 16614 3782 16628 3834
rect 16652 3782 16666 3834
rect 16666 3782 16678 3834
rect 16678 3782 16708 3834
rect 16732 3782 16742 3834
rect 16742 3782 16788 3834
rect 16492 3780 16548 3782
rect 16572 3780 16628 3782
rect 16652 3780 16708 3782
rect 16732 3780 16788 3782
rect 16854 2896 16910 2952
rect 16492 2746 16548 2748
rect 16572 2746 16628 2748
rect 16652 2746 16708 2748
rect 16732 2746 16788 2748
rect 16492 2694 16538 2746
rect 16538 2694 16548 2746
rect 16572 2694 16602 2746
rect 16602 2694 16614 2746
rect 16614 2694 16628 2746
rect 16652 2694 16666 2746
rect 16666 2694 16678 2746
rect 16678 2694 16708 2746
rect 16732 2694 16742 2746
rect 16742 2694 16788 2746
rect 16492 2692 16548 2694
rect 16572 2692 16628 2694
rect 16652 2692 16708 2694
rect 16732 2692 16788 2694
rect 18711 4378 18767 4380
rect 18791 4378 18847 4380
rect 18871 4378 18927 4380
rect 18951 4378 19007 4380
rect 18711 4326 18757 4378
rect 18757 4326 18767 4378
rect 18791 4326 18821 4378
rect 18821 4326 18833 4378
rect 18833 4326 18847 4378
rect 18871 4326 18885 4378
rect 18885 4326 18897 4378
rect 18897 4326 18927 4378
rect 18951 4326 18961 4378
rect 18961 4326 19007 4378
rect 18711 4324 18767 4326
rect 18791 4324 18847 4326
rect 18871 4324 18927 4326
rect 18951 4324 19007 4326
rect 18711 3290 18767 3292
rect 18791 3290 18847 3292
rect 18871 3290 18927 3292
rect 18951 3290 19007 3292
rect 18711 3238 18757 3290
rect 18757 3238 18767 3290
rect 18791 3238 18821 3290
rect 18821 3238 18833 3290
rect 18833 3238 18847 3290
rect 18871 3238 18885 3290
rect 18885 3238 18897 3290
rect 18897 3238 18927 3290
rect 18951 3238 18961 3290
rect 18961 3238 19007 3290
rect 18711 3236 18767 3238
rect 18791 3236 18847 3238
rect 18871 3236 18927 3238
rect 18951 3236 19007 3238
rect 14272 2202 14328 2204
rect 14352 2202 14408 2204
rect 14432 2202 14488 2204
rect 14512 2202 14568 2204
rect 14272 2150 14318 2202
rect 14318 2150 14328 2202
rect 14352 2150 14382 2202
rect 14382 2150 14394 2202
rect 14394 2150 14408 2202
rect 14432 2150 14446 2202
rect 14446 2150 14458 2202
rect 14458 2150 14488 2202
rect 14512 2150 14522 2202
rect 14522 2150 14568 2202
rect 14272 2148 14328 2150
rect 14352 2148 14408 2150
rect 14432 2148 14488 2150
rect 14512 2148 14568 2150
rect 18711 2202 18767 2204
rect 18791 2202 18847 2204
rect 18871 2202 18927 2204
rect 18951 2202 19007 2204
rect 18711 2150 18757 2202
rect 18757 2150 18767 2202
rect 18791 2150 18821 2202
rect 18821 2150 18833 2202
rect 18833 2150 18847 2202
rect 18871 2150 18885 2202
rect 18885 2150 18897 2202
rect 18897 2150 18927 2202
rect 18951 2150 18961 2202
rect 18961 2150 19007 2202
rect 18711 2148 18767 2150
rect 18791 2148 18847 2150
rect 18871 2148 18927 2150
rect 18951 2148 19007 2150
<< metal3 >>
rect 5384 7648 5700 7649
rect 5384 7584 5390 7648
rect 5454 7584 5470 7648
rect 5534 7584 5550 7648
rect 5614 7584 5630 7648
rect 5694 7584 5700 7648
rect 5384 7583 5700 7584
rect 9823 7648 10139 7649
rect 9823 7584 9829 7648
rect 9893 7584 9909 7648
rect 9973 7584 9989 7648
rect 10053 7584 10069 7648
rect 10133 7584 10139 7648
rect 9823 7583 10139 7584
rect 14262 7648 14578 7649
rect 14262 7584 14268 7648
rect 14332 7584 14348 7648
rect 14412 7584 14428 7648
rect 14492 7584 14508 7648
rect 14572 7584 14578 7648
rect 14262 7583 14578 7584
rect 18701 7648 19017 7649
rect 18701 7584 18707 7648
rect 18771 7584 18787 7648
rect 18851 7584 18867 7648
rect 18931 7584 18947 7648
rect 19011 7584 19017 7648
rect 18701 7583 19017 7584
rect 3165 7104 3481 7105
rect 3165 7040 3171 7104
rect 3235 7040 3251 7104
rect 3315 7040 3331 7104
rect 3395 7040 3411 7104
rect 3475 7040 3481 7104
rect 3165 7039 3481 7040
rect 7604 7104 7920 7105
rect 7604 7040 7610 7104
rect 7674 7040 7690 7104
rect 7754 7040 7770 7104
rect 7834 7040 7850 7104
rect 7914 7040 7920 7104
rect 7604 7039 7920 7040
rect 12043 7104 12359 7105
rect 12043 7040 12049 7104
rect 12113 7040 12129 7104
rect 12193 7040 12209 7104
rect 12273 7040 12289 7104
rect 12353 7040 12359 7104
rect 12043 7039 12359 7040
rect 16482 7104 16798 7105
rect 16482 7040 16488 7104
rect 16552 7040 16568 7104
rect 16632 7040 16648 7104
rect 16712 7040 16728 7104
rect 16792 7040 16798 7104
rect 16482 7039 16798 7040
rect 5384 6560 5700 6561
rect 5384 6496 5390 6560
rect 5454 6496 5470 6560
rect 5534 6496 5550 6560
rect 5614 6496 5630 6560
rect 5694 6496 5700 6560
rect 5384 6495 5700 6496
rect 9823 6560 10139 6561
rect 9823 6496 9829 6560
rect 9893 6496 9909 6560
rect 9973 6496 9989 6560
rect 10053 6496 10069 6560
rect 10133 6496 10139 6560
rect 9823 6495 10139 6496
rect 14262 6560 14578 6561
rect 14262 6496 14268 6560
rect 14332 6496 14348 6560
rect 14412 6496 14428 6560
rect 14492 6496 14508 6560
rect 14572 6496 14578 6560
rect 14262 6495 14578 6496
rect 18701 6560 19017 6561
rect 18701 6496 18707 6560
rect 18771 6496 18787 6560
rect 18851 6496 18867 6560
rect 18931 6496 18947 6560
rect 19011 6496 19017 6560
rect 18701 6495 19017 6496
rect 3165 6016 3481 6017
rect 3165 5952 3171 6016
rect 3235 5952 3251 6016
rect 3315 5952 3331 6016
rect 3395 5952 3411 6016
rect 3475 5952 3481 6016
rect 3165 5951 3481 5952
rect 7604 6016 7920 6017
rect 7604 5952 7610 6016
rect 7674 5952 7690 6016
rect 7754 5952 7770 6016
rect 7834 5952 7850 6016
rect 7914 5952 7920 6016
rect 7604 5951 7920 5952
rect 12043 6016 12359 6017
rect 12043 5952 12049 6016
rect 12113 5952 12129 6016
rect 12193 5952 12209 6016
rect 12273 5952 12289 6016
rect 12353 5952 12359 6016
rect 12043 5951 12359 5952
rect 16482 6016 16798 6017
rect 16482 5952 16488 6016
rect 16552 5952 16568 6016
rect 16632 5952 16648 6016
rect 16712 5952 16728 6016
rect 16792 5952 16798 6016
rect 16482 5951 16798 5952
rect 5384 5472 5700 5473
rect 5384 5408 5390 5472
rect 5454 5408 5470 5472
rect 5534 5408 5550 5472
rect 5614 5408 5630 5472
rect 5694 5408 5700 5472
rect 5384 5407 5700 5408
rect 9823 5472 10139 5473
rect 9823 5408 9829 5472
rect 9893 5408 9909 5472
rect 9973 5408 9989 5472
rect 10053 5408 10069 5472
rect 10133 5408 10139 5472
rect 9823 5407 10139 5408
rect 14262 5472 14578 5473
rect 14262 5408 14268 5472
rect 14332 5408 14348 5472
rect 14412 5408 14428 5472
rect 14492 5408 14508 5472
rect 14572 5408 14578 5472
rect 14262 5407 14578 5408
rect 18701 5472 19017 5473
rect 18701 5408 18707 5472
rect 18771 5408 18787 5472
rect 18851 5408 18867 5472
rect 18931 5408 18947 5472
rect 19011 5408 19017 5472
rect 18701 5407 19017 5408
rect 3165 4928 3481 4929
rect 3165 4864 3171 4928
rect 3235 4864 3251 4928
rect 3315 4864 3331 4928
rect 3395 4864 3411 4928
rect 3475 4864 3481 4928
rect 3165 4863 3481 4864
rect 7604 4928 7920 4929
rect 7604 4864 7610 4928
rect 7674 4864 7690 4928
rect 7754 4864 7770 4928
rect 7834 4864 7850 4928
rect 7914 4864 7920 4928
rect 7604 4863 7920 4864
rect 12043 4928 12359 4929
rect 12043 4864 12049 4928
rect 12113 4864 12129 4928
rect 12193 4864 12209 4928
rect 12273 4864 12289 4928
rect 12353 4864 12359 4928
rect 12043 4863 12359 4864
rect 16482 4928 16798 4929
rect 16482 4864 16488 4928
rect 16552 4864 16568 4928
rect 16632 4864 16648 4928
rect 16712 4864 16728 4928
rect 16792 4864 16798 4928
rect 16482 4863 16798 4864
rect 4337 4722 4403 4725
rect 6269 4722 6335 4725
rect 7281 4722 7347 4725
rect 4337 4720 7347 4722
rect 4337 4664 4342 4720
rect 4398 4664 6274 4720
rect 6330 4664 7286 4720
rect 7342 4664 7347 4720
rect 4337 4662 7347 4664
rect 4337 4659 4403 4662
rect 6269 4659 6335 4662
rect 7281 4659 7347 4662
rect 5073 4586 5139 4589
rect 6085 4586 6151 4589
rect 5073 4584 6151 4586
rect 5073 4528 5078 4584
rect 5134 4528 6090 4584
rect 6146 4528 6151 4584
rect 5073 4526 6151 4528
rect 5073 4523 5139 4526
rect 6085 4523 6151 4526
rect 5384 4384 5700 4385
rect 5384 4320 5390 4384
rect 5454 4320 5470 4384
rect 5534 4320 5550 4384
rect 5614 4320 5630 4384
rect 5694 4320 5700 4384
rect 5384 4319 5700 4320
rect 9823 4384 10139 4385
rect 9823 4320 9829 4384
rect 9893 4320 9909 4384
rect 9973 4320 9989 4384
rect 10053 4320 10069 4384
rect 10133 4320 10139 4384
rect 9823 4319 10139 4320
rect 14262 4384 14578 4385
rect 14262 4320 14268 4384
rect 14332 4320 14348 4384
rect 14412 4320 14428 4384
rect 14492 4320 14508 4384
rect 14572 4320 14578 4384
rect 14262 4319 14578 4320
rect 18701 4384 19017 4385
rect 18701 4320 18707 4384
rect 18771 4320 18787 4384
rect 18851 4320 18867 4384
rect 18931 4320 18947 4384
rect 19011 4320 19017 4384
rect 18701 4319 19017 4320
rect 7189 4178 7255 4181
rect 9305 4178 9371 4181
rect 7189 4176 9371 4178
rect 7189 4120 7194 4176
rect 7250 4120 9310 4176
rect 9366 4120 9371 4176
rect 7189 4118 9371 4120
rect 7189 4115 7255 4118
rect 9305 4115 9371 4118
rect 3165 3840 3481 3841
rect 3165 3776 3171 3840
rect 3235 3776 3251 3840
rect 3315 3776 3331 3840
rect 3395 3776 3411 3840
rect 3475 3776 3481 3840
rect 3165 3775 3481 3776
rect 7604 3840 7920 3841
rect 7604 3776 7610 3840
rect 7674 3776 7690 3840
rect 7754 3776 7770 3840
rect 7834 3776 7850 3840
rect 7914 3776 7920 3840
rect 7604 3775 7920 3776
rect 12043 3840 12359 3841
rect 12043 3776 12049 3840
rect 12113 3776 12129 3840
rect 12193 3776 12209 3840
rect 12273 3776 12289 3840
rect 12353 3776 12359 3840
rect 12043 3775 12359 3776
rect 16482 3840 16798 3841
rect 16482 3776 16488 3840
rect 16552 3776 16568 3840
rect 16632 3776 16648 3840
rect 16712 3776 16728 3840
rect 16792 3776 16798 3840
rect 16482 3775 16798 3776
rect 5384 3296 5700 3297
rect 5384 3232 5390 3296
rect 5454 3232 5470 3296
rect 5534 3232 5550 3296
rect 5614 3232 5630 3296
rect 5694 3232 5700 3296
rect 5384 3231 5700 3232
rect 9823 3296 10139 3297
rect 9823 3232 9829 3296
rect 9893 3232 9909 3296
rect 9973 3232 9989 3296
rect 10053 3232 10069 3296
rect 10133 3232 10139 3296
rect 9823 3231 10139 3232
rect 14262 3296 14578 3297
rect 14262 3232 14268 3296
rect 14332 3232 14348 3296
rect 14412 3232 14428 3296
rect 14492 3232 14508 3296
rect 14572 3232 14578 3296
rect 14262 3231 14578 3232
rect 18701 3296 19017 3297
rect 18701 3232 18707 3296
rect 18771 3232 18787 3296
rect 18851 3232 18867 3296
rect 18931 3232 18947 3296
rect 19011 3232 19017 3296
rect 18701 3231 19017 3232
rect 11697 2954 11763 2957
rect 16849 2954 16915 2957
rect 11697 2952 16915 2954
rect 11697 2896 11702 2952
rect 11758 2896 16854 2952
rect 16910 2896 16915 2952
rect 11697 2894 16915 2896
rect 11697 2891 11763 2894
rect 16849 2891 16915 2894
rect 3165 2752 3481 2753
rect 3165 2688 3171 2752
rect 3235 2688 3251 2752
rect 3315 2688 3331 2752
rect 3395 2688 3411 2752
rect 3475 2688 3481 2752
rect 3165 2687 3481 2688
rect 7604 2752 7920 2753
rect 7604 2688 7610 2752
rect 7674 2688 7690 2752
rect 7754 2688 7770 2752
rect 7834 2688 7850 2752
rect 7914 2688 7920 2752
rect 7604 2687 7920 2688
rect 12043 2752 12359 2753
rect 12043 2688 12049 2752
rect 12113 2688 12129 2752
rect 12193 2688 12209 2752
rect 12273 2688 12289 2752
rect 12353 2688 12359 2752
rect 12043 2687 12359 2688
rect 16482 2752 16798 2753
rect 16482 2688 16488 2752
rect 16552 2688 16568 2752
rect 16632 2688 16648 2752
rect 16712 2688 16728 2752
rect 16792 2688 16798 2752
rect 16482 2687 16798 2688
rect 5384 2208 5700 2209
rect 5384 2144 5390 2208
rect 5454 2144 5470 2208
rect 5534 2144 5550 2208
rect 5614 2144 5630 2208
rect 5694 2144 5700 2208
rect 5384 2143 5700 2144
rect 9823 2208 10139 2209
rect 9823 2144 9829 2208
rect 9893 2144 9909 2208
rect 9973 2144 9989 2208
rect 10053 2144 10069 2208
rect 10133 2144 10139 2208
rect 9823 2143 10139 2144
rect 14262 2208 14578 2209
rect 14262 2144 14268 2208
rect 14332 2144 14348 2208
rect 14412 2144 14428 2208
rect 14492 2144 14508 2208
rect 14572 2144 14578 2208
rect 14262 2143 14578 2144
rect 18701 2208 19017 2209
rect 18701 2144 18707 2208
rect 18771 2144 18787 2208
rect 18851 2144 18867 2208
rect 18931 2144 18947 2208
rect 19011 2144 19017 2208
rect 18701 2143 19017 2144
<< via3 >>
rect 5390 7644 5454 7648
rect 5390 7588 5394 7644
rect 5394 7588 5450 7644
rect 5450 7588 5454 7644
rect 5390 7584 5454 7588
rect 5470 7644 5534 7648
rect 5470 7588 5474 7644
rect 5474 7588 5530 7644
rect 5530 7588 5534 7644
rect 5470 7584 5534 7588
rect 5550 7644 5614 7648
rect 5550 7588 5554 7644
rect 5554 7588 5610 7644
rect 5610 7588 5614 7644
rect 5550 7584 5614 7588
rect 5630 7644 5694 7648
rect 5630 7588 5634 7644
rect 5634 7588 5690 7644
rect 5690 7588 5694 7644
rect 5630 7584 5694 7588
rect 9829 7644 9893 7648
rect 9829 7588 9833 7644
rect 9833 7588 9889 7644
rect 9889 7588 9893 7644
rect 9829 7584 9893 7588
rect 9909 7644 9973 7648
rect 9909 7588 9913 7644
rect 9913 7588 9969 7644
rect 9969 7588 9973 7644
rect 9909 7584 9973 7588
rect 9989 7644 10053 7648
rect 9989 7588 9993 7644
rect 9993 7588 10049 7644
rect 10049 7588 10053 7644
rect 9989 7584 10053 7588
rect 10069 7644 10133 7648
rect 10069 7588 10073 7644
rect 10073 7588 10129 7644
rect 10129 7588 10133 7644
rect 10069 7584 10133 7588
rect 14268 7644 14332 7648
rect 14268 7588 14272 7644
rect 14272 7588 14328 7644
rect 14328 7588 14332 7644
rect 14268 7584 14332 7588
rect 14348 7644 14412 7648
rect 14348 7588 14352 7644
rect 14352 7588 14408 7644
rect 14408 7588 14412 7644
rect 14348 7584 14412 7588
rect 14428 7644 14492 7648
rect 14428 7588 14432 7644
rect 14432 7588 14488 7644
rect 14488 7588 14492 7644
rect 14428 7584 14492 7588
rect 14508 7644 14572 7648
rect 14508 7588 14512 7644
rect 14512 7588 14568 7644
rect 14568 7588 14572 7644
rect 14508 7584 14572 7588
rect 18707 7644 18771 7648
rect 18707 7588 18711 7644
rect 18711 7588 18767 7644
rect 18767 7588 18771 7644
rect 18707 7584 18771 7588
rect 18787 7644 18851 7648
rect 18787 7588 18791 7644
rect 18791 7588 18847 7644
rect 18847 7588 18851 7644
rect 18787 7584 18851 7588
rect 18867 7644 18931 7648
rect 18867 7588 18871 7644
rect 18871 7588 18927 7644
rect 18927 7588 18931 7644
rect 18867 7584 18931 7588
rect 18947 7644 19011 7648
rect 18947 7588 18951 7644
rect 18951 7588 19007 7644
rect 19007 7588 19011 7644
rect 18947 7584 19011 7588
rect 3171 7100 3235 7104
rect 3171 7044 3175 7100
rect 3175 7044 3231 7100
rect 3231 7044 3235 7100
rect 3171 7040 3235 7044
rect 3251 7100 3315 7104
rect 3251 7044 3255 7100
rect 3255 7044 3311 7100
rect 3311 7044 3315 7100
rect 3251 7040 3315 7044
rect 3331 7100 3395 7104
rect 3331 7044 3335 7100
rect 3335 7044 3391 7100
rect 3391 7044 3395 7100
rect 3331 7040 3395 7044
rect 3411 7100 3475 7104
rect 3411 7044 3415 7100
rect 3415 7044 3471 7100
rect 3471 7044 3475 7100
rect 3411 7040 3475 7044
rect 7610 7100 7674 7104
rect 7610 7044 7614 7100
rect 7614 7044 7670 7100
rect 7670 7044 7674 7100
rect 7610 7040 7674 7044
rect 7690 7100 7754 7104
rect 7690 7044 7694 7100
rect 7694 7044 7750 7100
rect 7750 7044 7754 7100
rect 7690 7040 7754 7044
rect 7770 7100 7834 7104
rect 7770 7044 7774 7100
rect 7774 7044 7830 7100
rect 7830 7044 7834 7100
rect 7770 7040 7834 7044
rect 7850 7100 7914 7104
rect 7850 7044 7854 7100
rect 7854 7044 7910 7100
rect 7910 7044 7914 7100
rect 7850 7040 7914 7044
rect 12049 7100 12113 7104
rect 12049 7044 12053 7100
rect 12053 7044 12109 7100
rect 12109 7044 12113 7100
rect 12049 7040 12113 7044
rect 12129 7100 12193 7104
rect 12129 7044 12133 7100
rect 12133 7044 12189 7100
rect 12189 7044 12193 7100
rect 12129 7040 12193 7044
rect 12209 7100 12273 7104
rect 12209 7044 12213 7100
rect 12213 7044 12269 7100
rect 12269 7044 12273 7100
rect 12209 7040 12273 7044
rect 12289 7100 12353 7104
rect 12289 7044 12293 7100
rect 12293 7044 12349 7100
rect 12349 7044 12353 7100
rect 12289 7040 12353 7044
rect 16488 7100 16552 7104
rect 16488 7044 16492 7100
rect 16492 7044 16548 7100
rect 16548 7044 16552 7100
rect 16488 7040 16552 7044
rect 16568 7100 16632 7104
rect 16568 7044 16572 7100
rect 16572 7044 16628 7100
rect 16628 7044 16632 7100
rect 16568 7040 16632 7044
rect 16648 7100 16712 7104
rect 16648 7044 16652 7100
rect 16652 7044 16708 7100
rect 16708 7044 16712 7100
rect 16648 7040 16712 7044
rect 16728 7100 16792 7104
rect 16728 7044 16732 7100
rect 16732 7044 16788 7100
rect 16788 7044 16792 7100
rect 16728 7040 16792 7044
rect 5390 6556 5454 6560
rect 5390 6500 5394 6556
rect 5394 6500 5450 6556
rect 5450 6500 5454 6556
rect 5390 6496 5454 6500
rect 5470 6556 5534 6560
rect 5470 6500 5474 6556
rect 5474 6500 5530 6556
rect 5530 6500 5534 6556
rect 5470 6496 5534 6500
rect 5550 6556 5614 6560
rect 5550 6500 5554 6556
rect 5554 6500 5610 6556
rect 5610 6500 5614 6556
rect 5550 6496 5614 6500
rect 5630 6556 5694 6560
rect 5630 6500 5634 6556
rect 5634 6500 5690 6556
rect 5690 6500 5694 6556
rect 5630 6496 5694 6500
rect 9829 6556 9893 6560
rect 9829 6500 9833 6556
rect 9833 6500 9889 6556
rect 9889 6500 9893 6556
rect 9829 6496 9893 6500
rect 9909 6556 9973 6560
rect 9909 6500 9913 6556
rect 9913 6500 9969 6556
rect 9969 6500 9973 6556
rect 9909 6496 9973 6500
rect 9989 6556 10053 6560
rect 9989 6500 9993 6556
rect 9993 6500 10049 6556
rect 10049 6500 10053 6556
rect 9989 6496 10053 6500
rect 10069 6556 10133 6560
rect 10069 6500 10073 6556
rect 10073 6500 10129 6556
rect 10129 6500 10133 6556
rect 10069 6496 10133 6500
rect 14268 6556 14332 6560
rect 14268 6500 14272 6556
rect 14272 6500 14328 6556
rect 14328 6500 14332 6556
rect 14268 6496 14332 6500
rect 14348 6556 14412 6560
rect 14348 6500 14352 6556
rect 14352 6500 14408 6556
rect 14408 6500 14412 6556
rect 14348 6496 14412 6500
rect 14428 6556 14492 6560
rect 14428 6500 14432 6556
rect 14432 6500 14488 6556
rect 14488 6500 14492 6556
rect 14428 6496 14492 6500
rect 14508 6556 14572 6560
rect 14508 6500 14512 6556
rect 14512 6500 14568 6556
rect 14568 6500 14572 6556
rect 14508 6496 14572 6500
rect 18707 6556 18771 6560
rect 18707 6500 18711 6556
rect 18711 6500 18767 6556
rect 18767 6500 18771 6556
rect 18707 6496 18771 6500
rect 18787 6556 18851 6560
rect 18787 6500 18791 6556
rect 18791 6500 18847 6556
rect 18847 6500 18851 6556
rect 18787 6496 18851 6500
rect 18867 6556 18931 6560
rect 18867 6500 18871 6556
rect 18871 6500 18927 6556
rect 18927 6500 18931 6556
rect 18867 6496 18931 6500
rect 18947 6556 19011 6560
rect 18947 6500 18951 6556
rect 18951 6500 19007 6556
rect 19007 6500 19011 6556
rect 18947 6496 19011 6500
rect 3171 6012 3235 6016
rect 3171 5956 3175 6012
rect 3175 5956 3231 6012
rect 3231 5956 3235 6012
rect 3171 5952 3235 5956
rect 3251 6012 3315 6016
rect 3251 5956 3255 6012
rect 3255 5956 3311 6012
rect 3311 5956 3315 6012
rect 3251 5952 3315 5956
rect 3331 6012 3395 6016
rect 3331 5956 3335 6012
rect 3335 5956 3391 6012
rect 3391 5956 3395 6012
rect 3331 5952 3395 5956
rect 3411 6012 3475 6016
rect 3411 5956 3415 6012
rect 3415 5956 3471 6012
rect 3471 5956 3475 6012
rect 3411 5952 3475 5956
rect 7610 6012 7674 6016
rect 7610 5956 7614 6012
rect 7614 5956 7670 6012
rect 7670 5956 7674 6012
rect 7610 5952 7674 5956
rect 7690 6012 7754 6016
rect 7690 5956 7694 6012
rect 7694 5956 7750 6012
rect 7750 5956 7754 6012
rect 7690 5952 7754 5956
rect 7770 6012 7834 6016
rect 7770 5956 7774 6012
rect 7774 5956 7830 6012
rect 7830 5956 7834 6012
rect 7770 5952 7834 5956
rect 7850 6012 7914 6016
rect 7850 5956 7854 6012
rect 7854 5956 7910 6012
rect 7910 5956 7914 6012
rect 7850 5952 7914 5956
rect 12049 6012 12113 6016
rect 12049 5956 12053 6012
rect 12053 5956 12109 6012
rect 12109 5956 12113 6012
rect 12049 5952 12113 5956
rect 12129 6012 12193 6016
rect 12129 5956 12133 6012
rect 12133 5956 12189 6012
rect 12189 5956 12193 6012
rect 12129 5952 12193 5956
rect 12209 6012 12273 6016
rect 12209 5956 12213 6012
rect 12213 5956 12269 6012
rect 12269 5956 12273 6012
rect 12209 5952 12273 5956
rect 12289 6012 12353 6016
rect 12289 5956 12293 6012
rect 12293 5956 12349 6012
rect 12349 5956 12353 6012
rect 12289 5952 12353 5956
rect 16488 6012 16552 6016
rect 16488 5956 16492 6012
rect 16492 5956 16548 6012
rect 16548 5956 16552 6012
rect 16488 5952 16552 5956
rect 16568 6012 16632 6016
rect 16568 5956 16572 6012
rect 16572 5956 16628 6012
rect 16628 5956 16632 6012
rect 16568 5952 16632 5956
rect 16648 6012 16712 6016
rect 16648 5956 16652 6012
rect 16652 5956 16708 6012
rect 16708 5956 16712 6012
rect 16648 5952 16712 5956
rect 16728 6012 16792 6016
rect 16728 5956 16732 6012
rect 16732 5956 16788 6012
rect 16788 5956 16792 6012
rect 16728 5952 16792 5956
rect 5390 5468 5454 5472
rect 5390 5412 5394 5468
rect 5394 5412 5450 5468
rect 5450 5412 5454 5468
rect 5390 5408 5454 5412
rect 5470 5468 5534 5472
rect 5470 5412 5474 5468
rect 5474 5412 5530 5468
rect 5530 5412 5534 5468
rect 5470 5408 5534 5412
rect 5550 5468 5614 5472
rect 5550 5412 5554 5468
rect 5554 5412 5610 5468
rect 5610 5412 5614 5468
rect 5550 5408 5614 5412
rect 5630 5468 5694 5472
rect 5630 5412 5634 5468
rect 5634 5412 5690 5468
rect 5690 5412 5694 5468
rect 5630 5408 5694 5412
rect 9829 5468 9893 5472
rect 9829 5412 9833 5468
rect 9833 5412 9889 5468
rect 9889 5412 9893 5468
rect 9829 5408 9893 5412
rect 9909 5468 9973 5472
rect 9909 5412 9913 5468
rect 9913 5412 9969 5468
rect 9969 5412 9973 5468
rect 9909 5408 9973 5412
rect 9989 5468 10053 5472
rect 9989 5412 9993 5468
rect 9993 5412 10049 5468
rect 10049 5412 10053 5468
rect 9989 5408 10053 5412
rect 10069 5468 10133 5472
rect 10069 5412 10073 5468
rect 10073 5412 10129 5468
rect 10129 5412 10133 5468
rect 10069 5408 10133 5412
rect 14268 5468 14332 5472
rect 14268 5412 14272 5468
rect 14272 5412 14328 5468
rect 14328 5412 14332 5468
rect 14268 5408 14332 5412
rect 14348 5468 14412 5472
rect 14348 5412 14352 5468
rect 14352 5412 14408 5468
rect 14408 5412 14412 5468
rect 14348 5408 14412 5412
rect 14428 5468 14492 5472
rect 14428 5412 14432 5468
rect 14432 5412 14488 5468
rect 14488 5412 14492 5468
rect 14428 5408 14492 5412
rect 14508 5468 14572 5472
rect 14508 5412 14512 5468
rect 14512 5412 14568 5468
rect 14568 5412 14572 5468
rect 14508 5408 14572 5412
rect 18707 5468 18771 5472
rect 18707 5412 18711 5468
rect 18711 5412 18767 5468
rect 18767 5412 18771 5468
rect 18707 5408 18771 5412
rect 18787 5468 18851 5472
rect 18787 5412 18791 5468
rect 18791 5412 18847 5468
rect 18847 5412 18851 5468
rect 18787 5408 18851 5412
rect 18867 5468 18931 5472
rect 18867 5412 18871 5468
rect 18871 5412 18927 5468
rect 18927 5412 18931 5468
rect 18867 5408 18931 5412
rect 18947 5468 19011 5472
rect 18947 5412 18951 5468
rect 18951 5412 19007 5468
rect 19007 5412 19011 5468
rect 18947 5408 19011 5412
rect 3171 4924 3235 4928
rect 3171 4868 3175 4924
rect 3175 4868 3231 4924
rect 3231 4868 3235 4924
rect 3171 4864 3235 4868
rect 3251 4924 3315 4928
rect 3251 4868 3255 4924
rect 3255 4868 3311 4924
rect 3311 4868 3315 4924
rect 3251 4864 3315 4868
rect 3331 4924 3395 4928
rect 3331 4868 3335 4924
rect 3335 4868 3391 4924
rect 3391 4868 3395 4924
rect 3331 4864 3395 4868
rect 3411 4924 3475 4928
rect 3411 4868 3415 4924
rect 3415 4868 3471 4924
rect 3471 4868 3475 4924
rect 3411 4864 3475 4868
rect 7610 4924 7674 4928
rect 7610 4868 7614 4924
rect 7614 4868 7670 4924
rect 7670 4868 7674 4924
rect 7610 4864 7674 4868
rect 7690 4924 7754 4928
rect 7690 4868 7694 4924
rect 7694 4868 7750 4924
rect 7750 4868 7754 4924
rect 7690 4864 7754 4868
rect 7770 4924 7834 4928
rect 7770 4868 7774 4924
rect 7774 4868 7830 4924
rect 7830 4868 7834 4924
rect 7770 4864 7834 4868
rect 7850 4924 7914 4928
rect 7850 4868 7854 4924
rect 7854 4868 7910 4924
rect 7910 4868 7914 4924
rect 7850 4864 7914 4868
rect 12049 4924 12113 4928
rect 12049 4868 12053 4924
rect 12053 4868 12109 4924
rect 12109 4868 12113 4924
rect 12049 4864 12113 4868
rect 12129 4924 12193 4928
rect 12129 4868 12133 4924
rect 12133 4868 12189 4924
rect 12189 4868 12193 4924
rect 12129 4864 12193 4868
rect 12209 4924 12273 4928
rect 12209 4868 12213 4924
rect 12213 4868 12269 4924
rect 12269 4868 12273 4924
rect 12209 4864 12273 4868
rect 12289 4924 12353 4928
rect 12289 4868 12293 4924
rect 12293 4868 12349 4924
rect 12349 4868 12353 4924
rect 12289 4864 12353 4868
rect 16488 4924 16552 4928
rect 16488 4868 16492 4924
rect 16492 4868 16548 4924
rect 16548 4868 16552 4924
rect 16488 4864 16552 4868
rect 16568 4924 16632 4928
rect 16568 4868 16572 4924
rect 16572 4868 16628 4924
rect 16628 4868 16632 4924
rect 16568 4864 16632 4868
rect 16648 4924 16712 4928
rect 16648 4868 16652 4924
rect 16652 4868 16708 4924
rect 16708 4868 16712 4924
rect 16648 4864 16712 4868
rect 16728 4924 16792 4928
rect 16728 4868 16732 4924
rect 16732 4868 16788 4924
rect 16788 4868 16792 4924
rect 16728 4864 16792 4868
rect 5390 4380 5454 4384
rect 5390 4324 5394 4380
rect 5394 4324 5450 4380
rect 5450 4324 5454 4380
rect 5390 4320 5454 4324
rect 5470 4380 5534 4384
rect 5470 4324 5474 4380
rect 5474 4324 5530 4380
rect 5530 4324 5534 4380
rect 5470 4320 5534 4324
rect 5550 4380 5614 4384
rect 5550 4324 5554 4380
rect 5554 4324 5610 4380
rect 5610 4324 5614 4380
rect 5550 4320 5614 4324
rect 5630 4380 5694 4384
rect 5630 4324 5634 4380
rect 5634 4324 5690 4380
rect 5690 4324 5694 4380
rect 5630 4320 5694 4324
rect 9829 4380 9893 4384
rect 9829 4324 9833 4380
rect 9833 4324 9889 4380
rect 9889 4324 9893 4380
rect 9829 4320 9893 4324
rect 9909 4380 9973 4384
rect 9909 4324 9913 4380
rect 9913 4324 9969 4380
rect 9969 4324 9973 4380
rect 9909 4320 9973 4324
rect 9989 4380 10053 4384
rect 9989 4324 9993 4380
rect 9993 4324 10049 4380
rect 10049 4324 10053 4380
rect 9989 4320 10053 4324
rect 10069 4380 10133 4384
rect 10069 4324 10073 4380
rect 10073 4324 10129 4380
rect 10129 4324 10133 4380
rect 10069 4320 10133 4324
rect 14268 4380 14332 4384
rect 14268 4324 14272 4380
rect 14272 4324 14328 4380
rect 14328 4324 14332 4380
rect 14268 4320 14332 4324
rect 14348 4380 14412 4384
rect 14348 4324 14352 4380
rect 14352 4324 14408 4380
rect 14408 4324 14412 4380
rect 14348 4320 14412 4324
rect 14428 4380 14492 4384
rect 14428 4324 14432 4380
rect 14432 4324 14488 4380
rect 14488 4324 14492 4380
rect 14428 4320 14492 4324
rect 14508 4380 14572 4384
rect 14508 4324 14512 4380
rect 14512 4324 14568 4380
rect 14568 4324 14572 4380
rect 14508 4320 14572 4324
rect 18707 4380 18771 4384
rect 18707 4324 18711 4380
rect 18711 4324 18767 4380
rect 18767 4324 18771 4380
rect 18707 4320 18771 4324
rect 18787 4380 18851 4384
rect 18787 4324 18791 4380
rect 18791 4324 18847 4380
rect 18847 4324 18851 4380
rect 18787 4320 18851 4324
rect 18867 4380 18931 4384
rect 18867 4324 18871 4380
rect 18871 4324 18927 4380
rect 18927 4324 18931 4380
rect 18867 4320 18931 4324
rect 18947 4380 19011 4384
rect 18947 4324 18951 4380
rect 18951 4324 19007 4380
rect 19007 4324 19011 4380
rect 18947 4320 19011 4324
rect 3171 3836 3235 3840
rect 3171 3780 3175 3836
rect 3175 3780 3231 3836
rect 3231 3780 3235 3836
rect 3171 3776 3235 3780
rect 3251 3836 3315 3840
rect 3251 3780 3255 3836
rect 3255 3780 3311 3836
rect 3311 3780 3315 3836
rect 3251 3776 3315 3780
rect 3331 3836 3395 3840
rect 3331 3780 3335 3836
rect 3335 3780 3391 3836
rect 3391 3780 3395 3836
rect 3331 3776 3395 3780
rect 3411 3836 3475 3840
rect 3411 3780 3415 3836
rect 3415 3780 3471 3836
rect 3471 3780 3475 3836
rect 3411 3776 3475 3780
rect 7610 3836 7674 3840
rect 7610 3780 7614 3836
rect 7614 3780 7670 3836
rect 7670 3780 7674 3836
rect 7610 3776 7674 3780
rect 7690 3836 7754 3840
rect 7690 3780 7694 3836
rect 7694 3780 7750 3836
rect 7750 3780 7754 3836
rect 7690 3776 7754 3780
rect 7770 3836 7834 3840
rect 7770 3780 7774 3836
rect 7774 3780 7830 3836
rect 7830 3780 7834 3836
rect 7770 3776 7834 3780
rect 7850 3836 7914 3840
rect 7850 3780 7854 3836
rect 7854 3780 7910 3836
rect 7910 3780 7914 3836
rect 7850 3776 7914 3780
rect 12049 3836 12113 3840
rect 12049 3780 12053 3836
rect 12053 3780 12109 3836
rect 12109 3780 12113 3836
rect 12049 3776 12113 3780
rect 12129 3836 12193 3840
rect 12129 3780 12133 3836
rect 12133 3780 12189 3836
rect 12189 3780 12193 3836
rect 12129 3776 12193 3780
rect 12209 3836 12273 3840
rect 12209 3780 12213 3836
rect 12213 3780 12269 3836
rect 12269 3780 12273 3836
rect 12209 3776 12273 3780
rect 12289 3836 12353 3840
rect 12289 3780 12293 3836
rect 12293 3780 12349 3836
rect 12349 3780 12353 3836
rect 12289 3776 12353 3780
rect 16488 3836 16552 3840
rect 16488 3780 16492 3836
rect 16492 3780 16548 3836
rect 16548 3780 16552 3836
rect 16488 3776 16552 3780
rect 16568 3836 16632 3840
rect 16568 3780 16572 3836
rect 16572 3780 16628 3836
rect 16628 3780 16632 3836
rect 16568 3776 16632 3780
rect 16648 3836 16712 3840
rect 16648 3780 16652 3836
rect 16652 3780 16708 3836
rect 16708 3780 16712 3836
rect 16648 3776 16712 3780
rect 16728 3836 16792 3840
rect 16728 3780 16732 3836
rect 16732 3780 16788 3836
rect 16788 3780 16792 3836
rect 16728 3776 16792 3780
rect 5390 3292 5454 3296
rect 5390 3236 5394 3292
rect 5394 3236 5450 3292
rect 5450 3236 5454 3292
rect 5390 3232 5454 3236
rect 5470 3292 5534 3296
rect 5470 3236 5474 3292
rect 5474 3236 5530 3292
rect 5530 3236 5534 3292
rect 5470 3232 5534 3236
rect 5550 3292 5614 3296
rect 5550 3236 5554 3292
rect 5554 3236 5610 3292
rect 5610 3236 5614 3292
rect 5550 3232 5614 3236
rect 5630 3292 5694 3296
rect 5630 3236 5634 3292
rect 5634 3236 5690 3292
rect 5690 3236 5694 3292
rect 5630 3232 5694 3236
rect 9829 3292 9893 3296
rect 9829 3236 9833 3292
rect 9833 3236 9889 3292
rect 9889 3236 9893 3292
rect 9829 3232 9893 3236
rect 9909 3292 9973 3296
rect 9909 3236 9913 3292
rect 9913 3236 9969 3292
rect 9969 3236 9973 3292
rect 9909 3232 9973 3236
rect 9989 3292 10053 3296
rect 9989 3236 9993 3292
rect 9993 3236 10049 3292
rect 10049 3236 10053 3292
rect 9989 3232 10053 3236
rect 10069 3292 10133 3296
rect 10069 3236 10073 3292
rect 10073 3236 10129 3292
rect 10129 3236 10133 3292
rect 10069 3232 10133 3236
rect 14268 3292 14332 3296
rect 14268 3236 14272 3292
rect 14272 3236 14328 3292
rect 14328 3236 14332 3292
rect 14268 3232 14332 3236
rect 14348 3292 14412 3296
rect 14348 3236 14352 3292
rect 14352 3236 14408 3292
rect 14408 3236 14412 3292
rect 14348 3232 14412 3236
rect 14428 3292 14492 3296
rect 14428 3236 14432 3292
rect 14432 3236 14488 3292
rect 14488 3236 14492 3292
rect 14428 3232 14492 3236
rect 14508 3292 14572 3296
rect 14508 3236 14512 3292
rect 14512 3236 14568 3292
rect 14568 3236 14572 3292
rect 14508 3232 14572 3236
rect 18707 3292 18771 3296
rect 18707 3236 18711 3292
rect 18711 3236 18767 3292
rect 18767 3236 18771 3292
rect 18707 3232 18771 3236
rect 18787 3292 18851 3296
rect 18787 3236 18791 3292
rect 18791 3236 18847 3292
rect 18847 3236 18851 3292
rect 18787 3232 18851 3236
rect 18867 3292 18931 3296
rect 18867 3236 18871 3292
rect 18871 3236 18927 3292
rect 18927 3236 18931 3292
rect 18867 3232 18931 3236
rect 18947 3292 19011 3296
rect 18947 3236 18951 3292
rect 18951 3236 19007 3292
rect 19007 3236 19011 3292
rect 18947 3232 19011 3236
rect 3171 2748 3235 2752
rect 3171 2692 3175 2748
rect 3175 2692 3231 2748
rect 3231 2692 3235 2748
rect 3171 2688 3235 2692
rect 3251 2748 3315 2752
rect 3251 2692 3255 2748
rect 3255 2692 3311 2748
rect 3311 2692 3315 2748
rect 3251 2688 3315 2692
rect 3331 2748 3395 2752
rect 3331 2692 3335 2748
rect 3335 2692 3391 2748
rect 3391 2692 3395 2748
rect 3331 2688 3395 2692
rect 3411 2748 3475 2752
rect 3411 2692 3415 2748
rect 3415 2692 3471 2748
rect 3471 2692 3475 2748
rect 3411 2688 3475 2692
rect 7610 2748 7674 2752
rect 7610 2692 7614 2748
rect 7614 2692 7670 2748
rect 7670 2692 7674 2748
rect 7610 2688 7674 2692
rect 7690 2748 7754 2752
rect 7690 2692 7694 2748
rect 7694 2692 7750 2748
rect 7750 2692 7754 2748
rect 7690 2688 7754 2692
rect 7770 2748 7834 2752
rect 7770 2692 7774 2748
rect 7774 2692 7830 2748
rect 7830 2692 7834 2748
rect 7770 2688 7834 2692
rect 7850 2748 7914 2752
rect 7850 2692 7854 2748
rect 7854 2692 7910 2748
rect 7910 2692 7914 2748
rect 7850 2688 7914 2692
rect 12049 2748 12113 2752
rect 12049 2692 12053 2748
rect 12053 2692 12109 2748
rect 12109 2692 12113 2748
rect 12049 2688 12113 2692
rect 12129 2748 12193 2752
rect 12129 2692 12133 2748
rect 12133 2692 12189 2748
rect 12189 2692 12193 2748
rect 12129 2688 12193 2692
rect 12209 2748 12273 2752
rect 12209 2692 12213 2748
rect 12213 2692 12269 2748
rect 12269 2692 12273 2748
rect 12209 2688 12273 2692
rect 12289 2748 12353 2752
rect 12289 2692 12293 2748
rect 12293 2692 12349 2748
rect 12349 2692 12353 2748
rect 12289 2688 12353 2692
rect 16488 2748 16552 2752
rect 16488 2692 16492 2748
rect 16492 2692 16548 2748
rect 16548 2692 16552 2748
rect 16488 2688 16552 2692
rect 16568 2748 16632 2752
rect 16568 2692 16572 2748
rect 16572 2692 16628 2748
rect 16628 2692 16632 2748
rect 16568 2688 16632 2692
rect 16648 2748 16712 2752
rect 16648 2692 16652 2748
rect 16652 2692 16708 2748
rect 16708 2692 16712 2748
rect 16648 2688 16712 2692
rect 16728 2748 16792 2752
rect 16728 2692 16732 2748
rect 16732 2692 16788 2748
rect 16788 2692 16792 2748
rect 16728 2688 16792 2692
rect 5390 2204 5454 2208
rect 5390 2148 5394 2204
rect 5394 2148 5450 2204
rect 5450 2148 5454 2204
rect 5390 2144 5454 2148
rect 5470 2204 5534 2208
rect 5470 2148 5474 2204
rect 5474 2148 5530 2204
rect 5530 2148 5534 2204
rect 5470 2144 5534 2148
rect 5550 2204 5614 2208
rect 5550 2148 5554 2204
rect 5554 2148 5610 2204
rect 5610 2148 5614 2204
rect 5550 2144 5614 2148
rect 5630 2204 5694 2208
rect 5630 2148 5634 2204
rect 5634 2148 5690 2204
rect 5690 2148 5694 2204
rect 5630 2144 5694 2148
rect 9829 2204 9893 2208
rect 9829 2148 9833 2204
rect 9833 2148 9889 2204
rect 9889 2148 9893 2204
rect 9829 2144 9893 2148
rect 9909 2204 9973 2208
rect 9909 2148 9913 2204
rect 9913 2148 9969 2204
rect 9969 2148 9973 2204
rect 9909 2144 9973 2148
rect 9989 2204 10053 2208
rect 9989 2148 9993 2204
rect 9993 2148 10049 2204
rect 10049 2148 10053 2204
rect 9989 2144 10053 2148
rect 10069 2204 10133 2208
rect 10069 2148 10073 2204
rect 10073 2148 10129 2204
rect 10129 2148 10133 2204
rect 10069 2144 10133 2148
rect 14268 2204 14332 2208
rect 14268 2148 14272 2204
rect 14272 2148 14328 2204
rect 14328 2148 14332 2204
rect 14268 2144 14332 2148
rect 14348 2204 14412 2208
rect 14348 2148 14352 2204
rect 14352 2148 14408 2204
rect 14408 2148 14412 2204
rect 14348 2144 14412 2148
rect 14428 2204 14492 2208
rect 14428 2148 14432 2204
rect 14432 2148 14488 2204
rect 14488 2148 14492 2204
rect 14428 2144 14492 2148
rect 14508 2204 14572 2208
rect 14508 2148 14512 2204
rect 14512 2148 14568 2204
rect 14568 2148 14572 2204
rect 14508 2144 14572 2148
rect 18707 2204 18771 2208
rect 18707 2148 18711 2204
rect 18711 2148 18767 2204
rect 18767 2148 18771 2204
rect 18707 2144 18771 2148
rect 18787 2204 18851 2208
rect 18787 2148 18791 2204
rect 18791 2148 18847 2204
rect 18847 2148 18851 2204
rect 18787 2144 18851 2148
rect 18867 2204 18931 2208
rect 18867 2148 18871 2204
rect 18871 2148 18927 2204
rect 18927 2148 18931 2204
rect 18867 2144 18931 2148
rect 18947 2204 19011 2208
rect 18947 2148 18951 2204
rect 18951 2148 19007 2204
rect 19007 2148 19011 2204
rect 18947 2144 19011 2148
<< metal4 >>
rect 3163 7104 3483 7664
rect 3163 7040 3171 7104
rect 3235 7040 3251 7104
rect 3315 7040 3331 7104
rect 3395 7040 3411 7104
rect 3475 7040 3483 7104
rect 3163 6016 3483 7040
rect 3163 5952 3171 6016
rect 3235 5952 3251 6016
rect 3315 5952 3331 6016
rect 3395 5952 3411 6016
rect 3475 5952 3483 6016
rect 3163 4928 3483 5952
rect 3163 4864 3171 4928
rect 3235 4864 3251 4928
rect 3315 4864 3331 4928
rect 3395 4864 3411 4928
rect 3475 4864 3483 4928
rect 3163 3840 3483 4864
rect 3163 3776 3171 3840
rect 3235 3776 3251 3840
rect 3315 3776 3331 3840
rect 3395 3776 3411 3840
rect 3475 3776 3483 3840
rect 3163 2752 3483 3776
rect 3163 2688 3171 2752
rect 3235 2688 3251 2752
rect 3315 2688 3331 2752
rect 3395 2688 3411 2752
rect 3475 2688 3483 2752
rect 3163 2128 3483 2688
rect 5382 7648 5702 7664
rect 5382 7584 5390 7648
rect 5454 7584 5470 7648
rect 5534 7584 5550 7648
rect 5614 7584 5630 7648
rect 5694 7584 5702 7648
rect 5382 6560 5702 7584
rect 5382 6496 5390 6560
rect 5454 6496 5470 6560
rect 5534 6496 5550 6560
rect 5614 6496 5630 6560
rect 5694 6496 5702 6560
rect 5382 5472 5702 6496
rect 5382 5408 5390 5472
rect 5454 5408 5470 5472
rect 5534 5408 5550 5472
rect 5614 5408 5630 5472
rect 5694 5408 5702 5472
rect 5382 4384 5702 5408
rect 5382 4320 5390 4384
rect 5454 4320 5470 4384
rect 5534 4320 5550 4384
rect 5614 4320 5630 4384
rect 5694 4320 5702 4384
rect 5382 3296 5702 4320
rect 5382 3232 5390 3296
rect 5454 3232 5470 3296
rect 5534 3232 5550 3296
rect 5614 3232 5630 3296
rect 5694 3232 5702 3296
rect 5382 2208 5702 3232
rect 5382 2144 5390 2208
rect 5454 2144 5470 2208
rect 5534 2144 5550 2208
rect 5614 2144 5630 2208
rect 5694 2144 5702 2208
rect 5382 2128 5702 2144
rect 7602 7104 7922 7664
rect 7602 7040 7610 7104
rect 7674 7040 7690 7104
rect 7754 7040 7770 7104
rect 7834 7040 7850 7104
rect 7914 7040 7922 7104
rect 7602 6016 7922 7040
rect 7602 5952 7610 6016
rect 7674 5952 7690 6016
rect 7754 5952 7770 6016
rect 7834 5952 7850 6016
rect 7914 5952 7922 6016
rect 7602 4928 7922 5952
rect 7602 4864 7610 4928
rect 7674 4864 7690 4928
rect 7754 4864 7770 4928
rect 7834 4864 7850 4928
rect 7914 4864 7922 4928
rect 7602 3840 7922 4864
rect 7602 3776 7610 3840
rect 7674 3776 7690 3840
rect 7754 3776 7770 3840
rect 7834 3776 7850 3840
rect 7914 3776 7922 3840
rect 7602 2752 7922 3776
rect 7602 2688 7610 2752
rect 7674 2688 7690 2752
rect 7754 2688 7770 2752
rect 7834 2688 7850 2752
rect 7914 2688 7922 2752
rect 7602 2128 7922 2688
rect 9821 7648 10141 7664
rect 9821 7584 9829 7648
rect 9893 7584 9909 7648
rect 9973 7584 9989 7648
rect 10053 7584 10069 7648
rect 10133 7584 10141 7648
rect 9821 6560 10141 7584
rect 9821 6496 9829 6560
rect 9893 6496 9909 6560
rect 9973 6496 9989 6560
rect 10053 6496 10069 6560
rect 10133 6496 10141 6560
rect 9821 5472 10141 6496
rect 9821 5408 9829 5472
rect 9893 5408 9909 5472
rect 9973 5408 9989 5472
rect 10053 5408 10069 5472
rect 10133 5408 10141 5472
rect 9821 4384 10141 5408
rect 9821 4320 9829 4384
rect 9893 4320 9909 4384
rect 9973 4320 9989 4384
rect 10053 4320 10069 4384
rect 10133 4320 10141 4384
rect 9821 3296 10141 4320
rect 9821 3232 9829 3296
rect 9893 3232 9909 3296
rect 9973 3232 9989 3296
rect 10053 3232 10069 3296
rect 10133 3232 10141 3296
rect 9821 2208 10141 3232
rect 9821 2144 9829 2208
rect 9893 2144 9909 2208
rect 9973 2144 9989 2208
rect 10053 2144 10069 2208
rect 10133 2144 10141 2208
rect 9821 2128 10141 2144
rect 12041 7104 12361 7664
rect 12041 7040 12049 7104
rect 12113 7040 12129 7104
rect 12193 7040 12209 7104
rect 12273 7040 12289 7104
rect 12353 7040 12361 7104
rect 12041 6016 12361 7040
rect 12041 5952 12049 6016
rect 12113 5952 12129 6016
rect 12193 5952 12209 6016
rect 12273 5952 12289 6016
rect 12353 5952 12361 6016
rect 12041 4928 12361 5952
rect 12041 4864 12049 4928
rect 12113 4864 12129 4928
rect 12193 4864 12209 4928
rect 12273 4864 12289 4928
rect 12353 4864 12361 4928
rect 12041 3840 12361 4864
rect 12041 3776 12049 3840
rect 12113 3776 12129 3840
rect 12193 3776 12209 3840
rect 12273 3776 12289 3840
rect 12353 3776 12361 3840
rect 12041 2752 12361 3776
rect 12041 2688 12049 2752
rect 12113 2688 12129 2752
rect 12193 2688 12209 2752
rect 12273 2688 12289 2752
rect 12353 2688 12361 2752
rect 12041 2128 12361 2688
rect 14260 7648 14580 7664
rect 14260 7584 14268 7648
rect 14332 7584 14348 7648
rect 14412 7584 14428 7648
rect 14492 7584 14508 7648
rect 14572 7584 14580 7648
rect 14260 6560 14580 7584
rect 14260 6496 14268 6560
rect 14332 6496 14348 6560
rect 14412 6496 14428 6560
rect 14492 6496 14508 6560
rect 14572 6496 14580 6560
rect 14260 5472 14580 6496
rect 14260 5408 14268 5472
rect 14332 5408 14348 5472
rect 14412 5408 14428 5472
rect 14492 5408 14508 5472
rect 14572 5408 14580 5472
rect 14260 4384 14580 5408
rect 14260 4320 14268 4384
rect 14332 4320 14348 4384
rect 14412 4320 14428 4384
rect 14492 4320 14508 4384
rect 14572 4320 14580 4384
rect 14260 3296 14580 4320
rect 14260 3232 14268 3296
rect 14332 3232 14348 3296
rect 14412 3232 14428 3296
rect 14492 3232 14508 3296
rect 14572 3232 14580 3296
rect 14260 2208 14580 3232
rect 14260 2144 14268 2208
rect 14332 2144 14348 2208
rect 14412 2144 14428 2208
rect 14492 2144 14508 2208
rect 14572 2144 14580 2208
rect 14260 2128 14580 2144
rect 16480 7104 16800 7664
rect 16480 7040 16488 7104
rect 16552 7040 16568 7104
rect 16632 7040 16648 7104
rect 16712 7040 16728 7104
rect 16792 7040 16800 7104
rect 16480 6016 16800 7040
rect 16480 5952 16488 6016
rect 16552 5952 16568 6016
rect 16632 5952 16648 6016
rect 16712 5952 16728 6016
rect 16792 5952 16800 6016
rect 16480 4928 16800 5952
rect 16480 4864 16488 4928
rect 16552 4864 16568 4928
rect 16632 4864 16648 4928
rect 16712 4864 16728 4928
rect 16792 4864 16800 4928
rect 16480 3840 16800 4864
rect 16480 3776 16488 3840
rect 16552 3776 16568 3840
rect 16632 3776 16648 3840
rect 16712 3776 16728 3840
rect 16792 3776 16800 3840
rect 16480 2752 16800 3776
rect 16480 2688 16488 2752
rect 16552 2688 16568 2752
rect 16632 2688 16648 2752
rect 16712 2688 16728 2752
rect 16792 2688 16800 2752
rect 16480 2128 16800 2688
rect 18699 7648 19019 7664
rect 18699 7584 18707 7648
rect 18771 7584 18787 7648
rect 18851 7584 18867 7648
rect 18931 7584 18947 7648
rect 19011 7584 19019 7648
rect 18699 6560 19019 7584
rect 18699 6496 18707 6560
rect 18771 6496 18787 6560
rect 18851 6496 18867 6560
rect 18931 6496 18947 6560
rect 19011 6496 19019 6560
rect 18699 5472 19019 6496
rect 18699 5408 18707 5472
rect 18771 5408 18787 5472
rect 18851 5408 18867 5472
rect 18931 5408 18947 5472
rect 19011 5408 19019 5472
rect 18699 4384 19019 5408
rect 18699 4320 18707 4384
rect 18771 4320 18787 4384
rect 18851 4320 18867 4384
rect 18931 4320 18947 4384
rect 19011 4320 19019 4384
rect 18699 3296 19019 4320
rect 18699 3232 18707 3296
rect 18771 3232 18787 3296
rect 18851 3232 18867 3296
rect 18931 3232 18947 3296
rect 19011 3232 19019 3296
rect 18699 2208 19019 3232
rect 18699 2144 18707 2208
rect 18771 2144 18787 2208
rect 18851 2144 18867 2208
rect 18931 2144 18947 2208
rect 19011 2144 19019 2208
rect 18699 2128 19019 2144
<< labels >>
rlabel metal1 s 9982 7072 9982 7072 4 vccd1
rlabel metal2 s 10061 7616 10061 7616 4 vssd1
rlabel metal1 s 11760 3094 11760 3094 4 _00_
rlabel metal2 s 14766 2584 14766 2584 4 _01_
rlabel metal2 s 10069 2346 10069 2346 4 _02_
rlabel metal2 s 12001 4182 12001 4182 4 _03_
rlabel metal2 s 12466 3978 12466 3978 4 _04_
rlabel metal1 s 10299 3502 10299 3502 4 _05_
rlabel metal1 s 8321 3502 8321 3502 4 _06_
rlabel metal2 s 4273 3502 4273 3502 4 _07_
rlabel metal1 s 4319 3434 4319 3434 4 _08_
rlabel metal2 s 5754 4114 5754 4114 4 _09_
rlabel metal1 s 5070 2414 5070 2414 4 _10_
rlabel metal2 s 3082 5066 3082 5066 4 _11_
rlabel metal2 s 7038 5202 7038 5202 4 _12_
rlabel metal1 s 4722 2346 4722 2346 4 _13_
rlabel metal1 s 3782 4114 3782 4114 4 _14_
rlabel metal2 s 16882 2771 16882 2771 4 _15_
rlabel metal1 s 9169 2346 9169 2346 4 _16_
rlabel metal2 s 9338 4692 9338 4692 4 _17_
rlabel metal2 s 17066 3196 17066 3196 4 _18_
rlabel metal2 s 15686 4284 15686 4284 4 _19_
rlabel metal2 s 13110 4896 13110 4896 4 _20_
rlabel metal1 s 13478 4658 13478 4658 4 _21_
rlabel metal2 s 10902 4896 10902 4896 4 _22_
rlabel metal1 s 9614 5202 9614 5202 4 _23_
rlabel metal1 s 5658 4794 5658 4794 4 _24_
rlabel metal2 s 6670 4352 6670 4352 4 _25_
rlabel metal1 s 6394 4794 6394 4794 4 _26_
rlabel metal1 s 8280 4114 8280 4114 4 _27_
rlabel metal2 s 4002 5236 4002 5236 4 _28_
rlabel metal2 s 2898 5508 2898 5508 4 _29_
rlabel metal2 s 1978 4556 1978 4556 4 _30_
rlabel metal1 s 6463 5202 6463 5202 4 _31_
rlabel metal1 s 17158 2414 17158 2414 4 _32_
rlabel metal1 s 16192 3502 16192 3502 4 _33_
rlabel metal1 s 7544 3026 7544 3026 4 clk
rlabel metal1 s 7636 4182 7636 4182 4 clknet_0_clk
rlabel metal1 s 4324 2482 4324 2482 4 clknet_1_0__leaf_clk
rlabel metal1 s 12512 2414 12512 2414 4 clknet_1_1__leaf_clk
rlabel metal1 s 10212 7446 10212 7446 4 comp
rlabel metal1 s 1426 7514 1426 7514 4 dq[0]
rlabel metal1 s 3726 7514 3726 7514 4 dq[1]
rlabel metal2 s 5750 8415 5750 8415 4 dq[2]
rlabel metal1 s 7912 7514 7912 7514 4 dq[3]
rlabel metal2 s 12374 8415 12374 8415 4 dq[4]
rlabel metal2 s 14674 8415 14674 8415 4 dq[5]
rlabel metal1 s 16836 7514 16836 7514 4 dq[6]
rlabel metal1 s 18354 7514 18354 7514 4 dq[7]
rlabel metal2 s 17434 1520 17434 1520 4 last_cycle
rlabel metal2 s 13570 5474 13570 5474 4 net1
rlabel metal1 s 18078 7344 18078 7344 4 net10
rlabel metal2 s 17526 2992 17526 2992 4 net11
rlabel metal2 s 12466 1792 12466 1792 4 net12
rlabel metal2 s 2162 4148 2162 4148 4 net2
rlabel metal1 s 1978 2618 1978 2618 4 net3
rlabel metal2 s 4646 5814 4646 5814 4 net4
rlabel metal1 s 6992 5338 6992 5338 4 net5
rlabel metal2 s 7130 4454 7130 4454 4 net6
rlabel metal1 s 10442 5678 10442 5678 4 net7
rlabel metal1 s 12604 5542 12604 5542 4 net8
rlabel metal2 s 14674 4624 14674 4624 4 net9
rlabel metal1 s 2254 3026 2254 3026 4 rst_n
rlabel metal3 s 6302 4675 6302 4675 4 sr\[1\]
rlabel metal1 s 6302 2618 6302 2618 4 sr\[2\]
rlabel metal1 s 10051 5746 10051 5746 4 sr\[3\]
rlabel metal1 s 10074 5134 10074 5134 4 sr\[4\]
rlabel metal1 s 8556 2278 8556 2278 4 sr\[5\]
rlabel metal1 s 16698 3468 16698 3468 4 sr\[6\]
rlabel metal1 s 13202 3162 13202 3162 4 sr\[7\]
rlabel metal1 s 11454 5134 11454 5134 4 sr_dly\[0\]
flabel metal2 s 7470 0 7526 800 0 FreeSans 280 90 0 0 clk
port 1 nsew
flabel metal2 s 9954 9200 10010 10000 0 FreeSans 280 90 0 0 comp
port 2 nsew
flabel metal2 s 1122 9200 1178 10000 0 FreeSans 280 90 0 0 dq[0]
port 3 nsew
flabel metal2 s 3330 9200 3386 10000 0 FreeSans 280 90 0 0 dq[1]
port 4 nsew
flabel metal2 s 5538 9200 5594 10000 0 FreeSans 280 90 0 0 dq[2]
port 5 nsew
flabel metal2 s 7746 9200 7802 10000 0 FreeSans 280 90 0 0 dq[3]
port 6 nsew
flabel metal2 s 12162 9200 12218 10000 0 FreeSans 280 90 0 0 dq[4]
port 7 nsew
flabel metal2 s 14370 9200 14426 10000 0 FreeSans 280 90 0 0 dq[5]
port 8 nsew
flabel metal2 s 16578 9200 16634 10000 0 FreeSans 280 90 0 0 dq[6]
port 9 nsew
flabel metal2 s 18786 9200 18842 10000 0 FreeSans 280 90 0 0 dq[7]
port 10 nsew
flabel metal2 s 17406 0 17462 800 0 FreeSans 280 90 0 0 last_cycle
port 11 nsew
flabel metal2 s 2502 0 2558 800 0 FreeSans 280 90 0 0 rst_n
port 12 nsew
flabel metal2 s 12438 0 12494 800 0 FreeSans 280 90 0 0 valid
port 13 nsew
flabel metal4 s 3163 2128 3483 7664 0 FreeSans 2400 90 0 0 vccd1
port 14 nsew
flabel metal4 s 7602 2128 7922 7664 0 FreeSans 2400 90 0 0 vccd1
port 14 nsew
flabel metal4 s 12041 2128 12361 7664 0 FreeSans 2400 90 0 0 vccd1
port 14 nsew
flabel metal4 s 16480 2128 16800 7664 0 FreeSans 2400 90 0 0 vccd1
port 14 nsew
flabel metal4 s 5382 2128 5702 7664 0 FreeSans 2400 90 0 0 vssd1
port 15 nsew
flabel metal4 s 9821 2128 10141 7664 0 FreeSans 2400 90 0 0 vssd1
port 15 nsew
flabel metal4 s 14260 2128 14580 7664 0 FreeSans 2400 90 0 0 vssd1
port 15 nsew
flabel metal4 s 18699 2128 19019 7664 0 FreeSans 2400 90 0 0 vssd1
port 15 nsew
<< end >>