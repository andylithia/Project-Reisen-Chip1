magic
tech sky130A
magscale 1 2
timestamp 1672464819
<< pwell >>
rect 4180 1431 5070 2657
rect 4180 1397 4216 1431
rect 5034 1397 5070 1431
rect 4180 1361 5070 1397
<< psubdiff >>
rect 4216 2587 4312 2621
rect 4518 2587 4676 2621
rect 4882 2587 5034 2621
rect 4216 2525 4250 2587
rect 4580 2525 4614 2587
rect 4944 1431 5034 2587
rect 4216 1397 5034 1431
<< psubdiffcont >>
rect 4312 2587 4518 2621
rect 4676 2587 4882 2621
rect 4216 1431 4250 2525
rect 4580 1431 4614 2525
<< xpolycontact >>
rect 4346 2059 4484 2491
rect 4346 1527 4484 1959
rect 4710 2059 4848 2491
rect 4710 1527 4848 1959
<< ppolyres >>
rect 4346 1959 4484 2059
rect 4710 1959 4848 2059
<< locali >>
rect 4216 2621 4287 2658
rect 4216 2587 4312 2621
rect 4518 2587 4676 2621
rect 4882 2587 4944 2621
rect 4216 2574 4287 2587
rect 4216 2525 4229 2574
rect 4274 1431 4287 2574
rect 4580 2525 4614 2587
rect 4216 1397 4287 1431
rect 4580 1397 4614 1431
<< viali >>
rect 4229 2525 4274 2574
rect 4229 1431 4250 2525
rect 4250 1431 4274 2525
rect 4362 2076 4468 2473
rect 4362 1545 4468 1942
rect 4726 2076 4832 2473
rect 4726 1545 4832 1942
<< metal1 >>
rect 4216 2574 4287 2658
rect 4216 1431 4225 2574
rect 4277 1431 4287 2574
rect 4356 2473 4474 2485
rect 4356 2076 4362 2473
rect 4468 2076 4474 2473
rect 4356 2064 4474 2076
rect 4710 2473 4848 2491
rect 4710 2076 4726 2473
rect 4832 2076 4848 2473
rect 4710 2059 4848 2076
rect 4346 1942 4484 1959
rect 4346 1545 4362 1942
rect 4468 1545 4484 1942
rect 4346 1527 4484 1545
rect 4720 1942 4838 1954
rect 4720 1545 4726 1942
rect 4832 1545 4838 1942
rect 4720 1533 4838 1545
rect 4216 1397 4287 1431
<< via1 >>
rect 4225 1431 4229 2574
rect 4229 1431 4274 2574
rect 4274 1431 4277 2574
rect 4362 2076 4468 2473
rect 4726 2076 4832 2473
rect 4362 1545 4468 1942
rect 4726 1545 4832 1942
<< metal2 >>
rect 4250 2658 4280 2670
rect 4216 2574 4287 2658
rect 4216 1431 4225 2574
rect 4277 1431 4287 2574
rect 4346 2473 4484 2491
rect 4346 2076 4362 2473
rect 4468 2250 4484 2473
rect 4710 2473 4848 2491
rect 4710 2250 4726 2473
rect 4468 2190 4726 2250
rect 4468 2150 4484 2190
rect 4710 2150 4726 2190
rect 4468 2090 4726 2150
rect 4468 2076 4484 2090
rect 4346 2059 4484 2076
rect 4710 2076 4726 2090
rect 4832 2076 4848 2473
rect 4710 2059 4848 2076
rect 4346 1942 4484 1959
rect 4346 1545 4362 1942
rect 4468 1940 4484 1942
rect 4710 1942 4848 1959
rect 4710 1940 4726 1942
rect 4468 1880 4726 1940
rect 4468 1840 4484 1880
rect 4710 1840 4726 1880
rect 4468 1780 4726 1840
rect 4468 1545 4484 1780
rect 4346 1527 4484 1545
rect 4710 1545 4726 1780
rect 4832 1545 4848 1942
rect 4710 1527 4848 1545
<< via2 >>
rect 4362 2076 4468 2473
rect 4726 1545 4832 1942
<< metal3 >>
rect 4346 2473 4484 2491
rect 4346 2440 4362 2473
rect 4190 2380 4362 2440
rect 4330 2340 4362 2380
rect 4346 2076 4362 2340
rect 4468 2076 4484 2473
rect 4346 2059 4484 2076
rect 4870 2340 5034 2440
rect 4870 1960 4930 2340
rect 4810 1959 4930 1960
rect 4710 1942 4930 1959
rect 4710 1545 4726 1942
rect 4832 1900 4930 1942
rect 4832 1545 4848 1900
rect 4710 1527 4848 1545
<< labels >>
rlabel metal2 4250 2660 4280 2670 5 VLO
port 2 s
rlabel metal3 5014 2340 5034 2440 1 IO2
port 1 n
rlabel metal3 4190 2380 4212 2440 1 IO1
port 4 n
<< end >>
