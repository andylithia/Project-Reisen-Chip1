magic
tech sky130B
magscale 1 2
timestamp 1668572718
<< nwell >>
rect 3166 -3954 6378 -2940
<< pwell >>
rect 3198 -4110 6346 -4072
rect 3198 -4144 3539 -4110
rect 3542 -4144 3600 -4110
rect 3605 -4144 5939 -4110
rect 5944 -4144 6002 -4110
rect 6005 -4144 6346 -4110
rect 3198 -4728 6346 -4144
<< nmos >>
rect 3269 -4582 3299 -4182
rect 3365 -4582 3395 -4182
rect 3461 -4582 3491 -4182
rect 3557 -4582 3587 -4182
rect 3653 -4582 3683 -4182
rect 3749 -4582 3779 -4182
rect 3845 -4582 3875 -4182
rect 3941 -4582 3971 -4182
rect 4037 -4582 4067 -4182
rect 4133 -4582 4163 -4182
rect 4229 -4582 4259 -4182
rect 4325 -4582 4355 -4182
rect 4421 -4582 4451 -4182
rect 4517 -4582 4547 -4182
rect 4613 -4582 4643 -4182
rect 4709 -4582 4739 -4182
rect 4805 -4582 4835 -4182
rect 4901 -4582 4931 -4182
rect 4997 -4582 5027 -4182
rect 5093 -4582 5123 -4182
rect 5189 -4582 5219 -4182
rect 5285 -4582 5315 -4182
rect 5381 -4582 5411 -4182
rect 5477 -4582 5507 -4182
rect 5573 -4582 5603 -4182
rect 5669 -4582 5699 -4182
rect 5765 -4582 5795 -4182
rect 5861 -4582 5891 -4182
rect 5957 -4582 5987 -4182
rect 6053 -4582 6083 -4182
rect 6149 -4582 6179 -4182
rect 6245 -4582 6275 -4182
<< pmos >>
rect 3269 -3827 3299 -3107
rect 3365 -3827 3395 -3107
rect 3461 -3827 3491 -3107
rect 3557 -3827 3587 -3107
rect 3653 -3827 3683 -3107
rect 3749 -3827 3779 -3107
rect 3845 -3827 3875 -3107
rect 3941 -3827 3971 -3107
rect 4037 -3827 4067 -3107
rect 4133 -3827 4163 -3107
rect 4229 -3827 4259 -3107
rect 4325 -3827 4355 -3107
rect 4421 -3827 4451 -3107
rect 4517 -3827 4547 -3107
rect 4613 -3827 4643 -3107
rect 4709 -3827 4739 -3107
rect 4805 -3827 4835 -3107
rect 4901 -3827 4931 -3107
rect 4997 -3827 5027 -3107
rect 5093 -3827 5123 -3107
rect 5189 -3827 5219 -3107
rect 5285 -3827 5315 -3107
rect 5381 -3827 5411 -3107
rect 5477 -3827 5507 -3107
rect 5573 -3827 5603 -3107
rect 5669 -3827 5699 -3107
rect 5765 -3827 5795 -3107
rect 5861 -3827 5891 -3107
rect 5957 -3827 5987 -3107
rect 6053 -3827 6083 -3107
rect 6149 -3827 6179 -3107
rect 6245 -3827 6275 -3107
<< ndiff >>
rect 3207 -4194 3269 -4182
rect 3207 -4570 3219 -4194
rect 3253 -4570 3269 -4194
rect 3207 -4582 3269 -4570
rect 3299 -4194 3365 -4182
rect 3299 -4570 3315 -4194
rect 3349 -4570 3365 -4194
rect 3299 -4582 3365 -4570
rect 3395 -4194 3461 -4182
rect 3395 -4570 3411 -4194
rect 3445 -4570 3461 -4194
rect 3395 -4582 3461 -4570
rect 3491 -4194 3557 -4182
rect 3491 -4570 3507 -4194
rect 3541 -4570 3557 -4194
rect 3491 -4582 3557 -4570
rect 3587 -4194 3653 -4182
rect 3587 -4570 3603 -4194
rect 3637 -4570 3653 -4194
rect 3587 -4582 3653 -4570
rect 3683 -4194 3749 -4182
rect 3683 -4570 3699 -4194
rect 3733 -4570 3749 -4194
rect 3683 -4582 3749 -4570
rect 3779 -4194 3845 -4182
rect 3779 -4570 3795 -4194
rect 3829 -4570 3845 -4194
rect 3779 -4582 3845 -4570
rect 3875 -4194 3941 -4182
rect 3875 -4570 3891 -4194
rect 3925 -4570 3941 -4194
rect 3875 -4582 3941 -4570
rect 3971 -4194 4037 -4182
rect 3971 -4570 3987 -4194
rect 4021 -4570 4037 -4194
rect 3971 -4582 4037 -4570
rect 4067 -4194 4133 -4182
rect 4067 -4570 4083 -4194
rect 4117 -4570 4133 -4194
rect 4067 -4582 4133 -4570
rect 4163 -4194 4229 -4182
rect 4163 -4570 4179 -4194
rect 4213 -4570 4229 -4194
rect 4163 -4582 4229 -4570
rect 4259 -4194 4325 -4182
rect 4259 -4570 4275 -4194
rect 4309 -4570 4325 -4194
rect 4259 -4582 4325 -4570
rect 4355 -4194 4421 -4182
rect 4355 -4570 4371 -4194
rect 4405 -4570 4421 -4194
rect 4355 -4582 4421 -4570
rect 4451 -4194 4517 -4182
rect 4451 -4570 4467 -4194
rect 4501 -4570 4517 -4194
rect 4451 -4582 4517 -4570
rect 4547 -4194 4613 -4182
rect 4547 -4570 4563 -4194
rect 4597 -4570 4613 -4194
rect 4547 -4582 4613 -4570
rect 4643 -4194 4709 -4182
rect 4643 -4570 4659 -4194
rect 4693 -4570 4709 -4194
rect 4643 -4582 4709 -4570
rect 4739 -4194 4805 -4182
rect 4739 -4570 4755 -4194
rect 4789 -4570 4805 -4194
rect 4739 -4582 4805 -4570
rect 4835 -4194 4901 -4182
rect 4835 -4570 4851 -4194
rect 4885 -4570 4901 -4194
rect 4835 -4582 4901 -4570
rect 4931 -4194 4997 -4182
rect 4931 -4570 4947 -4194
rect 4981 -4570 4997 -4194
rect 4931 -4582 4997 -4570
rect 5027 -4194 5093 -4182
rect 5027 -4570 5043 -4194
rect 5077 -4570 5093 -4194
rect 5027 -4582 5093 -4570
rect 5123 -4194 5189 -4182
rect 5123 -4570 5139 -4194
rect 5173 -4570 5189 -4194
rect 5123 -4582 5189 -4570
rect 5219 -4194 5285 -4182
rect 5219 -4570 5235 -4194
rect 5269 -4570 5285 -4194
rect 5219 -4582 5285 -4570
rect 5315 -4194 5381 -4182
rect 5315 -4570 5331 -4194
rect 5365 -4570 5381 -4194
rect 5315 -4582 5381 -4570
rect 5411 -4194 5477 -4182
rect 5411 -4570 5427 -4194
rect 5461 -4570 5477 -4194
rect 5411 -4582 5477 -4570
rect 5507 -4194 5573 -4182
rect 5507 -4570 5523 -4194
rect 5557 -4570 5573 -4194
rect 5507 -4582 5573 -4570
rect 5603 -4194 5669 -4182
rect 5603 -4570 5619 -4194
rect 5653 -4570 5669 -4194
rect 5603 -4582 5669 -4570
rect 5699 -4194 5765 -4182
rect 5699 -4570 5715 -4194
rect 5749 -4570 5765 -4194
rect 5699 -4582 5765 -4570
rect 5795 -4194 5861 -4182
rect 5795 -4570 5811 -4194
rect 5845 -4570 5861 -4194
rect 5795 -4582 5861 -4570
rect 5891 -4194 5957 -4182
rect 5891 -4570 5907 -4194
rect 5941 -4570 5957 -4194
rect 5891 -4582 5957 -4570
rect 5987 -4194 6053 -4182
rect 5987 -4570 6003 -4194
rect 6037 -4570 6053 -4194
rect 5987 -4582 6053 -4570
rect 6083 -4194 6149 -4182
rect 6083 -4570 6099 -4194
rect 6133 -4570 6149 -4194
rect 6083 -4582 6149 -4570
rect 6179 -4194 6245 -4182
rect 6179 -4570 6195 -4194
rect 6229 -4570 6245 -4194
rect 6179 -4582 6245 -4570
rect 6275 -4194 6337 -4182
rect 6275 -4570 6291 -4194
rect 6325 -4570 6337 -4194
rect 6275 -4582 6337 -4570
<< pdiff >>
rect 3207 -3119 3269 -3107
rect 3207 -3815 3219 -3119
rect 3253 -3815 3269 -3119
rect 3207 -3827 3269 -3815
rect 3299 -3119 3365 -3107
rect 3299 -3815 3315 -3119
rect 3349 -3815 3365 -3119
rect 3299 -3827 3365 -3815
rect 3395 -3119 3461 -3107
rect 3395 -3815 3411 -3119
rect 3445 -3815 3461 -3119
rect 3395 -3827 3461 -3815
rect 3491 -3119 3557 -3107
rect 3491 -3815 3507 -3119
rect 3541 -3815 3557 -3119
rect 3491 -3827 3557 -3815
rect 3587 -3119 3653 -3107
rect 3587 -3815 3603 -3119
rect 3637 -3815 3653 -3119
rect 3587 -3827 3653 -3815
rect 3683 -3119 3749 -3107
rect 3683 -3815 3699 -3119
rect 3733 -3815 3749 -3119
rect 3683 -3827 3749 -3815
rect 3779 -3119 3845 -3107
rect 3779 -3815 3795 -3119
rect 3829 -3815 3845 -3119
rect 3779 -3827 3845 -3815
rect 3875 -3119 3941 -3107
rect 3875 -3815 3891 -3119
rect 3925 -3815 3941 -3119
rect 3875 -3827 3941 -3815
rect 3971 -3119 4037 -3107
rect 3971 -3815 3987 -3119
rect 4021 -3815 4037 -3119
rect 3971 -3827 4037 -3815
rect 4067 -3119 4133 -3107
rect 4067 -3815 4083 -3119
rect 4117 -3815 4133 -3119
rect 4067 -3827 4133 -3815
rect 4163 -3119 4229 -3107
rect 4163 -3815 4179 -3119
rect 4213 -3815 4229 -3119
rect 4163 -3827 4229 -3815
rect 4259 -3119 4325 -3107
rect 4259 -3815 4275 -3119
rect 4309 -3815 4325 -3119
rect 4259 -3827 4325 -3815
rect 4355 -3119 4421 -3107
rect 4355 -3815 4371 -3119
rect 4405 -3815 4421 -3119
rect 4355 -3827 4421 -3815
rect 4451 -3119 4517 -3107
rect 4451 -3815 4467 -3119
rect 4501 -3815 4517 -3119
rect 4451 -3827 4517 -3815
rect 4547 -3119 4613 -3107
rect 4547 -3815 4563 -3119
rect 4597 -3815 4613 -3119
rect 4547 -3827 4613 -3815
rect 4643 -3119 4709 -3107
rect 4643 -3815 4659 -3119
rect 4693 -3815 4709 -3119
rect 4643 -3827 4709 -3815
rect 4739 -3119 4805 -3107
rect 4739 -3815 4755 -3119
rect 4789 -3815 4805 -3119
rect 4739 -3827 4805 -3815
rect 4835 -3119 4901 -3107
rect 4835 -3815 4851 -3119
rect 4885 -3815 4901 -3119
rect 4835 -3827 4901 -3815
rect 4931 -3119 4997 -3107
rect 4931 -3815 4947 -3119
rect 4981 -3815 4997 -3119
rect 4931 -3827 4997 -3815
rect 5027 -3119 5093 -3107
rect 5027 -3815 5043 -3119
rect 5077 -3815 5093 -3119
rect 5027 -3827 5093 -3815
rect 5123 -3119 5189 -3107
rect 5123 -3815 5139 -3119
rect 5173 -3815 5189 -3119
rect 5123 -3827 5189 -3815
rect 5219 -3119 5285 -3107
rect 5219 -3815 5235 -3119
rect 5269 -3815 5285 -3119
rect 5219 -3827 5285 -3815
rect 5315 -3119 5381 -3107
rect 5315 -3815 5331 -3119
rect 5365 -3815 5381 -3119
rect 5315 -3827 5381 -3815
rect 5411 -3119 5477 -3107
rect 5411 -3815 5427 -3119
rect 5461 -3815 5477 -3119
rect 5411 -3827 5477 -3815
rect 5507 -3119 5573 -3107
rect 5507 -3815 5523 -3119
rect 5557 -3815 5573 -3119
rect 5507 -3827 5573 -3815
rect 5603 -3119 5669 -3107
rect 5603 -3815 5619 -3119
rect 5653 -3815 5669 -3119
rect 5603 -3827 5669 -3815
rect 5699 -3119 5765 -3107
rect 5699 -3815 5715 -3119
rect 5749 -3815 5765 -3119
rect 5699 -3827 5765 -3815
rect 5795 -3119 5861 -3107
rect 5795 -3815 5811 -3119
rect 5845 -3815 5861 -3119
rect 5795 -3827 5861 -3815
rect 5891 -3119 5957 -3107
rect 5891 -3815 5907 -3119
rect 5941 -3815 5957 -3119
rect 5891 -3827 5957 -3815
rect 5987 -3119 6053 -3107
rect 5987 -3815 6003 -3119
rect 6037 -3815 6053 -3119
rect 5987 -3827 6053 -3815
rect 6083 -3119 6149 -3107
rect 6083 -3815 6099 -3119
rect 6133 -3815 6149 -3119
rect 6083 -3827 6149 -3815
rect 6179 -3119 6245 -3107
rect 6179 -3815 6195 -3119
rect 6229 -3815 6245 -3119
rect 6179 -3827 6245 -3815
rect 6275 -3119 6337 -3107
rect 6275 -3815 6291 -3119
rect 6325 -3815 6337 -3119
rect 6275 -3827 6337 -3815
<< ndiffc >>
rect 3219 -4570 3253 -4194
rect 3315 -4570 3349 -4194
rect 3411 -4570 3445 -4194
rect 3507 -4570 3541 -4194
rect 3603 -4570 3637 -4194
rect 3699 -4570 3733 -4194
rect 3795 -4570 3829 -4194
rect 3891 -4570 3925 -4194
rect 3987 -4570 4021 -4194
rect 4083 -4570 4117 -4194
rect 4179 -4570 4213 -4194
rect 4275 -4570 4309 -4194
rect 4371 -4570 4405 -4194
rect 4467 -4570 4501 -4194
rect 4563 -4570 4597 -4194
rect 4659 -4570 4693 -4194
rect 4755 -4570 4789 -4194
rect 4851 -4570 4885 -4194
rect 4947 -4570 4981 -4194
rect 5043 -4570 5077 -4194
rect 5139 -4570 5173 -4194
rect 5235 -4570 5269 -4194
rect 5331 -4570 5365 -4194
rect 5427 -4570 5461 -4194
rect 5523 -4570 5557 -4194
rect 5619 -4570 5653 -4194
rect 5715 -4570 5749 -4194
rect 5811 -4570 5845 -4194
rect 5907 -4570 5941 -4194
rect 6003 -4570 6037 -4194
rect 6099 -4570 6133 -4194
rect 6195 -4570 6229 -4194
rect 6291 -4570 6325 -4194
<< pdiffc >>
rect 3219 -3815 3253 -3119
rect 3315 -3815 3349 -3119
rect 3411 -3815 3445 -3119
rect 3507 -3815 3541 -3119
rect 3603 -3815 3637 -3119
rect 3699 -3815 3733 -3119
rect 3795 -3815 3829 -3119
rect 3891 -3815 3925 -3119
rect 3987 -3815 4021 -3119
rect 4083 -3815 4117 -3119
rect 4179 -3815 4213 -3119
rect 4275 -3815 4309 -3119
rect 4371 -3815 4405 -3119
rect 4467 -3815 4501 -3119
rect 4563 -3815 4597 -3119
rect 4659 -3815 4693 -3119
rect 4755 -3815 4789 -3119
rect 4851 -3815 4885 -3119
rect 4947 -3815 4981 -3119
rect 5043 -3815 5077 -3119
rect 5139 -3815 5173 -3119
rect 5235 -3815 5269 -3119
rect 5331 -3815 5365 -3119
rect 5427 -3815 5461 -3119
rect 5523 -3815 5557 -3119
rect 5619 -3815 5653 -3119
rect 5715 -3815 5749 -3119
rect 5811 -3815 5845 -3119
rect 5907 -3815 5941 -3119
rect 6003 -3815 6037 -3119
rect 6099 -3815 6133 -3119
rect 6195 -3815 6229 -3119
rect 6291 -3815 6325 -3119
<< psubdiff >>
rect 3212 -4712 3312 -4678
rect 6232 -4712 6332 -4678
<< nsubdiff >>
rect 3212 -3010 3312 -2976
rect 6232 -3010 6332 -2976
<< psubdiffcont >>
rect 3312 -4712 6232 -4678
<< nsubdiffcont >>
rect 3312 -3010 6232 -2976
<< poly >>
rect 3269 -3107 3299 -3076
rect 3365 -3107 3395 -3076
rect 3461 -3107 3491 -3076
rect 3557 -3107 3587 -3076
rect 3653 -3107 3683 -3076
rect 3749 -3107 3779 -3076
rect 3845 -3107 3875 -3076
rect 3941 -3107 3971 -3076
rect 4037 -3107 4067 -3076
rect 4133 -3107 4163 -3076
rect 4229 -3107 4259 -3076
rect 4325 -3107 4355 -3076
rect 4421 -3107 4451 -3076
rect 4517 -3107 4547 -3076
rect 4613 -3107 4643 -3076
rect 4709 -3107 4739 -3076
rect 4805 -3107 4835 -3076
rect 4901 -3107 4931 -3076
rect 4997 -3107 5027 -3076
rect 5093 -3107 5123 -3076
rect 5189 -3107 5219 -3076
rect 5285 -3107 5315 -3076
rect 5381 -3107 5411 -3076
rect 5477 -3107 5507 -3076
rect 5573 -3107 5603 -3076
rect 5669 -3107 5699 -3076
rect 5765 -3107 5795 -3076
rect 5861 -3107 5891 -3076
rect 5957 -3107 5987 -3076
rect 6053 -3107 6083 -3076
rect 6149 -3107 6179 -3076
rect 6245 -3107 6275 -3076
rect 3269 -3858 3299 -3827
rect 3365 -3858 3395 -3827
rect 3269 -3874 3395 -3858
rect 3269 -3908 3279 -3874
rect 3384 -3908 3395 -3874
rect 3269 -3924 3395 -3908
rect 3461 -3858 3491 -3827
rect 3557 -3858 3587 -3827
rect 3461 -3874 3587 -3858
rect 3461 -3908 3471 -3874
rect 3576 -3908 3587 -3874
rect 3461 -3924 3587 -3908
rect 3653 -3858 3683 -3827
rect 3749 -3858 3779 -3827
rect 3653 -3874 3779 -3858
rect 3653 -3908 3663 -3874
rect 3768 -3908 3779 -3874
rect 3653 -3924 3779 -3908
rect 3845 -3858 3875 -3827
rect 3941 -3858 3971 -3827
rect 3845 -3874 3971 -3858
rect 3845 -3908 3855 -3874
rect 3960 -3908 3971 -3874
rect 3845 -3924 3971 -3908
rect 4037 -3858 4067 -3827
rect 4133 -3858 4163 -3827
rect 4037 -3874 4163 -3858
rect 4037 -3908 4047 -3874
rect 4152 -3908 4163 -3874
rect 4037 -3924 4163 -3908
rect 4229 -3858 4259 -3827
rect 4325 -3858 4355 -3827
rect 4229 -3874 4355 -3858
rect 4229 -3908 4239 -3874
rect 4344 -3908 4355 -3874
rect 4229 -3924 4355 -3908
rect 4421 -3858 4451 -3827
rect 4517 -3858 4547 -3827
rect 4421 -3874 4547 -3858
rect 4421 -3908 4431 -3874
rect 4536 -3908 4547 -3874
rect 4421 -3924 4547 -3908
rect 4613 -3858 4643 -3827
rect 4709 -3858 4739 -3827
rect 4613 -3874 4739 -3858
rect 4613 -3908 4623 -3874
rect 4728 -3908 4739 -3874
rect 4613 -3924 4739 -3908
rect 4805 -3858 4835 -3827
rect 4901 -3858 4931 -3827
rect 4805 -3874 4931 -3858
rect 4805 -3908 4816 -3874
rect 4921 -3908 4931 -3874
rect 4805 -3924 4931 -3908
rect 4997 -3858 5027 -3827
rect 5093 -3858 5123 -3827
rect 4997 -3874 5123 -3858
rect 4997 -3908 5008 -3874
rect 5113 -3908 5123 -3874
rect 4997 -3924 5123 -3908
rect 5189 -3858 5219 -3827
rect 5285 -3858 5315 -3827
rect 5189 -3874 5315 -3858
rect 5189 -3908 5200 -3874
rect 5305 -3908 5315 -3874
rect 5189 -3924 5315 -3908
rect 5381 -3858 5411 -3827
rect 5477 -3858 5507 -3827
rect 5381 -3874 5507 -3858
rect 5381 -3908 5392 -3874
rect 5497 -3908 5507 -3874
rect 5381 -3924 5507 -3908
rect 5573 -3858 5603 -3827
rect 5669 -3858 5699 -3827
rect 5573 -3874 5699 -3858
rect 5573 -3908 5584 -3874
rect 5689 -3908 5699 -3874
rect 5573 -3924 5699 -3908
rect 5765 -3858 5795 -3827
rect 5861 -3858 5891 -3827
rect 5765 -3874 5891 -3858
rect 5765 -3908 5776 -3874
rect 5881 -3908 5891 -3874
rect 5765 -3924 5891 -3908
rect 5957 -3858 5987 -3827
rect 6053 -3858 6083 -3827
rect 5957 -3874 6083 -3858
rect 5957 -3908 5968 -3874
rect 6073 -3908 6083 -3874
rect 5957 -3924 6083 -3908
rect 6149 -3858 6179 -3827
rect 6245 -3858 6275 -3827
rect 6149 -3874 6275 -3858
rect 6149 -3908 6160 -3874
rect 6265 -3908 6275 -3874
rect 6149 -3924 6275 -3908
rect 3269 -4110 3491 -4094
rect 3269 -4144 3279 -4110
rect 3384 -4144 3491 -4110
rect 3269 -4160 3491 -4144
rect 3536 -4104 3608 -4094
rect 3536 -4138 3554 -4104
rect 3588 -4138 3608 -4104
rect 3536 -4160 3608 -4138
rect 3653 -4110 3779 -4094
rect 3653 -4144 3663 -4110
rect 3768 -4144 3779 -4110
rect 3653 -4160 3779 -4144
rect 3269 -4182 3299 -4160
rect 3365 -4182 3395 -4160
rect 3461 -4182 3491 -4160
rect 3557 -4182 3587 -4160
rect 3653 -4182 3683 -4160
rect 3749 -4182 3779 -4160
rect 3845 -4110 3971 -4094
rect 3845 -4144 3855 -4110
rect 3960 -4144 3971 -4110
rect 3845 -4160 3971 -4144
rect 3845 -4182 3875 -4160
rect 3941 -4182 3971 -4160
rect 4037 -4110 4163 -4094
rect 4037 -4144 4047 -4110
rect 4152 -4144 4163 -4110
rect 4037 -4160 4163 -4144
rect 4037 -4182 4067 -4160
rect 4133 -4182 4163 -4160
rect 4229 -4110 4355 -4094
rect 4229 -4144 4239 -4110
rect 4344 -4144 4355 -4110
rect 4229 -4160 4355 -4144
rect 4229 -4182 4259 -4160
rect 4325 -4182 4355 -4160
rect 4421 -4110 4547 -4094
rect 4421 -4144 4431 -4110
rect 4536 -4144 4547 -4110
rect 4421 -4160 4547 -4144
rect 4421 -4182 4451 -4160
rect 4517 -4182 4547 -4160
rect 4613 -4110 4739 -4094
rect 4613 -4144 4623 -4110
rect 4728 -4144 4739 -4110
rect 4613 -4160 4739 -4144
rect 4613 -4182 4643 -4160
rect 4709 -4182 4739 -4160
rect 4805 -4110 4931 -4094
rect 4805 -4144 4816 -4110
rect 4921 -4144 4931 -4110
rect 4805 -4160 4931 -4144
rect 4805 -4182 4835 -4160
rect 4901 -4182 4931 -4160
rect 4997 -4110 5123 -4094
rect 4997 -4144 5008 -4110
rect 5113 -4144 5123 -4110
rect 4997 -4160 5123 -4144
rect 4997 -4182 5027 -4160
rect 5093 -4182 5123 -4160
rect 5189 -4110 5315 -4094
rect 5189 -4144 5200 -4110
rect 5305 -4144 5315 -4110
rect 5189 -4160 5315 -4144
rect 5189 -4182 5219 -4160
rect 5285 -4182 5315 -4160
rect 5381 -4110 5507 -4094
rect 5381 -4144 5392 -4110
rect 5497 -4144 5507 -4110
rect 5381 -4160 5507 -4144
rect 5381 -4182 5411 -4160
rect 5477 -4182 5507 -4160
rect 5573 -4110 5699 -4094
rect 5573 -4144 5584 -4110
rect 5689 -4144 5699 -4110
rect 5573 -4160 5699 -4144
rect 5573 -4182 5603 -4160
rect 5669 -4182 5699 -4160
rect 5765 -4110 5891 -4094
rect 5765 -4144 5776 -4110
rect 5881 -4144 5891 -4110
rect 5765 -4160 5891 -4144
rect 5936 -4104 6008 -4094
rect 5936 -4138 5956 -4104
rect 5990 -4138 6008 -4104
rect 5936 -4160 6008 -4138
rect 6053 -4110 6275 -4094
rect 6053 -4144 6160 -4110
rect 6265 -4144 6275 -4110
rect 6053 -4160 6275 -4144
rect 5765 -4182 5795 -4160
rect 5861 -4182 5891 -4160
rect 5957 -4182 5987 -4160
rect 6053 -4182 6083 -4160
rect 6149 -4182 6179 -4160
rect 6245 -4182 6275 -4160
rect 3269 -4608 3299 -4582
rect 3365 -4608 3395 -4582
rect 3461 -4608 3491 -4582
rect 3557 -4608 3587 -4582
rect 3653 -4608 3683 -4582
rect 3749 -4608 3779 -4582
rect 3845 -4608 3875 -4582
rect 3941 -4608 3971 -4582
rect 4037 -4608 4067 -4582
rect 4133 -4608 4163 -4582
rect 4229 -4608 4259 -4582
rect 4325 -4608 4355 -4582
rect 4421 -4608 4451 -4582
rect 4517 -4608 4547 -4582
rect 4613 -4608 4643 -4582
rect 4709 -4608 4739 -4582
rect 4805 -4608 4835 -4582
rect 4901 -4608 4931 -4582
rect 4997 -4608 5027 -4582
rect 5093 -4608 5123 -4582
rect 5189 -4608 5219 -4582
rect 5285 -4608 5315 -4582
rect 5381 -4608 5411 -4582
rect 5477 -4608 5507 -4582
rect 5573 -4608 5603 -4582
rect 5669 -4608 5699 -4582
rect 5765 -4608 5795 -4582
rect 5861 -4608 5891 -4582
rect 5957 -4608 5987 -4582
rect 6053 -4608 6083 -4582
rect 6149 -4608 6179 -4582
rect 6245 -4608 6275 -4582
<< polycont >>
rect 3279 -3908 3384 -3874
rect 3471 -3908 3576 -3874
rect 3663 -3908 3768 -3874
rect 3855 -3908 3960 -3874
rect 4047 -3908 4152 -3874
rect 4239 -3908 4344 -3874
rect 4431 -3908 4536 -3874
rect 4623 -3908 4728 -3874
rect 4816 -3908 4921 -3874
rect 5008 -3908 5113 -3874
rect 5200 -3908 5305 -3874
rect 5392 -3908 5497 -3874
rect 5584 -3908 5689 -3874
rect 5776 -3908 5881 -3874
rect 5968 -3908 6073 -3874
rect 6160 -3908 6265 -3874
rect 3279 -4144 3384 -4110
rect 3554 -4138 3588 -4104
rect 3663 -4144 3768 -4110
rect 3855 -4144 3960 -4110
rect 4047 -4144 4152 -4110
rect 4239 -4144 4344 -4110
rect 4431 -4144 4536 -4110
rect 4623 -4144 4728 -4110
rect 4816 -4144 4921 -4110
rect 5008 -4144 5113 -4110
rect 5200 -4144 5305 -4110
rect 5392 -4144 5497 -4110
rect 5584 -4144 5689 -4110
rect 5776 -4144 5881 -4110
rect 5956 -4138 5990 -4104
rect 6160 -4144 6265 -4110
<< locali >>
rect 3212 -3010 3312 -2976
rect 6232 -3010 6332 -2976
rect 3219 -3119 3253 -3103
rect 3219 -3831 3253 -3815
rect 3315 -3119 3349 -3103
rect 3315 -3831 3349 -3815
rect 3411 -3119 3445 -3103
rect 3411 -3831 3445 -3815
rect 3507 -3119 3541 -3103
rect 3507 -3831 3541 -3815
rect 3603 -3119 3637 -3103
rect 3603 -3831 3637 -3815
rect 3699 -3119 3733 -3103
rect 3699 -3831 3733 -3815
rect 3795 -3119 3829 -3103
rect 3795 -3831 3829 -3815
rect 3891 -3119 3925 -3103
rect 3891 -3831 3925 -3815
rect 3987 -3119 4021 -3103
rect 3987 -3831 4021 -3815
rect 4083 -3119 4117 -3103
rect 4083 -3831 4117 -3815
rect 4179 -3119 4213 -3103
rect 4179 -3831 4213 -3815
rect 4275 -3119 4309 -3103
rect 4275 -3831 4309 -3815
rect 4371 -3119 4405 -3103
rect 4371 -3831 4405 -3815
rect 4467 -3119 4501 -3103
rect 4467 -3831 4501 -3815
rect 4563 -3119 4597 -3103
rect 4563 -3831 4597 -3815
rect 4659 -3119 4693 -3103
rect 4659 -3831 4693 -3815
rect 4755 -3119 4789 -3103
rect 4755 -3831 4789 -3815
rect 4851 -3119 4885 -3103
rect 4851 -3831 4885 -3815
rect 4947 -3119 4981 -3103
rect 4947 -3831 4981 -3815
rect 5043 -3119 5077 -3103
rect 5043 -3831 5077 -3815
rect 5139 -3119 5173 -3103
rect 5139 -3831 5173 -3815
rect 5235 -3119 5269 -3103
rect 5235 -3831 5269 -3815
rect 5331 -3119 5365 -3103
rect 5331 -3831 5365 -3815
rect 5427 -3119 5461 -3103
rect 5427 -3831 5461 -3815
rect 5523 -3119 5557 -3103
rect 5523 -3831 5557 -3815
rect 5619 -3119 5653 -3103
rect 5619 -3831 5653 -3815
rect 5715 -3119 5749 -3103
rect 5715 -3831 5749 -3815
rect 5811 -3119 5845 -3103
rect 5811 -3831 5845 -3815
rect 5907 -3119 5941 -3103
rect 5907 -3831 5941 -3815
rect 6003 -3119 6037 -3103
rect 6003 -3831 6037 -3815
rect 6099 -3119 6133 -3103
rect 6099 -3831 6133 -3815
rect 6195 -3119 6229 -3103
rect 6195 -3831 6229 -3815
rect 6291 -3119 6325 -3103
rect 6291 -3831 6325 -3815
rect 3263 -3908 3279 -3874
rect 3384 -3908 3400 -3874
rect 3455 -3908 3471 -3874
rect 3576 -3908 3592 -3874
rect 3647 -3908 3663 -3874
rect 3768 -3908 3784 -3874
rect 3839 -3908 3855 -3874
rect 3960 -3908 3976 -3874
rect 4031 -3908 4047 -3874
rect 4152 -3908 4168 -3874
rect 4223 -3908 4239 -3874
rect 4344 -3908 4360 -3874
rect 4415 -3908 4431 -3874
rect 4536 -3908 4552 -3874
rect 4607 -3908 4623 -3874
rect 4728 -3908 4744 -3874
rect 4800 -3908 4816 -3874
rect 4921 -3908 4937 -3874
rect 4992 -3908 5008 -3874
rect 5113 -3908 5129 -3874
rect 5184 -3908 5200 -3874
rect 5305 -3908 5321 -3874
rect 5376 -3908 5392 -3874
rect 5497 -3908 5513 -3874
rect 5568 -3908 5584 -3874
rect 5689 -3908 5705 -3874
rect 5760 -3908 5776 -3874
rect 5881 -3908 5897 -3874
rect 5952 -3908 5968 -3874
rect 6073 -3908 6089 -3874
rect 6144 -3908 6160 -3874
rect 6265 -3908 6281 -3874
rect 3302 -3914 3314 -3908
rect 3348 -3914 3360 -3908
rect 3302 -3924 3360 -3914
rect 3494 -3914 3506 -3908
rect 3540 -3914 3552 -3908
rect 3494 -3924 3552 -3914
rect 3686 -3914 3698 -3908
rect 3732 -3914 3744 -3908
rect 3686 -3952 3744 -3914
rect 3686 -3986 3698 -3952
rect 3732 -3986 3744 -3952
rect 3686 -3992 3744 -3986
rect 3878 -3914 3890 -3908
rect 3924 -3914 3936 -3908
rect 3878 -3952 3936 -3914
rect 3878 -3986 3890 -3952
rect 3924 -3986 3936 -3952
rect 3878 -3992 3936 -3986
rect 4070 -3914 4082 -3908
rect 4116 -3914 4128 -3908
rect 4070 -3952 4128 -3914
rect 4070 -3986 4082 -3952
rect 4116 -3986 4128 -3952
rect 4070 -3992 4128 -3986
rect 4262 -3914 4274 -3908
rect 4308 -3914 4320 -3908
rect 4262 -3952 4320 -3914
rect 4262 -3986 4274 -3952
rect 4308 -3986 4320 -3952
rect 4262 -3992 4320 -3986
rect 4454 -3914 4466 -3908
rect 4500 -3914 4512 -3908
rect 4454 -3952 4512 -3914
rect 4454 -3986 4466 -3952
rect 4500 -3986 4512 -3952
rect 4454 -3992 4512 -3986
rect 4646 -3914 4658 -3908
rect 4692 -3914 4704 -3908
rect 4646 -3952 4704 -3914
rect 4646 -3986 4658 -3952
rect 4692 -3986 4704 -3952
rect 4646 -3992 4704 -3986
rect 4840 -3914 4852 -3908
rect 4886 -3914 4898 -3908
rect 4840 -3952 4898 -3914
rect 4840 -3986 4852 -3952
rect 4886 -3986 4898 -3952
rect 4840 -3992 4898 -3986
rect 5032 -3914 5044 -3908
rect 5078 -3914 5090 -3908
rect 5032 -3952 5090 -3914
rect 5032 -3986 5044 -3952
rect 5078 -3986 5090 -3952
rect 5032 -3992 5090 -3986
rect 5224 -3914 5236 -3908
rect 5270 -3914 5282 -3908
rect 5224 -3952 5282 -3914
rect 5224 -3986 5236 -3952
rect 5270 -3986 5282 -3952
rect 5224 -3992 5282 -3986
rect 5416 -3914 5428 -3908
rect 5462 -3914 5474 -3908
rect 5416 -3952 5474 -3914
rect 5416 -3986 5428 -3952
rect 5462 -3986 5474 -3952
rect 5416 -3992 5474 -3986
rect 5608 -3914 5620 -3908
rect 5654 -3914 5666 -3908
rect 5608 -3952 5666 -3914
rect 5608 -3986 5620 -3952
rect 5654 -3986 5666 -3952
rect 5608 -3992 5666 -3986
rect 5800 -3914 5812 -3908
rect 5846 -3914 5858 -3908
rect 5800 -3952 5858 -3914
rect 5992 -3914 6004 -3908
rect 6038 -3914 6050 -3908
rect 5992 -3924 6050 -3914
rect 6184 -3914 6196 -3908
rect 6230 -3914 6242 -3908
rect 6184 -3924 6242 -3914
rect 5800 -3986 5812 -3952
rect 5846 -3986 5858 -3952
rect 5800 -3992 5858 -3986
rect 3536 -4032 3608 -4026
rect 3536 -4066 3554 -4032
rect 3588 -4066 3608 -4032
rect 3302 -4104 3360 -4094
rect 3302 -4110 3314 -4104
rect 3348 -4110 3360 -4104
rect 3536 -4104 3608 -4066
rect 3263 -4144 3279 -4110
rect 3384 -4144 3400 -4110
rect 3536 -4138 3554 -4104
rect 3588 -4138 3608 -4104
rect 3686 -4032 3744 -4026
rect 3686 -4066 3698 -4032
rect 3732 -4066 3744 -4032
rect 3686 -4104 3744 -4066
rect 3686 -4110 3698 -4104
rect 3732 -4110 3744 -4104
rect 3878 -4032 3936 -4026
rect 3878 -4066 3890 -4032
rect 3924 -4066 3936 -4032
rect 3878 -4104 3936 -4066
rect 3878 -4110 3890 -4104
rect 3924 -4110 3936 -4104
rect 4070 -4032 4128 -4026
rect 4070 -4066 4082 -4032
rect 4116 -4066 4128 -4032
rect 4070 -4104 4128 -4066
rect 4070 -4110 4082 -4104
rect 4116 -4110 4128 -4104
rect 4262 -4032 4320 -4026
rect 4262 -4066 4274 -4032
rect 4308 -4066 4320 -4032
rect 4262 -4104 4320 -4066
rect 4262 -4110 4274 -4104
rect 4308 -4110 4320 -4104
rect 4454 -4032 4512 -4026
rect 4454 -4066 4466 -4032
rect 4500 -4066 4512 -4032
rect 4454 -4104 4512 -4066
rect 4454 -4110 4466 -4104
rect 4500 -4110 4512 -4104
rect 4646 -4032 4704 -4026
rect 4646 -4066 4658 -4032
rect 4692 -4066 4704 -4032
rect 4646 -4104 4704 -4066
rect 4646 -4110 4658 -4104
rect 4692 -4110 4704 -4104
rect 4840 -4032 4898 -4026
rect 4840 -4066 4852 -4032
rect 4886 -4066 4898 -4032
rect 4840 -4104 4898 -4066
rect 4840 -4110 4852 -4104
rect 4886 -4110 4898 -4104
rect 5032 -4032 5090 -4026
rect 5032 -4066 5044 -4032
rect 5078 -4066 5090 -4032
rect 5032 -4104 5090 -4066
rect 5032 -4110 5044 -4104
rect 5078 -4110 5090 -4104
rect 5224 -4032 5282 -4026
rect 5224 -4066 5236 -4032
rect 5270 -4066 5282 -4032
rect 5224 -4104 5282 -4066
rect 5224 -4110 5236 -4104
rect 5270 -4110 5282 -4104
rect 5416 -4032 5474 -4026
rect 5416 -4066 5428 -4032
rect 5462 -4066 5474 -4032
rect 5416 -4104 5474 -4066
rect 5416 -4110 5428 -4104
rect 5462 -4110 5474 -4104
rect 5608 -4032 5666 -4026
rect 5608 -4066 5620 -4032
rect 5654 -4066 5666 -4032
rect 5608 -4104 5666 -4066
rect 5608 -4110 5620 -4104
rect 5654 -4110 5666 -4104
rect 5800 -4032 5858 -4026
rect 5800 -4066 5812 -4032
rect 5846 -4066 5858 -4032
rect 5800 -4104 5858 -4066
rect 5800 -4110 5812 -4104
rect 5846 -4110 5858 -4104
rect 5936 -4032 6008 -4026
rect 5936 -4066 5956 -4032
rect 5990 -4066 6008 -4032
rect 5936 -4104 6008 -4066
rect 3536 -4144 3608 -4138
rect 3647 -4144 3663 -4110
rect 3768 -4144 3784 -4110
rect 3839 -4144 3855 -4110
rect 3960 -4144 3976 -4110
rect 4031 -4144 4047 -4110
rect 4152 -4144 4168 -4110
rect 4223 -4144 4239 -4110
rect 4344 -4144 4360 -4110
rect 4415 -4144 4431 -4110
rect 4536 -4144 4552 -4110
rect 4607 -4144 4623 -4110
rect 4728 -4144 4744 -4110
rect 4800 -4144 4816 -4110
rect 4921 -4144 4937 -4110
rect 4992 -4144 5008 -4110
rect 5113 -4144 5129 -4110
rect 5184 -4144 5200 -4110
rect 5305 -4144 5321 -4110
rect 5376 -4144 5392 -4110
rect 5497 -4144 5513 -4110
rect 5568 -4144 5584 -4110
rect 5689 -4144 5705 -4110
rect 5760 -4144 5776 -4110
rect 5881 -4144 5897 -4110
rect 5936 -4138 5956 -4104
rect 5990 -4138 6008 -4104
rect 6184 -4104 6242 -4094
rect 6184 -4110 6196 -4104
rect 6230 -4110 6242 -4104
rect 5936 -4144 6008 -4138
rect 6144 -4144 6160 -4110
rect 6265 -4144 6281 -4110
rect 3219 -4194 3253 -4178
rect 3219 -4586 3253 -4570
rect 3315 -4194 3349 -4178
rect 3315 -4586 3349 -4570
rect 3411 -4194 3445 -4178
rect 3411 -4586 3445 -4570
rect 3507 -4194 3541 -4178
rect 3507 -4586 3541 -4570
rect 3603 -4194 3637 -4178
rect 3603 -4586 3637 -4570
rect 3699 -4194 3733 -4178
rect 3699 -4586 3733 -4570
rect 3795 -4194 3829 -4178
rect 3795 -4586 3829 -4570
rect 3891 -4194 3925 -4178
rect 3891 -4586 3925 -4570
rect 3987 -4194 4021 -4178
rect 3987 -4586 4021 -4570
rect 4083 -4194 4117 -4178
rect 4083 -4586 4117 -4570
rect 4179 -4194 4213 -4178
rect 4179 -4586 4213 -4570
rect 4275 -4194 4309 -4178
rect 4275 -4586 4309 -4570
rect 4371 -4194 4405 -4178
rect 4371 -4586 4405 -4570
rect 4467 -4194 4501 -4178
rect 4467 -4586 4501 -4570
rect 4563 -4194 4597 -4178
rect 4563 -4586 4597 -4570
rect 4659 -4194 4693 -4178
rect 4659 -4586 4693 -4570
rect 4755 -4194 4789 -4178
rect 4755 -4586 4789 -4570
rect 4851 -4194 4885 -4178
rect 4851 -4586 4885 -4570
rect 4947 -4194 4981 -4178
rect 4947 -4586 4981 -4570
rect 5043 -4194 5077 -4178
rect 5043 -4586 5077 -4570
rect 5139 -4194 5173 -4178
rect 5139 -4586 5173 -4570
rect 5235 -4194 5269 -4178
rect 5235 -4586 5269 -4570
rect 5331 -4194 5365 -4178
rect 5331 -4586 5365 -4570
rect 5427 -4194 5461 -4178
rect 5427 -4586 5461 -4570
rect 5523 -4194 5557 -4178
rect 5523 -4586 5557 -4570
rect 5619 -4194 5653 -4178
rect 5619 -4586 5653 -4570
rect 5715 -4194 5749 -4178
rect 5715 -4586 5749 -4570
rect 5811 -4194 5845 -4178
rect 5811 -4586 5845 -4570
rect 5907 -4194 5941 -4178
rect 5907 -4586 5941 -4570
rect 6003 -4194 6037 -4178
rect 6003 -4586 6037 -4570
rect 6099 -4194 6133 -4178
rect 6099 -4586 6133 -4570
rect 6195 -4194 6229 -4178
rect 6195 -4586 6229 -4570
rect 6291 -4194 6325 -4178
rect 6291 -4586 6325 -4570
rect 3212 -4712 3312 -4678
rect 6232 -4712 6332 -4678
<< viali >>
rect 3312 -3010 6232 -2976
rect 3219 -3815 3253 -3119
rect 3315 -3815 3349 -3119
rect 3411 -3815 3445 -3119
rect 3507 -3815 3541 -3119
rect 3603 -3815 3637 -3119
rect 3699 -3815 3733 -3119
rect 3795 -3815 3829 -3119
rect 3891 -3815 3925 -3119
rect 3987 -3815 4021 -3119
rect 4083 -3815 4117 -3119
rect 4179 -3815 4213 -3119
rect 4275 -3815 4309 -3119
rect 4371 -3815 4405 -3119
rect 4467 -3815 4501 -3119
rect 4563 -3815 4597 -3119
rect 4659 -3815 4693 -3119
rect 4755 -3815 4789 -3119
rect 4851 -3815 4885 -3119
rect 4947 -3815 4981 -3119
rect 5043 -3815 5077 -3119
rect 5139 -3815 5173 -3119
rect 5235 -3815 5269 -3119
rect 5331 -3815 5365 -3119
rect 5427 -3815 5461 -3119
rect 5523 -3815 5557 -3119
rect 5619 -3815 5653 -3119
rect 5715 -3815 5749 -3119
rect 5811 -3815 5845 -3119
rect 5907 -3815 5941 -3119
rect 6003 -3815 6037 -3119
rect 6099 -3815 6133 -3119
rect 6195 -3815 6229 -3119
rect 6291 -3815 6325 -3119
rect 3314 -3908 3348 -3880
rect 3506 -3908 3540 -3880
rect 3698 -3908 3732 -3880
rect 3890 -3908 3924 -3880
rect 4082 -3908 4116 -3880
rect 4274 -3908 4308 -3880
rect 4466 -3908 4500 -3880
rect 4658 -3908 4692 -3880
rect 4852 -3908 4886 -3880
rect 5044 -3908 5078 -3880
rect 5236 -3908 5270 -3880
rect 5428 -3908 5462 -3880
rect 5620 -3908 5654 -3880
rect 5812 -3908 5846 -3880
rect 6004 -3908 6038 -3880
rect 6196 -3908 6230 -3880
rect 3314 -3914 3348 -3908
rect 3506 -3914 3540 -3908
rect 3698 -3914 3732 -3908
rect 3698 -3986 3732 -3952
rect 3890 -3914 3924 -3908
rect 3890 -3986 3924 -3952
rect 4082 -3914 4116 -3908
rect 4082 -3986 4116 -3952
rect 4274 -3914 4308 -3908
rect 4274 -3986 4308 -3952
rect 4466 -3914 4500 -3908
rect 4466 -3986 4500 -3952
rect 4658 -3914 4692 -3908
rect 4658 -3986 4692 -3952
rect 4852 -3914 4886 -3908
rect 4852 -3986 4886 -3952
rect 5044 -3914 5078 -3908
rect 5044 -3986 5078 -3952
rect 5236 -3914 5270 -3908
rect 5236 -3986 5270 -3952
rect 5428 -3914 5462 -3908
rect 5428 -3986 5462 -3952
rect 5620 -3914 5654 -3908
rect 5620 -3986 5654 -3952
rect 5812 -3914 5846 -3908
rect 6004 -3914 6038 -3908
rect 6196 -3914 6230 -3908
rect 5812 -3986 5846 -3952
rect 3554 -4066 3588 -4032
rect 3314 -4110 3348 -4104
rect 3314 -4138 3348 -4110
rect 3554 -4138 3588 -4104
rect 3698 -4066 3732 -4032
rect 3698 -4110 3732 -4104
rect 3890 -4066 3924 -4032
rect 3890 -4110 3924 -4104
rect 4082 -4066 4116 -4032
rect 4082 -4110 4116 -4104
rect 4274 -4066 4308 -4032
rect 4274 -4110 4308 -4104
rect 4466 -4066 4500 -4032
rect 4466 -4110 4500 -4104
rect 4658 -4066 4692 -4032
rect 4658 -4110 4692 -4104
rect 4852 -4066 4886 -4032
rect 4852 -4110 4886 -4104
rect 5044 -4066 5078 -4032
rect 5044 -4110 5078 -4104
rect 5236 -4066 5270 -4032
rect 5236 -4110 5270 -4104
rect 5428 -4066 5462 -4032
rect 5428 -4110 5462 -4104
rect 5620 -4066 5654 -4032
rect 5620 -4110 5654 -4104
rect 5812 -4066 5846 -4032
rect 5812 -4110 5846 -4104
rect 5956 -4066 5990 -4032
rect 3698 -4138 3732 -4110
rect 3890 -4138 3924 -4110
rect 4082 -4138 4116 -4110
rect 4274 -4138 4308 -4110
rect 4466 -4138 4500 -4110
rect 4658 -4138 4692 -4110
rect 4852 -4138 4886 -4110
rect 5044 -4138 5078 -4110
rect 5236 -4138 5270 -4110
rect 5428 -4138 5462 -4110
rect 5620 -4138 5654 -4110
rect 5812 -4138 5846 -4110
rect 5956 -4138 5990 -4104
rect 6196 -4110 6230 -4104
rect 6196 -4138 6230 -4110
rect 3219 -4570 3253 -4194
rect 3315 -4570 3349 -4194
rect 3411 -4570 3445 -4194
rect 3507 -4570 3541 -4194
rect 3603 -4570 3637 -4194
rect 3699 -4570 3733 -4194
rect 3795 -4570 3829 -4194
rect 3891 -4570 3925 -4194
rect 3987 -4570 4021 -4194
rect 4083 -4570 4117 -4194
rect 4179 -4570 4213 -4194
rect 4275 -4570 4309 -4194
rect 4371 -4570 4405 -4194
rect 4467 -4570 4501 -4194
rect 4563 -4570 4597 -4194
rect 4659 -4570 4693 -4194
rect 4755 -4570 4789 -4194
rect 4851 -4570 4885 -4194
rect 4947 -4570 4981 -4194
rect 5043 -4570 5077 -4194
rect 5139 -4570 5173 -4194
rect 5235 -4570 5269 -4194
rect 5331 -4570 5365 -4194
rect 5427 -4570 5461 -4194
rect 5523 -4570 5557 -4194
rect 5619 -4570 5653 -4194
rect 5715 -4570 5749 -4194
rect 5811 -4570 5845 -4194
rect 5907 -4570 5941 -4194
rect 6003 -4570 6037 -4194
rect 6099 -4570 6133 -4194
rect 6195 -4570 6229 -4194
rect 6291 -4570 6325 -4194
rect 3312 -4712 6232 -4678
<< metal1 >>
rect 3212 -2976 6332 -2940
rect 3212 -3010 3312 -2976
rect 6232 -3010 6332 -2976
rect 3212 -3040 6332 -3010
rect 3212 -3119 3260 -3040
rect 3308 -3102 3356 -3040
rect 3212 -3815 3219 -3119
rect 3253 -3815 3260 -3119
rect 3212 -3858 3260 -3815
rect 3306 -3118 3358 -3102
rect 3306 -3830 3358 -3816
rect 3404 -3119 3452 -3040
rect 3500 -3102 3548 -3040
rect 3404 -3815 3411 -3119
rect 3445 -3815 3452 -3119
rect 3404 -3858 3452 -3815
rect 3498 -3118 3550 -3102
rect 3498 -3830 3550 -3816
rect 3596 -3119 3644 -3040
rect 3596 -3815 3603 -3119
rect 3637 -3815 3644 -3119
rect 3596 -3858 3644 -3815
rect 3690 -3118 3742 -3102
rect 3690 -3830 3742 -3816
rect 3788 -3119 3836 -3040
rect 3788 -3815 3795 -3119
rect 3829 -3815 3836 -3119
rect 3788 -3828 3836 -3815
rect 3882 -3118 3934 -3102
rect 3882 -3830 3934 -3816
rect 3980 -3119 4028 -3040
rect 3980 -3815 3987 -3119
rect 4021 -3815 4028 -3119
rect 3980 -3828 4028 -3815
rect 4074 -3118 4126 -3102
rect 4074 -3830 4126 -3816
rect 4172 -3119 4220 -3040
rect 4172 -3815 4179 -3119
rect 4213 -3815 4220 -3119
rect 4172 -3828 4220 -3815
rect 4266 -3118 4318 -3102
rect 4266 -3830 4318 -3816
rect 4364 -3119 4412 -3040
rect 4364 -3815 4371 -3119
rect 4405 -3815 4412 -3119
rect 4364 -3828 4412 -3815
rect 4458 -3118 4510 -3102
rect 4458 -3830 4510 -3816
rect 4556 -3119 4604 -3040
rect 4556 -3815 4563 -3119
rect 4597 -3815 4604 -3119
rect 4556 -3828 4604 -3815
rect 4650 -3118 4702 -3102
rect 4650 -3830 4702 -3816
rect 4748 -3119 4796 -3040
rect 4748 -3815 4755 -3119
rect 4789 -3815 4796 -3119
rect 4748 -3828 4796 -3815
rect 4842 -3119 4894 -3103
rect 4842 -3831 4894 -3817
rect 4940 -3119 4988 -3040
rect 4940 -3815 4947 -3119
rect 4981 -3815 4988 -3119
rect 4940 -3828 4988 -3815
rect 5034 -3119 5086 -3103
rect 5034 -3831 5086 -3817
rect 5132 -3119 5180 -3040
rect 5132 -3815 5139 -3119
rect 5173 -3815 5180 -3119
rect 5132 -3828 5180 -3815
rect 5226 -3119 5278 -3103
rect 5226 -3831 5278 -3817
rect 5324 -3119 5372 -3040
rect 5324 -3815 5331 -3119
rect 5365 -3815 5372 -3119
rect 5324 -3828 5372 -3815
rect 5418 -3119 5470 -3103
rect 5418 -3831 5470 -3817
rect 5516 -3119 5564 -3040
rect 5516 -3815 5523 -3119
rect 5557 -3815 5564 -3119
rect 5516 -3828 5564 -3815
rect 5610 -3119 5662 -3103
rect 5610 -3831 5662 -3817
rect 5708 -3119 5756 -3040
rect 5708 -3815 5715 -3119
rect 5749 -3815 5756 -3119
rect 5708 -3828 5756 -3815
rect 5802 -3119 5854 -3103
rect 5802 -3831 5854 -3817
rect 5900 -3119 5948 -3040
rect 5996 -3102 6044 -3040
rect 5900 -3815 5907 -3119
rect 5941 -3815 5948 -3119
rect 3212 -3880 3644 -3858
rect 5900 -3858 5948 -3815
rect 5994 -3118 6046 -3102
rect 5994 -3830 6046 -3816
rect 6092 -3119 6140 -3040
rect 6188 -3102 6236 -3040
rect 6092 -3815 6099 -3119
rect 6133 -3815 6140 -3119
rect 6092 -3858 6140 -3815
rect 6186 -3118 6238 -3102
rect 6186 -3830 6238 -3816
rect 6284 -3119 6332 -3040
rect 6284 -3815 6291 -3119
rect 6325 -3815 6332 -3119
rect 6284 -3858 6332 -3815
rect 3212 -3914 3314 -3880
rect 3348 -3914 3506 -3880
rect 3540 -3914 3644 -3880
rect 3212 -3924 3644 -3914
rect 3686 -3880 3744 -3874
rect 3686 -3914 3698 -3880
rect 3732 -3914 3744 -3880
rect 3686 -3952 3744 -3914
rect 3878 -3880 3936 -3874
rect 3878 -3914 3890 -3880
rect 3924 -3914 3936 -3880
rect 3878 -3952 3936 -3914
rect 4070 -3880 4128 -3874
rect 4070 -3914 4082 -3880
rect 4116 -3914 4128 -3880
rect 4070 -3952 4128 -3914
rect 4262 -3880 4320 -3874
rect 4262 -3914 4274 -3880
rect 4308 -3914 4320 -3880
rect 4262 -3952 4320 -3914
rect 4454 -3880 4512 -3874
rect 4454 -3914 4466 -3880
rect 4500 -3914 4512 -3880
rect 4454 -3952 4512 -3914
rect 4646 -3880 4704 -3874
rect 4646 -3914 4658 -3880
rect 4692 -3914 4704 -3880
rect 4646 -3952 4704 -3914
rect 3686 -3986 3698 -3952
rect 3732 -3986 3890 -3952
rect 3924 -3986 4082 -3952
rect 4116 -3986 4274 -3952
rect 4308 -3986 4320 -3952
rect 3536 -4006 3608 -4000
rect 3536 -4058 3544 -4006
rect 3596 -4058 3608 -4006
rect 3536 -4066 3554 -4058
rect 3588 -4066 3608 -4058
rect 3536 -4086 3608 -4066
rect 3212 -4104 3452 -4094
rect 3212 -4138 3314 -4104
rect 3348 -4138 3452 -4104
rect 3212 -4144 3452 -4138
rect 3536 -4138 3544 -4086
rect 3596 -4138 3608 -4086
rect 3536 -4144 3608 -4138
rect 3686 -4032 4320 -3986
rect 3686 -4066 3698 -4032
rect 3732 -4066 3890 -4032
rect 3924 -4066 4082 -4032
rect 4116 -4066 4274 -4032
rect 4308 -4066 4320 -4032
rect 4356 -3958 4466 -3952
rect 4356 -4028 4362 -3958
rect 4436 -3986 4466 -3958
rect 4500 -3986 4658 -3952
rect 4692 -3986 4704 -3952
rect 4436 -4028 4704 -3986
rect 4356 -4032 4704 -4028
rect 4356 -4034 4466 -4032
rect 3686 -4104 3744 -4066
rect 3686 -4138 3698 -4104
rect 3732 -4138 3744 -4104
rect 3686 -4144 3744 -4138
rect 3878 -4104 3936 -4066
rect 3878 -4138 3890 -4104
rect 3924 -4138 3936 -4104
rect 3878 -4144 3936 -4138
rect 4070 -4104 4128 -4066
rect 4070 -4138 4082 -4104
rect 4116 -4138 4128 -4104
rect 4070 -4144 4128 -4138
rect 4262 -4072 4320 -4066
rect 4454 -4066 4466 -4034
rect 4500 -4066 4658 -4032
rect 4692 -4066 4704 -4032
rect 4262 -4078 4420 -4072
rect 4262 -4104 4356 -4078
rect 4262 -4138 4274 -4104
rect 4308 -4138 4356 -4104
rect 4262 -4140 4356 -4138
rect 4262 -4144 4420 -4140
rect 4454 -4104 4512 -4066
rect 4454 -4138 4466 -4104
rect 4500 -4138 4512 -4104
rect 4454 -4144 4512 -4138
rect 4646 -4104 4704 -4066
rect 4646 -4138 4658 -4104
rect 4692 -4138 4704 -4104
rect 4646 -4144 4704 -4138
rect 4840 -3880 4898 -3874
rect 4840 -3914 4852 -3880
rect 4886 -3914 4898 -3880
rect 4840 -3952 4898 -3914
rect 5032 -3880 5090 -3874
rect 5032 -3914 5044 -3880
rect 5078 -3914 5090 -3880
rect 5032 -3952 5090 -3914
rect 5224 -3880 5282 -3874
rect 5224 -3914 5236 -3880
rect 5270 -3914 5282 -3880
rect 5224 -3952 5282 -3914
rect 5416 -3880 5474 -3874
rect 5416 -3914 5428 -3880
rect 5462 -3914 5474 -3880
rect 5416 -3952 5474 -3914
rect 5608 -3880 5666 -3874
rect 5608 -3914 5620 -3880
rect 5654 -3914 5666 -3880
rect 5608 -3952 5666 -3914
rect 5800 -3880 5858 -3874
rect 5800 -3914 5812 -3880
rect 5846 -3914 5858 -3880
rect 5800 -3952 5858 -3914
rect 5900 -3880 6332 -3858
rect 5900 -3914 6004 -3880
rect 6038 -3914 6196 -3880
rect 6230 -3914 6332 -3880
rect 5900 -3924 6332 -3914
rect 4840 -3986 4852 -3952
rect 4886 -3986 5044 -3952
rect 5078 -3958 5188 -3952
rect 5078 -3986 5108 -3958
rect 4840 -4028 5108 -3986
rect 5182 -4028 5188 -3958
rect 4840 -4032 5188 -4028
rect 4840 -4066 4852 -4032
rect 4886 -4066 5044 -4032
rect 5078 -4034 5188 -4032
rect 5224 -3986 5236 -3952
rect 5270 -3986 5428 -3952
rect 5462 -3986 5620 -3952
rect 5654 -3986 5812 -3952
rect 5846 -3986 5858 -3952
rect 5224 -4032 5858 -3986
rect 5078 -4066 5090 -4034
rect 4840 -4104 4898 -4066
rect 4840 -4138 4852 -4104
rect 4886 -4138 4898 -4104
rect 4840 -4144 4898 -4138
rect 5032 -4104 5090 -4066
rect 5224 -4066 5236 -4032
rect 5270 -4066 5428 -4032
rect 5462 -4066 5620 -4032
rect 5654 -4066 5812 -4032
rect 5846 -4066 5858 -4032
rect 5224 -4072 5282 -4066
rect 5032 -4138 5044 -4104
rect 5078 -4138 5090 -4104
rect 5032 -4144 5090 -4138
rect 5124 -4078 5282 -4072
rect 5188 -4104 5282 -4078
rect 5188 -4138 5236 -4104
rect 5270 -4138 5282 -4104
rect 5188 -4140 5282 -4138
rect 5124 -4144 5282 -4140
rect 5416 -4104 5474 -4066
rect 5416 -4138 5428 -4104
rect 5462 -4138 5474 -4104
rect 5416 -4144 5474 -4138
rect 5608 -4104 5666 -4066
rect 5608 -4138 5620 -4104
rect 5654 -4138 5666 -4104
rect 5608 -4144 5666 -4138
rect 5800 -4104 5858 -4066
rect 5800 -4138 5812 -4104
rect 5846 -4138 5858 -4104
rect 5800 -4144 5858 -4138
rect 5936 -4006 6008 -4000
rect 5936 -4058 5948 -4006
rect 6000 -4058 6008 -4006
rect 5936 -4066 5956 -4058
rect 5990 -4066 6008 -4058
rect 5936 -4086 6008 -4066
rect 5936 -4138 5948 -4086
rect 6000 -4138 6008 -4086
rect 5936 -4144 6008 -4138
rect 6092 -4104 6332 -4094
rect 6092 -4138 6196 -4104
rect 6230 -4138 6332 -4104
rect 6092 -4144 6332 -4138
rect 3212 -4194 3260 -4144
rect 3212 -4570 3219 -4194
rect 3253 -4570 3260 -4194
rect 3212 -4648 3260 -4570
rect 3306 -4194 3358 -4178
rect 3306 -4586 3358 -4572
rect 3404 -4194 3452 -4144
rect 4356 -4154 4420 -4144
rect 5124 -4146 5224 -4144
rect 3404 -4570 3411 -4194
rect 3445 -4570 3452 -4194
rect 3308 -4648 3356 -4586
rect 3404 -4648 3452 -4570
rect 3498 -4194 3550 -4178
rect 3498 -4586 3550 -4572
rect 3596 -4194 3644 -4182
rect 3596 -4570 3603 -4194
rect 3637 -4570 3644 -4194
rect 3596 -4648 3644 -4570
rect 3690 -4194 3742 -4178
rect 3690 -4586 3742 -4572
rect 3788 -4194 3836 -4182
rect 3788 -4570 3795 -4194
rect 3829 -4570 3836 -4194
rect 3788 -4648 3836 -4570
rect 3882 -4194 3934 -4178
rect 3882 -4586 3934 -4572
rect 3980 -4194 4028 -4182
rect 3980 -4570 3987 -4194
rect 4021 -4570 4028 -4194
rect 3980 -4648 4028 -4570
rect 4074 -4194 4126 -4178
rect 4074 -4586 4126 -4572
rect 4172 -4194 4220 -4182
rect 4172 -4570 4179 -4194
rect 4213 -4570 4220 -4194
rect 4172 -4648 4220 -4570
rect 4266 -4194 4318 -4178
rect 4266 -4586 4318 -4572
rect 4364 -4194 4412 -4182
rect 4364 -4570 4371 -4194
rect 4405 -4570 4412 -4194
rect 4364 -4648 4412 -4570
rect 4458 -4194 4510 -4178
rect 4458 -4586 4510 -4572
rect 4556 -4194 4604 -4182
rect 4556 -4570 4563 -4194
rect 4597 -4570 4604 -4194
rect 4556 -4648 4604 -4570
rect 4650 -4194 4702 -4178
rect 4650 -4586 4702 -4572
rect 4748 -4194 4796 -4182
rect 4748 -4570 4755 -4194
rect 4789 -4570 4796 -4194
rect 4748 -4648 4796 -4570
rect 4842 -4194 4894 -4178
rect 4842 -4586 4894 -4572
rect 4940 -4194 4988 -4182
rect 4940 -4570 4947 -4194
rect 4981 -4570 4988 -4194
rect 4940 -4648 4988 -4570
rect 5034 -4194 5086 -4178
rect 5034 -4586 5086 -4572
rect 5132 -4194 5180 -4182
rect 5132 -4570 5139 -4194
rect 5173 -4570 5180 -4194
rect 5132 -4648 5180 -4570
rect 5226 -4194 5278 -4178
rect 5226 -4586 5278 -4572
rect 5324 -4194 5372 -4182
rect 5324 -4570 5331 -4194
rect 5365 -4570 5372 -4194
rect 5324 -4648 5372 -4570
rect 5418 -4194 5470 -4178
rect 5418 -4586 5470 -4572
rect 5516 -4194 5564 -4182
rect 5516 -4570 5523 -4194
rect 5557 -4570 5564 -4194
rect 5516 -4648 5564 -4570
rect 5610 -4194 5662 -4178
rect 5610 -4586 5662 -4572
rect 5708 -4194 5756 -4182
rect 5708 -4570 5715 -4194
rect 5749 -4570 5756 -4194
rect 5708 -4648 5756 -4570
rect 5802 -4194 5854 -4178
rect 5802 -4586 5854 -4572
rect 5900 -4194 5948 -4182
rect 5900 -4570 5907 -4194
rect 5941 -4570 5948 -4194
rect 5900 -4648 5948 -4570
rect 5994 -4194 6046 -4178
rect 5994 -4586 6046 -4572
rect 6092 -4194 6140 -4144
rect 6092 -4570 6099 -4194
rect 6133 -4570 6140 -4194
rect 6092 -4648 6140 -4570
rect 6186 -4194 6238 -4178
rect 6186 -4586 6238 -4572
rect 6284 -4194 6332 -4144
rect 6284 -4570 6291 -4194
rect 6325 -4570 6332 -4194
rect 6188 -4648 6236 -4586
rect 6284 -4648 6332 -4570
rect 3212 -4678 6332 -4648
rect 3212 -4712 3312 -4678
rect 6232 -4712 6332 -4678
rect 3212 -4728 6332 -4712
<< via1 >>
rect 3306 -3119 3358 -3118
rect 3306 -3815 3315 -3119
rect 3315 -3815 3349 -3119
rect 3349 -3815 3358 -3119
rect 3306 -3816 3358 -3815
rect 3498 -3119 3550 -3118
rect 3498 -3815 3507 -3119
rect 3507 -3815 3541 -3119
rect 3541 -3815 3550 -3119
rect 3498 -3816 3550 -3815
rect 3690 -3119 3742 -3118
rect 3690 -3815 3699 -3119
rect 3699 -3815 3733 -3119
rect 3733 -3815 3742 -3119
rect 3690 -3816 3742 -3815
rect 3882 -3119 3934 -3118
rect 3882 -3815 3891 -3119
rect 3891 -3815 3925 -3119
rect 3925 -3815 3934 -3119
rect 3882 -3816 3934 -3815
rect 4074 -3119 4126 -3118
rect 4074 -3815 4083 -3119
rect 4083 -3815 4117 -3119
rect 4117 -3815 4126 -3119
rect 4074 -3816 4126 -3815
rect 4266 -3119 4318 -3118
rect 4266 -3815 4275 -3119
rect 4275 -3815 4309 -3119
rect 4309 -3815 4318 -3119
rect 4266 -3816 4318 -3815
rect 4458 -3119 4510 -3118
rect 4458 -3815 4467 -3119
rect 4467 -3815 4501 -3119
rect 4501 -3815 4510 -3119
rect 4458 -3816 4510 -3815
rect 4650 -3119 4702 -3118
rect 4650 -3815 4659 -3119
rect 4659 -3815 4693 -3119
rect 4693 -3815 4702 -3119
rect 4650 -3816 4702 -3815
rect 4842 -3815 4851 -3119
rect 4851 -3815 4885 -3119
rect 4885 -3815 4894 -3119
rect 4842 -3817 4894 -3815
rect 5034 -3815 5043 -3119
rect 5043 -3815 5077 -3119
rect 5077 -3815 5086 -3119
rect 5034 -3817 5086 -3815
rect 5226 -3815 5235 -3119
rect 5235 -3815 5269 -3119
rect 5269 -3815 5278 -3119
rect 5226 -3817 5278 -3815
rect 5418 -3815 5427 -3119
rect 5427 -3815 5461 -3119
rect 5461 -3815 5470 -3119
rect 5418 -3817 5470 -3815
rect 5610 -3815 5619 -3119
rect 5619 -3815 5653 -3119
rect 5653 -3815 5662 -3119
rect 5610 -3817 5662 -3815
rect 5802 -3815 5811 -3119
rect 5811 -3815 5845 -3119
rect 5845 -3815 5854 -3119
rect 5802 -3817 5854 -3815
rect 5994 -3119 6046 -3118
rect 5994 -3815 6003 -3119
rect 6003 -3815 6037 -3119
rect 6037 -3815 6046 -3119
rect 5994 -3816 6046 -3815
rect 6186 -3119 6238 -3118
rect 6186 -3815 6195 -3119
rect 6195 -3815 6229 -3119
rect 6229 -3815 6238 -3119
rect 6186 -3816 6238 -3815
rect 3544 -4032 3596 -4006
rect 3544 -4058 3554 -4032
rect 3554 -4058 3588 -4032
rect 3588 -4058 3596 -4032
rect 3544 -4104 3596 -4086
rect 3544 -4138 3554 -4104
rect 3554 -4138 3588 -4104
rect 3588 -4138 3596 -4104
rect 4362 -4028 4436 -3958
rect 4356 -4140 4420 -4078
rect 5108 -4028 5182 -3958
rect 5124 -4140 5188 -4078
rect 5948 -4032 6000 -4006
rect 5948 -4058 5956 -4032
rect 5956 -4058 5990 -4032
rect 5990 -4058 6000 -4032
rect 5948 -4104 6000 -4086
rect 5948 -4138 5956 -4104
rect 5956 -4138 5990 -4104
rect 5990 -4138 6000 -4104
rect 3306 -4570 3315 -4194
rect 3315 -4570 3349 -4194
rect 3349 -4570 3358 -4194
rect 3306 -4572 3358 -4570
rect 3498 -4570 3507 -4194
rect 3507 -4570 3541 -4194
rect 3541 -4570 3550 -4194
rect 3498 -4572 3550 -4570
rect 3690 -4570 3699 -4194
rect 3699 -4570 3733 -4194
rect 3733 -4570 3742 -4194
rect 3690 -4572 3742 -4570
rect 3882 -4570 3891 -4194
rect 3891 -4570 3925 -4194
rect 3925 -4570 3934 -4194
rect 3882 -4572 3934 -4570
rect 4074 -4570 4083 -4194
rect 4083 -4570 4117 -4194
rect 4117 -4570 4126 -4194
rect 4074 -4572 4126 -4570
rect 4266 -4570 4275 -4194
rect 4275 -4570 4309 -4194
rect 4309 -4570 4318 -4194
rect 4266 -4572 4318 -4570
rect 4458 -4570 4467 -4194
rect 4467 -4570 4501 -4194
rect 4501 -4570 4510 -4194
rect 4458 -4572 4510 -4570
rect 4650 -4570 4659 -4194
rect 4659 -4570 4693 -4194
rect 4693 -4570 4702 -4194
rect 4650 -4572 4702 -4570
rect 4842 -4570 4851 -4194
rect 4851 -4570 4885 -4194
rect 4885 -4570 4894 -4194
rect 4842 -4572 4894 -4570
rect 5034 -4570 5043 -4194
rect 5043 -4570 5077 -4194
rect 5077 -4570 5086 -4194
rect 5034 -4572 5086 -4570
rect 5226 -4570 5235 -4194
rect 5235 -4570 5269 -4194
rect 5269 -4570 5278 -4194
rect 5226 -4572 5278 -4570
rect 5418 -4570 5427 -4194
rect 5427 -4570 5461 -4194
rect 5461 -4570 5470 -4194
rect 5418 -4572 5470 -4570
rect 5610 -4570 5619 -4194
rect 5619 -4570 5653 -4194
rect 5653 -4570 5662 -4194
rect 5610 -4572 5662 -4570
rect 5802 -4570 5811 -4194
rect 5811 -4570 5845 -4194
rect 5845 -4570 5854 -4194
rect 5802 -4572 5854 -4570
rect 5994 -4570 6003 -4194
rect 6003 -4570 6037 -4194
rect 6037 -4570 6046 -4194
rect 5994 -4572 6046 -4570
rect 6186 -4570 6195 -4194
rect 6195 -4570 6229 -4194
rect 6229 -4570 6238 -4194
rect 6186 -4572 6238 -4570
<< metal2 >>
rect 3303 -3118 3360 -3102
rect 3303 -3830 3360 -3816
rect 3495 -3118 3552 -3102
rect 3495 -3830 3552 -3816
rect 3687 -3118 3744 -3102
rect 3687 -3830 3744 -3816
rect 3879 -3118 3936 -3102
rect 3879 -3830 3936 -3816
rect 4071 -3118 4128 -3102
rect 4071 -3830 4128 -3816
rect 4263 -3118 4320 -3102
rect 4263 -3830 4320 -3816
rect 4455 -3118 4512 -3102
rect 4455 -3830 4512 -3816
rect 4647 -3118 4704 -3102
rect 4647 -3830 4704 -3816
rect 4840 -3119 4897 -3103
rect 4840 -3831 4897 -3817
rect 5032 -3119 5089 -3103
rect 5032 -3831 5089 -3817
rect 5224 -3119 5281 -3103
rect 5224 -3831 5281 -3817
rect 5416 -3119 5473 -3103
rect 5416 -3831 5473 -3817
rect 5608 -3119 5665 -3103
rect 5608 -3831 5665 -3817
rect 5800 -3119 5857 -3103
rect 5800 -3831 5857 -3817
rect 5992 -3118 6049 -3102
rect 5992 -3830 6049 -3816
rect 6184 -3118 6241 -3102
rect 6184 -3830 6241 -3816
rect 4352 -3958 4446 -3948
rect 3536 -4006 3608 -4000
rect 3536 -4058 3544 -4006
rect 3596 -4058 3608 -4006
rect 4352 -4028 4362 -3958
rect 4436 -4028 4446 -3958
rect 4352 -4038 4446 -4028
rect 5098 -3958 5192 -3948
rect 5098 -4028 5108 -3958
rect 5182 -4028 5192 -3958
rect 5098 -4038 5192 -4028
rect 5936 -4006 6008 -4000
rect 3536 -4072 3608 -4058
rect 5936 -4058 5948 -4006
rect 6000 -4058 6008 -4006
rect 5936 -4072 6008 -4058
rect 3396 -4086 3608 -4072
rect 3396 -4138 3544 -4086
rect 3596 -4138 3608 -4086
rect 3396 -4140 3608 -4138
rect 3303 -4194 3360 -4178
rect 3303 -4586 3360 -4572
rect 3396 -4868 3460 -4140
rect 3495 -4144 3608 -4140
rect 4356 -4078 4420 -4072
rect 3495 -4194 3552 -4178
rect 3495 -4586 3552 -4572
rect 3687 -4194 3744 -4178
rect 3687 -4586 3744 -4572
rect 3879 -4194 3936 -4178
rect 3879 -4586 3936 -4572
rect 4071 -4194 4128 -4178
rect 4071 -4586 4128 -4572
rect 4263 -4194 4320 -4178
rect 4263 -4586 4320 -4572
rect 4356 -4868 4420 -4140
rect 5124 -4078 5188 -4072
rect 4455 -4194 4512 -4178
rect 4455 -4586 4512 -4572
rect 4647 -4194 4704 -4178
rect 4647 -4586 4704 -4572
rect 4840 -4194 4897 -4178
rect 4840 -4586 4897 -4572
rect 5032 -4194 5089 -4178
rect 5032 -4586 5089 -4572
rect 5124 -4868 5188 -4140
rect 5936 -4086 6148 -4072
rect 5936 -4138 5948 -4086
rect 6000 -4138 6148 -4086
rect 5936 -4140 6148 -4138
rect 5936 -4144 6049 -4140
rect 5224 -4194 5281 -4178
rect 5224 -4586 5281 -4572
rect 5416 -4194 5473 -4178
rect 5416 -4586 5473 -4572
rect 5608 -4194 5665 -4178
rect 5608 -4586 5665 -4572
rect 5800 -4194 5857 -4178
rect 5800 -4586 5857 -4572
rect 5992 -4194 6049 -4178
rect 5992 -4586 6049 -4572
rect 6084 -4868 6148 -4140
rect 6184 -4194 6241 -4178
rect 6184 -4586 6241 -4572
rect 3394 -4874 3462 -4868
rect 3394 -4930 3400 -4874
rect 3456 -4930 3462 -4874
rect 3394 -4956 3462 -4930
rect 3394 -5012 3400 -4956
rect 3456 -5012 3462 -4956
rect 3394 -5032 3462 -5012
rect 4354 -4874 4422 -4868
rect 4354 -4930 4360 -4874
rect 4416 -4930 4422 -4874
rect 4354 -4956 4422 -4930
rect 4354 -5012 4360 -4956
rect 4416 -5012 4422 -4956
rect 4354 -5032 4422 -5012
rect 5122 -4874 5190 -4868
rect 5122 -4930 5128 -4874
rect 5184 -4930 5190 -4874
rect 5122 -4956 5190 -4930
rect 5122 -5012 5128 -4956
rect 5184 -5012 5190 -4956
rect 5122 -5032 5190 -5012
rect 6082 -4874 6150 -4868
rect 6082 -4930 6088 -4874
rect 6144 -4930 6150 -4874
rect 6082 -4956 6150 -4930
rect 6082 -5012 6088 -4956
rect 6144 -5012 6150 -4956
rect 6082 -5032 6150 -5012
<< via2 >>
rect 3303 -3816 3306 -3118
rect 3306 -3816 3358 -3118
rect 3358 -3816 3360 -3118
rect 3495 -3816 3498 -3118
rect 3498 -3816 3550 -3118
rect 3550 -3816 3552 -3118
rect 3687 -3816 3690 -3118
rect 3690 -3816 3742 -3118
rect 3742 -3816 3744 -3118
rect 3879 -3816 3882 -3118
rect 3882 -3816 3934 -3118
rect 3934 -3816 3936 -3118
rect 4071 -3816 4074 -3118
rect 4074 -3816 4126 -3118
rect 4126 -3816 4128 -3118
rect 4263 -3816 4266 -3118
rect 4266 -3816 4318 -3118
rect 4318 -3816 4320 -3118
rect 4455 -3816 4458 -3118
rect 4458 -3816 4510 -3118
rect 4510 -3816 4512 -3118
rect 4647 -3816 4650 -3118
rect 4650 -3816 4702 -3118
rect 4702 -3816 4704 -3118
rect 4840 -3817 4842 -3119
rect 4842 -3817 4894 -3119
rect 4894 -3817 4897 -3119
rect 5032 -3817 5034 -3119
rect 5034 -3817 5086 -3119
rect 5086 -3817 5089 -3119
rect 5224 -3817 5226 -3119
rect 5226 -3817 5278 -3119
rect 5278 -3817 5281 -3119
rect 5416 -3817 5418 -3119
rect 5418 -3817 5470 -3119
rect 5470 -3817 5473 -3119
rect 5608 -3817 5610 -3119
rect 5610 -3817 5662 -3119
rect 5662 -3817 5665 -3119
rect 5800 -3817 5802 -3119
rect 5802 -3817 5854 -3119
rect 5854 -3817 5857 -3119
rect 5992 -3816 5994 -3118
rect 5994 -3816 6046 -3118
rect 6046 -3816 6049 -3118
rect 6184 -3816 6186 -3118
rect 6186 -3816 6238 -3118
rect 6238 -3816 6241 -3118
rect 4362 -4028 4436 -3958
rect 5108 -4028 5182 -3958
rect 3303 -4572 3306 -4194
rect 3306 -4572 3358 -4194
rect 3358 -4572 3360 -4194
rect 3495 -4572 3498 -4194
rect 3498 -4572 3550 -4194
rect 3550 -4572 3552 -4194
rect 3687 -4572 3690 -4194
rect 3690 -4572 3742 -4194
rect 3742 -4572 3744 -4194
rect 3879 -4572 3882 -4194
rect 3882 -4572 3934 -4194
rect 3934 -4572 3936 -4194
rect 4071 -4572 4074 -4194
rect 4074 -4572 4126 -4194
rect 4126 -4572 4128 -4194
rect 4263 -4572 4266 -4194
rect 4266 -4572 4318 -4194
rect 4318 -4572 4320 -4194
rect 4455 -4572 4458 -4194
rect 4458 -4572 4510 -4194
rect 4510 -4572 4512 -4194
rect 4647 -4572 4650 -4194
rect 4650 -4572 4702 -4194
rect 4702 -4572 4704 -4194
rect 4840 -4572 4842 -4194
rect 4842 -4572 4894 -4194
rect 4894 -4572 4897 -4194
rect 5032 -4572 5034 -4194
rect 5034 -4572 5086 -4194
rect 5086 -4572 5089 -4194
rect 5224 -4572 5226 -4194
rect 5226 -4572 5278 -4194
rect 5278 -4572 5281 -4194
rect 5416 -4572 5418 -4194
rect 5418 -4572 5470 -4194
rect 5470 -4572 5473 -4194
rect 5608 -4572 5610 -4194
rect 5610 -4572 5662 -4194
rect 5662 -4572 5665 -4194
rect 5800 -4572 5802 -4194
rect 5802 -4572 5854 -4194
rect 5854 -4572 5857 -4194
rect 5992 -4572 5994 -4194
rect 5994 -4572 6046 -4194
rect 6046 -4572 6049 -4194
rect 6184 -4572 6186 -4194
rect 6186 -4572 6238 -4194
rect 6238 -4572 6241 -4194
rect 3400 -4930 3456 -4874
rect 3400 -5012 3456 -4956
rect 4360 -4930 4416 -4874
rect 4360 -5012 4416 -4956
rect 5128 -4930 5184 -4874
rect 5128 -5012 5184 -4956
rect 6088 -4930 6144 -4874
rect 6088 -5012 6144 -4956
<< metal3 >>
rect 3298 -3118 3366 -3102
rect 3298 -3816 3303 -3118
rect 3360 -3816 3366 -3118
rect 3298 -3830 3366 -3816
rect 3490 -3118 3558 -3102
rect 3490 -3816 3495 -3118
rect 3552 -3816 3558 -3118
rect 3490 -3830 3558 -3816
rect 3682 -3118 3750 -3102
rect 3682 -3816 3687 -3118
rect 3744 -3816 3750 -3118
rect 3298 -4194 3366 -4178
rect 3298 -4572 3303 -4194
rect 3360 -4572 3366 -4194
rect 3298 -4586 3366 -4572
rect 3490 -4194 3558 -4178
rect 3490 -4572 3495 -4194
rect 3552 -4572 3558 -4194
rect 3490 -4748 3558 -4572
rect 3682 -4194 3750 -3816
rect 3682 -4572 3687 -4194
rect 3744 -4572 3750 -4194
rect 3490 -4808 3586 -4748
rect 3682 -4808 3750 -4572
rect 3874 -3118 3942 -3102
rect 3874 -3816 3879 -3118
rect 3936 -3816 3942 -3118
rect 3874 -4194 3942 -3816
rect 3874 -4572 3879 -4194
rect 3936 -4572 3942 -4194
rect 3874 -4808 3942 -4572
rect 4066 -3118 4134 -3102
rect 4066 -3816 4071 -3118
rect 4128 -3816 4134 -3118
rect 4066 -4194 4134 -3816
rect 4066 -4572 4071 -4194
rect 4128 -4572 4134 -4194
rect 4066 -4808 4134 -4572
rect 4258 -3118 4326 -3102
rect 4258 -3816 4263 -3118
rect 4320 -3816 4326 -3118
rect 4258 -3948 4326 -3816
rect 4450 -3118 4518 -3102
rect 4450 -3816 4455 -3118
rect 4512 -3776 4518 -3118
rect 4642 -3118 4710 -3102
rect 4512 -3816 4582 -3776
rect 4450 -3836 4582 -3816
rect 4258 -3958 4446 -3948
rect 4258 -4028 4362 -3958
rect 4436 -4028 4446 -3958
rect 4258 -4038 4446 -4028
rect 4258 -4194 4326 -4038
rect 4514 -4182 4582 -3836
rect 4258 -4572 4263 -4194
rect 4320 -4572 4326 -4194
rect 4258 -4748 4326 -4572
rect 4230 -4808 4326 -4748
rect 4450 -4194 4582 -4182
rect 4450 -4572 4455 -4194
rect 4512 -4244 4582 -4194
rect 4642 -3816 4647 -3118
rect 4704 -3816 4710 -3118
rect 4642 -4194 4710 -3816
rect 4512 -4572 4518 -4244
rect 4450 -4748 4518 -4572
rect 4642 -4572 4647 -4194
rect 4704 -4572 4710 -4194
rect 4450 -4808 4546 -4748
rect 4642 -4808 4710 -4572
rect 3390 -4874 3466 -4868
rect 3390 -4930 3400 -4874
rect 3456 -4930 3466 -4874
rect 3526 -4914 4290 -4808
rect 4350 -4874 4426 -4868
rect 3390 -4956 3466 -4930
rect 3390 -5012 3400 -4956
rect 3456 -5012 3466 -4956
rect 3390 -5032 3466 -5012
rect 4066 -5032 4134 -4914
rect 4350 -4930 4360 -4874
rect 4416 -4930 4426 -4874
rect 4486 -4914 4710 -4808
rect 4350 -4956 4426 -4930
rect 4350 -5012 4360 -4956
rect 4416 -5012 4426 -4956
rect 4350 -5032 4426 -5012
rect 4642 -5034 4710 -4914
rect 4834 -3119 4902 -3103
rect 4834 -3817 4840 -3119
rect 4897 -3817 4902 -3119
rect 5026 -3119 5094 -3103
rect 5026 -3776 5032 -3119
rect 4834 -4194 4902 -3817
rect 4834 -4572 4840 -4194
rect 4897 -4572 4902 -4194
rect 4962 -3817 5032 -3776
rect 5089 -3817 5094 -3119
rect 4962 -3836 5094 -3817
rect 5218 -3119 5286 -3103
rect 5218 -3817 5224 -3119
rect 5281 -3817 5286 -3119
rect 4962 -4182 5030 -3836
rect 5218 -3948 5286 -3817
rect 5098 -3958 5286 -3948
rect 5098 -4028 5108 -3958
rect 5182 -4028 5286 -3958
rect 5098 -4038 5286 -4028
rect 4962 -4194 5094 -4182
rect 4962 -4244 5032 -4194
rect 4834 -4808 4902 -4572
rect 5026 -4572 5032 -4244
rect 5089 -4572 5094 -4194
rect 5026 -4748 5094 -4572
rect 4998 -4808 5094 -4748
rect 5218 -4194 5286 -4038
rect 5218 -4572 5224 -4194
rect 5281 -4572 5286 -4194
rect 5218 -4748 5286 -4572
rect 5410 -3119 5478 -3103
rect 5410 -3817 5416 -3119
rect 5473 -3817 5478 -3119
rect 5410 -4194 5478 -3817
rect 5410 -4572 5416 -4194
rect 5473 -4572 5478 -4194
rect 5218 -4808 5314 -4748
rect 5410 -4808 5478 -4572
rect 5602 -3119 5670 -3103
rect 5602 -3817 5608 -3119
rect 5665 -3817 5670 -3119
rect 5602 -4194 5670 -3817
rect 5602 -4572 5608 -4194
rect 5665 -4572 5670 -4194
rect 5602 -4808 5670 -4572
rect 5794 -3119 5862 -3103
rect 5794 -3817 5800 -3119
rect 5857 -3817 5862 -3119
rect 5794 -4194 5862 -3817
rect 5986 -3118 6054 -3102
rect 5986 -3816 5992 -3118
rect 6049 -3816 6054 -3118
rect 5986 -3924 6054 -3816
rect 6178 -3118 6246 -3102
rect 6178 -3816 6184 -3118
rect 6241 -3816 6246 -3118
rect 6178 -3924 6246 -3816
rect 5794 -4572 5800 -4194
rect 5857 -4572 5862 -4194
rect 5794 -4808 5862 -4572
rect 5986 -4194 6054 -4178
rect 5986 -4572 5992 -4194
rect 6049 -4572 6054 -4194
rect 5986 -4748 6054 -4572
rect 6178 -4194 6246 -4178
rect 6178 -4572 6184 -4194
rect 6241 -4572 6246 -4194
rect 6178 -4586 6246 -4572
rect 5958 -4808 6054 -4748
rect 4834 -4914 5058 -4808
rect 5118 -4874 5194 -4868
rect 4834 -5034 4902 -4914
rect 5118 -4930 5128 -4874
rect 5184 -4930 5194 -4874
rect 5254 -4914 6018 -4808
rect 6078 -4874 6154 -4868
rect 5118 -4956 5194 -4930
rect 5118 -5012 5128 -4956
rect 5184 -5012 5194 -4956
rect 5118 -5032 5194 -5012
rect 5410 -5032 5478 -4914
rect 6078 -4930 6088 -4874
rect 6144 -4930 6154 -4874
rect 6078 -4956 6154 -4930
rect 6078 -5012 6088 -4956
rect 6144 -5012 6154 -4956
rect 6078 -5032 6154 -5012
<< comment >>
rect 3260 -3040 3274 -3010
rect 3452 -3040 3466 -3010
rect 6078 -3040 6092 -3010
rect 6270 -3040 6284 -3010
<< end >>
