magic
tech sky130A
timestamp 1671210538
<< pwell >>
rect -889 -467 889 467
<< psubdiff >>
rect -871 432 -823 449
rect 823 432 871 449
rect -871 401 -854 432
rect 854 401 871 432
rect -871 -432 -854 -401
rect 854 -432 871 -401
rect -871 -449 -823 -432
rect 823 -449 871 -432
<< psubdiffcont >>
rect -823 432 823 449
rect -871 -401 -854 401
rect 854 -401 871 401
rect -823 -449 823 -432
<< xpolycontact >>
rect -806 -384 -771 -168
rect 771 -384 806 -168
<< xpolyres >>
rect -806 349 -688 384
rect -806 -168 -771 349
rect -723 -81 -688 349
rect -640 349 -522 384
rect -640 -81 -605 349
rect -723 -116 -605 -81
rect -557 -81 -522 349
rect -474 349 -356 384
rect -474 -81 -439 349
rect -557 -116 -439 -81
rect -391 -81 -356 349
rect -308 349 -190 384
rect -308 -81 -273 349
rect -391 -116 -273 -81
rect -225 -81 -190 349
rect -142 349 -24 384
rect -142 -81 -107 349
rect -225 -116 -107 -81
rect -59 -81 -24 349
rect 24 349 142 384
rect 24 -81 59 349
rect -59 -116 59 -81
rect 107 -81 142 349
rect 190 349 308 384
rect 190 -81 225 349
rect 107 -116 225 -81
rect 273 -81 308 349
rect 356 349 474 384
rect 356 -81 391 349
rect 273 -116 391 -81
rect 439 -81 474 349
rect 522 349 640 384
rect 522 -81 557 349
rect 439 -116 557 -81
rect 605 -81 640 349
rect 688 349 806 384
rect 688 -81 723 349
rect 605 -116 723 -81
rect 771 -168 806 349
<< locali >>
rect -871 432 -823 449
rect 823 432 871 449
rect -871 401 -854 432
rect 854 401 871 432
rect -871 -432 -854 -401
rect 854 -432 871 -401
rect -871 -449 -823 -432
rect 823 -449 871 -432
<< properties >>
string FIXED_BBOX -862 -440 862 440
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.35 l 5 m 1 nx 20 wmin 0.350 lmin 0.50 rho 2000 val 610.504k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 1 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
