// This is the unpowered netlist.
module dac_con (clk,
    dummy,
    llsb,
    llsb_n,
    rst_n,
    test_mode,
    dac_in,
    lsb,
    lsb_n,
    msb,
    msb_n);
 input clk;
 input dummy;
 output llsb;
 output llsb_n;
 input rst_n;
 input test_mode;
 input [9:0] dac_in;
 output [5:0] lsb;
 output [5:0] lsb_n;
 output [15:0] msb;
 output [15:0] msb_n;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire \cnt_r[0] ;
 wire \cnt_r[1] ;
 wire \cnt_r[2] ;
 wire \cnt_r[3] ;
 wire \cnt_r[4] ;
 wire \cnt_r[5] ;
 wire \cnt_r[6] ;
 wire \cnt_r[7] ;
 wire \cnt_r[8] ;
 wire \cnt_r[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;

 sky130_fd_sc_hd__clkinv_2 _093_ (.A(net14),
    .Y(net15));
 sky130_fd_sc_hd__clkinv_2 _094_ (.A(net28),
    .Y(net44));
 sky130_fd_sc_hd__clkinv_2 _095_ (.A(net35),
    .Y(net51));
 sky130_fd_sc_hd__clkinv_2 _096_ (.A(net36),
    .Y(net52));
 sky130_fd_sc_hd__clkinv_2 _097_ (.A(net37),
    .Y(net53));
 sky130_fd_sc_hd__clkinv_2 _098_ (.A(net38),
    .Y(net54));
 sky130_fd_sc_hd__clkinv_2 _099_ (.A(net39),
    .Y(net55));
 sky130_fd_sc_hd__clkinv_2 _100_ (.A(net40),
    .Y(net56));
 sky130_fd_sc_hd__clkinv_2 _101_ (.A(net41),
    .Y(net57));
 sky130_fd_sc_hd__clkinv_2 _102_ (.A(net42),
    .Y(net58));
 sky130_fd_sc_hd__clkinv_2 _103_ (.A(net43),
    .Y(net59));
 sky130_fd_sc_hd__clkinv_2 _104_ (.A(net29),
    .Y(net45));
 sky130_fd_sc_hd__clkinv_2 _105_ (.A(net30),
    .Y(net46));
 sky130_fd_sc_hd__clkinv_2 _106_ (.A(net31),
    .Y(net47));
 sky130_fd_sc_hd__clkinv_2 _107_ (.A(net32),
    .Y(net48));
 sky130_fd_sc_hd__clkinv_2 _108_ (.A(net33),
    .Y(net49));
 sky130_fd_sc_hd__clkinv_2 _109_ (.A(net34),
    .Y(net50));
 sky130_fd_sc_hd__clkinv_2 _110_ (.A(net16),
    .Y(net22));
 sky130_fd_sc_hd__clkinv_2 _111_ (.A(net17),
    .Y(net23));
 sky130_fd_sc_hd__clkinv_2 _112_ (.A(net18),
    .Y(net24));
 sky130_fd_sc_hd__clkinv_2 _113_ (.A(net19),
    .Y(net25));
 sky130_fd_sc_hd__clkinv_2 _114_ (.A(net20),
    .Y(net26));
 sky130_fd_sc_hd__clkinv_2 _115_ (.A(net21),
    .Y(net27));
 sky130_fd_sc_hd__clkbuf_1 _116_ (.A(net12),
    .X(_033_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _117_ (.A(_033_),
    .X(_034_));
 sky130_fd_sc_hd__clkbuf_1 _118_ (.A(_034_),
    .X(_035_));
 sky130_fd_sc_hd__clkbuf_1 _119_ (.A(_035_),
    .X(_000_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _120_ (.A(\cnt_r[0] ),
    .X(_036_));
 sky130_fd_sc_hd__inv_2 _121_ (.A(net12),
    .Y(_037_));
 sky130_fd_sc_hd__nor2_1 _122_ (.A(_036_),
    .B(_037_),
    .Y(_001_));
 sky130_fd_sc_hd__clkbuf_1 _123_ (.A(\cnt_r[1] ),
    .X(_038_));
 sky130_fd_sc_hd__o21ai_1 _124_ (.A1(_036_),
    .A2(_038_),
    .B1(_034_),
    .Y(_039_));
 sky130_fd_sc_hd__a21oi_1 _125_ (.A1(_036_),
    .A2(_038_),
    .B1(_039_),
    .Y(_002_));
 sky130_fd_sc_hd__and3_1 _126_ (.A(\cnt_r[0] ),
    .B(_038_),
    .C(\cnt_r[2] ),
    .X(_040_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _127_ (.A(_033_),
    .X(_041_));
 sky130_fd_sc_hd__a21o_1 _128_ (.A1(_036_),
    .A2(_038_),
    .B1(\cnt_r[2] ),
    .X(_042_));
 sky130_fd_sc_hd__and3b_1 _129_ (.A_N(_040_),
    .B(_041_),
    .C(_042_),
    .X(_043_));
 sky130_fd_sc_hd__clkbuf_1 _130_ (.A(_043_),
    .X(_003_));
 sky130_fd_sc_hd__and4_1 _131_ (.A(\cnt_r[0] ),
    .B(\cnt_r[1] ),
    .C(\cnt_r[2] ),
    .D(\cnt_r[3] ),
    .X(_044_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _132_ (.A(_044_),
    .X(_045_));
 sky130_fd_sc_hd__nor2_1 _133_ (.A(_037_),
    .B(_045_),
    .Y(_046_));
 sky130_fd_sc_hd__o21a_1 _134_ (.A1(\cnt_r[3] ),
    .A2(_040_),
    .B1(_046_),
    .X(_004_));
 sky130_fd_sc_hd__clkbuf_1 _135_ (.A(\cnt_r[4] ),
    .X(_047_));
 sky130_fd_sc_hd__a21oi_1 _136_ (.A1(_047_),
    .A2(_045_),
    .B1(_037_),
    .Y(_048_));
 sky130_fd_sc_hd__o21a_1 _137_ (.A1(_047_),
    .A2(_045_),
    .B1(_048_),
    .X(_005_));
 sky130_fd_sc_hd__and3_1 _138_ (.A(_047_),
    .B(\cnt_r[5] ),
    .C(_045_),
    .X(_049_));
 sky130_fd_sc_hd__a21o_1 _139_ (.A1(_047_),
    .A2(_045_),
    .B1(\cnt_r[5] ),
    .X(_050_));
 sky130_fd_sc_hd__and3b_1 _140_ (.A_N(_049_),
    .B(_041_),
    .C(_050_),
    .X(_051_));
 sky130_fd_sc_hd__clkbuf_1 _141_ (.A(_051_),
    .X(_006_));
 sky130_fd_sc_hd__and4_1 _142_ (.A(\cnt_r[4] ),
    .B(\cnt_r[5] ),
    .C(\cnt_r[6] ),
    .D(_044_),
    .X(_052_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _143_ (.A(_052_),
    .X(_053_));
 sky130_fd_sc_hd__o21ai_1 _144_ (.A1(\cnt_r[6] ),
    .A2(_049_),
    .B1(_034_),
    .Y(_054_));
 sky130_fd_sc_hd__nor2_1 _145_ (.A(_053_),
    .B(_054_),
    .Y(_007_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _146_ (.A(\cnt_r[7] ),
    .X(_055_));
 sky130_fd_sc_hd__a21oi_1 _147_ (.A1(_055_),
    .A2(_053_),
    .B1(_037_),
    .Y(_056_));
 sky130_fd_sc_hd__o21a_1 _148_ (.A1(_055_),
    .A2(_053_),
    .B1(_056_),
    .X(_008_));
 sky130_fd_sc_hd__a21o_1 _149_ (.A1(_055_),
    .A2(_052_),
    .B1(\cnt_r[8] ),
    .X(_057_));
 sky130_fd_sc_hd__nand3_1 _150_ (.A(\cnt_r[8] ),
    .B(_055_),
    .C(_053_),
    .Y(_058_));
 sky130_fd_sc_hd__and3_1 _151_ (.A(_041_),
    .B(_057_),
    .C(_058_),
    .X(_059_));
 sky130_fd_sc_hd__clkbuf_1 _152_ (.A(_059_),
    .X(_009_));
 sky130_fd_sc_hd__inv_2 _153_ (.A(\cnt_r[9] ),
    .Y(_060_));
 sky130_fd_sc_hd__a41o_1 _154_ (.A1(\cnt_r[9] ),
    .A2(\cnt_r[8] ),
    .A3(_055_),
    .A4(_053_),
    .B1(_037_),
    .X(_061_));
 sky130_fd_sc_hd__a21oi_1 _155_ (.A1(_060_),
    .A2(_058_),
    .B1(_061_),
    .Y(_010_));
 sky130_fd_sc_hd__and2_1 _156_ (.A(_034_),
    .B(net11),
    .X(_062_));
 sky130_fd_sc_hd__clkbuf_1 _157_ (.A(_062_),
    .X(_011_));
 sky130_fd_sc_hd__clkbuf_1 _158_ (.A(_033_),
    .X(_063_));
 sky130_fd_sc_hd__clkbuf_2 _159_ (.A(net13),
    .X(_064_));
 sky130_fd_sc_hd__clkbuf_2 _160_ (.A(_064_),
    .X(_065_));
 sky130_fd_sc_hd__mux2_1 _161_ (.A0(net1),
    .A1(_036_),
    .S(_065_),
    .X(_066_));
 sky130_fd_sc_hd__and2_1 _162_ (.A(_063_),
    .B(_066_),
    .X(_067_));
 sky130_fd_sc_hd__clkbuf_1 _163_ (.A(_067_),
    .X(_012_));
 sky130_fd_sc_hd__mux2_1 _164_ (.A0(net2),
    .A1(_038_),
    .S(_065_),
    .X(_068_));
 sky130_fd_sc_hd__and2_1 _165_ (.A(_063_),
    .B(_068_),
    .X(_069_));
 sky130_fd_sc_hd__clkbuf_1 _166_ (.A(_069_),
    .X(_013_));
 sky130_fd_sc_hd__mux2_1 _167_ (.A0(net3),
    .A1(\cnt_r[2] ),
    .S(_065_),
    .X(_070_));
 sky130_fd_sc_hd__and2_1 _168_ (.A(_063_),
    .B(_070_),
    .X(_071_));
 sky130_fd_sc_hd__clkbuf_1 _169_ (.A(_071_),
    .X(_014_));
 sky130_fd_sc_hd__mux2_1 _170_ (.A0(net4),
    .A1(\cnt_r[3] ),
    .S(_065_),
    .X(_072_));
 sky130_fd_sc_hd__and2_1 _171_ (.A(_063_),
    .B(_072_),
    .X(_073_));
 sky130_fd_sc_hd__clkbuf_1 _172_ (.A(_073_),
    .X(_015_));
 sky130_fd_sc_hd__mux2_1 _173_ (.A0(net5),
    .A1(_047_),
    .S(_065_),
    .X(_074_));
 sky130_fd_sc_hd__and2_1 _174_ (.A(_063_),
    .B(_074_),
    .X(_075_));
 sky130_fd_sc_hd__clkbuf_1 _175_ (.A(_075_),
    .X(_016_));
 sky130_fd_sc_hd__mux2_1 _176_ (.A0(net6),
    .A1(\cnt_r[5] ),
    .S(_064_),
    .X(_076_));
 sky130_fd_sc_hd__and2_1 _177_ (.A(_041_),
    .B(_076_),
    .X(_077_));
 sky130_fd_sc_hd__clkbuf_1 _178_ (.A(_077_),
    .X(_017_));
 sky130_fd_sc_hd__mux2_1 _179_ (.A0(net10),
    .A1(\cnt_r[9] ),
    .S(net13),
    .X(_078_));
 sky130_fd_sc_hd__and2_1 _180_ (.A(_033_),
    .B(_078_),
    .X(_079_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _181_ (.A(_079_),
    .X(_032_));
 sky130_fd_sc_hd__mux2_1 _182_ (.A0(net7),
    .A1(\cnt_r[6] ),
    .S(_064_),
    .X(_080_));
 sky130_fd_sc_hd__mux2_1 _183_ (.A0(net8),
    .A1(\cnt_r[7] ),
    .S(_064_),
    .X(_081_));
 sky130_fd_sc_hd__or2_1 _184_ (.A(_080_),
    .B(_081_),
    .X(_082_));
 sky130_fd_sc_hd__mux2_1 _185_ (.A0(net9),
    .A1(\cnt_r[8] ),
    .S(_064_),
    .X(_083_));
 sky130_fd_sc_hd__and3_1 _186_ (.A(net12),
    .B(_078_),
    .C(_083_),
    .X(_084_));
 sky130_fd_sc_hd__clkbuf_1 _187_ (.A(_084_),
    .X(_021_));
 sky130_fd_sc_hd__a21o_1 _188_ (.A1(_032_),
    .A2(_082_),
    .B1(_021_),
    .X(_018_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _189_ (.A(_081_),
    .X(_085_));
 sky130_fd_sc_hd__a21o_1 _190_ (.A1(_032_),
    .A2(_085_),
    .B1(_021_),
    .X(_019_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _191_ (.A(_083_),
    .X(_086_));
 sky130_fd_sc_hd__and2_1 _192_ (.A(_080_),
    .B(_085_),
    .X(_087_));
 sky130_fd_sc_hd__o21a_1 _193_ (.A1(_086_),
    .A2(_087_),
    .B1(_032_),
    .X(_020_));
 sky130_fd_sc_hd__and2_1 _194_ (.A(_021_),
    .B(_082_),
    .X(_088_));
 sky130_fd_sc_hd__clkbuf_1 _195_ (.A(_088_),
    .X(_022_));
 sky130_fd_sc_hd__and2_1 _196_ (.A(_021_),
    .B(_085_),
    .X(_089_));
 sky130_fd_sc_hd__clkbuf_1 _197_ (.A(_089_),
    .X(_023_));
 sky130_fd_sc_hd__and2_1 _198_ (.A(_084_),
    .B(_087_),
    .X(_090_));
 sky130_fd_sc_hd__clkbuf_1 _199_ (.A(_090_),
    .X(_024_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _200_ (.A(_041_),
    .X(_091_));
 sky130_fd_sc_hd__o21a_1 _201_ (.A1(_078_),
    .A2(_086_),
    .B1(_033_),
    .X(_092_));
 sky130_fd_sc_hd__clkbuf_1 _202_ (.A(_092_),
    .X(_028_));
 sky130_fd_sc_hd__a21o_1 _203_ (.A1(_091_),
    .A2(_082_),
    .B1(_028_),
    .X(_025_));
 sky130_fd_sc_hd__a21o_1 _204_ (.A1(_091_),
    .A2(_085_),
    .B1(_028_),
    .X(_026_));
 sky130_fd_sc_hd__a21o_1 _205_ (.A1(_091_),
    .A2(_087_),
    .B1(_028_),
    .X(_027_));
 sky130_fd_sc_hd__a31o_1 _206_ (.A1(_091_),
    .A2(_086_),
    .A3(_082_),
    .B1(_032_),
    .X(_029_));
 sky130_fd_sc_hd__a31o_1 _207_ (.A1(_091_),
    .A2(_086_),
    .A3(_085_),
    .B1(_079_),
    .X(_030_));
 sky130_fd_sc_hd__a31o_1 _208_ (.A1(_034_),
    .A2(_086_),
    .A3(_087_),
    .B1(_079_),
    .X(_031_));
 sky130_fd_sc_hd__dfxtp_1 _209_ (.CLK(clknet_2_3__leaf_clk),
    .D(_000_),
    .Q(net28));
 sky130_fd_sc_hd__dfxtp_1 _210_ (.CLK(clknet_2_1__leaf_clk),
    .D(_001_),
    .Q(\cnt_r[0] ));
 sky130_fd_sc_hd__dfxtp_1 _211_ (.CLK(clknet_2_1__leaf_clk),
    .D(_002_),
    .Q(\cnt_r[1] ));
 sky130_fd_sc_hd__dfxtp_1 _212_ (.CLK(clknet_2_1__leaf_clk),
    .D(_003_),
    .Q(\cnt_r[2] ));
 sky130_fd_sc_hd__dfxtp_1 _213_ (.CLK(clknet_2_1__leaf_clk),
    .D(_004_),
    .Q(\cnt_r[3] ));
 sky130_fd_sc_hd__dfxtp_1 _214_ (.CLK(clknet_2_0__leaf_clk),
    .D(_005_),
    .Q(\cnt_r[4] ));
 sky130_fd_sc_hd__dfxtp_1 _215_ (.CLK(clknet_2_1__leaf_clk),
    .D(_006_),
    .Q(\cnt_r[5] ));
 sky130_fd_sc_hd__dfxtp_1 _216_ (.CLK(clknet_2_1__leaf_clk),
    .D(_007_),
    .Q(\cnt_r[6] ));
 sky130_fd_sc_hd__dfxtp_1 _217_ (.CLK(clknet_2_0__leaf_clk),
    .D(_008_),
    .Q(\cnt_r[7] ));
 sky130_fd_sc_hd__dfxtp_1 _218_ (.CLK(clknet_2_0__leaf_clk),
    .D(_009_),
    .Q(\cnt_r[8] ));
 sky130_fd_sc_hd__dfxtp_1 _219_ (.CLK(clknet_2_0__leaf_clk),
    .D(_010_),
    .Q(\cnt_r[9] ));
 sky130_fd_sc_hd__dfxtp_1 _220_ (.CLK(clknet_2_1__leaf_clk),
    .D(_011_),
    .Q(net14));
 sky130_fd_sc_hd__dfxtp_1 _221_ (.CLK(clknet_2_3__leaf_clk),
    .D(_012_),
    .Q(net16));
 sky130_fd_sc_hd__dfxtp_1 _222_ (.CLK(clknet_2_3__leaf_clk),
    .D(_013_),
    .Q(net17));
 sky130_fd_sc_hd__dfxtp_1 _223_ (.CLK(clknet_2_3__leaf_clk),
    .D(_014_),
    .Q(net18));
 sky130_fd_sc_hd__dfxtp_1 _224_ (.CLK(clknet_2_3__leaf_clk),
    .D(_015_),
    .Q(net19));
 sky130_fd_sc_hd__dfxtp_1 _225_ (.CLK(clknet_2_3__leaf_clk),
    .D(_016_),
    .Q(net20));
 sky130_fd_sc_hd__dfxtp_1 _226_ (.CLK(clknet_2_1__leaf_clk),
    .D(_017_),
    .Q(net21));
 sky130_fd_sc_hd__dfxtp_1 _227_ (.CLK(clknet_2_2__leaf_clk),
    .D(_018_),
    .Q(net43));
 sky130_fd_sc_hd__dfxtp_1 _228_ (.CLK(clknet_2_2__leaf_clk),
    .D(_019_),
    .Q(net29));
 sky130_fd_sc_hd__dfxtp_1 _229_ (.CLK(clknet_2_2__leaf_clk),
    .D(_020_),
    .Q(net30));
 sky130_fd_sc_hd__dfxtp_1 _230_ (.CLK(clknet_2_2__leaf_clk),
    .D(_021_),
    .Q(net31));
 sky130_fd_sc_hd__dfxtp_1 _231_ (.CLK(clknet_2_2__leaf_clk),
    .D(_022_),
    .Q(net32));
 sky130_fd_sc_hd__dfxtp_1 _232_ (.CLK(clknet_2_3__leaf_clk),
    .D(_023_),
    .Q(net33));
 sky130_fd_sc_hd__dfxtp_1 _233_ (.CLK(clknet_2_0__leaf_clk),
    .D(_024_),
    .Q(net34));
 sky130_fd_sc_hd__dfxtp_1 _234_ (.CLK(clknet_2_2__leaf_clk),
    .D(_025_),
    .Q(net35));
 sky130_fd_sc_hd__dfxtp_1 _235_ (.CLK(clknet_2_3__leaf_clk),
    .D(_026_),
    .Q(net36));
 sky130_fd_sc_hd__dfxtp_1 _236_ (.CLK(clknet_2_3__leaf_clk),
    .D(_027_),
    .Q(net37));
 sky130_fd_sc_hd__dfxtp_1 _237_ (.CLK(clknet_2_2__leaf_clk),
    .D(_028_),
    .Q(net38));
 sky130_fd_sc_hd__dfxtp_1 _238_ (.CLK(clknet_2_2__leaf_clk),
    .D(_029_),
    .Q(net39));
 sky130_fd_sc_hd__dfxtp_1 _239_ (.CLK(clknet_2_2__leaf_clk),
    .D(_030_),
    .Q(net40));
 sky130_fd_sc_hd__dfxtp_1 _240_ (.CLK(clknet_2_0__leaf_clk),
    .D(_031_),
    .Q(net41));
 sky130_fd_sc_hd__dfxtp_1 _241_ (.CLK(clknet_2_3__leaf_clk),
    .D(_032_),
    .Q(net42));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(dac_in[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(dac_in[1]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(dac_in[2]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(dac_in[3]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(dac_in[4]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(dac_in[5]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(dac_in[6]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(dac_in[7]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(dac_in[8]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(dac_in[9]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(dummy),
    .X(net11));
 sky130_fd_sc_hd__dlymetal6s2s_1 input12 (.A(rst_n),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(test_mode),
    .X(net13));
 sky130_fd_sc_hd__buf_2 output14 (.A(net14),
    .X(llsb));
 sky130_fd_sc_hd__buf_2 output15 (.A(net15),
    .X(llsb_n));
 sky130_fd_sc_hd__buf_2 output16 (.A(net16),
    .X(lsb[0]));
 sky130_fd_sc_hd__buf_2 output17 (.A(net17),
    .X(lsb[1]));
 sky130_fd_sc_hd__buf_2 output18 (.A(net18),
    .X(lsb[2]));
 sky130_fd_sc_hd__buf_2 output19 (.A(net19),
    .X(lsb[3]));
 sky130_fd_sc_hd__buf_2 output20 (.A(net20),
    .X(lsb[4]));
 sky130_fd_sc_hd__buf_2 output21 (.A(net21),
    .X(lsb[5]));
 sky130_fd_sc_hd__buf_2 output22 (.A(net22),
    .X(lsb_n[0]));
 sky130_fd_sc_hd__buf_2 output23 (.A(net23),
    .X(lsb_n[1]));
 sky130_fd_sc_hd__buf_2 output24 (.A(net24),
    .X(lsb_n[2]));
 sky130_fd_sc_hd__buf_2 output25 (.A(net25),
    .X(lsb_n[3]));
 sky130_fd_sc_hd__buf_2 output26 (.A(net26),
    .X(lsb_n[4]));
 sky130_fd_sc_hd__buf_2 output27 (.A(net27),
    .X(lsb_n[5]));
 sky130_fd_sc_hd__buf_2 output28 (.A(net28),
    .X(msb[0]));
 sky130_fd_sc_hd__buf_2 output29 (.A(net29),
    .X(msb[10]));
 sky130_fd_sc_hd__buf_2 output30 (.A(net30),
    .X(msb[11]));
 sky130_fd_sc_hd__buf_2 output31 (.A(net31),
    .X(msb[12]));
 sky130_fd_sc_hd__buf_2 output32 (.A(net32),
    .X(msb[13]));
 sky130_fd_sc_hd__buf_2 output33 (.A(net33),
    .X(msb[14]));
 sky130_fd_sc_hd__buf_2 output34 (.A(net34),
    .X(msb[15]));
 sky130_fd_sc_hd__buf_2 output35 (.A(net35),
    .X(msb[1]));
 sky130_fd_sc_hd__buf_2 output36 (.A(net36),
    .X(msb[2]));
 sky130_fd_sc_hd__buf_2 output37 (.A(net37),
    .X(msb[3]));
 sky130_fd_sc_hd__buf_2 output38 (.A(net38),
    .X(msb[4]));
 sky130_fd_sc_hd__buf_2 output39 (.A(net39),
    .X(msb[5]));
 sky130_fd_sc_hd__buf_2 output40 (.A(net40),
    .X(msb[6]));
 sky130_fd_sc_hd__buf_2 output41 (.A(net41),
    .X(msb[7]));
 sky130_fd_sc_hd__buf_2 output42 (.A(net42),
    .X(msb[8]));
 sky130_fd_sc_hd__buf_2 output43 (.A(net43),
    .X(msb[9]));
 sky130_fd_sc_hd__buf_2 output44 (.A(net44),
    .X(msb_n[0]));
 sky130_fd_sc_hd__buf_2 output45 (.A(net45),
    .X(msb_n[10]));
 sky130_fd_sc_hd__buf_2 output46 (.A(net46),
    .X(msb_n[11]));
 sky130_fd_sc_hd__buf_2 output47 (.A(net47),
    .X(msb_n[12]));
 sky130_fd_sc_hd__buf_2 output48 (.A(net48),
    .X(msb_n[13]));
 sky130_fd_sc_hd__buf_2 output49 (.A(net49),
    .X(msb_n[14]));
 sky130_fd_sc_hd__buf_2 output50 (.A(net50),
    .X(msb_n[15]));
 sky130_fd_sc_hd__buf_2 output51 (.A(net51),
    .X(msb_n[1]));
 sky130_fd_sc_hd__buf_2 output52 (.A(net52),
    .X(msb_n[2]));
 sky130_fd_sc_hd__buf_2 output53 (.A(net53),
    .X(msb_n[3]));
 sky130_fd_sc_hd__buf_2 output54 (.A(net54),
    .X(msb_n[4]));
 sky130_fd_sc_hd__buf_2 output55 (.A(net55),
    .X(msb_n[5]));
 sky130_fd_sc_hd__buf_2 output56 (.A(net56),
    .X(msb_n[6]));
 sky130_fd_sc_hd__buf_2 output57 (.A(net57),
    .X(msb_n[7]));
 sky130_fd_sc_hd__buf_2 output58 (.A(net58),
    .X(msb_n[8]));
 sky130_fd_sc_hd__buf_2 output59 (.A(net59),
    .X(msb_n[9]));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(dac_in[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(dac_in[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(dac_in[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(dac_in[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(dac_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(dac_in[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(dac_in[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(dac_in[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(dac_in[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(dac_in[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(dummy));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(rst_n));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(test_mode));
 sky130_fd_sc_hd__diode_2 ANTENNA_output14_A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__093__A (.DIODE(net14));
 sky130_fd_sc_hd__decap_6 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_84 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_30 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_145 ();
endmodule

