magic
tech sky130A
magscale 1 2
timestamp 1671152619
<< error_p >>
rect 1177 147 1235 153
rect 1295 147 1353 153
rect 1413 147 1471 153
rect 1531 147 1589 153
rect 1649 147 1707 153
rect 1767 147 1825 153
rect 1885 147 1943 153
rect 2003 147 2061 153
rect 2121 147 2179 153
rect 2239 147 2297 153
rect 2357 147 2415 153
rect 2475 147 2533 153
rect 2593 147 2651 153
rect 2711 147 2769 153
rect 2829 147 2887 153
rect 2947 147 3005 153
rect 3065 147 3123 153
rect 3183 147 3241 153
rect 3301 147 3359 153
rect 3419 147 3477 153
rect 3537 147 3595 153
rect 3655 147 3713 153
rect 3773 147 3831 153
rect 3891 147 3949 153
rect 4009 147 4067 153
rect 4127 147 4185 153
rect 4245 147 4303 153
rect 4363 147 4421 153
rect 4481 147 4539 153
rect 4599 147 4657 153
rect 4717 147 4775 153
rect 4835 147 4893 153
rect 4953 147 5011 153
rect 5071 147 5129 153
rect 5189 147 5247 153
rect 5307 147 5365 153
rect 5425 147 5483 153
rect 5543 147 5601 153
rect 5661 147 5719 153
rect 5779 147 5837 153
rect 5897 147 5955 153
rect 6015 147 6073 153
rect 6133 147 6191 153
rect 6251 147 6309 153
rect 6369 147 6427 153
rect 6487 147 6545 153
rect 1177 113 1189 147
rect 1295 113 1307 147
rect 1413 113 1425 147
rect 1531 113 1543 147
rect 1649 113 1661 147
rect 1767 113 1779 147
rect 1885 113 1897 147
rect 2003 113 2015 147
rect 2121 113 2133 147
rect 2239 113 2251 147
rect 2357 113 2369 147
rect 2475 113 2487 147
rect 2593 113 2605 147
rect 2711 113 2723 147
rect 2829 113 2841 147
rect 2947 113 2959 147
rect 3065 113 3077 147
rect 3183 113 3195 147
rect 3301 113 3313 147
rect 3419 113 3431 147
rect 3537 113 3549 147
rect 3655 113 3667 147
rect 3773 113 3785 147
rect 3891 113 3903 147
rect 4009 113 4021 147
rect 4127 113 4139 147
rect 4245 113 4257 147
rect 4363 113 4375 147
rect 4481 113 4493 147
rect 4599 113 4611 147
rect 4717 113 4729 147
rect 4835 113 4847 147
rect 4953 113 4965 147
rect 5071 113 5083 147
rect 5189 113 5201 147
rect 5307 113 5319 147
rect 5425 113 5437 147
rect 5543 113 5555 147
rect 5661 113 5673 147
rect 5779 113 5791 147
rect 5897 113 5909 147
rect 6015 113 6027 147
rect 6133 113 6145 147
rect 6251 113 6263 147
rect 6369 113 6381 147
rect 6487 113 6499 147
rect 1177 107 1235 113
rect 1295 107 1353 113
rect 1413 107 1471 113
rect 1531 107 1589 113
rect 1649 107 1707 113
rect 1767 107 1825 113
rect 1885 107 1943 113
rect 2003 107 2061 113
rect 2121 107 2179 113
rect 2239 107 2297 113
rect 2357 107 2415 113
rect 2475 107 2533 113
rect 2593 107 2651 113
rect 2711 107 2769 113
rect 2829 107 2887 113
rect 2947 107 3005 113
rect 3065 107 3123 113
rect 3183 107 3241 113
rect 3301 107 3359 113
rect 3419 107 3477 113
rect 3537 107 3595 113
rect 3655 107 3713 113
rect 3773 107 3831 113
rect 3891 107 3949 113
rect 4009 107 4067 113
rect 4127 107 4185 113
rect 4245 107 4303 113
rect 4363 107 4421 113
rect 4481 107 4539 113
rect 4599 107 4657 113
rect 4717 107 4775 113
rect 4835 107 4893 113
rect 4953 107 5011 113
rect 5071 107 5129 113
rect 5189 107 5247 113
rect 5307 107 5365 113
rect 5425 107 5483 113
rect 5543 107 5601 113
rect 5661 107 5719 113
rect 5779 107 5837 113
rect 5897 107 5955 113
rect 6015 107 6073 113
rect 6133 107 6191 113
rect 6251 107 6309 113
rect 6369 107 6427 113
rect 6487 107 6545 113
<< error_s >>
rect 1177 -1981 1235 -1975
rect 1295 -1981 1353 -1975
rect 1413 -1981 1471 -1975
rect 1531 -1981 1589 -1975
rect 1649 -1981 1707 -1975
rect 1767 -1981 1825 -1975
rect 1885 -1981 1943 -1975
rect 2003 -1981 2061 -1975
rect 2121 -1981 2179 -1975
rect 2239 -1981 2297 -1975
rect 2357 -1981 2415 -1975
rect 2475 -1981 2533 -1975
rect 2593 -1981 2651 -1975
rect 2711 -1981 2769 -1975
rect 2829 -1981 2887 -1975
rect 2947 -1981 3005 -1975
rect 3065 -1981 3123 -1975
rect 3183 -1981 3241 -1975
rect 3301 -1981 3359 -1975
rect 3419 -1981 3477 -1975
rect 3537 -1981 3595 -1975
rect 3655 -1981 3713 -1975
rect 3773 -1981 3831 -1975
rect 3891 -1981 3949 -1975
rect 4009 -1981 4067 -1975
rect 4127 -1981 4185 -1975
rect 4245 -1981 4303 -1975
rect 4363 -1981 4421 -1975
rect 4481 -1981 4539 -1975
rect 4599 -1981 4657 -1975
rect 4717 -1981 4775 -1975
rect 4835 -1981 4893 -1975
rect 4953 -1981 5011 -1975
rect 5071 -1981 5129 -1975
rect 5189 -1981 5247 -1975
rect 5307 -1981 5365 -1975
rect 5425 -1981 5483 -1975
rect 5543 -1981 5601 -1975
rect 5661 -1981 5719 -1975
rect 5779 -1981 5837 -1975
rect 5897 -1981 5955 -1975
rect 6015 -1981 6073 -1975
rect 6133 -1981 6191 -1975
rect 6251 -1981 6309 -1975
rect 6369 -1981 6427 -1975
rect 6487 -1981 6545 -1975
rect 1177 -2015 1189 -1981
rect 1295 -2015 1307 -1981
rect 1413 -2015 1425 -1981
rect 1531 -2015 1543 -1981
rect 1649 -2015 1661 -1981
rect 1767 -2015 1779 -1981
rect 1885 -2015 1897 -1981
rect 2003 -2015 2015 -1981
rect 2121 -2015 2133 -1981
rect 2239 -2015 2251 -1981
rect 2357 -2015 2369 -1981
rect 2475 -2015 2487 -1981
rect 2593 -2015 2605 -1981
rect 2711 -2015 2723 -1981
rect 2829 -2015 2841 -1981
rect 2947 -2015 2959 -1981
rect 3065 -2015 3077 -1981
rect 3183 -2015 3195 -1981
rect 3301 -2015 3313 -1981
rect 3419 -2015 3431 -1981
rect 3537 -2015 3549 -1981
rect 3655 -2015 3667 -1981
rect 3773 -2015 3785 -1981
rect 3891 -2015 3903 -1981
rect 4009 -2015 4021 -1981
rect 4127 -2015 4139 -1981
rect 4245 -2015 4257 -1981
rect 4363 -2015 4375 -1981
rect 4481 -2015 4493 -1981
rect 4599 -2015 4611 -1981
rect 4717 -2015 4729 -1981
rect 4835 -2015 4847 -1981
rect 4953 -2015 4965 -1981
rect 5071 -2015 5083 -1981
rect 5189 -2015 5201 -1981
rect 5307 -2015 5319 -1981
rect 5425 -2015 5437 -1981
rect 5543 -2015 5555 -1981
rect 5661 -2015 5673 -1981
rect 5779 -2015 5791 -1981
rect 5897 -2015 5909 -1981
rect 6015 -2015 6027 -1981
rect 6133 -2015 6145 -1981
rect 6251 -2015 6263 -1981
rect 6369 -2015 6381 -1981
rect 6487 -2015 6499 -1981
rect 1177 -2021 1235 -2015
rect 1295 -2021 1353 -2015
rect 1413 -2021 1471 -2015
rect 1531 -2021 1589 -2015
rect 1649 -2021 1707 -2015
rect 1767 -2021 1825 -2015
rect 1885 -2021 1943 -2015
rect 2003 -2021 2061 -2015
rect 2121 -2021 2179 -2015
rect 2239 -2021 2297 -2015
rect 2357 -2021 2415 -2015
rect 2475 -2021 2533 -2015
rect 2593 -2021 2651 -2015
rect 2711 -2021 2769 -2015
rect 2829 -2021 2887 -2015
rect 2947 -2021 3005 -2015
rect 3065 -2021 3123 -2015
rect 3183 -2021 3241 -2015
rect 3301 -2021 3359 -2015
rect 3419 -2021 3477 -2015
rect 3537 -2021 3595 -2015
rect 3655 -2021 3713 -2015
rect 3773 -2021 3831 -2015
rect 3891 -2021 3949 -2015
rect 4009 -2021 4067 -2015
rect 4127 -2021 4185 -2015
rect 4245 -2021 4303 -2015
rect 4363 -2021 4421 -2015
rect 4481 -2021 4539 -2015
rect 4599 -2021 4657 -2015
rect 4717 -2021 4775 -2015
rect 4835 -2021 4893 -2015
rect 4953 -2021 5011 -2015
rect 5071 -2021 5129 -2015
rect 5189 -2021 5247 -2015
rect 5307 -2021 5365 -2015
rect 5425 -2021 5483 -2015
rect 5543 -2021 5601 -2015
rect 5661 -2021 5719 -2015
rect 5779 -2021 5837 -2015
rect 5897 -2021 5955 -2015
rect 6015 -2021 6073 -2015
rect 6133 -2021 6191 -2015
rect 6251 -2021 6309 -2015
rect 6369 -2021 6427 -2015
rect 6487 -2021 6545 -2015
rect 1177 -2292 1235 -2286
rect 1295 -2292 1353 -2286
rect 1413 -2292 1471 -2286
rect 1531 -2292 1589 -2286
rect 1649 -2292 1707 -2286
rect 1767 -2292 1825 -2286
rect 1885 -2292 1943 -2286
rect 2003 -2292 2061 -2286
rect 5662 -2291 5720 -2285
rect 5780 -2291 5838 -2285
rect 5898 -2291 5956 -2285
rect 6016 -2291 6074 -2285
rect 6134 -2291 6192 -2285
rect 6252 -2291 6310 -2285
rect 6370 -2291 6428 -2285
rect 6488 -2291 6546 -2285
rect 1177 -2326 1189 -2292
rect 1295 -2326 1307 -2292
rect 1413 -2326 1425 -2292
rect 1531 -2326 1543 -2292
rect 1649 -2326 1661 -2292
rect 1767 -2326 1779 -2292
rect 1885 -2326 1897 -2292
rect 2003 -2326 2015 -2292
rect 5662 -2325 5674 -2291
rect 5780 -2325 5792 -2291
rect 5898 -2325 5910 -2291
rect 6016 -2325 6028 -2291
rect 6134 -2325 6146 -2291
rect 6252 -2325 6264 -2291
rect 6370 -2325 6382 -2291
rect 6488 -2325 6500 -2291
rect 1177 -2332 1235 -2326
rect 1295 -2332 1353 -2326
rect 1413 -2332 1471 -2326
rect 1531 -2332 1589 -2326
rect 1649 -2332 1707 -2326
rect 1767 -2332 1825 -2326
rect 1885 -2332 1943 -2326
rect 2003 -2332 2061 -2326
rect 5662 -2331 5720 -2325
rect 5780 -2331 5838 -2325
rect 5898 -2331 5956 -2325
rect 6016 -2331 6074 -2325
rect 6134 -2331 6192 -2325
rect 6252 -2331 6310 -2325
rect 6370 -2331 6428 -2325
rect 6488 -2331 6546 -2325
rect 1177 -4402 1235 -4396
rect 1295 -4402 1353 -4396
rect 1413 -4402 1471 -4396
rect 1531 -4402 1589 -4396
rect 1649 -4402 1707 -4396
rect 1767 -4402 1825 -4396
rect 1885 -4402 1943 -4396
rect 2003 -4402 2061 -4396
rect 5662 -4401 5720 -4395
rect 5780 -4401 5838 -4395
rect 5898 -4401 5956 -4395
rect 6016 -4401 6074 -4395
rect 6134 -4401 6192 -4395
rect 6252 -4401 6310 -4395
rect 6370 -4401 6428 -4395
rect 6488 -4401 6546 -4395
rect 1177 -4436 1189 -4402
rect 1295 -4436 1307 -4402
rect 1413 -4436 1425 -4402
rect 1531 -4436 1543 -4402
rect 1649 -4436 1661 -4402
rect 1767 -4436 1779 -4402
rect 1885 -4436 1897 -4402
rect 2003 -4436 2015 -4402
rect 5662 -4435 5674 -4401
rect 5780 -4435 5792 -4401
rect 5898 -4435 5910 -4401
rect 6016 -4435 6028 -4401
rect 6134 -4435 6146 -4401
rect 6252 -4435 6264 -4401
rect 6370 -4435 6382 -4401
rect 6488 -4435 6500 -4401
rect 1177 -4442 1235 -4436
rect 1295 -4442 1353 -4436
rect 1413 -4442 1471 -4436
rect 1531 -4442 1589 -4436
rect 1649 -4442 1707 -4436
rect 1767 -4442 1825 -4436
rect 1885 -4442 1943 -4436
rect 2003 -4442 2061 -4436
rect 5662 -4441 5720 -4435
rect 5780 -4441 5838 -4435
rect 5898 -4441 5956 -4435
rect 6016 -4441 6074 -4435
rect 6134 -4441 6192 -4435
rect 6252 -4441 6310 -4435
rect 6370 -4441 6428 -4435
rect 6488 -4441 6546 -4435
<< metal1 >>
rect 3396 -2426 4038 -2376
rect 4164 -2426 4268 -2376
rect 4222 -2464 4268 -2426
rect 3252 -3464 3258 -2464
rect 3312 -3464 3318 -2464
rect 3348 -3464 3354 -2464
rect 3408 -3464 3414 -2464
rect 3444 -3464 3450 -2464
rect 3504 -3464 3510 -2464
rect 3540 -3464 3546 -2464
rect 3600 -3464 3606 -2464
rect 3636 -3464 3642 -2464
rect 3696 -3464 3702 -2464
rect 3732 -3464 3738 -2464
rect 3792 -3464 3798 -2464
rect 3828 -3464 3834 -2464
rect 3888 -3464 3894 -2464
rect 3924 -3464 3930 -2464
rect 3984 -3464 3990 -2464
rect 4020 -3464 4026 -2464
rect 4080 -3464 4086 -2464
rect 4116 -3464 4122 -2464
rect 4176 -3464 4182 -2464
rect 4212 -3464 4218 -2464
rect 4272 -3464 4278 -2464
rect 3268 -3502 3308 -3464
rect 3268 -3542 3366 -3502
rect 3492 -3552 4134 -3502
<< via1 >>
rect 3258 -3464 3312 -2464
rect 3354 -3464 3408 -2464
rect 3450 -3464 3504 -2464
rect 3546 -3464 3600 -2464
rect 3642 -3464 3696 -2464
rect 3738 -3464 3792 -2464
rect 3834 -3464 3888 -2464
rect 3930 -3464 3984 -2464
rect 4026 -3464 4080 -2464
rect 4122 -3464 4176 -2464
rect 4218 -3464 4272 -2464
<< metal2 >>
rect 3348 -2464 3414 -2350
rect 3252 -3464 3258 -2464
rect 3312 -3464 3318 -2464
rect 3348 -3464 3354 -2464
rect 3408 -3464 3414 -2464
rect 3444 -3464 3450 -2464
rect 3504 -3464 3510 -2464
rect 3540 -3464 3546 -2464
rect 3600 -3464 3606 -2464
rect 3636 -3464 3642 -2464
rect 3696 -3464 3702 -2464
rect 3732 -3464 3738 -2464
rect 3792 -3464 3798 -2464
rect 3828 -3464 3834 -2464
rect 3888 -3464 3894 -2464
rect 3924 -3464 3930 -2464
rect 3984 -3464 3990 -2464
rect 4020 -3464 4026 -2464
rect 4080 -3464 4086 -2464
rect 4116 -3464 4122 -2464
rect 4176 -3464 4182 -2464
rect 4212 -3464 4218 -2464
rect 4272 -3464 4278 -2464
rect 3444 -3674 3510 -3464
rect 3636 -3674 3702 -3464
rect 3828 -3674 3894 -3464
rect 4020 -3674 4086 -3464
use sky130_fd_pr__nfet_01v8_P4JNYZ  sky130_fd_pr__nfet_01v8_P4JNYZ_0
timestamp 1671152619
transform 1 0 3765 0 1 -2964
box -647 -710 647 710
use sky130_fd_pr__nfet_01v8_RSFWNV  sky130_fd_pr__nfet_01v8_RSFWNV_0
timestamp 1671152619
transform 1 0 6104 0 1 -3363
box -639 -1210 639 1210
use sky130_fd_pr__nfet_01v8_RSFWNV  sky130_fd_pr__nfet_01v8_RSFWNV_2
timestamp 1671152619
transform 1 0 1619 0 1 -3364
box -639 -1210 639 1210
use sky130_fd_pr__nfet_01v8_U52XAY  sky130_fd_pr__nfet_01v8_U52XAY_0
timestamp 1671152619
transform 1 0 4141 0 1 -5644
box -1999 -710 1999 710
use sky130_fd_pr__pfet_01v8_4D836H  sky130_fd_pr__pfet_01v8_4D836H_0
timestamp 1671152619
transform 1 0 3861 0 1 -934
box -2881 -1219 2881 1219
<< end >>
