magic
tech sky130A
magscale 1 2
timestamp 1671985581
<< locali >>
rect 220 1107 285 1174
rect -774 1072 -710 1081
rect -1051 1049 -987 1058
rect -1051 1015 -1036 1049
rect -1002 1015 -987 1049
rect -774 1038 -759 1072
rect -725 1038 -710 1072
rect -774 1029 -710 1038
rect -660 1074 -596 1083
rect -660 1040 -645 1074
rect -611 1040 -596 1074
rect -660 1031 -596 1040
rect -267 1061 -203 1070
rect -267 1027 -252 1061
rect -218 1027 -203 1061
rect 220 1040 455 1107
rect 902 1046 966 1055
rect -267 1018 -203 1027
rect -1051 1006 -987 1015
rect 902 1012 917 1046
rect 951 1012 966 1046
rect 4267 1046 4403 1055
rect 902 1003 966 1012
rect 2981 1014 3045 1023
rect 2981 980 2996 1014
rect 3030 980 3045 1014
rect 4267 1012 4282 1046
rect 4316 1012 4354 1046
rect 4388 1012 4403 1046
rect 4267 1003 4403 1012
rect 4654 1046 4790 1055
rect 4654 1012 4669 1046
rect 4703 1012 4741 1046
rect 4775 1012 4790 1046
rect 4654 1003 4790 1012
rect 2981 971 3045 980
rect 4865 970 4965 1050
rect 3671 943 3723 958
rect 3671 909 3680 943
rect 3714 909 3723 943
rect -375 887 -311 896
rect -375 853 -360 887
rect -326 853 -311 887
rect -375 844 -311 853
rect 3671 871 3723 909
rect 3671 837 3680 871
rect 3714 837 3723 871
rect -167 815 -115 830
rect 3671 822 3723 837
rect -167 781 -158 815
rect -124 781 -115 815
rect -167 766 -115 781
rect 3265 490 3317 505
rect 3265 456 3274 490
rect 3308 456 3317 490
rect 3265 418 3317 456
rect 3265 384 3274 418
rect 3308 384 3317 418
rect 3265 369 3317 384
rect 3674 486 3726 501
rect 3674 452 3683 486
rect 3717 452 3726 486
rect 3674 414 3726 452
rect 3674 380 3683 414
rect 3717 380 3726 414
rect 3674 365 3726 380
rect 2983 353 3047 362
rect 490 342 554 351
rect 490 308 505 342
rect 539 308 554 342
rect 490 299 554 308
rect 906 320 970 329
rect 217 225 452 292
rect 906 286 921 320
rect 955 286 970 320
rect 2983 319 2998 353
rect 3032 319 3047 353
rect 2983 310 3047 319
rect 4245 341 4311 356
rect 4245 307 4262 341
rect 4296 307 4311 341
rect 4245 290 4311 307
rect 4372 334 4450 343
rect 4372 300 4387 334
rect 4421 300 4450 334
rect 4916 327 4974 345
rect 4372 291 4450 300
rect 4757 287 4974 327
rect 906 277 970 286
rect 4916 265 4974 287
rect 220 191 286 225
<< viali >>
rect -1036 1015 -1002 1049
rect -759 1038 -725 1072
rect -645 1040 -611 1074
rect -252 1027 -218 1061
rect 509 991 543 1025
rect 917 1012 951 1046
rect 2996 980 3030 1014
rect 4282 1012 4316 1046
rect 4354 1012 4388 1046
rect 4669 1012 4703 1046
rect 4741 1012 4775 1046
rect 3680 909 3714 943
rect -360 853 -326 887
rect 3680 837 3714 871
rect -158 781 -124 815
rect 3274 456 3308 490
rect 3274 384 3308 418
rect 3683 452 3717 486
rect 3683 380 3717 414
rect 505 308 539 342
rect 921 286 955 320
rect 2998 319 3032 353
rect 4262 307 4296 341
rect 4387 300 4421 334
<< metal1 >>
rect -1051 1006 -1045 1058
rect -993 1006 -987 1058
rect -774 1029 -768 1081
rect -716 1029 -710 1081
rect -660 1031 -654 1083
rect -602 1031 -596 1083
rect -267 1018 -261 1070
rect -209 1018 -203 1070
rect 497 1025 555 1034
rect 497 991 509 1025
rect 543 991 555 1025
rect 902 1003 908 1055
rect 960 1003 966 1055
rect 497 982 555 991
rect -375 844 -369 896
rect -317 844 -311 896
rect -167 824 -115 830
rect -167 766 -115 772
rect 501 715 547 982
rect 2632 700 2660 1013
rect 2981 971 2987 1023
rect 3039 971 3045 1023
rect 4267 1003 4273 1055
rect 4325 1003 4345 1055
rect 4397 1003 4403 1055
rect 4654 1003 4660 1055
rect 4712 1003 4732 1055
rect 4784 1003 4790 1055
rect 3671 952 3723 958
rect 3671 880 3723 900
rect 3671 822 3723 828
rect 2632 640 2640 700
rect 490 299 496 351
rect 548 299 554 351
rect 906 277 912 329
rect 964 277 970 329
rect 2632 319 2660 640
rect 3265 499 3317 505
rect 3265 427 3317 447
rect 3265 369 3317 375
rect 3674 495 3726 501
rect 3674 423 3726 443
rect 3674 365 3726 371
rect 2983 310 2989 362
rect 3041 310 3047 362
rect 4245 350 4311 356
rect 4245 298 4253 350
rect 4305 298 4311 350
rect 4245 290 4311 298
rect 4372 291 4378 343
rect 4430 291 4450 343
<< via1 >>
rect 240 1960 660 2040
rect 1440 1960 1860 2040
rect 2640 1960 3060 2040
rect 3840 1960 4260 2040
rect -460 1300 -40 1380
rect 840 1300 1260 1360
rect 2040 1300 2460 1360
rect 3240 1300 3660 1360
rect 4440 1300 4860 1360
rect -1045 1049 -993 1058
rect -1045 1015 -1036 1049
rect -1036 1015 -1002 1049
rect -1002 1015 -993 1049
rect -1045 1006 -993 1015
rect -768 1072 -716 1081
rect -768 1038 -759 1072
rect -759 1038 -725 1072
rect -725 1038 -716 1072
rect -768 1029 -716 1038
rect -654 1074 -602 1083
rect -654 1040 -645 1074
rect -645 1040 -611 1074
rect -611 1040 -602 1074
rect -654 1031 -602 1040
rect -261 1061 -209 1070
rect -261 1027 -252 1061
rect -252 1027 -218 1061
rect -218 1027 -209 1061
rect -261 1018 -209 1027
rect 908 1046 960 1055
rect 908 1012 917 1046
rect 917 1012 951 1046
rect 951 1012 960 1046
rect 908 1003 960 1012
rect -369 887 -317 896
rect -369 853 -360 887
rect -360 853 -326 887
rect -326 853 -317 887
rect -369 844 -317 853
rect -167 815 -115 824
rect -167 781 -158 815
rect -158 781 -124 815
rect -124 781 -115 815
rect -167 772 -115 781
rect 2987 1014 3039 1023
rect 2987 980 2996 1014
rect 2996 980 3030 1014
rect 3030 980 3039 1014
rect 2987 971 3039 980
rect 4273 1046 4325 1055
rect 4273 1012 4282 1046
rect 4282 1012 4316 1046
rect 4316 1012 4325 1046
rect 4273 1003 4325 1012
rect 4345 1046 4397 1055
rect 4345 1012 4354 1046
rect 4354 1012 4388 1046
rect 4388 1012 4397 1046
rect 4345 1003 4397 1012
rect 4660 1046 4712 1055
rect 4660 1012 4669 1046
rect 4669 1012 4703 1046
rect 4703 1012 4712 1046
rect 4660 1003 4712 1012
rect 4732 1046 4784 1055
rect 4732 1012 4741 1046
rect 4741 1012 4775 1046
rect 4775 1012 4784 1046
rect 4732 1003 4784 1012
rect 3671 943 3723 952
rect 3671 909 3680 943
rect 3680 909 3714 943
rect 3714 909 3723 943
rect 3671 900 3723 909
rect 3671 871 3723 880
rect 3671 837 3680 871
rect 3680 837 3714 871
rect 3714 837 3723 871
rect 3671 828 3723 837
rect 240 640 660 700
rect 1440 640 1860 700
rect 2640 640 3060 700
rect 3840 640 4260 700
rect 496 342 548 351
rect 496 308 505 342
rect 505 308 539 342
rect 539 308 548 342
rect 496 299 548 308
rect 912 320 964 329
rect 912 286 921 320
rect 921 286 955 320
rect 955 286 964 320
rect 912 277 964 286
rect 3265 490 3317 499
rect 3265 456 3274 490
rect 3274 456 3308 490
rect 3308 456 3317 490
rect 3265 447 3317 456
rect 3265 418 3317 427
rect 3265 384 3274 418
rect 3274 384 3308 418
rect 3308 384 3317 418
rect 3265 375 3317 384
rect 3674 486 3726 495
rect 3674 452 3683 486
rect 3683 452 3717 486
rect 3717 452 3726 486
rect 3674 443 3726 452
rect 3674 414 3726 423
rect 3674 380 3683 414
rect 3683 380 3717 414
rect 3717 380 3726 414
rect 3674 371 3726 380
rect 2989 353 3041 362
rect 2989 319 2998 353
rect 2998 319 3032 353
rect 3032 319 3041 353
rect 2989 310 3041 319
rect 4253 341 4305 350
rect 4253 307 4262 341
rect 4262 307 4296 341
rect 4296 307 4305 341
rect 4253 298 4305 307
rect 4378 334 4430 343
rect 4378 300 4387 334
rect 4387 300 4421 334
rect 4421 300 4430 334
rect 4378 291 4430 300
rect 840 -40 1260 20
rect 2040 -40 2460 20
rect 3240 -40 3660 20
rect 4440 -40 4860 20
<< metal2 >>
rect -2280 2960 -996 3040
rect -2920 1580 -2820 1660
rect -2940 1000 -2840 1080
rect -2280 180 -2200 2960
rect -2320 160 -2200 180
rect -2320 80 -2300 160
rect -2220 80 -2200 160
rect -2320 60 -2200 80
rect -2280 -1460 -2200 60
rect -2140 2246 -986 2326
rect -2140 0 -2060 2246
rect 220 2040 680 2060
rect 220 1960 240 2040
rect 660 1960 680 2040
rect 220 1940 680 1960
rect 1420 2040 1880 2060
rect 1420 1960 1440 2040
rect 1860 1960 1880 2040
rect 1420 1940 1880 1960
rect 2620 2040 3080 2060
rect 2620 1960 2640 2040
rect 3060 1960 3080 2040
rect 2620 1940 3080 1960
rect 3820 2040 4280 2060
rect 3820 1960 3840 2040
rect 4260 1960 4280 2040
rect 3820 1940 4280 1960
rect -1204 1439 -1141 1461
rect -1204 1409 -613 1439
rect -1204 1238 -1141 1249
rect -1204 1208 -726 1238
rect -1204 1197 -1141 1208
rect -1144 1128 -910 1165
rect -1493 550 -1441 552
rect -1144 550 -1107 1128
rect -1051 1006 -1045 1058
rect -993 1006 -987 1058
rect -1045 970 -993 1006
rect -947 977 -910 1128
rect -756 1081 -726 1208
rect -643 1083 -613 1409
rect -480 1380 -20 1400
rect -480 1300 -460 1380
rect -40 1300 -20 1380
rect -480 1280 -20 1300
rect 820 1360 1280 1380
rect 820 1280 840 1360
rect 1260 1280 1280 1360
rect 820 1260 1280 1280
rect 2020 1360 2480 1380
rect 2020 1280 2040 1360
rect 2460 1280 2480 1360
rect 2020 1260 2480 1280
rect 3220 1360 3680 1380
rect 3220 1280 3240 1360
rect 3660 1280 3680 1360
rect 3220 1260 3680 1280
rect 4420 1360 4880 1380
rect 4420 1280 4440 1360
rect 4860 1280 4880 1360
rect 4420 1260 4880 1280
rect 767 1101 3033 1141
rect -774 1029 -768 1081
rect -716 1029 -710 1081
rect -660 1031 -654 1083
rect -602 1031 -596 1083
rect -267 1018 -261 1070
rect -209 1018 -203 1070
rect -259 977 -222 1018
rect -1038 581 -997 970
rect -947 940 -222 977
rect 767 908 807 1101
rect 902 1041 908 1055
rect -375 896 807 908
rect -375 844 -369 896
rect -317 868 807 896
rect 856 1003 908 1041
rect 960 1003 966 1055
rect 2993 1023 3033 1101
rect 4049 1107 4714 1144
rect -317 844 -310 868
rect 856 830 894 1003
rect 2981 971 2987 1023
rect 3039 971 3045 1023
rect -167 824 894 830
rect -115 792 894 824
rect 3671 952 3723 958
rect 3723 943 3740 952
rect 4049 943 4086 1107
rect 4677 1055 4714 1107
rect 4267 1003 4273 1055
rect 4325 1003 4345 1055
rect 4397 1003 4403 1055
rect 4654 1003 4660 1055
rect 4712 1003 4732 1055
rect 4784 1003 4790 1055
rect 3723 906 4086 943
rect 3723 900 3740 906
rect 3671 880 3723 900
rect 3671 822 3723 828
rect -167 766 -115 772
rect 220 720 680 740
rect 220 640 240 720
rect 660 640 680 720
rect 220 620 680 640
rect 1420 720 1880 740
rect 1420 640 1440 720
rect 1860 640 1880 720
rect 1420 620 1880 640
rect 2620 720 3080 740
rect 2620 640 2640 720
rect 3060 640 3080 720
rect 2620 620 3080 640
rect 3820 720 4280 740
rect 3820 640 3840 720
rect 4260 640 4280 720
rect 3820 620 4280 640
rect -1493 498 -1100 550
rect -1038 540 3370 581
rect -1980 340 -1860 360
rect -1980 260 -1960 340
rect -1880 260 -1640 340
rect -1493 319 -1441 498
rect -1572 267 -1441 319
rect -820 400 -400 420
rect -1980 240 -1860 260
rect -820 160 -800 400
rect -420 160 -400 400
rect 502 351 543 540
rect 3265 499 3370 540
rect 3317 447 3370 499
rect 3265 427 3370 447
rect 3317 416 3370 427
rect 3674 495 3726 501
rect 3674 423 3726 443
rect 4330 423 4363 1003
rect 3317 375 3594 416
rect 3265 369 3317 375
rect 490 299 496 351
rect 548 299 554 351
rect 906 325 912 329
rect -820 140 -400 160
rect 784 277 912 325
rect 964 277 970 329
rect 2983 310 2989 362
rect 3041 310 3047 362
rect 784 131 832 277
rect 2983 274 3047 310
rect 3549 327 3590 375
rect 3726 390 4363 423
rect 3726 371 3759 390
rect 3674 365 3726 371
rect 4205 350 4311 356
rect 4205 327 4253 350
rect 3549 298 4253 327
rect 4305 298 4311 350
rect 4700 343 4733 1003
rect 3549 290 4311 298
rect 4372 291 4378 343
rect 4430 291 4733 343
rect 3549 286 4205 290
rect -52 83 832 131
rect 820 20 1280 40
rect -2140 -20 -2020 0
rect -2140 -100 -2120 -20
rect -2040 -100 -2020 -20
rect 820 -60 840 20
rect 1260 -60 1280 20
rect 820 -80 1280 -60
rect 2020 20 2480 40
rect 2020 -60 2040 20
rect 2460 -60 2480 20
rect 2020 -80 2480 -60
rect 3220 20 3680 40
rect 3220 -60 3240 20
rect 3660 -60 3680 20
rect 3220 -80 3680 -60
rect 4420 20 4880 40
rect 4420 -60 4440 20
rect 4860 -60 4880 20
rect 4420 -80 4880 -60
rect -2140 -120 -2020 -100
rect -2140 -740 -2060 -120
rect -2140 -820 -1440 -740
rect -2280 -1540 -1380 -1460
<< via2 >>
rect -2300 80 -2220 160
rect 240 1960 660 2040
rect 1440 1960 1860 2040
rect 2640 1960 3060 2040
rect 3840 1960 4260 2040
rect -1960 1500 -1580 1720
rect -1960 940 -1580 1160
rect -460 1300 -40 1380
rect 840 1300 1260 1360
rect 840 1280 1260 1300
rect 2040 1300 2460 1360
rect 2040 1280 2460 1300
rect 3240 1300 3660 1360
rect 3240 1280 3660 1300
rect 4440 1300 4860 1360
rect 4440 1280 4860 1300
rect 240 700 660 720
rect 240 640 660 700
rect 1440 700 1860 720
rect 1440 640 1860 700
rect 2640 700 3060 720
rect 2640 640 3060 700
rect 3840 700 4260 720
rect 3840 640 4260 700
rect -1960 260 -1880 340
rect -800 160 -420 400
rect -2120 -100 -2040 -20
rect 840 -40 1260 20
rect 840 -60 1260 -40
rect 2040 -40 2460 20
rect 2040 -60 2460 -40
rect 3240 -40 3660 20
rect 3240 -60 3660 -40
rect 4440 -40 4860 20
rect 4440 -60 4860 -40
<< metal3 >>
rect -1980 1720 -1560 1740
rect -1980 1500 -1960 1720
rect -1580 1500 -1560 1720
rect -1980 1480 -1560 1500
rect -1420 1420 -1260 3460
rect 220 2040 4280 2060
rect 220 1960 240 2040
rect 660 1960 1440 2040
rect 1860 1960 2640 2040
rect 3060 1960 3840 2040
rect 4260 1960 4280 2040
rect 220 1940 4280 1960
rect -1420 1380 40 1420
rect -1420 1300 -460 1380
rect -40 1300 40 1380
rect -1420 1260 40 1300
rect -1980 1160 -1560 1180
rect -1980 940 -1960 1160
rect -1580 940 -1560 1160
rect -1980 920 -1560 940
rect -1420 820 -1260 1260
rect -1780 660 -1260 820
rect 220 740 340 1940
rect 560 740 680 1940
rect 220 720 680 740
rect -2480 340 -1860 360
rect -2480 260 -1960 340
rect -1880 260 -1860 340
rect -2480 240 -1860 260
rect -2480 160 -2200 180
rect -2480 80 -2300 160
rect -2220 80 -2200 160
rect -2480 60 -2200 80
rect -1780 40 -1620 660
rect 220 640 240 720
rect 660 640 680 720
rect 220 620 680 640
rect 820 1360 1280 1380
rect 820 1280 840 1360
rect 1260 1280 1280 1360
rect 820 1260 1280 1280
rect -820 400 -400 420
rect -820 160 -800 400
rect -420 160 -400 400
rect -820 140 -400 160
rect 820 40 940 1260
rect 1160 40 1280 1260
rect 1420 740 1540 1940
rect 1760 740 1880 1940
rect 1420 720 1880 740
rect 1420 640 1440 720
rect 1860 640 1880 720
rect 1420 620 1880 640
rect 2020 1360 2480 1380
rect 2020 1280 2040 1360
rect 2460 1280 2480 1360
rect 2020 1260 2480 1280
rect 2020 40 2140 1260
rect 2360 40 2480 1260
rect 2620 740 2740 1940
rect 2960 740 3080 1940
rect 2620 720 3080 740
rect 2620 640 2640 720
rect 3060 640 3080 720
rect 2620 620 3080 640
rect 3220 1360 3680 1380
rect 3220 1280 3240 1360
rect 3660 1280 3680 1360
rect 3220 1260 3680 1280
rect 3220 40 3340 1260
rect 3560 40 3680 1260
rect 3820 740 3940 1940
rect 4160 740 4280 1940
rect 3820 720 4280 740
rect 3820 640 3840 720
rect 4260 640 4280 720
rect 3820 620 4280 640
rect 4420 1360 4880 1380
rect 4420 1280 4440 1360
rect 4860 1280 4880 1360
rect 4420 1260 4880 1280
rect 4420 40 4540 1260
rect 4760 40 4880 1260
rect -1780 20 4880 40
rect -2480 -20 -2020 0
rect -2480 -100 -2120 -20
rect -2040 -100 -2020 -20
rect -2480 -120 -2020 -100
rect -1780 -60 840 20
rect 1260 -60 2040 20
rect 2460 -60 3240 20
rect 3660 -60 4440 20
rect 4860 -60 4880 20
rect -1780 -80 4880 -60
rect -1780 -1580 -1620 -80
<< via3 >>
rect -1960 1500 -1580 1720
rect -1960 940 -1580 1160
rect -800 160 -420 400
<< metal4 >>
rect -2500 1200 -2300 3400
rect -360 1760 -160 3460
rect -2000 1720 -160 1760
rect -2000 1500 -1960 1720
rect -1580 1560 -160 1720
rect -1580 1500 -1500 1560
rect -2000 1460 -1500 1500
rect -2500 1160 -1500 1200
rect -2500 1000 -1960 1160
rect -2000 940 -1960 1000
rect -1580 940 -1500 1160
rect -2000 900 -1500 940
rect -820 400 -400 420
rect -820 160 -800 400
rect -420 160 -400 400
rect -820 140 -400 160
rect -680 -1400 -480 140
use sky130_fd_sc_hs__and2_4  sky130_fd_sc_hs__and2_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1670771148
transform -1 0 4896 0 1 0
box -38 -49 902 715
use sky130_fd_sc_hs__decap_4  sky130_fd_sc_hs__decap_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1670771148
transform 1 0 4224 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_0 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1670771148
transform 1 0 -1152 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_2
timestamp 1670771148
transform 1 0 192 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_3
timestamp 1670771148
transform 1 0 864 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_4
timestamp 1670771148
transform 1 0 1536 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_6
timestamp 1670771148
transform 1 0 2880 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__decap_8  sky130_fd_sc_hs__decap_8_7
timestamp 1670771148
transform 1 0 3552 0 1 1332
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1670771148
transform 1 0 -96 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  sky130_fd_sc_hs__fill_1_1
timestamp 1670771148
transform 1 0 4800 0 1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  sky130_fd_sc_hs__fill_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1670771148
transform 1 0 4608 0 1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1670771148
transform 1 0 -480 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_1
timestamp 1670771148
transform 1 0 2112 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__fill_4  sky130_fd_sc_hs__fill_4_3
timestamp 1670771148
transform 1 0 2496 0 1 1332
box -38 -49 422 715
use sky130_fd_sc_hs__fill_diode_2  sky130_fd_sc_hs__fill_diode_2_1 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1670771148
transform 1 0 3840 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__fill_diode_2  sky130_fd_sc_hs__fill_diode_2_3
timestamp 1670771148
transform 1 0 3840 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__inv_2  sky130_fd_sc_hs__inv_2_1 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1670771148
transform 1 0 -288 0 -1 1332
box -38 -49 326 715
use sky130_fd_sc_hs__mux2_1  sky130_fd_sc_hs__mux2_1_1 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1670771148
transform 1 0 -1152 0 -1 1332
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_4  sky130_fd_sc_hs__nand2_4_3 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1670771148
transform 1 0 4032 0 -1 1332
box -38 -49 902 715
use sky130_fd_sc_hs__sdfbbn_2  sky130_fd_sc_hs__sdfbbn_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1670771148
transform 1 0 192 0 -1 1332
box -38 -49 3686 715
use sky130_fd_sc_hs__sdfbbn_2  sky130_fd_sc_hs__sdfbbn_2_1
timestamp 1670771148
transform 1 0 192 0 1 0
box -38 -49 3686 715
use sky130_fd_sc_hs__tapmet1_2  sky130_fd_sc_hs__tapmet1_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1670771148
transform 1 0 0 0 1 0
box -38 -49 230 715
use sky130_fd_sc_hs__tapmet1_2  sky130_fd_sc_hs__tapmet1_2_1
timestamp 1670771148
transform 1 0 0 0 -1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__tapmet1_2  sky130_fd_sc_hs__tapmet1_2_2
timestamp 1670771148
transform 1 0 0 0 1 1332
box -38 -49 230 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1670771148
transform 1 0 4896 0 1 0
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_2
timestamp 1670771148
transform 1 0 4896 0 -1 1332
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_3
timestamp 1670771148
transform 1 0 4896 0 1 1332
box -38 -49 134 715
use tcap_50f  tcap_50f_0
timestamp 1671378086
transform -1 0 -1519 0 1 2915
box -233 -53 2220 767
use tcap_50f  tcap_50f_2
timestamp 1671378086
transform 1 0 -1486 0 1 -855
box -233 -53 2220 767
use tcap_50f  tcap_50f_3
timestamp 1671378086
transform 1 0 -1053 0 1 2915
box -233 -53 2220 767
use tcap_100f  tcap_100f_0
timestamp 1671378102
transform -1 0 -1519 0 1 2201
box -233 -53 3790 767
use tcap_100f  tcap_100f_2
timestamp 1671378102
transform 1 0 -1486 0 1 -1569
box -233 -53 3790 767
use tcap_100f  tcap_100f_3
timestamp 1671378102
transform 1 0 -1053 0 1 2201
box -233 -53 3790 767
use twcon_tdly  twcon_tdly_0
timestamp 1671673121
transform 1 0 1365 0 1 216
box -3131 -265 -1327 499
use twcon_tdly  twcon_tdly_1
timestamp 1671673121
transform 1 0 213 0 -1 1116
box -3131 -265 -1327 499
use twcon_tdly  twcon_tdly_2
timestamp 1671673121
transform 1 0 213 0 1 1548
box -3131 -265 -1327 499
<< labels >>
rlabel metal2 3720 371 3759 423 1 UPDN
port 1 n
rlabel metal3 -2480 240 -2420 360 1 CLKIN
port 2 n
rlabel metal2 -2940 1000 -2840 1080 1 A0
port 3 n
rlabel metal2 -2920 1580 -2820 1660 1 A1
port 4 n
rlabel metal2 2983 274 3047 362 1 RSTB
port 5 n
rlabel metal3 720 2037 788 2060 1 VHI
port 6 n
rlabel metal3 -439 1396 -371 1419 1 VLO
port 7 n
rlabel metal3 -2480 60 -2420 180 1 C100
port 8 n
rlabel metal3 -2480 -120 -2420 0 1 C50
port 9 n
rlabel metal2 2 870 32 906 1 MUX_OUT
port 10 n
rlabel metal2 180 792 210 828 1 ENCLK
port 11 n
rlabel locali 4934 265 4974 345 1 GN
port 12 n
rlabel locali 4925 970 4965 1050 1 GP
port 13 n
<< end >>
