magic
tech sky130A
magscale 1 2
timestamp 1671166957
<< error_p >>
rect -560 1072 -502 1078
rect -442 1072 -384 1078
rect -324 1072 -266 1078
rect -206 1072 -148 1078
rect -88 1072 -30 1078
rect 30 1072 88 1078
rect 148 1072 206 1078
rect 266 1072 324 1078
rect 384 1072 442 1078
rect 502 1072 560 1078
rect -560 1038 -548 1072
rect -442 1038 -430 1072
rect -324 1038 -312 1072
rect -206 1038 -194 1072
rect -88 1038 -76 1072
rect 30 1038 42 1072
rect 148 1038 160 1072
rect 266 1038 278 1072
rect 384 1038 396 1072
rect 502 1038 514 1072
rect -560 1032 -502 1038
rect -442 1032 -384 1038
rect -324 1032 -266 1038
rect -206 1032 -148 1038
rect -88 1032 -30 1038
rect 30 1032 88 1038
rect 148 1032 206 1038
rect 266 1032 324 1038
rect 384 1032 442 1038
rect 502 1032 560 1038
rect -560 -1038 -502 -1032
rect -442 -1038 -384 -1032
rect -324 -1038 -266 -1032
rect -206 -1038 -148 -1032
rect -88 -1038 -30 -1032
rect 30 -1038 88 -1032
rect 148 -1038 206 -1032
rect 266 -1038 324 -1032
rect 384 -1038 442 -1032
rect 502 -1038 560 -1032
rect -560 -1072 -548 -1038
rect -442 -1072 -430 -1038
rect -324 -1072 -312 -1038
rect -206 -1072 -194 -1038
rect -88 -1072 -76 -1038
rect 30 -1072 42 -1038
rect 148 -1072 160 -1038
rect 266 -1072 278 -1038
rect 384 -1072 396 -1038
rect 502 -1072 514 -1038
rect -560 -1078 -502 -1072
rect -442 -1078 -384 -1072
rect -324 -1078 -266 -1072
rect -206 -1078 -148 -1072
rect -88 -1078 -30 -1072
rect 30 -1078 88 -1072
rect 148 -1078 206 -1072
rect 266 -1078 324 -1072
rect 384 -1078 442 -1072
rect 502 -1078 560 -1072
<< pwell >>
rect -757 -1210 757 1210
<< nmos >>
rect -561 -1000 -501 1000
rect -443 -1000 -383 1000
rect -325 -1000 -265 1000
rect -207 -1000 -147 1000
rect -89 -1000 -29 1000
rect 29 -1000 89 1000
rect 147 -1000 207 1000
rect 265 -1000 325 1000
rect 383 -1000 443 1000
rect 501 -1000 561 1000
<< ndiff >>
rect -619 988 -561 1000
rect -619 -988 -607 988
rect -573 -988 -561 988
rect -619 -1000 -561 -988
rect -501 988 -443 1000
rect -501 -988 -489 988
rect -455 -988 -443 988
rect -501 -1000 -443 -988
rect -383 988 -325 1000
rect -383 -988 -371 988
rect -337 -988 -325 988
rect -383 -1000 -325 -988
rect -265 988 -207 1000
rect -265 -988 -253 988
rect -219 -988 -207 988
rect -265 -1000 -207 -988
rect -147 988 -89 1000
rect -147 -988 -135 988
rect -101 -988 -89 988
rect -147 -1000 -89 -988
rect -29 988 29 1000
rect -29 -988 -17 988
rect 17 -988 29 988
rect -29 -1000 29 -988
rect 89 988 147 1000
rect 89 -988 101 988
rect 135 -988 147 988
rect 89 -1000 147 -988
rect 207 988 265 1000
rect 207 -988 219 988
rect 253 -988 265 988
rect 207 -1000 265 -988
rect 325 988 383 1000
rect 325 -988 337 988
rect 371 -988 383 988
rect 325 -1000 383 -988
rect 443 988 501 1000
rect 443 -988 455 988
rect 489 -988 501 988
rect 443 -1000 501 -988
rect 561 988 619 1000
rect 561 -988 573 988
rect 607 -988 619 988
rect 561 -1000 619 -988
<< ndiffc >>
rect -607 -988 -573 988
rect -489 -988 -455 988
rect -371 -988 -337 988
rect -253 -988 -219 988
rect -135 -988 -101 988
rect -17 -988 17 988
rect 101 -988 135 988
rect 219 -988 253 988
rect 337 -988 371 988
rect 455 -988 489 988
rect 573 -988 607 988
<< psubdiff >>
rect -721 1140 -625 1174
rect 625 1140 721 1174
rect -721 1078 -687 1140
rect 687 1078 721 1140
rect -721 -1140 -687 -1078
rect 687 -1140 721 -1078
rect -721 -1174 -625 -1140
rect 625 -1174 721 -1140
<< psubdiffcont >>
rect -625 1140 625 1174
rect -721 -1078 -687 1078
rect 687 -1078 721 1078
rect -625 -1174 625 -1140
<< poly >>
rect -564 1072 -498 1088
rect -564 1038 -548 1072
rect -514 1038 -498 1072
rect -564 1022 -498 1038
rect -446 1072 -380 1088
rect -446 1038 -430 1072
rect -396 1038 -380 1072
rect -446 1022 -380 1038
rect -328 1072 -262 1088
rect -328 1038 -312 1072
rect -278 1038 -262 1072
rect -328 1022 -262 1038
rect -210 1072 -144 1088
rect -210 1038 -194 1072
rect -160 1038 -144 1072
rect -210 1022 -144 1038
rect -92 1072 -26 1088
rect -92 1038 -76 1072
rect -42 1038 -26 1072
rect -92 1022 -26 1038
rect 26 1072 92 1088
rect 26 1038 42 1072
rect 76 1038 92 1072
rect 26 1022 92 1038
rect 144 1072 210 1088
rect 144 1038 160 1072
rect 194 1038 210 1072
rect 144 1022 210 1038
rect 262 1072 328 1088
rect 262 1038 278 1072
rect 312 1038 328 1072
rect 262 1022 328 1038
rect 380 1072 446 1088
rect 380 1038 396 1072
rect 430 1038 446 1072
rect 380 1022 446 1038
rect 498 1072 564 1088
rect 498 1038 514 1072
rect 548 1038 564 1072
rect 498 1022 564 1038
rect -561 1000 -501 1022
rect -443 1000 -383 1022
rect -325 1000 -265 1022
rect -207 1000 -147 1022
rect -89 1000 -29 1022
rect 29 1000 89 1022
rect 147 1000 207 1022
rect 265 1000 325 1022
rect 383 1000 443 1022
rect 501 1000 561 1022
rect -561 -1022 -501 -1000
rect -443 -1022 -383 -1000
rect -325 -1022 -265 -1000
rect -207 -1022 -147 -1000
rect -89 -1022 -29 -1000
rect 29 -1022 89 -1000
rect 147 -1022 207 -1000
rect 265 -1022 325 -1000
rect 383 -1022 443 -1000
rect 501 -1022 561 -1000
rect -564 -1038 -498 -1022
rect -564 -1072 -548 -1038
rect -514 -1072 -498 -1038
rect -564 -1088 -498 -1072
rect -446 -1038 -380 -1022
rect -446 -1072 -430 -1038
rect -396 -1072 -380 -1038
rect -446 -1088 -380 -1072
rect -328 -1038 -262 -1022
rect -328 -1072 -312 -1038
rect -278 -1072 -262 -1038
rect -328 -1088 -262 -1072
rect -210 -1038 -144 -1022
rect -210 -1072 -194 -1038
rect -160 -1072 -144 -1038
rect -210 -1088 -144 -1072
rect -92 -1038 -26 -1022
rect -92 -1072 -76 -1038
rect -42 -1072 -26 -1038
rect -92 -1088 -26 -1072
rect 26 -1038 92 -1022
rect 26 -1072 42 -1038
rect 76 -1072 92 -1038
rect 26 -1088 92 -1072
rect 144 -1038 210 -1022
rect 144 -1072 160 -1038
rect 194 -1072 210 -1038
rect 144 -1088 210 -1072
rect 262 -1038 328 -1022
rect 262 -1072 278 -1038
rect 312 -1072 328 -1038
rect 262 -1088 328 -1072
rect 380 -1038 446 -1022
rect 380 -1072 396 -1038
rect 430 -1072 446 -1038
rect 380 -1088 446 -1072
rect 498 -1038 564 -1022
rect 498 -1072 514 -1038
rect 548 -1072 564 -1038
rect 498 -1088 564 -1072
<< polycont >>
rect -548 1038 -514 1072
rect -430 1038 -396 1072
rect -312 1038 -278 1072
rect -194 1038 -160 1072
rect -76 1038 -42 1072
rect 42 1038 76 1072
rect 160 1038 194 1072
rect 278 1038 312 1072
rect 396 1038 430 1072
rect 514 1038 548 1072
rect -548 -1072 -514 -1038
rect -430 -1072 -396 -1038
rect -312 -1072 -278 -1038
rect -194 -1072 -160 -1038
rect -76 -1072 -42 -1038
rect 42 -1072 76 -1038
rect 160 -1072 194 -1038
rect 278 -1072 312 -1038
rect 396 -1072 430 -1038
rect 514 -1072 548 -1038
<< locali >>
rect -721 1140 -625 1174
rect 625 1140 721 1174
rect -721 1078 -687 1140
rect 687 1078 721 1140
rect -564 1038 -548 1072
rect -514 1038 -498 1072
rect -446 1038 -430 1072
rect -396 1038 -380 1072
rect -328 1038 -312 1072
rect -278 1038 -262 1072
rect -210 1038 -194 1072
rect -160 1038 -144 1072
rect -92 1038 -76 1072
rect -42 1038 -26 1072
rect 26 1038 42 1072
rect 76 1038 92 1072
rect 144 1038 160 1072
rect 194 1038 210 1072
rect 262 1038 278 1072
rect 312 1038 328 1072
rect 380 1038 396 1072
rect 430 1038 446 1072
rect 498 1038 514 1072
rect 548 1038 564 1072
rect -607 988 -573 1004
rect -607 -1004 -573 -988
rect -489 988 -455 1004
rect -489 -1004 -455 -988
rect -371 988 -337 1004
rect -371 -1004 -337 -988
rect -253 988 -219 1004
rect -253 -1004 -219 -988
rect -135 988 -101 1004
rect -135 -1004 -101 -988
rect -17 988 17 1004
rect -17 -1004 17 -988
rect 101 988 135 1004
rect 101 -1004 135 -988
rect 219 988 253 1004
rect 219 -1004 253 -988
rect 337 988 371 1004
rect 337 -1004 371 -988
rect 455 988 489 1004
rect 455 -1004 489 -988
rect 573 988 607 1004
rect 573 -1004 607 -988
rect -564 -1072 -548 -1038
rect -514 -1072 -498 -1038
rect -446 -1072 -430 -1038
rect -396 -1072 -380 -1038
rect -328 -1072 -312 -1038
rect -278 -1072 -262 -1038
rect -210 -1072 -194 -1038
rect -160 -1072 -144 -1038
rect -92 -1072 -76 -1038
rect -42 -1072 -26 -1038
rect 26 -1072 42 -1038
rect 76 -1072 92 -1038
rect 144 -1072 160 -1038
rect 194 -1072 210 -1038
rect 262 -1072 278 -1038
rect 312 -1072 328 -1038
rect 380 -1072 396 -1038
rect 430 -1072 446 -1038
rect 498 -1072 514 -1038
rect 548 -1072 564 -1038
rect -721 -1140 -687 -1078
rect 687 -1140 721 -1078
rect -721 -1174 -625 -1140
rect 625 -1174 721 -1140
<< viali >>
rect -548 1038 -514 1072
rect -430 1038 -396 1072
rect -312 1038 -278 1072
rect -194 1038 -160 1072
rect -76 1038 -42 1072
rect 42 1038 76 1072
rect 160 1038 194 1072
rect 278 1038 312 1072
rect 396 1038 430 1072
rect 514 1038 548 1072
rect -607 -988 -573 988
rect -489 -988 -455 988
rect -371 -988 -337 988
rect -253 -988 -219 988
rect -135 -988 -101 988
rect -17 -988 17 988
rect 101 -988 135 988
rect 219 -988 253 988
rect 337 -988 371 988
rect 455 -988 489 988
rect 573 -988 607 988
rect -548 -1072 -514 -1038
rect -430 -1072 -396 -1038
rect -312 -1072 -278 -1038
rect -194 -1072 -160 -1038
rect -76 -1072 -42 -1038
rect 42 -1072 76 -1038
rect 160 -1072 194 -1038
rect 278 -1072 312 -1038
rect 396 -1072 430 -1038
rect 514 -1072 548 -1038
<< metal1 >>
rect -560 1072 -502 1078
rect -560 1038 -548 1072
rect -514 1038 -502 1072
rect -560 1032 -502 1038
rect -442 1072 -384 1078
rect -442 1038 -430 1072
rect -396 1038 -384 1072
rect -442 1032 -384 1038
rect -324 1072 -266 1078
rect -324 1038 -312 1072
rect -278 1038 -266 1072
rect -324 1032 -266 1038
rect -206 1072 -148 1078
rect -206 1038 -194 1072
rect -160 1038 -148 1072
rect -206 1032 -148 1038
rect -88 1072 -30 1078
rect -88 1038 -76 1072
rect -42 1038 -30 1072
rect -88 1032 -30 1038
rect 30 1072 88 1078
rect 30 1038 42 1072
rect 76 1038 88 1072
rect 30 1032 88 1038
rect 148 1072 206 1078
rect 148 1038 160 1072
rect 194 1038 206 1072
rect 148 1032 206 1038
rect 266 1072 324 1078
rect 266 1038 278 1072
rect 312 1038 324 1072
rect 266 1032 324 1038
rect 384 1072 442 1078
rect 384 1038 396 1072
rect 430 1038 442 1072
rect 384 1032 442 1038
rect 502 1072 560 1078
rect 502 1038 514 1072
rect 548 1038 560 1072
rect 502 1032 560 1038
rect -613 988 -567 1000
rect -613 -988 -607 988
rect -573 -988 -567 988
rect -613 -1000 -567 -988
rect -495 988 -449 1000
rect -495 -988 -489 988
rect -455 -988 -449 988
rect -495 -1000 -449 -988
rect -377 988 -331 1000
rect -377 -988 -371 988
rect -337 -988 -331 988
rect -377 -1000 -331 -988
rect -259 988 -213 1000
rect -259 -988 -253 988
rect -219 -988 -213 988
rect -259 -1000 -213 -988
rect -141 988 -95 1000
rect -141 -988 -135 988
rect -101 -988 -95 988
rect -141 -1000 -95 -988
rect -23 988 23 1000
rect -23 -988 -17 988
rect 17 -988 23 988
rect -23 -1000 23 -988
rect 95 988 141 1000
rect 95 -988 101 988
rect 135 -988 141 988
rect 95 -1000 141 -988
rect 213 988 259 1000
rect 213 -988 219 988
rect 253 -988 259 988
rect 213 -1000 259 -988
rect 331 988 377 1000
rect 331 -988 337 988
rect 371 -988 377 988
rect 331 -1000 377 -988
rect 449 988 495 1000
rect 449 -988 455 988
rect 489 -988 495 988
rect 449 -1000 495 -988
rect 567 988 613 1000
rect 567 -988 573 988
rect 607 -988 613 988
rect 567 -1000 613 -988
rect -560 -1038 -502 -1032
rect -560 -1072 -548 -1038
rect -514 -1072 -502 -1038
rect -560 -1078 -502 -1072
rect -442 -1038 -384 -1032
rect -442 -1072 -430 -1038
rect -396 -1072 -384 -1038
rect -442 -1078 -384 -1072
rect -324 -1038 -266 -1032
rect -324 -1072 -312 -1038
rect -278 -1072 -266 -1038
rect -324 -1078 -266 -1072
rect -206 -1038 -148 -1032
rect -206 -1072 -194 -1038
rect -160 -1072 -148 -1038
rect -206 -1078 -148 -1072
rect -88 -1038 -30 -1032
rect -88 -1072 -76 -1038
rect -42 -1072 -30 -1038
rect -88 -1078 -30 -1072
rect 30 -1038 88 -1032
rect 30 -1072 42 -1038
rect 76 -1072 88 -1038
rect 30 -1078 88 -1072
rect 148 -1038 206 -1032
rect 148 -1072 160 -1038
rect 194 -1072 206 -1038
rect 148 -1078 206 -1072
rect 266 -1038 324 -1032
rect 266 -1072 278 -1038
rect 312 -1072 324 -1038
rect 266 -1078 324 -1072
rect 384 -1038 442 -1032
rect 384 -1072 396 -1038
rect 430 -1072 442 -1038
rect 384 -1078 442 -1072
rect 502 -1038 560 -1032
rect 502 -1072 514 -1038
rect 548 -1072 560 -1038
rect 502 -1078 560 -1072
<< properties >>
string FIXED_BBOX -704 -1157 704 1157
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 10 l 0.3 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
