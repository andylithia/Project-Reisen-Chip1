VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_pr__res_xhigh_po_0p35_FE9J4G
  CLASS BLOCK ;
  FOREIGN sky130_fd_pr__res_xhigh_po_0p35_FE9J4G ;
  ORIGIN 0.740 52.725 ;
  SIZE 1.480 BY 105.450 ;
  OBS
      LAYER pwell ;
        RECT -0.955 52.510 0.955 52.940 ;
        RECT -0.955 -52.510 -0.525 52.510 ;
        RECT 0.525 -52.510 0.955 52.510 ;
        RECT -0.955 -52.940 0.955 -52.510 ;
      LAYER li1 ;
        RECT -0.825 52.640 0.825 52.810 ;
        RECT -0.825 -52.640 -0.655 52.640 ;
        RECT -0.175 50.000 0.175 52.160 ;
        RECT -0.175 -52.160 0.175 -50.000 ;
        RECT 0.655 -52.640 0.825 52.640 ;
        RECT -0.825 -52.810 0.825 -52.640 ;
      LAYER mcon ;
        RECT -0.085 51.890 0.085 52.060 ;
        RECT -0.085 51.530 0.085 51.700 ;
        RECT -0.085 51.170 0.085 51.340 ;
        RECT -0.085 50.810 0.085 50.980 ;
        RECT -0.085 50.450 0.085 50.620 ;
        RECT -0.085 50.090 0.085 50.260 ;
        RECT -0.085 -50.265 0.085 -50.095 ;
        RECT -0.085 -50.625 0.085 -50.455 ;
        RECT -0.085 -50.985 0.085 -50.815 ;
        RECT -0.085 -51.345 0.085 -51.175 ;
        RECT -0.085 -51.705 0.085 -51.535 ;
        RECT -0.085 -52.065 0.085 -51.895 ;
      LAYER met1 ;
        RECT -0.125 50.025 0.125 52.130 ;
        RECT -0.125 -52.130 0.125 -50.025 ;
  END
END sky130_fd_pr__res_xhigh_po_0p35_FE9J4G
MACRO largecap1
  CLASS BLOCK ;
  FOREIGN largecap1 ;
  ORIGIN -219.000 -26.000 ;
  SIZE 1211.000 BY 208.000 ;
  PIN A
    PORT
      LAYER met5 ;
        RECT 219.000 128.000 219.950 133.000 ;
    END
  END A
  PIN VLO
    PORT
      LAYER met4 ;
        RECT 225.200 78.750 225.800 83.750 ;
    END
  END VLO
  PIN B
    PORT
      LAYER met5 ;
        RECT 219.000 27.000 219.950 32.000 ;
    END
  END B
  OBS
      LAYER pwell ;
        RECT 226.050 132.500 227.960 132.930 ;
        RECT 226.050 27.480 226.480 132.500 ;
        RECT 227.530 27.480 227.960 132.500 ;
        RECT 226.050 27.050 227.960 27.480 ;
      LAYER li1 ;
        RECT 226.180 132.630 227.830 132.800 ;
        RECT 226.180 83.750 226.350 132.630 ;
        RECT 226.830 129.990 227.180 132.150 ;
        RECT 225.700 78.750 226.350 83.750 ;
        RECT 226.180 27.350 226.350 78.750 ;
        RECT 226.830 27.830 227.180 29.990 ;
        RECT 227.660 27.350 227.830 132.630 ;
        RECT 226.180 27.180 227.830 27.350 ;
      LAYER mcon ;
        RECT 226.920 131.885 227.090 132.055 ;
        RECT 226.920 131.525 227.090 131.695 ;
        RECT 226.920 131.165 227.090 131.335 ;
        RECT 226.920 130.805 227.090 130.975 ;
        RECT 226.920 130.445 227.090 130.615 ;
        RECT 226.920 130.085 227.090 130.255 ;
        RECT 225.915 83.325 226.085 83.495 ;
        RECT 225.915 82.965 226.085 83.135 ;
        RECT 225.915 82.605 226.085 82.775 ;
        RECT 225.915 82.245 226.085 82.415 ;
        RECT 225.915 81.885 226.085 82.055 ;
        RECT 225.915 81.525 226.085 81.695 ;
        RECT 225.915 81.165 226.085 81.335 ;
        RECT 225.915 80.805 226.085 80.975 ;
        RECT 225.915 80.445 226.085 80.615 ;
        RECT 225.915 80.085 226.085 80.255 ;
        RECT 225.915 79.725 226.085 79.895 ;
        RECT 225.915 79.365 226.085 79.535 ;
        RECT 225.915 79.005 226.085 79.175 ;
        RECT 226.920 29.730 227.090 29.900 ;
        RECT 226.920 29.370 227.090 29.540 ;
        RECT 226.920 29.010 227.090 29.180 ;
        RECT 226.920 28.650 227.090 28.820 ;
        RECT 226.920 28.290 227.090 28.460 ;
        RECT 226.920 27.930 227.090 28.100 ;
      LAYER met1 ;
        RECT 226.800 130.000 227.200 132.200 ;
        RECT 225.700 78.750 226.300 83.750 ;
        RECT 226.800 27.800 227.200 30.000 ;
      LAYER via ;
        RECT 226.870 131.770 227.130 132.030 ;
        RECT 226.870 131.450 227.130 131.710 ;
        RECT 226.870 131.130 227.130 131.390 ;
        RECT 226.870 130.810 227.130 131.070 ;
        RECT 226.870 130.490 227.130 130.750 ;
        RECT 226.870 130.170 227.130 130.430 ;
        RECT 225.870 83.360 226.130 83.620 ;
        RECT 225.870 83.040 226.130 83.300 ;
        RECT 225.870 82.720 226.130 82.980 ;
        RECT 225.870 82.400 226.130 82.660 ;
        RECT 225.870 82.080 226.130 82.340 ;
        RECT 225.870 81.760 226.130 82.020 ;
        RECT 225.870 81.440 226.130 81.700 ;
        RECT 225.870 81.120 226.130 81.380 ;
        RECT 225.870 80.800 226.130 81.060 ;
        RECT 225.870 80.480 226.130 80.740 ;
        RECT 225.870 80.160 226.130 80.420 ;
        RECT 225.870 79.840 226.130 80.100 ;
        RECT 225.870 79.520 226.130 79.780 ;
        RECT 225.870 79.200 226.130 79.460 ;
        RECT 225.870 78.880 226.130 79.140 ;
        RECT 226.870 29.570 227.130 29.830 ;
        RECT 226.870 29.250 227.130 29.510 ;
        RECT 226.870 28.930 227.130 29.190 ;
        RECT 226.870 28.610 227.130 28.870 ;
        RECT 226.870 28.290 227.130 28.550 ;
        RECT 226.870 27.970 227.130 28.230 ;
      LAYER met2 ;
        RECT 226.650 130.000 227.350 132.200 ;
        RECT 225.700 78.750 226.300 83.750 ;
        RECT 226.650 27.800 227.350 30.000 ;
      LAYER via2 ;
        RECT 226.860 131.760 227.140 132.040 ;
        RECT 226.860 131.360 227.140 131.640 ;
        RECT 226.860 130.960 227.140 131.240 ;
        RECT 226.860 130.560 227.140 130.840 ;
        RECT 226.860 130.160 227.140 130.440 ;
        RECT 225.860 83.310 226.140 83.590 ;
        RECT 225.860 82.910 226.140 83.190 ;
        RECT 225.860 82.510 226.140 82.790 ;
        RECT 225.860 82.110 226.140 82.390 ;
        RECT 225.860 81.710 226.140 81.990 ;
        RECT 225.860 81.310 226.140 81.590 ;
        RECT 225.860 80.910 226.140 81.190 ;
        RECT 225.860 80.510 226.140 80.790 ;
        RECT 225.860 80.110 226.140 80.390 ;
        RECT 225.860 79.710 226.140 79.990 ;
        RECT 225.860 79.310 226.140 79.590 ;
        RECT 225.860 78.910 226.140 79.190 ;
        RECT 226.860 29.560 227.140 29.840 ;
        RECT 226.860 29.160 227.140 29.440 ;
        RECT 226.860 28.760 227.140 29.040 ;
        RECT 226.860 28.360 227.140 28.640 ;
        RECT 226.860 27.960 227.140 28.240 ;
      LAYER met3 ;
        RECT 230.000 230.000 1430.000 234.000 ;
        RECT 226.650 130.000 227.350 132.200 ;
        RECT 230.000 131.000 272.000 230.000 ;
        RECT 280.000 131.000 322.000 230.000 ;
        RECT 330.000 131.000 372.000 230.000 ;
        RECT 380.000 131.000 422.000 230.000 ;
        RECT 430.000 131.000 472.000 230.000 ;
        RECT 480.000 131.000 522.000 230.000 ;
        RECT 530.000 131.000 572.000 230.000 ;
        RECT 580.000 131.000 622.000 230.000 ;
        RECT 630.000 131.000 672.000 230.000 ;
        RECT 680.000 131.000 722.000 230.000 ;
        RECT 730.000 131.000 772.000 230.000 ;
        RECT 780.000 131.000 822.000 230.000 ;
        RECT 830.000 131.000 872.000 230.000 ;
        RECT 880.000 131.000 922.000 230.000 ;
        RECT 930.000 131.000 972.000 230.000 ;
        RECT 980.000 131.000 1022.000 230.000 ;
        RECT 1030.000 131.000 1072.000 230.000 ;
        RECT 1080.000 131.000 1122.000 230.000 ;
        RECT 1130.000 131.000 1172.000 230.000 ;
        RECT 1180.000 131.000 1222.000 230.000 ;
        RECT 1230.000 131.000 1272.000 230.000 ;
        RECT 1280.000 131.000 1322.000 230.000 ;
        RECT 1330.000 131.000 1372.000 230.000 ;
        RECT 1380.000 131.000 1422.000 230.000 ;
        RECT 238.000 129.000 272.000 131.000 ;
        RECT 288.000 129.000 322.000 131.000 ;
        RECT 338.000 129.000 372.000 131.000 ;
        RECT 388.000 129.000 422.000 131.000 ;
        RECT 438.000 129.000 472.000 131.000 ;
        RECT 488.000 129.000 522.000 131.000 ;
        RECT 538.000 129.000 572.000 131.000 ;
        RECT 588.000 129.000 622.000 131.000 ;
        RECT 638.000 129.000 672.000 131.000 ;
        RECT 688.000 129.000 722.000 131.000 ;
        RECT 738.000 129.000 772.000 131.000 ;
        RECT 788.000 129.000 822.000 131.000 ;
        RECT 838.000 129.000 872.000 131.000 ;
        RECT 888.000 129.000 922.000 131.000 ;
        RECT 938.000 129.000 972.000 131.000 ;
        RECT 988.000 129.000 1022.000 131.000 ;
        RECT 1038.000 129.000 1072.000 131.000 ;
        RECT 1088.000 129.000 1122.000 131.000 ;
        RECT 1138.000 129.000 1172.000 131.000 ;
        RECT 1188.000 129.000 1222.000 131.000 ;
        RECT 1238.000 129.000 1272.000 131.000 ;
        RECT 1288.000 129.000 1322.000 131.000 ;
        RECT 1338.000 129.000 1372.000 131.000 ;
        RECT 1388.000 129.000 1422.000 131.000 ;
        RECT 225.700 78.750 226.300 83.750 ;
        RECT 238.000 30.000 280.000 129.000 ;
        RECT 288.000 30.000 330.000 129.000 ;
        RECT 338.000 30.000 380.000 129.000 ;
        RECT 388.000 30.000 430.000 129.000 ;
        RECT 438.000 30.000 480.000 129.000 ;
        RECT 488.000 30.000 530.000 129.000 ;
        RECT 538.000 30.000 580.000 129.000 ;
        RECT 588.000 30.000 630.000 129.000 ;
        RECT 638.000 30.000 680.000 129.000 ;
        RECT 688.000 30.000 730.000 129.000 ;
        RECT 738.000 30.000 780.000 129.000 ;
        RECT 788.000 30.000 830.000 129.000 ;
        RECT 838.000 30.000 880.000 129.000 ;
        RECT 888.000 30.000 930.000 129.000 ;
        RECT 938.000 30.000 980.000 129.000 ;
        RECT 988.000 30.000 1030.000 129.000 ;
        RECT 1038.000 30.000 1080.000 129.000 ;
        RECT 1088.000 30.000 1130.000 129.000 ;
        RECT 1138.000 30.000 1180.000 129.000 ;
        RECT 1188.000 30.000 1230.000 129.000 ;
        RECT 1238.000 30.000 1280.000 129.000 ;
        RECT 1288.000 30.000 1330.000 129.000 ;
        RECT 1338.000 30.000 1380.000 129.000 ;
        RECT 1388.000 30.000 1430.000 129.000 ;
        RECT 226.650 27.800 227.350 30.000 ;
        RECT 230.000 26.000 1430.000 30.000 ;
      LAYER via3 ;
        RECT 235.040 232.240 274.960 233.760 ;
        RECT 285.040 232.240 324.960 233.760 ;
        RECT 335.040 232.240 374.960 233.760 ;
        RECT 385.040 232.240 424.960 233.760 ;
        RECT 435.040 232.240 474.960 233.760 ;
        RECT 485.040 232.240 524.960 233.760 ;
        RECT 535.040 232.240 574.960 233.760 ;
        RECT 585.040 232.240 624.960 233.760 ;
        RECT 635.040 232.240 674.960 233.760 ;
        RECT 685.040 232.240 724.960 233.760 ;
        RECT 735.040 232.240 774.960 233.760 ;
        RECT 785.040 232.240 824.960 233.760 ;
        RECT 835.040 232.240 874.960 233.760 ;
        RECT 885.040 232.240 924.960 233.760 ;
        RECT 935.040 232.240 974.960 233.760 ;
        RECT 985.040 232.240 1024.960 233.760 ;
        RECT 1035.040 232.240 1074.960 233.760 ;
        RECT 1085.040 232.240 1124.960 233.760 ;
        RECT 1135.040 232.240 1174.960 233.760 ;
        RECT 1185.040 232.240 1224.960 233.760 ;
        RECT 1235.040 232.240 1274.960 233.760 ;
        RECT 1285.040 232.240 1324.960 233.760 ;
        RECT 1335.040 232.240 1374.960 233.760 ;
        RECT 1385.040 232.240 1424.960 233.760 ;
        RECT 226.840 131.740 227.160 132.060 ;
        RECT 226.840 131.340 227.160 131.660 ;
        RECT 226.840 130.940 227.160 131.260 ;
        RECT 226.840 130.540 227.160 130.860 ;
        RECT 226.840 130.140 227.160 130.460 ;
        RECT 225.840 83.290 226.160 83.610 ;
        RECT 225.840 82.890 226.160 83.210 ;
        RECT 225.840 82.490 226.160 82.810 ;
        RECT 225.840 82.090 226.160 82.410 ;
        RECT 225.840 81.690 226.160 82.010 ;
        RECT 225.840 81.290 226.160 81.610 ;
        RECT 225.840 80.890 226.160 81.210 ;
        RECT 225.840 80.490 226.160 80.810 ;
        RECT 225.840 80.090 226.160 80.410 ;
        RECT 225.840 79.690 226.160 80.010 ;
        RECT 225.840 79.290 226.160 79.610 ;
        RECT 225.840 78.890 226.160 79.210 ;
        RECT 226.840 29.540 227.160 29.860 ;
        RECT 226.840 29.140 227.160 29.460 ;
        RECT 226.840 28.740 227.160 29.060 ;
        RECT 226.840 28.340 227.160 28.660 ;
        RECT 226.840 27.940 227.160 28.260 ;
        RECT 235.040 26.240 279.760 27.760 ;
        RECT 285.040 26.240 329.760 27.760 ;
        RECT 335.040 26.240 379.760 27.760 ;
        RECT 385.040 26.240 429.760 27.760 ;
        RECT 435.040 26.240 479.760 27.760 ;
        RECT 485.040 26.240 529.760 27.760 ;
        RECT 535.040 26.240 579.760 27.760 ;
        RECT 585.040 26.240 629.760 27.760 ;
        RECT 635.040 26.240 679.760 27.760 ;
        RECT 685.040 26.240 729.760 27.760 ;
        RECT 735.040 26.240 779.760 27.760 ;
        RECT 785.040 26.240 829.760 27.760 ;
        RECT 835.040 26.240 879.760 27.760 ;
        RECT 885.040 26.240 929.760 27.760 ;
        RECT 935.040 26.240 979.760 27.760 ;
        RECT 985.040 26.240 1029.760 27.760 ;
        RECT 1035.040 26.240 1079.760 27.760 ;
        RECT 1085.040 26.240 1129.760 27.760 ;
        RECT 1135.040 26.240 1179.760 27.760 ;
        RECT 1185.040 26.240 1229.760 27.760 ;
        RECT 1235.040 26.240 1279.760 27.760 ;
        RECT 1285.040 26.240 1329.760 27.760 ;
        RECT 1335.040 26.240 1379.760 27.760 ;
        RECT 1385.040 26.240 1429.760 27.760 ;
      LAYER met4 ;
        RECT 230.000 232.000 1430.000 234.000 ;
        RECT 230.000 228.000 1422.000 230.000 ;
        RECT 219.000 132.000 228.000 133.000 ;
        RECT 230.000 132.000 272.000 228.000 ;
        RECT 280.000 132.000 322.000 228.000 ;
        RECT 330.000 132.000 372.000 228.000 ;
        RECT 380.000 132.000 422.000 228.000 ;
        RECT 430.000 132.000 472.000 228.000 ;
        RECT 480.000 132.000 522.000 228.000 ;
        RECT 530.000 132.000 572.000 228.000 ;
        RECT 580.000 132.000 622.000 228.000 ;
        RECT 630.000 132.000 672.000 228.000 ;
        RECT 680.000 132.000 722.000 228.000 ;
        RECT 730.000 132.000 772.000 228.000 ;
        RECT 780.000 132.000 822.000 228.000 ;
        RECT 830.000 132.000 872.000 228.000 ;
        RECT 880.000 132.000 922.000 228.000 ;
        RECT 930.000 132.000 972.000 228.000 ;
        RECT 980.000 132.000 1022.000 228.000 ;
        RECT 1030.000 132.000 1072.000 228.000 ;
        RECT 1080.000 132.000 1122.000 228.000 ;
        RECT 1130.000 132.000 1172.000 228.000 ;
        RECT 1180.000 132.000 1222.000 228.000 ;
        RECT 1230.000 132.000 1272.000 228.000 ;
        RECT 1280.000 132.000 1322.000 228.000 ;
        RECT 1330.000 132.000 1372.000 228.000 ;
        RECT 1380.000 132.000 1422.000 228.000 ;
        RECT 219.000 129.000 1422.000 132.000 ;
        RECT 219.000 128.000 1430.000 129.000 ;
        RECT 225.800 78.750 226.300 83.750 ;
        RECT 238.000 32.000 280.000 128.000 ;
        RECT 288.000 32.000 330.000 128.000 ;
        RECT 338.000 32.000 380.000 128.000 ;
        RECT 388.000 32.000 430.000 128.000 ;
        RECT 438.000 32.000 480.000 128.000 ;
        RECT 488.000 32.000 530.000 128.000 ;
        RECT 538.000 32.000 580.000 128.000 ;
        RECT 588.000 32.000 630.000 128.000 ;
        RECT 638.000 32.000 680.000 128.000 ;
        RECT 688.000 32.000 730.000 128.000 ;
        RECT 738.000 32.000 780.000 128.000 ;
        RECT 788.000 32.000 830.000 128.000 ;
        RECT 838.000 32.000 880.000 128.000 ;
        RECT 888.000 32.000 930.000 128.000 ;
        RECT 938.000 32.000 980.000 128.000 ;
        RECT 988.000 32.000 1030.000 128.000 ;
        RECT 1038.000 32.000 1080.000 128.000 ;
        RECT 1088.000 32.000 1130.000 128.000 ;
        RECT 1138.000 32.000 1180.000 128.000 ;
        RECT 1188.000 32.000 1230.000 128.000 ;
        RECT 1238.000 32.000 1280.000 128.000 ;
        RECT 1288.000 32.000 1330.000 128.000 ;
        RECT 1338.000 32.000 1380.000 128.000 ;
        RECT 1388.000 32.000 1430.000 128.000 ;
        RECT 219.000 29.000 228.000 32.000 ;
        RECT 238.000 30.000 1430.000 32.000 ;
        RECT 219.000 28.000 230.000 29.000 ;
        RECT 219.000 27.000 1430.000 28.000 ;
        RECT 230.000 26.000 1430.000 27.000 ;
      LAYER via4 ;
        RECT 235.210 232.410 236.390 233.590 ;
        RECT 236.810 232.410 237.990 233.590 ;
        RECT 238.410 232.410 239.590 233.590 ;
        RECT 240.010 232.410 241.190 233.590 ;
        RECT 241.610 232.410 242.790 233.590 ;
        RECT 243.210 232.410 244.390 233.590 ;
        RECT 244.810 232.410 245.990 233.590 ;
        RECT 246.410 232.410 247.590 233.590 ;
        RECT 248.010 232.410 249.190 233.590 ;
        RECT 249.610 232.410 250.790 233.590 ;
        RECT 251.210 232.410 252.390 233.590 ;
        RECT 252.810 232.410 253.990 233.590 ;
        RECT 254.410 232.410 255.590 233.590 ;
        RECT 256.010 232.410 257.190 233.590 ;
        RECT 257.610 232.410 258.790 233.590 ;
        RECT 259.210 232.410 260.390 233.590 ;
        RECT 260.810 232.410 261.990 233.590 ;
        RECT 262.410 232.410 263.590 233.590 ;
        RECT 264.010 232.410 265.190 233.590 ;
        RECT 265.610 232.410 266.790 233.590 ;
        RECT 267.210 232.410 268.390 233.590 ;
        RECT 268.810 232.410 269.990 233.590 ;
        RECT 270.410 232.410 271.590 233.590 ;
        RECT 272.010 232.410 273.190 233.590 ;
        RECT 273.610 232.410 274.790 233.590 ;
        RECT 285.210 232.410 286.390 233.590 ;
        RECT 286.810 232.410 287.990 233.590 ;
        RECT 288.410 232.410 289.590 233.590 ;
        RECT 290.010 232.410 291.190 233.590 ;
        RECT 291.610 232.410 292.790 233.590 ;
        RECT 293.210 232.410 294.390 233.590 ;
        RECT 294.810 232.410 295.990 233.590 ;
        RECT 296.410 232.410 297.590 233.590 ;
        RECT 298.010 232.410 299.190 233.590 ;
        RECT 299.610 232.410 300.790 233.590 ;
        RECT 301.210 232.410 302.390 233.590 ;
        RECT 302.810 232.410 303.990 233.590 ;
        RECT 304.410 232.410 305.590 233.590 ;
        RECT 306.010 232.410 307.190 233.590 ;
        RECT 307.610 232.410 308.790 233.590 ;
        RECT 309.210 232.410 310.390 233.590 ;
        RECT 310.810 232.410 311.990 233.590 ;
        RECT 312.410 232.410 313.590 233.590 ;
        RECT 314.010 232.410 315.190 233.590 ;
        RECT 315.610 232.410 316.790 233.590 ;
        RECT 317.210 232.410 318.390 233.590 ;
        RECT 318.810 232.410 319.990 233.590 ;
        RECT 320.410 232.410 321.590 233.590 ;
        RECT 322.010 232.410 323.190 233.590 ;
        RECT 323.610 232.410 324.790 233.590 ;
        RECT 335.210 232.410 336.390 233.590 ;
        RECT 336.810 232.410 337.990 233.590 ;
        RECT 338.410 232.410 339.590 233.590 ;
        RECT 340.010 232.410 341.190 233.590 ;
        RECT 341.610 232.410 342.790 233.590 ;
        RECT 343.210 232.410 344.390 233.590 ;
        RECT 344.810 232.410 345.990 233.590 ;
        RECT 346.410 232.410 347.590 233.590 ;
        RECT 348.010 232.410 349.190 233.590 ;
        RECT 349.610 232.410 350.790 233.590 ;
        RECT 351.210 232.410 352.390 233.590 ;
        RECT 352.810 232.410 353.990 233.590 ;
        RECT 354.410 232.410 355.590 233.590 ;
        RECT 356.010 232.410 357.190 233.590 ;
        RECT 357.610 232.410 358.790 233.590 ;
        RECT 359.210 232.410 360.390 233.590 ;
        RECT 360.810 232.410 361.990 233.590 ;
        RECT 362.410 232.410 363.590 233.590 ;
        RECT 364.010 232.410 365.190 233.590 ;
        RECT 365.610 232.410 366.790 233.590 ;
        RECT 367.210 232.410 368.390 233.590 ;
        RECT 368.810 232.410 369.990 233.590 ;
        RECT 370.410 232.410 371.590 233.590 ;
        RECT 372.010 232.410 373.190 233.590 ;
        RECT 373.610 232.410 374.790 233.590 ;
        RECT 385.210 232.410 386.390 233.590 ;
        RECT 386.810 232.410 387.990 233.590 ;
        RECT 388.410 232.410 389.590 233.590 ;
        RECT 390.010 232.410 391.190 233.590 ;
        RECT 391.610 232.410 392.790 233.590 ;
        RECT 393.210 232.410 394.390 233.590 ;
        RECT 394.810 232.410 395.990 233.590 ;
        RECT 396.410 232.410 397.590 233.590 ;
        RECT 398.010 232.410 399.190 233.590 ;
        RECT 399.610 232.410 400.790 233.590 ;
        RECT 401.210 232.410 402.390 233.590 ;
        RECT 402.810 232.410 403.990 233.590 ;
        RECT 404.410 232.410 405.590 233.590 ;
        RECT 406.010 232.410 407.190 233.590 ;
        RECT 407.610 232.410 408.790 233.590 ;
        RECT 409.210 232.410 410.390 233.590 ;
        RECT 410.810 232.410 411.990 233.590 ;
        RECT 412.410 232.410 413.590 233.590 ;
        RECT 414.010 232.410 415.190 233.590 ;
        RECT 415.610 232.410 416.790 233.590 ;
        RECT 417.210 232.410 418.390 233.590 ;
        RECT 418.810 232.410 419.990 233.590 ;
        RECT 420.410 232.410 421.590 233.590 ;
        RECT 422.010 232.410 423.190 233.590 ;
        RECT 423.610 232.410 424.790 233.590 ;
        RECT 435.210 232.410 436.390 233.590 ;
        RECT 436.810 232.410 437.990 233.590 ;
        RECT 438.410 232.410 439.590 233.590 ;
        RECT 440.010 232.410 441.190 233.590 ;
        RECT 441.610 232.410 442.790 233.590 ;
        RECT 443.210 232.410 444.390 233.590 ;
        RECT 444.810 232.410 445.990 233.590 ;
        RECT 446.410 232.410 447.590 233.590 ;
        RECT 448.010 232.410 449.190 233.590 ;
        RECT 449.610 232.410 450.790 233.590 ;
        RECT 451.210 232.410 452.390 233.590 ;
        RECT 452.810 232.410 453.990 233.590 ;
        RECT 454.410 232.410 455.590 233.590 ;
        RECT 456.010 232.410 457.190 233.590 ;
        RECT 457.610 232.410 458.790 233.590 ;
        RECT 459.210 232.410 460.390 233.590 ;
        RECT 460.810 232.410 461.990 233.590 ;
        RECT 462.410 232.410 463.590 233.590 ;
        RECT 464.010 232.410 465.190 233.590 ;
        RECT 465.610 232.410 466.790 233.590 ;
        RECT 467.210 232.410 468.390 233.590 ;
        RECT 468.810 232.410 469.990 233.590 ;
        RECT 470.410 232.410 471.590 233.590 ;
        RECT 472.010 232.410 473.190 233.590 ;
        RECT 473.610 232.410 474.790 233.590 ;
        RECT 485.210 232.410 486.390 233.590 ;
        RECT 486.810 232.410 487.990 233.590 ;
        RECT 488.410 232.410 489.590 233.590 ;
        RECT 490.010 232.410 491.190 233.590 ;
        RECT 491.610 232.410 492.790 233.590 ;
        RECT 493.210 232.410 494.390 233.590 ;
        RECT 494.810 232.410 495.990 233.590 ;
        RECT 496.410 232.410 497.590 233.590 ;
        RECT 498.010 232.410 499.190 233.590 ;
        RECT 499.610 232.410 500.790 233.590 ;
        RECT 501.210 232.410 502.390 233.590 ;
        RECT 502.810 232.410 503.990 233.590 ;
        RECT 504.410 232.410 505.590 233.590 ;
        RECT 506.010 232.410 507.190 233.590 ;
        RECT 507.610 232.410 508.790 233.590 ;
        RECT 509.210 232.410 510.390 233.590 ;
        RECT 510.810 232.410 511.990 233.590 ;
        RECT 512.410 232.410 513.590 233.590 ;
        RECT 514.010 232.410 515.190 233.590 ;
        RECT 515.610 232.410 516.790 233.590 ;
        RECT 517.210 232.410 518.390 233.590 ;
        RECT 518.810 232.410 519.990 233.590 ;
        RECT 520.410 232.410 521.590 233.590 ;
        RECT 522.010 232.410 523.190 233.590 ;
        RECT 523.610 232.410 524.790 233.590 ;
        RECT 535.210 232.410 536.390 233.590 ;
        RECT 536.810 232.410 537.990 233.590 ;
        RECT 538.410 232.410 539.590 233.590 ;
        RECT 540.010 232.410 541.190 233.590 ;
        RECT 541.610 232.410 542.790 233.590 ;
        RECT 543.210 232.410 544.390 233.590 ;
        RECT 544.810 232.410 545.990 233.590 ;
        RECT 546.410 232.410 547.590 233.590 ;
        RECT 548.010 232.410 549.190 233.590 ;
        RECT 549.610 232.410 550.790 233.590 ;
        RECT 551.210 232.410 552.390 233.590 ;
        RECT 552.810 232.410 553.990 233.590 ;
        RECT 554.410 232.410 555.590 233.590 ;
        RECT 556.010 232.410 557.190 233.590 ;
        RECT 557.610 232.410 558.790 233.590 ;
        RECT 559.210 232.410 560.390 233.590 ;
        RECT 560.810 232.410 561.990 233.590 ;
        RECT 562.410 232.410 563.590 233.590 ;
        RECT 564.010 232.410 565.190 233.590 ;
        RECT 565.610 232.410 566.790 233.590 ;
        RECT 567.210 232.410 568.390 233.590 ;
        RECT 568.810 232.410 569.990 233.590 ;
        RECT 570.410 232.410 571.590 233.590 ;
        RECT 572.010 232.410 573.190 233.590 ;
        RECT 573.610 232.410 574.790 233.590 ;
        RECT 585.210 232.410 586.390 233.590 ;
        RECT 586.810 232.410 587.990 233.590 ;
        RECT 588.410 232.410 589.590 233.590 ;
        RECT 590.010 232.410 591.190 233.590 ;
        RECT 591.610 232.410 592.790 233.590 ;
        RECT 593.210 232.410 594.390 233.590 ;
        RECT 594.810 232.410 595.990 233.590 ;
        RECT 596.410 232.410 597.590 233.590 ;
        RECT 598.010 232.410 599.190 233.590 ;
        RECT 599.610 232.410 600.790 233.590 ;
        RECT 601.210 232.410 602.390 233.590 ;
        RECT 602.810 232.410 603.990 233.590 ;
        RECT 604.410 232.410 605.590 233.590 ;
        RECT 606.010 232.410 607.190 233.590 ;
        RECT 607.610 232.410 608.790 233.590 ;
        RECT 609.210 232.410 610.390 233.590 ;
        RECT 610.810 232.410 611.990 233.590 ;
        RECT 612.410 232.410 613.590 233.590 ;
        RECT 614.010 232.410 615.190 233.590 ;
        RECT 615.610 232.410 616.790 233.590 ;
        RECT 617.210 232.410 618.390 233.590 ;
        RECT 618.810 232.410 619.990 233.590 ;
        RECT 620.410 232.410 621.590 233.590 ;
        RECT 622.010 232.410 623.190 233.590 ;
        RECT 623.610 232.410 624.790 233.590 ;
        RECT 635.210 232.410 636.390 233.590 ;
        RECT 636.810 232.410 637.990 233.590 ;
        RECT 638.410 232.410 639.590 233.590 ;
        RECT 640.010 232.410 641.190 233.590 ;
        RECT 641.610 232.410 642.790 233.590 ;
        RECT 643.210 232.410 644.390 233.590 ;
        RECT 644.810 232.410 645.990 233.590 ;
        RECT 646.410 232.410 647.590 233.590 ;
        RECT 648.010 232.410 649.190 233.590 ;
        RECT 649.610 232.410 650.790 233.590 ;
        RECT 651.210 232.410 652.390 233.590 ;
        RECT 652.810 232.410 653.990 233.590 ;
        RECT 654.410 232.410 655.590 233.590 ;
        RECT 656.010 232.410 657.190 233.590 ;
        RECT 657.610 232.410 658.790 233.590 ;
        RECT 659.210 232.410 660.390 233.590 ;
        RECT 660.810 232.410 661.990 233.590 ;
        RECT 662.410 232.410 663.590 233.590 ;
        RECT 664.010 232.410 665.190 233.590 ;
        RECT 665.610 232.410 666.790 233.590 ;
        RECT 667.210 232.410 668.390 233.590 ;
        RECT 668.810 232.410 669.990 233.590 ;
        RECT 670.410 232.410 671.590 233.590 ;
        RECT 672.010 232.410 673.190 233.590 ;
        RECT 673.610 232.410 674.790 233.590 ;
        RECT 685.210 232.410 686.390 233.590 ;
        RECT 686.810 232.410 687.990 233.590 ;
        RECT 688.410 232.410 689.590 233.590 ;
        RECT 690.010 232.410 691.190 233.590 ;
        RECT 691.610 232.410 692.790 233.590 ;
        RECT 693.210 232.410 694.390 233.590 ;
        RECT 694.810 232.410 695.990 233.590 ;
        RECT 696.410 232.410 697.590 233.590 ;
        RECT 698.010 232.410 699.190 233.590 ;
        RECT 699.610 232.410 700.790 233.590 ;
        RECT 701.210 232.410 702.390 233.590 ;
        RECT 702.810 232.410 703.990 233.590 ;
        RECT 704.410 232.410 705.590 233.590 ;
        RECT 706.010 232.410 707.190 233.590 ;
        RECT 707.610 232.410 708.790 233.590 ;
        RECT 709.210 232.410 710.390 233.590 ;
        RECT 710.810 232.410 711.990 233.590 ;
        RECT 712.410 232.410 713.590 233.590 ;
        RECT 714.010 232.410 715.190 233.590 ;
        RECT 715.610 232.410 716.790 233.590 ;
        RECT 717.210 232.410 718.390 233.590 ;
        RECT 718.810 232.410 719.990 233.590 ;
        RECT 720.410 232.410 721.590 233.590 ;
        RECT 722.010 232.410 723.190 233.590 ;
        RECT 723.610 232.410 724.790 233.590 ;
        RECT 735.210 232.410 736.390 233.590 ;
        RECT 736.810 232.410 737.990 233.590 ;
        RECT 738.410 232.410 739.590 233.590 ;
        RECT 740.010 232.410 741.190 233.590 ;
        RECT 741.610 232.410 742.790 233.590 ;
        RECT 743.210 232.410 744.390 233.590 ;
        RECT 744.810 232.410 745.990 233.590 ;
        RECT 746.410 232.410 747.590 233.590 ;
        RECT 748.010 232.410 749.190 233.590 ;
        RECT 749.610 232.410 750.790 233.590 ;
        RECT 751.210 232.410 752.390 233.590 ;
        RECT 752.810 232.410 753.990 233.590 ;
        RECT 754.410 232.410 755.590 233.590 ;
        RECT 756.010 232.410 757.190 233.590 ;
        RECT 757.610 232.410 758.790 233.590 ;
        RECT 759.210 232.410 760.390 233.590 ;
        RECT 760.810 232.410 761.990 233.590 ;
        RECT 762.410 232.410 763.590 233.590 ;
        RECT 764.010 232.410 765.190 233.590 ;
        RECT 765.610 232.410 766.790 233.590 ;
        RECT 767.210 232.410 768.390 233.590 ;
        RECT 768.810 232.410 769.990 233.590 ;
        RECT 770.410 232.410 771.590 233.590 ;
        RECT 772.010 232.410 773.190 233.590 ;
        RECT 773.610 232.410 774.790 233.590 ;
        RECT 785.210 232.410 786.390 233.590 ;
        RECT 786.810 232.410 787.990 233.590 ;
        RECT 788.410 232.410 789.590 233.590 ;
        RECT 790.010 232.410 791.190 233.590 ;
        RECT 791.610 232.410 792.790 233.590 ;
        RECT 793.210 232.410 794.390 233.590 ;
        RECT 794.810 232.410 795.990 233.590 ;
        RECT 796.410 232.410 797.590 233.590 ;
        RECT 798.010 232.410 799.190 233.590 ;
        RECT 799.610 232.410 800.790 233.590 ;
        RECT 801.210 232.410 802.390 233.590 ;
        RECT 802.810 232.410 803.990 233.590 ;
        RECT 804.410 232.410 805.590 233.590 ;
        RECT 806.010 232.410 807.190 233.590 ;
        RECT 807.610 232.410 808.790 233.590 ;
        RECT 809.210 232.410 810.390 233.590 ;
        RECT 810.810 232.410 811.990 233.590 ;
        RECT 812.410 232.410 813.590 233.590 ;
        RECT 814.010 232.410 815.190 233.590 ;
        RECT 815.610 232.410 816.790 233.590 ;
        RECT 817.210 232.410 818.390 233.590 ;
        RECT 818.810 232.410 819.990 233.590 ;
        RECT 820.410 232.410 821.590 233.590 ;
        RECT 822.010 232.410 823.190 233.590 ;
        RECT 823.610 232.410 824.790 233.590 ;
        RECT 835.210 232.410 836.390 233.590 ;
        RECT 836.810 232.410 837.990 233.590 ;
        RECT 838.410 232.410 839.590 233.590 ;
        RECT 840.010 232.410 841.190 233.590 ;
        RECT 841.610 232.410 842.790 233.590 ;
        RECT 843.210 232.410 844.390 233.590 ;
        RECT 844.810 232.410 845.990 233.590 ;
        RECT 846.410 232.410 847.590 233.590 ;
        RECT 848.010 232.410 849.190 233.590 ;
        RECT 849.610 232.410 850.790 233.590 ;
        RECT 851.210 232.410 852.390 233.590 ;
        RECT 852.810 232.410 853.990 233.590 ;
        RECT 854.410 232.410 855.590 233.590 ;
        RECT 856.010 232.410 857.190 233.590 ;
        RECT 857.610 232.410 858.790 233.590 ;
        RECT 859.210 232.410 860.390 233.590 ;
        RECT 860.810 232.410 861.990 233.590 ;
        RECT 862.410 232.410 863.590 233.590 ;
        RECT 864.010 232.410 865.190 233.590 ;
        RECT 865.610 232.410 866.790 233.590 ;
        RECT 867.210 232.410 868.390 233.590 ;
        RECT 868.810 232.410 869.990 233.590 ;
        RECT 870.410 232.410 871.590 233.590 ;
        RECT 872.010 232.410 873.190 233.590 ;
        RECT 873.610 232.410 874.790 233.590 ;
        RECT 885.210 232.410 886.390 233.590 ;
        RECT 886.810 232.410 887.990 233.590 ;
        RECT 888.410 232.410 889.590 233.590 ;
        RECT 890.010 232.410 891.190 233.590 ;
        RECT 891.610 232.410 892.790 233.590 ;
        RECT 893.210 232.410 894.390 233.590 ;
        RECT 894.810 232.410 895.990 233.590 ;
        RECT 896.410 232.410 897.590 233.590 ;
        RECT 898.010 232.410 899.190 233.590 ;
        RECT 899.610 232.410 900.790 233.590 ;
        RECT 901.210 232.410 902.390 233.590 ;
        RECT 902.810 232.410 903.990 233.590 ;
        RECT 904.410 232.410 905.590 233.590 ;
        RECT 906.010 232.410 907.190 233.590 ;
        RECT 907.610 232.410 908.790 233.590 ;
        RECT 909.210 232.410 910.390 233.590 ;
        RECT 910.810 232.410 911.990 233.590 ;
        RECT 912.410 232.410 913.590 233.590 ;
        RECT 914.010 232.410 915.190 233.590 ;
        RECT 915.610 232.410 916.790 233.590 ;
        RECT 917.210 232.410 918.390 233.590 ;
        RECT 918.810 232.410 919.990 233.590 ;
        RECT 920.410 232.410 921.590 233.590 ;
        RECT 922.010 232.410 923.190 233.590 ;
        RECT 923.610 232.410 924.790 233.590 ;
        RECT 935.210 232.410 936.390 233.590 ;
        RECT 936.810 232.410 937.990 233.590 ;
        RECT 938.410 232.410 939.590 233.590 ;
        RECT 940.010 232.410 941.190 233.590 ;
        RECT 941.610 232.410 942.790 233.590 ;
        RECT 943.210 232.410 944.390 233.590 ;
        RECT 944.810 232.410 945.990 233.590 ;
        RECT 946.410 232.410 947.590 233.590 ;
        RECT 948.010 232.410 949.190 233.590 ;
        RECT 949.610 232.410 950.790 233.590 ;
        RECT 951.210 232.410 952.390 233.590 ;
        RECT 952.810 232.410 953.990 233.590 ;
        RECT 954.410 232.410 955.590 233.590 ;
        RECT 956.010 232.410 957.190 233.590 ;
        RECT 957.610 232.410 958.790 233.590 ;
        RECT 959.210 232.410 960.390 233.590 ;
        RECT 960.810 232.410 961.990 233.590 ;
        RECT 962.410 232.410 963.590 233.590 ;
        RECT 964.010 232.410 965.190 233.590 ;
        RECT 965.610 232.410 966.790 233.590 ;
        RECT 967.210 232.410 968.390 233.590 ;
        RECT 968.810 232.410 969.990 233.590 ;
        RECT 970.410 232.410 971.590 233.590 ;
        RECT 972.010 232.410 973.190 233.590 ;
        RECT 973.610 232.410 974.790 233.590 ;
        RECT 985.210 232.410 986.390 233.590 ;
        RECT 986.810 232.410 987.990 233.590 ;
        RECT 988.410 232.410 989.590 233.590 ;
        RECT 990.010 232.410 991.190 233.590 ;
        RECT 991.610 232.410 992.790 233.590 ;
        RECT 993.210 232.410 994.390 233.590 ;
        RECT 994.810 232.410 995.990 233.590 ;
        RECT 996.410 232.410 997.590 233.590 ;
        RECT 998.010 232.410 999.190 233.590 ;
        RECT 999.610 232.410 1000.790 233.590 ;
        RECT 1001.210 232.410 1002.390 233.590 ;
        RECT 1002.810 232.410 1003.990 233.590 ;
        RECT 1004.410 232.410 1005.590 233.590 ;
        RECT 1006.010 232.410 1007.190 233.590 ;
        RECT 1007.610 232.410 1008.790 233.590 ;
        RECT 1009.210 232.410 1010.390 233.590 ;
        RECT 1010.810 232.410 1011.990 233.590 ;
        RECT 1012.410 232.410 1013.590 233.590 ;
        RECT 1014.010 232.410 1015.190 233.590 ;
        RECT 1015.610 232.410 1016.790 233.590 ;
        RECT 1017.210 232.410 1018.390 233.590 ;
        RECT 1018.810 232.410 1019.990 233.590 ;
        RECT 1020.410 232.410 1021.590 233.590 ;
        RECT 1022.010 232.410 1023.190 233.590 ;
        RECT 1023.610 232.410 1024.790 233.590 ;
        RECT 1035.210 232.410 1036.390 233.590 ;
        RECT 1036.810 232.410 1037.990 233.590 ;
        RECT 1038.410 232.410 1039.590 233.590 ;
        RECT 1040.010 232.410 1041.190 233.590 ;
        RECT 1041.610 232.410 1042.790 233.590 ;
        RECT 1043.210 232.410 1044.390 233.590 ;
        RECT 1044.810 232.410 1045.990 233.590 ;
        RECT 1046.410 232.410 1047.590 233.590 ;
        RECT 1048.010 232.410 1049.190 233.590 ;
        RECT 1049.610 232.410 1050.790 233.590 ;
        RECT 1051.210 232.410 1052.390 233.590 ;
        RECT 1052.810 232.410 1053.990 233.590 ;
        RECT 1054.410 232.410 1055.590 233.590 ;
        RECT 1056.010 232.410 1057.190 233.590 ;
        RECT 1057.610 232.410 1058.790 233.590 ;
        RECT 1059.210 232.410 1060.390 233.590 ;
        RECT 1060.810 232.410 1061.990 233.590 ;
        RECT 1062.410 232.410 1063.590 233.590 ;
        RECT 1064.010 232.410 1065.190 233.590 ;
        RECT 1065.610 232.410 1066.790 233.590 ;
        RECT 1067.210 232.410 1068.390 233.590 ;
        RECT 1068.810 232.410 1069.990 233.590 ;
        RECT 1070.410 232.410 1071.590 233.590 ;
        RECT 1072.010 232.410 1073.190 233.590 ;
        RECT 1073.610 232.410 1074.790 233.590 ;
        RECT 1085.210 232.410 1086.390 233.590 ;
        RECT 1086.810 232.410 1087.990 233.590 ;
        RECT 1088.410 232.410 1089.590 233.590 ;
        RECT 1090.010 232.410 1091.190 233.590 ;
        RECT 1091.610 232.410 1092.790 233.590 ;
        RECT 1093.210 232.410 1094.390 233.590 ;
        RECT 1094.810 232.410 1095.990 233.590 ;
        RECT 1096.410 232.410 1097.590 233.590 ;
        RECT 1098.010 232.410 1099.190 233.590 ;
        RECT 1099.610 232.410 1100.790 233.590 ;
        RECT 1101.210 232.410 1102.390 233.590 ;
        RECT 1102.810 232.410 1103.990 233.590 ;
        RECT 1104.410 232.410 1105.590 233.590 ;
        RECT 1106.010 232.410 1107.190 233.590 ;
        RECT 1107.610 232.410 1108.790 233.590 ;
        RECT 1109.210 232.410 1110.390 233.590 ;
        RECT 1110.810 232.410 1111.990 233.590 ;
        RECT 1112.410 232.410 1113.590 233.590 ;
        RECT 1114.010 232.410 1115.190 233.590 ;
        RECT 1115.610 232.410 1116.790 233.590 ;
        RECT 1117.210 232.410 1118.390 233.590 ;
        RECT 1118.810 232.410 1119.990 233.590 ;
        RECT 1120.410 232.410 1121.590 233.590 ;
        RECT 1122.010 232.410 1123.190 233.590 ;
        RECT 1123.610 232.410 1124.790 233.590 ;
        RECT 1135.210 232.410 1136.390 233.590 ;
        RECT 1136.810 232.410 1137.990 233.590 ;
        RECT 1138.410 232.410 1139.590 233.590 ;
        RECT 1140.010 232.410 1141.190 233.590 ;
        RECT 1141.610 232.410 1142.790 233.590 ;
        RECT 1143.210 232.410 1144.390 233.590 ;
        RECT 1144.810 232.410 1145.990 233.590 ;
        RECT 1146.410 232.410 1147.590 233.590 ;
        RECT 1148.010 232.410 1149.190 233.590 ;
        RECT 1149.610 232.410 1150.790 233.590 ;
        RECT 1151.210 232.410 1152.390 233.590 ;
        RECT 1152.810 232.410 1153.990 233.590 ;
        RECT 1154.410 232.410 1155.590 233.590 ;
        RECT 1156.010 232.410 1157.190 233.590 ;
        RECT 1157.610 232.410 1158.790 233.590 ;
        RECT 1159.210 232.410 1160.390 233.590 ;
        RECT 1160.810 232.410 1161.990 233.590 ;
        RECT 1162.410 232.410 1163.590 233.590 ;
        RECT 1164.010 232.410 1165.190 233.590 ;
        RECT 1165.610 232.410 1166.790 233.590 ;
        RECT 1167.210 232.410 1168.390 233.590 ;
        RECT 1168.810 232.410 1169.990 233.590 ;
        RECT 1170.410 232.410 1171.590 233.590 ;
        RECT 1172.010 232.410 1173.190 233.590 ;
        RECT 1173.610 232.410 1174.790 233.590 ;
        RECT 1185.210 232.410 1186.390 233.590 ;
        RECT 1186.810 232.410 1187.990 233.590 ;
        RECT 1188.410 232.410 1189.590 233.590 ;
        RECT 1190.010 232.410 1191.190 233.590 ;
        RECT 1191.610 232.410 1192.790 233.590 ;
        RECT 1193.210 232.410 1194.390 233.590 ;
        RECT 1194.810 232.410 1195.990 233.590 ;
        RECT 1196.410 232.410 1197.590 233.590 ;
        RECT 1198.010 232.410 1199.190 233.590 ;
        RECT 1199.610 232.410 1200.790 233.590 ;
        RECT 1201.210 232.410 1202.390 233.590 ;
        RECT 1202.810 232.410 1203.990 233.590 ;
        RECT 1204.410 232.410 1205.590 233.590 ;
        RECT 1206.010 232.410 1207.190 233.590 ;
        RECT 1207.610 232.410 1208.790 233.590 ;
        RECT 1209.210 232.410 1210.390 233.590 ;
        RECT 1210.810 232.410 1211.990 233.590 ;
        RECT 1212.410 232.410 1213.590 233.590 ;
        RECT 1214.010 232.410 1215.190 233.590 ;
        RECT 1215.610 232.410 1216.790 233.590 ;
        RECT 1217.210 232.410 1218.390 233.590 ;
        RECT 1218.810 232.410 1219.990 233.590 ;
        RECT 1220.410 232.410 1221.590 233.590 ;
        RECT 1222.010 232.410 1223.190 233.590 ;
        RECT 1223.610 232.410 1224.790 233.590 ;
        RECT 1235.210 232.410 1236.390 233.590 ;
        RECT 1236.810 232.410 1237.990 233.590 ;
        RECT 1238.410 232.410 1239.590 233.590 ;
        RECT 1240.010 232.410 1241.190 233.590 ;
        RECT 1241.610 232.410 1242.790 233.590 ;
        RECT 1243.210 232.410 1244.390 233.590 ;
        RECT 1244.810 232.410 1245.990 233.590 ;
        RECT 1246.410 232.410 1247.590 233.590 ;
        RECT 1248.010 232.410 1249.190 233.590 ;
        RECT 1249.610 232.410 1250.790 233.590 ;
        RECT 1251.210 232.410 1252.390 233.590 ;
        RECT 1252.810 232.410 1253.990 233.590 ;
        RECT 1254.410 232.410 1255.590 233.590 ;
        RECT 1256.010 232.410 1257.190 233.590 ;
        RECT 1257.610 232.410 1258.790 233.590 ;
        RECT 1259.210 232.410 1260.390 233.590 ;
        RECT 1260.810 232.410 1261.990 233.590 ;
        RECT 1262.410 232.410 1263.590 233.590 ;
        RECT 1264.010 232.410 1265.190 233.590 ;
        RECT 1265.610 232.410 1266.790 233.590 ;
        RECT 1267.210 232.410 1268.390 233.590 ;
        RECT 1268.810 232.410 1269.990 233.590 ;
        RECT 1270.410 232.410 1271.590 233.590 ;
        RECT 1272.010 232.410 1273.190 233.590 ;
        RECT 1273.610 232.410 1274.790 233.590 ;
        RECT 1285.210 232.410 1286.390 233.590 ;
        RECT 1286.810 232.410 1287.990 233.590 ;
        RECT 1288.410 232.410 1289.590 233.590 ;
        RECT 1290.010 232.410 1291.190 233.590 ;
        RECT 1291.610 232.410 1292.790 233.590 ;
        RECT 1293.210 232.410 1294.390 233.590 ;
        RECT 1294.810 232.410 1295.990 233.590 ;
        RECT 1296.410 232.410 1297.590 233.590 ;
        RECT 1298.010 232.410 1299.190 233.590 ;
        RECT 1299.610 232.410 1300.790 233.590 ;
        RECT 1301.210 232.410 1302.390 233.590 ;
        RECT 1302.810 232.410 1303.990 233.590 ;
        RECT 1304.410 232.410 1305.590 233.590 ;
        RECT 1306.010 232.410 1307.190 233.590 ;
        RECT 1307.610 232.410 1308.790 233.590 ;
        RECT 1309.210 232.410 1310.390 233.590 ;
        RECT 1310.810 232.410 1311.990 233.590 ;
        RECT 1312.410 232.410 1313.590 233.590 ;
        RECT 1314.010 232.410 1315.190 233.590 ;
        RECT 1315.610 232.410 1316.790 233.590 ;
        RECT 1317.210 232.410 1318.390 233.590 ;
        RECT 1318.810 232.410 1319.990 233.590 ;
        RECT 1320.410 232.410 1321.590 233.590 ;
        RECT 1322.010 232.410 1323.190 233.590 ;
        RECT 1323.610 232.410 1324.790 233.590 ;
        RECT 1335.210 232.410 1336.390 233.590 ;
        RECT 1336.810 232.410 1337.990 233.590 ;
        RECT 1338.410 232.410 1339.590 233.590 ;
        RECT 1340.010 232.410 1341.190 233.590 ;
        RECT 1341.610 232.410 1342.790 233.590 ;
        RECT 1343.210 232.410 1344.390 233.590 ;
        RECT 1344.810 232.410 1345.990 233.590 ;
        RECT 1346.410 232.410 1347.590 233.590 ;
        RECT 1348.010 232.410 1349.190 233.590 ;
        RECT 1349.610 232.410 1350.790 233.590 ;
        RECT 1351.210 232.410 1352.390 233.590 ;
        RECT 1352.810 232.410 1353.990 233.590 ;
        RECT 1354.410 232.410 1355.590 233.590 ;
        RECT 1356.010 232.410 1357.190 233.590 ;
        RECT 1357.610 232.410 1358.790 233.590 ;
        RECT 1359.210 232.410 1360.390 233.590 ;
        RECT 1360.810 232.410 1361.990 233.590 ;
        RECT 1362.410 232.410 1363.590 233.590 ;
        RECT 1364.010 232.410 1365.190 233.590 ;
        RECT 1365.610 232.410 1366.790 233.590 ;
        RECT 1367.210 232.410 1368.390 233.590 ;
        RECT 1368.810 232.410 1369.990 233.590 ;
        RECT 1370.410 232.410 1371.590 233.590 ;
        RECT 1372.010 232.410 1373.190 233.590 ;
        RECT 1373.610 232.410 1374.790 233.590 ;
        RECT 1385.210 232.410 1386.390 233.590 ;
        RECT 1386.810 232.410 1387.990 233.590 ;
        RECT 1388.410 232.410 1389.590 233.590 ;
        RECT 1390.010 232.410 1391.190 233.590 ;
        RECT 1391.610 232.410 1392.790 233.590 ;
        RECT 1393.210 232.410 1394.390 233.590 ;
        RECT 1394.810 232.410 1395.990 233.590 ;
        RECT 1396.410 232.410 1397.590 233.590 ;
        RECT 1398.010 232.410 1399.190 233.590 ;
        RECT 1399.610 232.410 1400.790 233.590 ;
        RECT 1401.210 232.410 1402.390 233.590 ;
        RECT 1402.810 232.410 1403.990 233.590 ;
        RECT 1404.410 232.410 1405.590 233.590 ;
        RECT 1406.010 232.410 1407.190 233.590 ;
        RECT 1407.610 232.410 1408.790 233.590 ;
        RECT 1409.210 232.410 1410.390 233.590 ;
        RECT 1410.810 232.410 1411.990 233.590 ;
        RECT 1412.410 232.410 1413.590 233.590 ;
        RECT 1414.010 232.410 1415.190 233.590 ;
        RECT 1415.610 232.410 1416.790 233.590 ;
        RECT 1417.210 232.410 1418.390 233.590 ;
        RECT 1418.810 232.410 1419.990 233.590 ;
        RECT 1420.410 232.410 1421.590 233.590 ;
        RECT 1422.010 232.410 1423.190 233.590 ;
        RECT 1423.610 232.410 1424.790 233.590 ;
        RECT 220.310 129.110 224.690 131.890 ;
        RECT 220.310 28.110 224.690 30.890 ;
        RECT 235.210 26.410 236.390 27.590 ;
        RECT 236.810 26.410 237.990 27.590 ;
        RECT 238.410 26.410 239.590 27.590 ;
        RECT 240.010 26.410 241.190 27.590 ;
        RECT 241.610 26.410 242.790 27.590 ;
        RECT 243.210 26.410 244.390 27.590 ;
        RECT 244.810 26.410 245.990 27.590 ;
        RECT 246.410 26.410 247.590 27.590 ;
        RECT 248.010 26.410 249.190 27.590 ;
        RECT 249.610 26.410 250.790 27.590 ;
        RECT 251.210 26.410 252.390 27.590 ;
        RECT 252.810 26.410 253.990 27.590 ;
        RECT 254.410 26.410 255.590 27.590 ;
        RECT 256.010 26.410 257.190 27.590 ;
        RECT 257.610 26.410 258.790 27.590 ;
        RECT 259.210 26.410 260.390 27.590 ;
        RECT 260.810 26.410 261.990 27.590 ;
        RECT 262.410 26.410 263.590 27.590 ;
        RECT 264.010 26.410 265.190 27.590 ;
        RECT 265.610 26.410 266.790 27.590 ;
        RECT 267.210 26.410 268.390 27.590 ;
        RECT 268.810 26.410 269.990 27.590 ;
        RECT 270.410 26.410 271.590 27.590 ;
        RECT 272.010 26.410 273.190 27.590 ;
        RECT 273.610 26.410 274.790 27.590 ;
        RECT 285.210 26.410 286.390 27.590 ;
        RECT 286.810 26.410 287.990 27.590 ;
        RECT 288.410 26.410 289.590 27.590 ;
        RECT 290.010 26.410 291.190 27.590 ;
        RECT 291.610 26.410 292.790 27.590 ;
        RECT 293.210 26.410 294.390 27.590 ;
        RECT 294.810 26.410 295.990 27.590 ;
        RECT 296.410 26.410 297.590 27.590 ;
        RECT 298.010 26.410 299.190 27.590 ;
        RECT 299.610 26.410 300.790 27.590 ;
        RECT 301.210 26.410 302.390 27.590 ;
        RECT 302.810 26.410 303.990 27.590 ;
        RECT 304.410 26.410 305.590 27.590 ;
        RECT 306.010 26.410 307.190 27.590 ;
        RECT 307.610 26.410 308.790 27.590 ;
        RECT 309.210 26.410 310.390 27.590 ;
        RECT 310.810 26.410 311.990 27.590 ;
        RECT 312.410 26.410 313.590 27.590 ;
        RECT 314.010 26.410 315.190 27.590 ;
        RECT 315.610 26.410 316.790 27.590 ;
        RECT 317.210 26.410 318.390 27.590 ;
        RECT 318.810 26.410 319.990 27.590 ;
        RECT 320.410 26.410 321.590 27.590 ;
        RECT 322.010 26.410 323.190 27.590 ;
        RECT 323.610 26.410 324.790 27.590 ;
        RECT 335.210 26.410 336.390 27.590 ;
        RECT 336.810 26.410 337.990 27.590 ;
        RECT 338.410 26.410 339.590 27.590 ;
        RECT 340.010 26.410 341.190 27.590 ;
        RECT 341.610 26.410 342.790 27.590 ;
        RECT 343.210 26.410 344.390 27.590 ;
        RECT 344.810 26.410 345.990 27.590 ;
        RECT 346.410 26.410 347.590 27.590 ;
        RECT 348.010 26.410 349.190 27.590 ;
        RECT 349.610 26.410 350.790 27.590 ;
        RECT 351.210 26.410 352.390 27.590 ;
        RECT 352.810 26.410 353.990 27.590 ;
        RECT 354.410 26.410 355.590 27.590 ;
        RECT 356.010 26.410 357.190 27.590 ;
        RECT 357.610 26.410 358.790 27.590 ;
        RECT 359.210 26.410 360.390 27.590 ;
        RECT 360.810 26.410 361.990 27.590 ;
        RECT 362.410 26.410 363.590 27.590 ;
        RECT 364.010 26.410 365.190 27.590 ;
        RECT 365.610 26.410 366.790 27.590 ;
        RECT 367.210 26.410 368.390 27.590 ;
        RECT 368.810 26.410 369.990 27.590 ;
        RECT 370.410 26.410 371.590 27.590 ;
        RECT 372.010 26.410 373.190 27.590 ;
        RECT 373.610 26.410 374.790 27.590 ;
        RECT 385.210 26.410 386.390 27.590 ;
        RECT 386.810 26.410 387.990 27.590 ;
        RECT 388.410 26.410 389.590 27.590 ;
        RECT 390.010 26.410 391.190 27.590 ;
        RECT 391.610 26.410 392.790 27.590 ;
        RECT 393.210 26.410 394.390 27.590 ;
        RECT 394.810 26.410 395.990 27.590 ;
        RECT 396.410 26.410 397.590 27.590 ;
        RECT 398.010 26.410 399.190 27.590 ;
        RECT 399.610 26.410 400.790 27.590 ;
        RECT 401.210 26.410 402.390 27.590 ;
        RECT 402.810 26.410 403.990 27.590 ;
        RECT 404.410 26.410 405.590 27.590 ;
        RECT 406.010 26.410 407.190 27.590 ;
        RECT 407.610 26.410 408.790 27.590 ;
        RECT 409.210 26.410 410.390 27.590 ;
        RECT 410.810 26.410 411.990 27.590 ;
        RECT 412.410 26.410 413.590 27.590 ;
        RECT 414.010 26.410 415.190 27.590 ;
        RECT 415.610 26.410 416.790 27.590 ;
        RECT 417.210 26.410 418.390 27.590 ;
        RECT 418.810 26.410 419.990 27.590 ;
        RECT 420.410 26.410 421.590 27.590 ;
        RECT 422.010 26.410 423.190 27.590 ;
        RECT 423.610 26.410 424.790 27.590 ;
        RECT 435.210 26.410 436.390 27.590 ;
        RECT 436.810 26.410 437.990 27.590 ;
        RECT 438.410 26.410 439.590 27.590 ;
        RECT 440.010 26.410 441.190 27.590 ;
        RECT 441.610 26.410 442.790 27.590 ;
        RECT 443.210 26.410 444.390 27.590 ;
        RECT 444.810 26.410 445.990 27.590 ;
        RECT 446.410 26.410 447.590 27.590 ;
        RECT 448.010 26.410 449.190 27.590 ;
        RECT 449.610 26.410 450.790 27.590 ;
        RECT 451.210 26.410 452.390 27.590 ;
        RECT 452.810 26.410 453.990 27.590 ;
        RECT 454.410 26.410 455.590 27.590 ;
        RECT 456.010 26.410 457.190 27.590 ;
        RECT 457.610 26.410 458.790 27.590 ;
        RECT 459.210 26.410 460.390 27.590 ;
        RECT 460.810 26.410 461.990 27.590 ;
        RECT 462.410 26.410 463.590 27.590 ;
        RECT 464.010 26.410 465.190 27.590 ;
        RECT 465.610 26.410 466.790 27.590 ;
        RECT 467.210 26.410 468.390 27.590 ;
        RECT 468.810 26.410 469.990 27.590 ;
        RECT 470.410 26.410 471.590 27.590 ;
        RECT 472.010 26.410 473.190 27.590 ;
        RECT 473.610 26.410 474.790 27.590 ;
        RECT 485.210 26.410 486.390 27.590 ;
        RECT 486.810 26.410 487.990 27.590 ;
        RECT 488.410 26.410 489.590 27.590 ;
        RECT 490.010 26.410 491.190 27.590 ;
        RECT 491.610 26.410 492.790 27.590 ;
        RECT 493.210 26.410 494.390 27.590 ;
        RECT 494.810 26.410 495.990 27.590 ;
        RECT 496.410 26.410 497.590 27.590 ;
        RECT 498.010 26.410 499.190 27.590 ;
        RECT 499.610 26.410 500.790 27.590 ;
        RECT 501.210 26.410 502.390 27.590 ;
        RECT 502.810 26.410 503.990 27.590 ;
        RECT 504.410 26.410 505.590 27.590 ;
        RECT 506.010 26.410 507.190 27.590 ;
        RECT 507.610 26.410 508.790 27.590 ;
        RECT 509.210 26.410 510.390 27.590 ;
        RECT 510.810 26.410 511.990 27.590 ;
        RECT 512.410 26.410 513.590 27.590 ;
        RECT 514.010 26.410 515.190 27.590 ;
        RECT 515.610 26.410 516.790 27.590 ;
        RECT 517.210 26.410 518.390 27.590 ;
        RECT 518.810 26.410 519.990 27.590 ;
        RECT 520.410 26.410 521.590 27.590 ;
        RECT 522.010 26.410 523.190 27.590 ;
        RECT 523.610 26.410 524.790 27.590 ;
        RECT 535.210 26.410 536.390 27.590 ;
        RECT 536.810 26.410 537.990 27.590 ;
        RECT 538.410 26.410 539.590 27.590 ;
        RECT 540.010 26.410 541.190 27.590 ;
        RECT 541.610 26.410 542.790 27.590 ;
        RECT 543.210 26.410 544.390 27.590 ;
        RECT 544.810 26.410 545.990 27.590 ;
        RECT 546.410 26.410 547.590 27.590 ;
        RECT 548.010 26.410 549.190 27.590 ;
        RECT 549.610 26.410 550.790 27.590 ;
        RECT 551.210 26.410 552.390 27.590 ;
        RECT 552.810 26.410 553.990 27.590 ;
        RECT 554.410 26.410 555.590 27.590 ;
        RECT 556.010 26.410 557.190 27.590 ;
        RECT 557.610 26.410 558.790 27.590 ;
        RECT 559.210 26.410 560.390 27.590 ;
        RECT 560.810 26.410 561.990 27.590 ;
        RECT 562.410 26.410 563.590 27.590 ;
        RECT 564.010 26.410 565.190 27.590 ;
        RECT 565.610 26.410 566.790 27.590 ;
        RECT 567.210 26.410 568.390 27.590 ;
        RECT 568.810 26.410 569.990 27.590 ;
        RECT 570.410 26.410 571.590 27.590 ;
        RECT 572.010 26.410 573.190 27.590 ;
        RECT 573.610 26.410 574.790 27.590 ;
        RECT 585.210 26.410 586.390 27.590 ;
        RECT 586.810 26.410 587.990 27.590 ;
        RECT 588.410 26.410 589.590 27.590 ;
        RECT 590.010 26.410 591.190 27.590 ;
        RECT 591.610 26.410 592.790 27.590 ;
        RECT 593.210 26.410 594.390 27.590 ;
        RECT 594.810 26.410 595.990 27.590 ;
        RECT 596.410 26.410 597.590 27.590 ;
        RECT 598.010 26.410 599.190 27.590 ;
        RECT 599.610 26.410 600.790 27.590 ;
        RECT 601.210 26.410 602.390 27.590 ;
        RECT 602.810 26.410 603.990 27.590 ;
        RECT 604.410 26.410 605.590 27.590 ;
        RECT 606.010 26.410 607.190 27.590 ;
        RECT 607.610 26.410 608.790 27.590 ;
        RECT 609.210 26.410 610.390 27.590 ;
        RECT 610.810 26.410 611.990 27.590 ;
        RECT 612.410 26.410 613.590 27.590 ;
        RECT 614.010 26.410 615.190 27.590 ;
        RECT 615.610 26.410 616.790 27.590 ;
        RECT 617.210 26.410 618.390 27.590 ;
        RECT 618.810 26.410 619.990 27.590 ;
        RECT 620.410 26.410 621.590 27.590 ;
        RECT 622.010 26.410 623.190 27.590 ;
        RECT 623.610 26.410 624.790 27.590 ;
        RECT 635.210 26.410 636.390 27.590 ;
        RECT 636.810 26.410 637.990 27.590 ;
        RECT 638.410 26.410 639.590 27.590 ;
        RECT 640.010 26.410 641.190 27.590 ;
        RECT 641.610 26.410 642.790 27.590 ;
        RECT 643.210 26.410 644.390 27.590 ;
        RECT 644.810 26.410 645.990 27.590 ;
        RECT 646.410 26.410 647.590 27.590 ;
        RECT 648.010 26.410 649.190 27.590 ;
        RECT 649.610 26.410 650.790 27.590 ;
        RECT 651.210 26.410 652.390 27.590 ;
        RECT 652.810 26.410 653.990 27.590 ;
        RECT 654.410 26.410 655.590 27.590 ;
        RECT 656.010 26.410 657.190 27.590 ;
        RECT 657.610 26.410 658.790 27.590 ;
        RECT 659.210 26.410 660.390 27.590 ;
        RECT 660.810 26.410 661.990 27.590 ;
        RECT 662.410 26.410 663.590 27.590 ;
        RECT 664.010 26.410 665.190 27.590 ;
        RECT 665.610 26.410 666.790 27.590 ;
        RECT 667.210 26.410 668.390 27.590 ;
        RECT 668.810 26.410 669.990 27.590 ;
        RECT 670.410 26.410 671.590 27.590 ;
        RECT 672.010 26.410 673.190 27.590 ;
        RECT 673.610 26.410 674.790 27.590 ;
        RECT 685.210 26.410 686.390 27.590 ;
        RECT 686.810 26.410 687.990 27.590 ;
        RECT 688.410 26.410 689.590 27.590 ;
        RECT 690.010 26.410 691.190 27.590 ;
        RECT 691.610 26.410 692.790 27.590 ;
        RECT 693.210 26.410 694.390 27.590 ;
        RECT 694.810 26.410 695.990 27.590 ;
        RECT 696.410 26.410 697.590 27.590 ;
        RECT 698.010 26.410 699.190 27.590 ;
        RECT 699.610 26.410 700.790 27.590 ;
        RECT 701.210 26.410 702.390 27.590 ;
        RECT 702.810 26.410 703.990 27.590 ;
        RECT 704.410 26.410 705.590 27.590 ;
        RECT 706.010 26.410 707.190 27.590 ;
        RECT 707.610 26.410 708.790 27.590 ;
        RECT 709.210 26.410 710.390 27.590 ;
        RECT 710.810 26.410 711.990 27.590 ;
        RECT 712.410 26.410 713.590 27.590 ;
        RECT 714.010 26.410 715.190 27.590 ;
        RECT 715.610 26.410 716.790 27.590 ;
        RECT 717.210 26.410 718.390 27.590 ;
        RECT 718.810 26.410 719.990 27.590 ;
        RECT 720.410 26.410 721.590 27.590 ;
        RECT 722.010 26.410 723.190 27.590 ;
        RECT 723.610 26.410 724.790 27.590 ;
        RECT 735.210 26.410 736.390 27.590 ;
        RECT 736.810 26.410 737.990 27.590 ;
        RECT 738.410 26.410 739.590 27.590 ;
        RECT 740.010 26.410 741.190 27.590 ;
        RECT 741.610 26.410 742.790 27.590 ;
        RECT 743.210 26.410 744.390 27.590 ;
        RECT 744.810 26.410 745.990 27.590 ;
        RECT 746.410 26.410 747.590 27.590 ;
        RECT 748.010 26.410 749.190 27.590 ;
        RECT 749.610 26.410 750.790 27.590 ;
        RECT 751.210 26.410 752.390 27.590 ;
        RECT 752.810 26.410 753.990 27.590 ;
        RECT 754.410 26.410 755.590 27.590 ;
        RECT 756.010 26.410 757.190 27.590 ;
        RECT 757.610 26.410 758.790 27.590 ;
        RECT 759.210 26.410 760.390 27.590 ;
        RECT 760.810 26.410 761.990 27.590 ;
        RECT 762.410 26.410 763.590 27.590 ;
        RECT 764.010 26.410 765.190 27.590 ;
        RECT 765.610 26.410 766.790 27.590 ;
        RECT 767.210 26.410 768.390 27.590 ;
        RECT 768.810 26.410 769.990 27.590 ;
        RECT 770.410 26.410 771.590 27.590 ;
        RECT 772.010 26.410 773.190 27.590 ;
        RECT 773.610 26.410 774.790 27.590 ;
        RECT 785.210 26.410 786.390 27.590 ;
        RECT 786.810 26.410 787.990 27.590 ;
        RECT 788.410 26.410 789.590 27.590 ;
        RECT 790.010 26.410 791.190 27.590 ;
        RECT 791.610 26.410 792.790 27.590 ;
        RECT 793.210 26.410 794.390 27.590 ;
        RECT 794.810 26.410 795.990 27.590 ;
        RECT 796.410 26.410 797.590 27.590 ;
        RECT 798.010 26.410 799.190 27.590 ;
        RECT 799.610 26.410 800.790 27.590 ;
        RECT 801.210 26.410 802.390 27.590 ;
        RECT 802.810 26.410 803.990 27.590 ;
        RECT 804.410 26.410 805.590 27.590 ;
        RECT 806.010 26.410 807.190 27.590 ;
        RECT 807.610 26.410 808.790 27.590 ;
        RECT 809.210 26.410 810.390 27.590 ;
        RECT 810.810 26.410 811.990 27.590 ;
        RECT 812.410 26.410 813.590 27.590 ;
        RECT 814.010 26.410 815.190 27.590 ;
        RECT 815.610 26.410 816.790 27.590 ;
        RECT 817.210 26.410 818.390 27.590 ;
        RECT 818.810 26.410 819.990 27.590 ;
        RECT 820.410 26.410 821.590 27.590 ;
        RECT 822.010 26.410 823.190 27.590 ;
        RECT 823.610 26.410 824.790 27.590 ;
        RECT 835.210 26.410 836.390 27.590 ;
        RECT 836.810 26.410 837.990 27.590 ;
        RECT 838.410 26.410 839.590 27.590 ;
        RECT 840.010 26.410 841.190 27.590 ;
        RECT 841.610 26.410 842.790 27.590 ;
        RECT 843.210 26.410 844.390 27.590 ;
        RECT 844.810 26.410 845.990 27.590 ;
        RECT 846.410 26.410 847.590 27.590 ;
        RECT 848.010 26.410 849.190 27.590 ;
        RECT 849.610 26.410 850.790 27.590 ;
        RECT 851.210 26.410 852.390 27.590 ;
        RECT 852.810 26.410 853.990 27.590 ;
        RECT 854.410 26.410 855.590 27.590 ;
        RECT 856.010 26.410 857.190 27.590 ;
        RECT 857.610 26.410 858.790 27.590 ;
        RECT 859.210 26.410 860.390 27.590 ;
        RECT 860.810 26.410 861.990 27.590 ;
        RECT 862.410 26.410 863.590 27.590 ;
        RECT 864.010 26.410 865.190 27.590 ;
        RECT 865.610 26.410 866.790 27.590 ;
        RECT 867.210 26.410 868.390 27.590 ;
        RECT 868.810 26.410 869.990 27.590 ;
        RECT 870.410 26.410 871.590 27.590 ;
        RECT 872.010 26.410 873.190 27.590 ;
        RECT 873.610 26.410 874.790 27.590 ;
        RECT 885.210 26.410 886.390 27.590 ;
        RECT 886.810 26.410 887.990 27.590 ;
        RECT 888.410 26.410 889.590 27.590 ;
        RECT 890.010 26.410 891.190 27.590 ;
        RECT 891.610 26.410 892.790 27.590 ;
        RECT 893.210 26.410 894.390 27.590 ;
        RECT 894.810 26.410 895.990 27.590 ;
        RECT 896.410 26.410 897.590 27.590 ;
        RECT 898.010 26.410 899.190 27.590 ;
        RECT 899.610 26.410 900.790 27.590 ;
        RECT 901.210 26.410 902.390 27.590 ;
        RECT 902.810 26.410 903.990 27.590 ;
        RECT 904.410 26.410 905.590 27.590 ;
        RECT 906.010 26.410 907.190 27.590 ;
        RECT 907.610 26.410 908.790 27.590 ;
        RECT 909.210 26.410 910.390 27.590 ;
        RECT 910.810 26.410 911.990 27.590 ;
        RECT 912.410 26.410 913.590 27.590 ;
        RECT 914.010 26.410 915.190 27.590 ;
        RECT 915.610 26.410 916.790 27.590 ;
        RECT 917.210 26.410 918.390 27.590 ;
        RECT 918.810 26.410 919.990 27.590 ;
        RECT 920.410 26.410 921.590 27.590 ;
        RECT 922.010 26.410 923.190 27.590 ;
        RECT 923.610 26.410 924.790 27.590 ;
        RECT 935.210 26.410 936.390 27.590 ;
        RECT 936.810 26.410 937.990 27.590 ;
        RECT 938.410 26.410 939.590 27.590 ;
        RECT 940.010 26.410 941.190 27.590 ;
        RECT 941.610 26.410 942.790 27.590 ;
        RECT 943.210 26.410 944.390 27.590 ;
        RECT 944.810 26.410 945.990 27.590 ;
        RECT 946.410 26.410 947.590 27.590 ;
        RECT 948.010 26.410 949.190 27.590 ;
        RECT 949.610 26.410 950.790 27.590 ;
        RECT 951.210 26.410 952.390 27.590 ;
        RECT 952.810 26.410 953.990 27.590 ;
        RECT 954.410 26.410 955.590 27.590 ;
        RECT 956.010 26.410 957.190 27.590 ;
        RECT 957.610 26.410 958.790 27.590 ;
        RECT 959.210 26.410 960.390 27.590 ;
        RECT 960.810 26.410 961.990 27.590 ;
        RECT 962.410 26.410 963.590 27.590 ;
        RECT 964.010 26.410 965.190 27.590 ;
        RECT 965.610 26.410 966.790 27.590 ;
        RECT 967.210 26.410 968.390 27.590 ;
        RECT 968.810 26.410 969.990 27.590 ;
        RECT 970.410 26.410 971.590 27.590 ;
        RECT 972.010 26.410 973.190 27.590 ;
        RECT 973.610 26.410 974.790 27.590 ;
        RECT 985.210 26.410 986.390 27.590 ;
        RECT 986.810 26.410 987.990 27.590 ;
        RECT 988.410 26.410 989.590 27.590 ;
        RECT 990.010 26.410 991.190 27.590 ;
        RECT 991.610 26.410 992.790 27.590 ;
        RECT 993.210 26.410 994.390 27.590 ;
        RECT 994.810 26.410 995.990 27.590 ;
        RECT 996.410 26.410 997.590 27.590 ;
        RECT 998.010 26.410 999.190 27.590 ;
        RECT 999.610 26.410 1000.790 27.590 ;
        RECT 1001.210 26.410 1002.390 27.590 ;
        RECT 1002.810 26.410 1003.990 27.590 ;
        RECT 1004.410 26.410 1005.590 27.590 ;
        RECT 1006.010 26.410 1007.190 27.590 ;
        RECT 1007.610 26.410 1008.790 27.590 ;
        RECT 1009.210 26.410 1010.390 27.590 ;
        RECT 1010.810 26.410 1011.990 27.590 ;
        RECT 1012.410 26.410 1013.590 27.590 ;
        RECT 1014.010 26.410 1015.190 27.590 ;
        RECT 1015.610 26.410 1016.790 27.590 ;
        RECT 1017.210 26.410 1018.390 27.590 ;
        RECT 1018.810 26.410 1019.990 27.590 ;
        RECT 1020.410 26.410 1021.590 27.590 ;
        RECT 1022.010 26.410 1023.190 27.590 ;
        RECT 1023.610 26.410 1024.790 27.590 ;
        RECT 1035.210 26.410 1036.390 27.590 ;
        RECT 1036.810 26.410 1037.990 27.590 ;
        RECT 1038.410 26.410 1039.590 27.590 ;
        RECT 1040.010 26.410 1041.190 27.590 ;
        RECT 1041.610 26.410 1042.790 27.590 ;
        RECT 1043.210 26.410 1044.390 27.590 ;
        RECT 1044.810 26.410 1045.990 27.590 ;
        RECT 1046.410 26.410 1047.590 27.590 ;
        RECT 1048.010 26.410 1049.190 27.590 ;
        RECT 1049.610 26.410 1050.790 27.590 ;
        RECT 1051.210 26.410 1052.390 27.590 ;
        RECT 1052.810 26.410 1053.990 27.590 ;
        RECT 1054.410 26.410 1055.590 27.590 ;
        RECT 1056.010 26.410 1057.190 27.590 ;
        RECT 1057.610 26.410 1058.790 27.590 ;
        RECT 1059.210 26.410 1060.390 27.590 ;
        RECT 1060.810 26.410 1061.990 27.590 ;
        RECT 1062.410 26.410 1063.590 27.590 ;
        RECT 1064.010 26.410 1065.190 27.590 ;
        RECT 1065.610 26.410 1066.790 27.590 ;
        RECT 1067.210 26.410 1068.390 27.590 ;
        RECT 1068.810 26.410 1069.990 27.590 ;
        RECT 1070.410 26.410 1071.590 27.590 ;
        RECT 1072.010 26.410 1073.190 27.590 ;
        RECT 1073.610 26.410 1074.790 27.590 ;
        RECT 1085.210 26.410 1086.390 27.590 ;
        RECT 1086.810 26.410 1087.990 27.590 ;
        RECT 1088.410 26.410 1089.590 27.590 ;
        RECT 1090.010 26.410 1091.190 27.590 ;
        RECT 1091.610 26.410 1092.790 27.590 ;
        RECT 1093.210 26.410 1094.390 27.590 ;
        RECT 1094.810 26.410 1095.990 27.590 ;
        RECT 1096.410 26.410 1097.590 27.590 ;
        RECT 1098.010 26.410 1099.190 27.590 ;
        RECT 1099.610 26.410 1100.790 27.590 ;
        RECT 1101.210 26.410 1102.390 27.590 ;
        RECT 1102.810 26.410 1103.990 27.590 ;
        RECT 1104.410 26.410 1105.590 27.590 ;
        RECT 1106.010 26.410 1107.190 27.590 ;
        RECT 1107.610 26.410 1108.790 27.590 ;
        RECT 1109.210 26.410 1110.390 27.590 ;
        RECT 1110.810 26.410 1111.990 27.590 ;
        RECT 1112.410 26.410 1113.590 27.590 ;
        RECT 1114.010 26.410 1115.190 27.590 ;
        RECT 1115.610 26.410 1116.790 27.590 ;
        RECT 1117.210 26.410 1118.390 27.590 ;
        RECT 1118.810 26.410 1119.990 27.590 ;
        RECT 1120.410 26.410 1121.590 27.590 ;
        RECT 1122.010 26.410 1123.190 27.590 ;
        RECT 1123.610 26.410 1124.790 27.590 ;
        RECT 1135.210 26.410 1136.390 27.590 ;
        RECT 1136.810 26.410 1137.990 27.590 ;
        RECT 1138.410 26.410 1139.590 27.590 ;
        RECT 1140.010 26.410 1141.190 27.590 ;
        RECT 1141.610 26.410 1142.790 27.590 ;
        RECT 1143.210 26.410 1144.390 27.590 ;
        RECT 1144.810 26.410 1145.990 27.590 ;
        RECT 1146.410 26.410 1147.590 27.590 ;
        RECT 1148.010 26.410 1149.190 27.590 ;
        RECT 1149.610 26.410 1150.790 27.590 ;
        RECT 1151.210 26.410 1152.390 27.590 ;
        RECT 1152.810 26.410 1153.990 27.590 ;
        RECT 1154.410 26.410 1155.590 27.590 ;
        RECT 1156.010 26.410 1157.190 27.590 ;
        RECT 1157.610 26.410 1158.790 27.590 ;
        RECT 1159.210 26.410 1160.390 27.590 ;
        RECT 1160.810 26.410 1161.990 27.590 ;
        RECT 1162.410 26.410 1163.590 27.590 ;
        RECT 1164.010 26.410 1165.190 27.590 ;
        RECT 1165.610 26.410 1166.790 27.590 ;
        RECT 1167.210 26.410 1168.390 27.590 ;
        RECT 1168.810 26.410 1169.990 27.590 ;
        RECT 1170.410 26.410 1171.590 27.590 ;
        RECT 1172.010 26.410 1173.190 27.590 ;
        RECT 1173.610 26.410 1174.790 27.590 ;
        RECT 1185.210 26.410 1186.390 27.590 ;
        RECT 1186.810 26.410 1187.990 27.590 ;
        RECT 1188.410 26.410 1189.590 27.590 ;
        RECT 1190.010 26.410 1191.190 27.590 ;
        RECT 1191.610 26.410 1192.790 27.590 ;
        RECT 1193.210 26.410 1194.390 27.590 ;
        RECT 1194.810 26.410 1195.990 27.590 ;
        RECT 1196.410 26.410 1197.590 27.590 ;
        RECT 1198.010 26.410 1199.190 27.590 ;
        RECT 1199.610 26.410 1200.790 27.590 ;
        RECT 1201.210 26.410 1202.390 27.590 ;
        RECT 1202.810 26.410 1203.990 27.590 ;
        RECT 1204.410 26.410 1205.590 27.590 ;
        RECT 1206.010 26.410 1207.190 27.590 ;
        RECT 1207.610 26.410 1208.790 27.590 ;
        RECT 1209.210 26.410 1210.390 27.590 ;
        RECT 1210.810 26.410 1211.990 27.590 ;
        RECT 1212.410 26.410 1213.590 27.590 ;
        RECT 1214.010 26.410 1215.190 27.590 ;
        RECT 1215.610 26.410 1216.790 27.590 ;
        RECT 1217.210 26.410 1218.390 27.590 ;
        RECT 1218.810 26.410 1219.990 27.590 ;
        RECT 1220.410 26.410 1221.590 27.590 ;
        RECT 1222.010 26.410 1223.190 27.590 ;
        RECT 1223.610 26.410 1224.790 27.590 ;
        RECT 1235.210 26.410 1236.390 27.590 ;
        RECT 1236.810 26.410 1237.990 27.590 ;
        RECT 1238.410 26.410 1239.590 27.590 ;
        RECT 1240.010 26.410 1241.190 27.590 ;
        RECT 1241.610 26.410 1242.790 27.590 ;
        RECT 1243.210 26.410 1244.390 27.590 ;
        RECT 1244.810 26.410 1245.990 27.590 ;
        RECT 1246.410 26.410 1247.590 27.590 ;
        RECT 1248.010 26.410 1249.190 27.590 ;
        RECT 1249.610 26.410 1250.790 27.590 ;
        RECT 1251.210 26.410 1252.390 27.590 ;
        RECT 1252.810 26.410 1253.990 27.590 ;
        RECT 1254.410 26.410 1255.590 27.590 ;
        RECT 1256.010 26.410 1257.190 27.590 ;
        RECT 1257.610 26.410 1258.790 27.590 ;
        RECT 1259.210 26.410 1260.390 27.590 ;
        RECT 1260.810 26.410 1261.990 27.590 ;
        RECT 1262.410 26.410 1263.590 27.590 ;
        RECT 1264.010 26.410 1265.190 27.590 ;
        RECT 1265.610 26.410 1266.790 27.590 ;
        RECT 1267.210 26.410 1268.390 27.590 ;
        RECT 1268.810 26.410 1269.990 27.590 ;
        RECT 1270.410 26.410 1271.590 27.590 ;
        RECT 1272.010 26.410 1273.190 27.590 ;
        RECT 1273.610 26.410 1274.790 27.590 ;
        RECT 1285.210 26.410 1286.390 27.590 ;
        RECT 1286.810 26.410 1287.990 27.590 ;
        RECT 1288.410 26.410 1289.590 27.590 ;
        RECT 1290.010 26.410 1291.190 27.590 ;
        RECT 1291.610 26.410 1292.790 27.590 ;
        RECT 1293.210 26.410 1294.390 27.590 ;
        RECT 1294.810 26.410 1295.990 27.590 ;
        RECT 1296.410 26.410 1297.590 27.590 ;
        RECT 1298.010 26.410 1299.190 27.590 ;
        RECT 1299.610 26.410 1300.790 27.590 ;
        RECT 1301.210 26.410 1302.390 27.590 ;
        RECT 1302.810 26.410 1303.990 27.590 ;
        RECT 1304.410 26.410 1305.590 27.590 ;
        RECT 1306.010 26.410 1307.190 27.590 ;
        RECT 1307.610 26.410 1308.790 27.590 ;
        RECT 1309.210 26.410 1310.390 27.590 ;
        RECT 1310.810 26.410 1311.990 27.590 ;
        RECT 1312.410 26.410 1313.590 27.590 ;
        RECT 1314.010 26.410 1315.190 27.590 ;
        RECT 1315.610 26.410 1316.790 27.590 ;
        RECT 1317.210 26.410 1318.390 27.590 ;
        RECT 1318.810 26.410 1319.990 27.590 ;
        RECT 1320.410 26.410 1321.590 27.590 ;
        RECT 1322.010 26.410 1323.190 27.590 ;
        RECT 1323.610 26.410 1324.790 27.590 ;
        RECT 1335.210 26.410 1336.390 27.590 ;
        RECT 1336.810 26.410 1337.990 27.590 ;
        RECT 1338.410 26.410 1339.590 27.590 ;
        RECT 1340.010 26.410 1341.190 27.590 ;
        RECT 1341.610 26.410 1342.790 27.590 ;
        RECT 1343.210 26.410 1344.390 27.590 ;
        RECT 1344.810 26.410 1345.990 27.590 ;
        RECT 1346.410 26.410 1347.590 27.590 ;
        RECT 1348.010 26.410 1349.190 27.590 ;
        RECT 1349.610 26.410 1350.790 27.590 ;
        RECT 1351.210 26.410 1352.390 27.590 ;
        RECT 1352.810 26.410 1353.990 27.590 ;
        RECT 1354.410 26.410 1355.590 27.590 ;
        RECT 1356.010 26.410 1357.190 27.590 ;
        RECT 1357.610 26.410 1358.790 27.590 ;
        RECT 1359.210 26.410 1360.390 27.590 ;
        RECT 1360.810 26.410 1361.990 27.590 ;
        RECT 1362.410 26.410 1363.590 27.590 ;
        RECT 1364.010 26.410 1365.190 27.590 ;
        RECT 1365.610 26.410 1366.790 27.590 ;
        RECT 1367.210 26.410 1368.390 27.590 ;
        RECT 1368.810 26.410 1369.990 27.590 ;
        RECT 1370.410 26.410 1371.590 27.590 ;
        RECT 1372.010 26.410 1373.190 27.590 ;
        RECT 1373.610 26.410 1374.790 27.590 ;
        RECT 1385.210 26.410 1386.390 27.590 ;
        RECT 1386.810 26.410 1387.990 27.590 ;
        RECT 1388.410 26.410 1389.590 27.590 ;
        RECT 1390.010 26.410 1391.190 27.590 ;
        RECT 1391.610 26.410 1392.790 27.590 ;
        RECT 1393.210 26.410 1394.390 27.590 ;
        RECT 1394.810 26.410 1395.990 27.590 ;
        RECT 1396.410 26.410 1397.590 27.590 ;
        RECT 1398.010 26.410 1399.190 27.590 ;
        RECT 1399.610 26.410 1400.790 27.590 ;
        RECT 1401.210 26.410 1402.390 27.590 ;
        RECT 1402.810 26.410 1403.990 27.590 ;
        RECT 1404.410 26.410 1405.590 27.590 ;
        RECT 1406.010 26.410 1407.190 27.590 ;
        RECT 1407.610 26.410 1408.790 27.590 ;
        RECT 1409.210 26.410 1410.390 27.590 ;
        RECT 1410.810 26.410 1411.990 27.590 ;
        RECT 1412.410 26.410 1413.590 27.590 ;
        RECT 1414.010 26.410 1415.190 27.590 ;
        RECT 1415.610 26.410 1416.790 27.590 ;
        RECT 1417.210 26.410 1418.390 27.590 ;
        RECT 1418.810 26.410 1419.990 27.590 ;
        RECT 1420.410 26.410 1421.590 27.590 ;
        RECT 1422.010 26.410 1423.190 27.590 ;
        RECT 1423.610 26.410 1424.790 27.590 ;
      LAYER met5 ;
        RECT 230.000 230.000 1430.000 234.000 ;
        RECT 219.950 128.000 226.000 133.000 ;
        RECT 230.000 131.000 272.000 230.000 ;
        RECT 280.000 131.000 322.000 230.000 ;
        RECT 330.000 131.000 372.000 230.000 ;
        RECT 380.000 131.000 422.000 230.000 ;
        RECT 430.000 131.000 472.000 230.000 ;
        RECT 480.000 131.000 522.000 230.000 ;
        RECT 530.000 131.000 572.000 230.000 ;
        RECT 580.000 131.000 622.000 230.000 ;
        RECT 630.000 131.000 672.000 230.000 ;
        RECT 680.000 131.000 722.000 230.000 ;
        RECT 730.000 131.000 772.000 230.000 ;
        RECT 780.000 131.000 822.000 230.000 ;
        RECT 830.000 131.000 872.000 230.000 ;
        RECT 880.000 131.000 922.000 230.000 ;
        RECT 930.000 131.000 972.000 230.000 ;
        RECT 980.000 131.000 1022.000 230.000 ;
        RECT 1030.000 131.000 1072.000 230.000 ;
        RECT 1080.000 131.000 1122.000 230.000 ;
        RECT 1130.000 131.000 1172.000 230.000 ;
        RECT 1180.000 131.000 1222.000 230.000 ;
        RECT 1230.000 131.000 1272.000 230.000 ;
        RECT 1280.000 131.000 1322.000 230.000 ;
        RECT 1330.000 131.000 1372.000 230.000 ;
        RECT 1380.000 131.000 1422.000 230.000 ;
        RECT 238.000 129.000 272.000 131.000 ;
        RECT 288.000 129.000 322.000 131.000 ;
        RECT 338.000 129.000 372.000 131.000 ;
        RECT 388.000 129.000 422.000 131.000 ;
        RECT 438.000 129.000 472.000 131.000 ;
        RECT 488.000 129.000 522.000 131.000 ;
        RECT 538.000 129.000 572.000 131.000 ;
        RECT 588.000 129.000 622.000 131.000 ;
        RECT 638.000 129.000 672.000 131.000 ;
        RECT 688.000 129.000 722.000 131.000 ;
        RECT 738.000 129.000 772.000 131.000 ;
        RECT 788.000 129.000 822.000 131.000 ;
        RECT 838.000 129.000 872.000 131.000 ;
        RECT 888.000 129.000 922.000 131.000 ;
        RECT 938.000 129.000 972.000 131.000 ;
        RECT 988.000 129.000 1022.000 131.000 ;
        RECT 1038.000 129.000 1072.000 131.000 ;
        RECT 1088.000 129.000 1122.000 131.000 ;
        RECT 1138.000 129.000 1172.000 131.000 ;
        RECT 1188.000 129.000 1222.000 131.000 ;
        RECT 1238.000 129.000 1272.000 131.000 ;
        RECT 1288.000 129.000 1322.000 131.000 ;
        RECT 1338.000 129.000 1372.000 131.000 ;
        RECT 1388.000 129.000 1422.000 131.000 ;
        RECT 219.950 27.000 226.000 32.000 ;
        RECT 238.000 30.000 280.000 129.000 ;
        RECT 288.000 30.000 330.000 129.000 ;
        RECT 338.000 30.000 380.000 129.000 ;
        RECT 388.000 30.000 430.000 129.000 ;
        RECT 438.000 30.000 480.000 129.000 ;
        RECT 488.000 30.000 530.000 129.000 ;
        RECT 538.000 30.000 580.000 129.000 ;
        RECT 588.000 30.000 630.000 129.000 ;
        RECT 638.000 30.000 680.000 129.000 ;
        RECT 688.000 30.000 730.000 129.000 ;
        RECT 738.000 30.000 780.000 129.000 ;
        RECT 788.000 30.000 830.000 129.000 ;
        RECT 838.000 30.000 880.000 129.000 ;
        RECT 888.000 30.000 930.000 129.000 ;
        RECT 938.000 30.000 980.000 129.000 ;
        RECT 988.000 30.000 1030.000 129.000 ;
        RECT 1038.000 30.000 1080.000 129.000 ;
        RECT 1088.000 30.000 1130.000 129.000 ;
        RECT 1138.000 30.000 1180.000 129.000 ;
        RECT 1188.000 30.000 1230.000 129.000 ;
        RECT 1238.000 30.000 1280.000 129.000 ;
        RECT 1288.000 30.000 1330.000 129.000 ;
        RECT 1338.000 30.000 1380.000 129.000 ;
        RECT 1388.000 30.000 1430.000 129.000 ;
        RECT 230.000 26.000 1430.000 30.000 ;
  END
END largecap1
END LIBRARY

