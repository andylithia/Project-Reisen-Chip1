magic
tech sky130A
timestamp 1672105061
<< metal4 >>
rect 0 -3950 400 0
rect 500 -3400 900 0
rect 1000 -2850 1400 0
rect 1500 -1450 2150 0
rect 2250 -50 2900 0
rect 2250 -1150 2300 -50
rect 2850 -1150 2900 -50
rect 2250 -1200 2900 -1150
rect 3100 -50 3750 0
rect 3100 -1150 3150 -50
rect 3700 -1150 3750 -50
rect 3100 -1200 3750 -1150
rect 1500 -2550 1550 -1450
rect 2100 -2550 2150 -1450
rect 1500 -2600 2150 -2550
rect 1000 -3100 1050 -2850
rect 1350 -3100 1400 -2850
rect 1000 -3150 1400 -3100
rect 500 -3650 550 -3400
rect 850 -3650 900 -3400
rect 500 -3700 900 -3650
rect 0 -4200 50 -3950
rect 350 -4200 400 -3950
rect 0 -4250 400 -4200
<< via4 >>
rect 2300 -1150 2850 -50
rect 3150 -1150 3700 -50
rect 1550 -2550 2100 -1450
rect 1050 -3100 1350 -2850
rect 550 -3650 850 -3400
rect 50 -4200 350 -3950
<< metal5 >>
rect 2250 -50 131100 0
rect 2250 -1150 2300 -50
rect 2850 -1150 3150 -50
rect 3700 -1150 131100 -50
rect 2250 -1200 131100 -1150
rect 1500 -1450 129500 -1400
rect 1500 -2550 1550 -1450
rect 2100 -2550 129500 -1450
rect 1500 -2600 129500 -2550
rect 1000 -2850 131000 -2800
rect 1000 -3100 1050 -2850
rect 1350 -3100 131000 -2850
rect 1000 -3150 131000 -3100
rect 500 -3400 130500 -3350
rect 500 -3650 550 -3400
rect 850 -3650 130500 -3400
rect 500 -3700 130500 -3650
rect 0 -3950 130000 -3900
rect 0 -4200 50 -3950
rect 350 -4200 130000 -3950
rect 0 -4250 130000 -4200
<< end >>
