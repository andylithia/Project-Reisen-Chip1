** sch_path:
*+ /home/andylithia/openmpw/Project-Yatsuhashi-Chip1/xschem/2stack_res_matching_newbias_PEX.sch
**.subckt 2stack_res_matching_newbias_PEX
V3 net1 GND 3.3
L1 net3 voi 2n m=1
L6 vout net4 1.3n m=1
C7 net4 voi 1.6p m=1
C1 voi GND 0.6p m=1
R7 net1 net2 1m m=1
R12 net2 net3 5 m=1
R10 vout GND 50 m=1
V1 bias_cascode GND 1.2
I1 GND net5 100u
V9 VDD GND 1.8
C3 VGATE vin 1.6p m=1
V2 vin GND SIN(0 0.9 5G)
XM1 net6 net5 GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 net5 net5 GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
R1 vref0 net6 0.1 m=1
x3 VDD VDD VDD GND GND vref0 vbiasl VDD GND pmirror_tunable_64x_PEX
**** begin user architecture code
.lib /home/andylithia/openmpw/pdk_1/sky130B/libs.tech/ngspice/sky130.lib.spice tt
* .include
*+ /home/andylithia/openmpw/pdk_1/sky130B/libs.ref/sky130_fd_sc_hvl/spice/sky130_fd_sc_hvl.spice


.subckt DUT IREF_L GND VBIAS_CAS INPUT OUTPUT

.subckt sky130_fd_pr__nfet_01v8_6H2JGK a_63_n800# a_n225_n800# a_111_822# a_n321_n800#  a_207_n888#
+ a_n369_n888# a_n33_n800# a_303_822# a_15_n888# a_n81_822# a_n177_n888#  a_159_n800# a_n515_n974# a_n273_822#
+ a_255_n800# a_n413_n800# a_351_n800# a_n129_n800#
X0 a_n129_n800# a_n177_n888# a_n225_n800# a_n515_n974# sky130_fd_pr__nfet_01v8 ad=2.64e+12p
+ pd=1.666e+07u as=2.64e+12p ps=1.666e+07u w=8e+06u l=150000u
X1 a_351_n800# a_303_822# a_255_n800# a_n515_n974# sky130_fd_pr__nfet_01v8 ad=2.48e+12p
+ pd=1.662e+07u as=2.64e+12p ps=1.666e+07u w=8e+06u l=150000u
X2 a_n33_n800# a_n81_822# a_n129_n800# a_n515_n974# sky130_fd_pr__nfet_01v8 ad=2.64e+12p
+ pd=1.666e+07u as=0p ps=0u w=8e+06u l=150000u
X3 a_255_n800# a_207_n888# a_159_n800# a_n515_n974# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.64e+12p
+ ps=1.666e+07u w=8e+06u l=150000u
X4 a_n321_n800# a_n369_n888# a_n413_n800# a_n515_n974# sky130_fd_pr__nfet_01v8 ad=2.64e+12p
+ pd=1.666e+07u as=2.48e+12p ps=1.662e+07u w=8e+06u l=150000u
X5 a_159_n800# a_111_822# a_63_n800# a_n515_n974# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.64e+12p
+ ps=1.666e+07u w=8e+06u l=150000u
X6 a_n225_n800# a_n273_822# a_n321_n800# a_n515_n974# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p
+ ps=0u w=8e+06u l=150000u
X7 a_63_n800# a_15_n888# a_n33_n800# a_n515_n974# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u
+ w=8e+06u l=150000u
.ends

.subckt sky130_fd_pr__res_high_po_0p35_ZE2H5K a_n35_300# a_n165_n862# a_n35_n732#
X0 a_n35_n732# a_n35_300# a_n165_n862# sky130_fd_pr__res_high_po_0p35 l=3e+06u
.ends

.subckt sky130_fd_pr__nfet_03v3_nvt_EV757D a_977_n997# a_n1135_1127# a_603_n1927#  a_n2557_n909#
+ a_n1551_21# a_2241_n2015# a_n445_n997# a_2183_109# a_1235_109# a_n2083_109#  a_n977_1127# a_819_1039#
+ a_n1709_n997# a_n1135_109# a_n2025_n997# a_n1767_n909#  a_1235_n1927# a_n2557_1127# a_n1077_1039# a_n2083_n909#
+ a_n2499_n2015# a_1709_n1927#  a_2399_n997# a_n1235_n997# a_345_1039# a_n503_n909# a_n1767_1127# a_n1293_n909#
+  a_129_n909# a_2083_n2015# a_445_n1927# a_977_21# a_n2083_1127# a_n2499_1039# a_503_n997#  a_919_n1927#
+ a_187_21# a_n503_1127# a_n919_1039# a_1077_n1927# a_129_1127# a_n1293_1127#  a_1609_n997# a_1077_109#
+ a_n977_109# a_977_1039# a_29_n2015# a_n1867_n997# a_1609_21#  a_n445_1039# a_287_n1927# a_n2183_n997#
+ a_n1709_1039# a_2399_n2015# a_1551_n1927#  a_n603_n997# a_1451_21# a_n2025_1039# a_1135_n997# a_n661_n909#
+ a_n1393_n997# a_287_n909#  a_129_109# a_2399_1039# a_n1925_n909# a_n445_21# a_n1235_1039# a_n2241_n909#
+ a_n29_n1927#  a_761_n1927# a_661_n997# a_n661_1127# a_503_1039# a_1393_n1927# a_n2183_21# a_287_1127#
+  a_n1925_1127# a_n1451_n909# a_n2241_1127# a_1867_n1927# a_1767_n997# a_2083_n997#  a_1709_109# a_n2557_109#
+ a_n1609_109# a_1609_1039# a_n1867_21# a_n1451_1127# a_n1867_1039#  a_n2183_1039# a_n761_n997# a_1293_n997#
+ a_n1077_21# a_n2341_n997# a_n603_1039# a_919_n909#  a_1135_1039# a_n29_109# a_n1393_1039# a_n1135_n1927#
+ a_1551_109# a_n1451_109# a_345_21#  a_29_21# a_661_1039# a_n1609_n1927# a_n1551_n997# a_919_1127# a_445_n909#
+ a_n503_n1927#  a_n129_n2015# a_2499_109# a_n503_109# a_n2399_109# a_603_109# a_445_1127# a_1767_1039#
+  a_n1235_n2015# a_2083_21# a_2083_1039# a_n1709_n2015# a_1925_n997# a_n603_n2015#  a_2241_n997# a_n761_1039#
+ a_n345_n1927# a_1767_21# a_1293_1039# a_n603_21# a_1077_n909#  a_n819_n1927# a_2025_n1927# a_n2341_1039#
+ a_1451_n997# a_1393_109# a_n1293_109#  a_n1077_n2015# a_n1451_n1927# a_n2341_21# a_n1925_n1927# a_1077_1127#
+ a_n1551_1039#  a_2499_n909# a_n445_n2015# a_503_n2015# a_n2691_n2149# a_n187_n1927# a_n345_109#  a_n2499_21#
+ a_n919_n2015# a_445_109# a_603_n909# a_n1551_n2015# a_1135_n2015# a_2499_1127#  a_n1293_n1927# a_n1235_21#
+ a_1609_n2015# a_n1767_n1927# a_1925_1039# a_603_1127#  a_1709_n909# a_345_n2015# a_n661_n1927# a_2241_1039#
+ a_n287_n2015# a_2341_n1927#  a_2025_n909# a_819_n2015# a_n1925_109# a_503_21# a_n1393_n2015# a_1451_1039#
+ a_1709_1127#  a_1235_n909# a_n1867_n2015# a_2025_1127# a_2025_109# a_n187_109# a_n761_n2015# a_2241_21#
+  a_761_n909# a_187_n2015# a_287_109# a_2183_n1927# a_1235_1127# a_1451_n2015# a_n977_n1927#  a_2399_21#
+ a_1925_n2015# a_1925_21# a_761_1127# a_1867_n909# a_2183_n909# a_661_n2015#  a_1135_21# a_1867_109# a_n1767_109#
+ a_n29_n909# a_n919_21# a_1867_1127# a_1293_n2015#  a_n761_21# a_2183_1127# a_1393_n909# a_2499_n1927#
+ a_n129_21# a_1767_n2015# a_29_n997#  a_n819_109# a_n29_1127# a_919_109# a_1393_1127# a_n129_n997# a_977_n2015#
+ a_n187_n909#  a_n2025_n2015# a_187_n997# a_n661_109# a_n1393_21# a_n187_1127# a_761_109# a_819_21#  a_2341_n909#
+ a_661_21# a_n2241_n1927# a_29_1039# a_1551_n909# a_n2399_n909# a_2341_1127#  a_n287_n997# a_n819_n909#
+ a_n129_1039# a_1551_1127# a_n2399_1127# a_n2341_n2015#  a_819_n997# a_n2083_n1927# a_2341_109# a_n2241_109#
+ a_n819_1127# a_187_1039# a_n345_n909#  a_n2557_n1927# a_n1077_n997# a_n1609_n909# a_345_n997# a_1293_21#
+ a_n2499_n997#  a_n345_1127# a_129_n1927# a_n2025_21# a_n1609_1127# a_n2183_n2015# a_n1135_n909#  a_n919_n997#
+ a_n287_21# a_n977_n909# a_n2399_n1927# a_n287_1039# a_n1709_21#
X0 a_n29_1127# a_n129_1039# a_n187_1127# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=1.16e+12p
+ pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X1 a_603_1127# a_503_1039# a_445_1127# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=1.16e+12p
+ pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X2 a_n661_109# a_n761_21# a_n819_109# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=1.16e+12p
+ pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X3 a_n1293_n1927# a_n1393_n2015# a_n1451_n1927# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt
+ ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X4 a_n661_n909# a_n761_n997# a_n819_n909# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=1.16e+12p
+ pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X5 a_n29_n1927# a_n129_n2015# a_n187_n1927# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=1.16e+12p
+ pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X6 a_129_109# a_29_21# a_n29_109# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=1.16e+12p
+ pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X7 a_1551_n1927# a_1451_n2015# a_1393_n1927# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=1.16e+12p
+ pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X8 a_n1609_n1927# a_n1709_n2015# a_n1767_n1927# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt
+ ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X9 a_2183_n1927# a_2083_n2015# a_2025_n1927# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=1.16e+12p
+ pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X10 a_n187_109# a_n287_21# a_n345_109# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=1.16e+12p
+ pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X11 a_919_n909# a_819_n997# a_761_n909# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=1.16e+12p
+ pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X12 a_n187_n1927# a_n287_n2015# a_n345_n1927# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u
+ as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X13 a_n1767_n1927# a_n1867_n2015# a_n1925_n1927# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p
+ pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X14 a_2025_n909# a_1925_n997# a_1867_n909# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=1.16e+12p
+ pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X15 a_1235_1127# a_1135_1039# a_1077_1127# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=1.16e+12p
+ pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X16 a_n2399_n1927# a_n2499_n2015# a_n2557_n1927# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt
+ ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X17 a_761_n909# a_661_n997# a_603_n909# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u
+ as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X18 a_n187_n909# a_n287_n997# a_n345_n909# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=1.16e+12p
+ pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X19 a_n1135_1127# a_n1235_1039# a_n1293_1127# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt
+ ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X20 a_2025_n1927# a_1925_n2015# a_1867_n1927# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u
+ as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X21 a_n819_109# a_n919_21# a_n977_109# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u
+ as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X22 a_2341_n909# a_2241_n997# a_2183_n909# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=1.16e+12p
+ pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X23 a_n2241_n909# a_n2341_n997# a_n2399_n909# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt
+ ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X24 a_n345_109# a_n445_21# a_n503_109# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u
+ as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X25 a_287_n909# a_187_n997# a_129_n909# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=1.16e+12p
+ pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X26 a_129_n1927# a_29_n2015# a_n29_n1927# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=1.16e+12p
+ pd=8.58e+06u as=0p ps=0u w=4e+06u l=500000u
X27 a_n503_109# a_n603_21# a_n661_109# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p
+ ps=0u w=4e+06u l=500000u
X28 a_1393_n909# a_1293_n997# a_1235_n909# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=1.16e+12p
+ pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X29 a_n1293_n909# a_n1393_n997# a_n1451_n909# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt
+ ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X30 a_1867_1127# a_1767_1039# a_1709_1127# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=1.16e+12p
+ pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X31 a_n1767_1127# a_n1867_1039# a_n1925_1127# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt
+ ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X32 a_n29_109# a_n129_21# a_n187_109# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p
+ ps=0u w=4e+06u l=500000u
X33 a_n2399_109# a_n2499_21# a_n2557_109# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=1.16e+12p
+ pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X34 a_445_n1927# a_345_n2015# a_287_n1927# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=1.16e+12p
+ pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X35 a_n2083_1127# a_n2183_1039# a_n2241_1127# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt
+ ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X36 a_2183_1127# a_2083_1039# a_2025_1127# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=1.16e+12p
+ pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X37 a_1867_109# a_1767_21# a_1709_109# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=1.16e+12p
+ pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X38 a_1393_109# a_1293_21# a_1235_109# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=1.16e+12p
+ pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X39 a_n345_n909# a_n445_n997# a_n503_n909# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u
+ as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X40 a_1077_109# a_977_21# a_919_109# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=1.16e+12p
+ pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X41 a_2499_n909# a_2399_n997# a_2341_n909# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=1.16e+12p
+ pd=8.58e+06u as=0p ps=0u w=4e+06u l=500000u
X42 a_n2083_109# a_n2183_21# a_n2241_109# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=1.16e+12p
+ pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X43 a_919_n1927# a_819_n2015# a_761_n1927# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=1.16e+12p
+ pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X44 a_n2399_n909# a_n2499_n997# a_n2557_n909# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u
+ as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X45 a_2025_109# a_1925_21# a_1867_109# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=1.16e+12p
+ pd=8.58e+06u as=0p ps=0u w=4e+06u l=500000u
X46 a_n819_1127# a_n919_1039# a_n977_1127# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=1.16e+12p
+ pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X47 a_n1925_n1927# a_n2025_n2015# a_n2083_n1927# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p
+ pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X48 a_1551_109# a_1451_21# a_1393_109# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=1.16e+12p
+ pd=8.58e+06u as=0p ps=0u w=4e+06u l=500000u
X49 a_129_n909# a_29_n997# a_n29_n909# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u
+ as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X50 a_n661_1127# a_n761_1039# a_n819_1127# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=1.16e+12p
+ pd=8.58e+06u as=0p ps=0u w=4e+06u l=500000u
X51 a_1077_n1927# a_977_n2015# a_919_n1927# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=1.16e+12p
+ pd=8.58e+06u as=0p ps=0u w=4e+06u l=500000u
X52 a_1709_n909# a_1609_n997# a_1551_n909# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=1.16e+12p
+ pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X53 a_n1451_n1927# a_n1551_n2015# a_n1609_n1927# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p
+ pd=0u as=0p ps=0u w=4e+06u l=500000u
X54 a_n1609_n909# a_n1709_n997# a_n1767_n909# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt
+ ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X55 a_n2083_n1927# a_n2183_n2015# a_n2241_n1927# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p
+ pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X56 a_445_n909# a_345_n997# a_287_n909# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=1.16e+12p
+ pd=8.58e+06u as=0p ps=0u w=4e+06u l=500000u
X57 a_n2241_109# a_n2341_21# a_n2399_109# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u
+ as=0p ps=0u w=4e+06u l=500000u
X58 a_761_109# a_661_21# a_603_109# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=1.16e+12p
+ pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X59 a_2341_n1927# a_2241_n2015# a_2183_n1927# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt
+ ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=500000u
X60 a_1551_n909# a_1451_n997# a_1393_n909# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u
+ as=0p ps=0u w=4e+06u l=500000u
X61 a_n1451_n909# a_n1551_n997# a_n1609_n909# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u
+ as=0p ps=0u w=4e+06u l=500000u
X62 a_n1925_n909# a_n2025_n997# a_n2083_n909# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt
+ ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X63 a_919_1127# a_819_1039# a_761_1127# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=1.16e+12p
+ pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X64 a_2025_1127# a_1925_1039# a_1867_1127# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u
+ as=0p ps=0u w=4e+06u l=500000u
X65 a_n345_n1927# a_n445_n2015# a_n503_n1927# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u
+ as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X66 a_1709_109# a_1609_21# a_1551_109# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p
+ ps=0u w=4e+06u l=500000u
X67 a_287_109# a_187_21# a_129_109# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=1.16e+12p
+ pd=8.58e+06u as=0p ps=0u w=4e+06u l=500000u
X68 a_n187_1127# a_n287_1039# a_n345_1127# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u
+ as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X69 a_761_1127# a_661_1039# a_603_1127# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p
+ ps=0u w=4e+06u l=500000u
X70 a_1235_109# a_1135_21# a_1077_109# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p
+ ps=0u w=4e+06u l=500000u
X71 a_2341_1127# a_2241_1039# a_2183_1127# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=1.16e+12p
+ pd=8.58e+06u as=0p ps=0u w=4e+06u l=500000u
X72 a_n2241_1127# a_n2341_1039# a_n2399_1127# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u
+ as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X73 a_n977_n909# a_n1077_n997# a_n1135_n909# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=1.16e+12p
+ pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X74 a_919_109# a_819_21# a_761_109# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p
+ ps=0u w=4e+06u l=500000u
X75 a_n1925_109# a_n2025_21# a_n2083_109# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=1.16e+12p
+ pd=8.58e+06u as=0p ps=0u w=4e+06u l=500000u
X76 a_n819_n1927# a_n919_n2015# a_n977_n1927# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt
+ ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X77 a_1077_n909# a_977_n997# a_919_n909# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=1.16e+12p
+ pd=8.58e+06u as=0p ps=0u w=4e+06u l=500000u
X78 a_445_109# a_345_21# a_287_109# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=1.16e+12p
+ pd=8.58e+06u as=0p ps=0u w=4e+06u l=500000u
X79 a_n503_n909# a_n603_n997# a_n661_n909# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u
+ as=0p ps=0u w=4e+06u l=500000u
X80 a_287_1127# a_187_1039# a_129_1127# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=1.16e+12p
+ pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X81 a_n977_n1927# a_n1077_n2015# a_n1135_n1927# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p
+ pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X82 a_1393_1127# a_1293_1039# a_1235_1127# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=1.16e+12p
+ pd=8.58e+06u as=0p ps=0u w=4e+06u l=500000u
X83 a_n1293_1127# a_n1393_1039# a_n1451_1127# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u
+ as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X84 a_1235_n1927# a_1135_n2015# a_1077_n1927# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt
+ ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=500000u
X85 a_603_109# a_503_21# a_445_109# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p
+ ps=0u w=4e+06u l=500000u
X86 a_603_n909# a_503_n997# a_445_n909# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p
+ ps=0u w=4e+06u l=500000u
X87 a_n29_n909# a_n129_n997# a_n187_n909# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u
+ as=0p ps=0u w=4e+06u l=500000u
X88 a_1393_n1927# a_1293_n2015# a_1235_n1927# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u
+ as=0p ps=0u w=4e+06u l=500000u
X89 a_603_n1927# a_503_n2015# a_445_n1927# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=1.16e+12p
+ pd=8.58e+06u as=0p ps=0u w=4e+06u l=500000u
X90 a_1709_n1927# a_1609_n2015# a_1551_n1927# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt
+ ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=500000u
X91 a_n345_1127# a_n445_1039# a_n503_1127# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u
+ as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X92 a_761_n1927# a_661_n2015# a_603_n1927# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u
+ as=0p ps=0u w=4e+06u l=500000u
X93 a_n2399_1127# a_n2499_1039# a_n2557_1127# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u
+ as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X94 a_2499_1127# a_2399_1039# a_2341_1127# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=1.16e+12p
+ pd=8.58e+06u as=0p ps=0u w=4e+06u l=500000u
X95 a_n1767_109# a_n1867_21# a_n1925_109# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=1.16e+12p
+ pd=8.58e+06u as=0p ps=0u w=4e+06u l=500000u
X96 a_1867_n1927# a_1767_n2015# a_1709_n1927# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u
+ as=0p ps=0u w=4e+06u l=500000u
X97 a_n1293_109# a_n1393_21# a_n1451_109# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=1.16e+12p
+ pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X98 a_2499_n1927# a_2399_n2015# a_2341_n1927# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt
+ ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=500000u
X99 a_1235_n909# a_1135_n997# a_1077_n909# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u
+ as=0p ps=0u w=4e+06u l=500000u
X100 a_n1135_n909# a_n1235_n997# a_n1293_n909# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p
+ pd=0u as=0p ps=0u w=4e+06u l=500000u
X101 a_129_1127# a_29_1039# a_n29_1127# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p
+ ps=0u w=4e+06u l=500000u
X102 a_n1609_1127# a_n1709_1039# a_n1767_1127# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt
+ ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=500000u
X103 a_1709_1127# a_1609_1039# a_1551_1127# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u
+ as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X104 a_445_1127# a_345_1039# a_287_1127# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u
+ as=0p ps=0u w=4e+06u l=500000u
X105 a_n1451_109# a_n1551_21# a_n1609_109# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u
+ as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X106 a_n2241_n1927# a_n2341_n2015# a_n2399_n1927# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p
+ pd=0u as=0p ps=0u w=4e+06u l=500000u
X107 a_n1925_1127# a_n2025_1039# a_n2083_1127# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p
+ pd=0u as=0p ps=0u w=4e+06u l=500000u
X108 a_n1451_1127# a_n1551_1039# a_n1609_1127# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p
+ pd=0u as=0p ps=0u w=4e+06u l=500000u
X109 a_1551_1127# a_1451_1039# a_1393_1127# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u
+ as=0p ps=0u w=4e+06u l=500000u
X110 a_2499_109# a_2399_21# a_2341_109# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=1.16e+12p
+ pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X111 a_n977_109# a_n1077_21# a_n1135_109# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u
+ as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X112 a_n503_n1927# a_n603_n2015# a_n661_n1927# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p
+ pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
X113 a_1867_n909# a_1767_n997# a_1709_n909# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u
+ as=0p ps=0u w=4e+06u l=500000u
X114 a_n1767_n909# a_n1867_n997# a_n1925_n909# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p
+ pd=0u as=0p ps=0u w=4e+06u l=500000u
X115 a_287_n1927# a_187_n2015# a_129_n1927# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u
+ as=0p ps=0u w=4e+06u l=500000u
X116 a_n977_1127# a_n1077_1039# a_n1135_1127# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u
+ as=0p ps=0u w=4e+06u l=500000u
X117 a_2183_n909# a_2083_n997# a_2025_n909# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u
+ as=0p ps=0u w=4e+06u l=500000u
X118 a_n1609_109# a_n1709_21# a_n1767_109# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u
+ as=0p ps=0u w=4e+06u l=500000u
X119 a_1077_1127# a_977_1039# a_919_1127# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u
+ as=0p ps=0u w=4e+06u l=500000u
X120 a_n661_n1927# a_n761_n2015# a_n819_n1927# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p
+ pd=0u as=0p ps=0u w=4e+06u l=500000u
X121 a_n2083_n909# a_n2183_n997# a_n2241_n909# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p
+ pd=0u as=0p ps=0u w=4e+06u l=500000u
X122 a_2183_109# a_2083_21# a_2025_109# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=1.16e+12p
+ pd=8.58e+06u as=0p ps=0u w=4e+06u l=500000u
X123 a_n1135_109# a_n1235_21# a_n1293_109# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u
+ as=0p ps=0u w=4e+06u l=500000u
X124 a_n503_1127# a_n603_1039# a_n661_1127# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u
+ as=0p ps=0u w=4e+06u l=500000u
X125 a_n1135_n1927# a_n1235_n2015# a_n1293_n1927# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p
+ pd=0u as=0p ps=0u w=4e+06u l=500000u
X126 a_2341_109# a_2241_21# a_2183_109# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p
+ ps=0u w=4e+06u l=500000u
X127 a_n819_n909# a_n919_n997# a_n977_n909# a_n2691_n2149# sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u
+ as=0p ps=0u w=4e+06u l=500000u
.ends

.subckt RF_nfet_3v_dnwell_cascode D G2 G1 SB DNW VSUBS
Xsky130_fd_pr__nfet_03v3_nvt_EV757D_0 G1 D SB SB G2 G1 G2 SB SB D SB G1 G2 D G2 D  SB SB G2 D G2 D
+ G1 G2 G1 D D SB D G1 D G1 D G2 G1 SB G1 D G2 D D SB G1 D SB G1 G1  G2 G1 G2 SB G2 G2 G1 SB G2 G1 G2 G1
+ SB G2 SB D G1 SB G2 G2 SB SB D G1 SB G1 D G2  SB SB D SB SB G1 G1 D SB SB G1 G2 D G2 G2 G2 G1 G2 G2 G2
+ SB G1 SB G2 D SB D G1 G1  G1 SB G2 SB D D G2 SB D D SB D G1 G2 G1 G1 G2 G1 G2 G1 G2 SB G1 G1 G2 D D D
+ G2 G1  D SB G2 D G2 SB D G2 SB G2 G1 SB D SB G2 G2 D SB G2 G1 SB SB G2 G1 D G1 SB D G1  SB G1 G2 D D
+ G1 SB G1 G2 G1 D SB G2 D D D G2 G1 D G1 SB SB SB G1 SB G1 G1 G1 D SB  SB G1 G1 SB D SB G2 SB G1 G2 SB
+ D SB G2 G1 G1 D SB SB D G2 G1 D G2 G1 SB G2 D D  G1 D G1 SB G1 SB D D G2 D G2 SB D G2 G1 D D SB D G1
+ SB SB G2 SB G1 G1 G2 SB D G2  SB G2 D G2 G2 SB D G2 G2 sky130_fd_pr__nfet_03v3_nvt_EV757D
C0 D SB 132.51fF
C1 G1 SB 25.45fF
C2 G2 DNW 3.39fF
C3 D G1 19.92fF
C4 DNW SB 92.93fF
C5 G2 SB 27.04fF
C6 G1 DNW 2.85fF
C7 D G2 19.94fF
C8 SB VSUBS -3.31fF
C9 DNW VSUBS 112.06fF
C10 D VSUBS -2.56fF
C11 G1 VSUBS 3.47fF
C12 G2 VSUBS 3.41fF
.ends

.subckt sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap G D S VSUBS
X0 D G S VSUBS sky130_fd_pr__nfet_01v8 ad=4.242e+12p pd=3.198e+07u as=2.828e+12p ps=2.132e+07u
+ w=5.05e+06u l=150000u
X1 D G S VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X2 S G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X3 S G D VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
C0 S D 6.34fF
.ends

.subckt RF_nfet_8xW5p0L0p15 G S SD
Xsky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0 G S SD S
+ sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap
Xsky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_1 G S SD S
+ sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap
Xsky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_2 G S SD S
+ sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap
C0 G 0 2.12fF
.ends

.subckt RF_nfet_driver_64x8 G D SG
XRF_nfet_8xW5p0L0p15_9 G SG D RF_nfet_8xW5p0L0p15
XRF_nfet_8xW5p0L0p15_10 G SG D RF_nfet_8xW5p0L0p15
XRF_nfet_8xW5p0L0p15_11 G SG D RF_nfet_8xW5p0L0p15
XRF_nfet_8xW5p0L0p15_0 G SG D RF_nfet_8xW5p0L0p15
XRF_nfet_8xW5p0L0p15_1 G SG D RF_nfet_8xW5p0L0p15
XRF_nfet_8xW5p0L0p15_2 G SG D RF_nfet_8xW5p0L0p15
XRF_nfet_8xW5p0L0p15_3 G SG D RF_nfet_8xW5p0L0p15
XRF_nfet_8xW5p0L0p15_4 G SG D RF_nfet_8xW5p0L0p15
XRF_nfet_8xW5p0L0p15_5 G SG D RF_nfet_8xW5p0L0p15
XRF_nfet_8xW5p0L0p15_6 G SG D RF_nfet_8xW5p0L0p15
XRF_nfet_8xW5p0L0p15_7 G SG D RF_nfet_8xW5p0L0p15
XRF_nfet_8xW5p0L0p15_8 G SG D RF_nfet_8xW5p0L0p15
C0 D G 18.33fF
C1 D SG 24.68fF
C2 G SG 14.51fF
C3 D 0 -3.92fF
C4 SG 0 -25.16fF
C5 G 0 17.76fF
.ends

.subckt PA_core_1 DRAIN TOPBIAS_R GATE TOPBIAS_L MID VSUB
XRF_nfet_3v_dnwell_cascode_0 DRAIN RF_nfet_3v_dnwell_cascode_0/G2 RF_nfet_3v_dnwell_cascode_0/G1
+  MID VSUB VSUB RF_nfet_3v_dnwell_cascode
XRF_nfet_driver_64x8_0 GATE MID VSUB RF_nfet_driver_64x8
Xsky130_fd_pr__res_high_po_0p35_ZE2H5K_0 RF_nfet_3v_dnwell_cascode_0/G2 VSUB TOPBIAS_L
+  sky130_fd_pr__res_high_po_0p35_ZE2H5K
Xsky130_fd_pr__res_high_po_0p35_ZE2H5K_1 TOPBIAS_R VSUB RF_nfet_3v_dnwell_cascode_0/G1
+  sky130_fd_pr__res_high_po_0p35_ZE2H5K
C0 VSUB DRAIN 2.00fF
C1 VSUB MID 6.73fF
C2 VSUB 0 85.58fF
C3 GATE 0 17.76fF
C4 MID 0 -11.48fF
C5 DRAIN 0 -2.02fF
C6 RF_nfet_3v_dnwell_cascode_0/G1 0 4.12fF
C7 RF_nfet_3v_dnwell_cascode_0/G2 0 4.07fF
.ends

* PORTS:
* IREF_L, GND, INPUT, OUTPUT, VGATE_CAS


Xsky130_fd_pr__nfet_01v8_6H2JGK_0 IREF_L GND IREF_L IREF_L IREF_L IREF_L GND IREF_L  IREF_L IREF_L
+ IREF_L GND GND IREF_L IREF_L GND GND IREF_L sky130_fd_pr__nfet_01v8_6H2JGK
Xsky130_fd_pr__res_high_po_0p35_ZE2H5K_0 IREF_L GND INPUT sky130_fd_pr__res_high_po_0p35_ZE2H5K
XPA_core_1_0 OUTPUT VGATE_CAS INPUT VGATE_CAS PA_core_1_0/MID GND PA_core_1
X0 VGATE_CAS GND sky130_fd_pr__cap_mim_m3_2 l=1.6e+07u w=1.9e+07u
X1 GND VGATE_CAS sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.9e+07u
X2 IREF_L GND sky130_fd_pr__cap_mim_m3_2 l=1.55e+07u w=2.25e+07u
X3 GND IREF_L sky130_fd_pr__cap_mim_m3_1 l=1.55e+07u w=2.25e+07u
C0 m5_n1000_18400# IREF_L 7.66fF
C1 VGATE_CAS GND 57.37fF
C2 GND IREF_L 84.58fF
C3 OUTPUT VGATE_CAS 4.71fF
C4 INPUT IREF_L 2.32fF
C8 VGATE_CAS 0 11.90fF
C10 INPUT 0 32.79fF
C12 OUTPUT 0 67.83fF
C13 PA_core_1_0/RF_nfet_3v_dnwell_cascode_0/G1 0 4.12fF
C14 PA_core_1_0/RF_nfet_3v_dnwell_cascode_0/G2 0 4.07fF
C15 IREF_L 0 16.35fF
.ends

XDUT vbiasl GND bias_cascode VGATE voi DUT

.options savecurrents
* XMU_0 gu voi mid mid rf_nfet_6xaM02_extracted
* XMU_1 gu voi mid mid rf_nfet_6xaM02_extracted
* XMU_2 gu voi mid mid rf_nfet_6xaM02_extracted
* XMU_3 gu voi mid mid rf_nfet_6xaM02_extracted
* XMU_4 gu voi mid mid rf_nfet_6xaM02_extracted
* XMU_5 gu voi mid mid rf_nfet_6xaM02_extracted
* XMD_0 gd mid gnd gnd rf_nfet_6xaM02_extracted
* XMD_1 gd mid gnd gnd rf_nfet_6xaM02_extracted
* XMD_2 gd mid gnd gnd rf_nfet_6xaM02_extracted
* XMD_3 gd mid gnd gnd rf_nfet_6xaM02_extracted
* XMD_4 gd mid gnd gnd rf_nfet_6xaM02_extracted
* XMD_5 gd mid gnd gnd rf_nfet_6xaM02_extracted
.tran 10ps 40ns
* .sp dec 1000 1e9 10e9 1
* .dc I1 0 10m 0.1m
.control
run
display
* plot @r5[i]
* let zout=@rload[r]
* let zin=50
* plot voi
* plot vout
* plot @c1[i]

plot vbiasl
plot @l1[i]


* meas TRAN vout_rms rms v(vout)
* meas TRAN isp_hi_avg  avg @r7[i]
* meas TRAN isp_mid_avg avg @r9[i]
* meas TRAN vin_rms rms v(vin)
* meas TRAN isp_1p8_avg avg @rsense2[i]
* let psp_rms  = isp_hi_avg*3.6 + isp_mid_avg*2.2
* let pout_rms = vout_rms^2/zout
* let pin_rms  = vin_rms^2/zin
* print psp_rms
* print ((pout_rms-pin_rms)/psp_rms)*100
* print 10*log10(pout_rms*1000)

* plot gd vmid voi vout

* let pout = mag(@rload[i]*vout)
* let poutdbm = log10((pout/(1e-3))*10
* plot pout

.endc


**** end user architecture code
**.ends

* expanding   symbol:  pmirror_tunable_64x_PEX.sym # of pins=9
** sym_path: /home/andylithia/openmpw/Project-Yatsuhashi-Chip1/xschem/pmirror_tunable_64x_PEX.sym
** sch_path: /home/andylithia/openmpw/Project-Yatsuhashi-Chip1/xschem/pmirror_tunable_64x_PEX.sch
.subckt pmirror_tunable_64x_PEX  VHI G2 G4 VSUBS G8 IREF IOUT G16 G32
*.ipin G2
*.ipin G4
*.ipin G8
*.ipin G16
*.ipin G32
*.iopin VHI
*.iopin VSUBS
*.iopin IREF
*.iopin IOUT
**** begin user architecture code

* SPICE3 file created from pmirror_pfet_64x_complete.ext - technology: sky130B
X0 pmirror_pfet_64x_flat_0/G32 IREF VSUBS sky130_fd_pr__res_xhigh_po_0p35 l=500000u
X1 pmirror_pfet_64x_flat_0/G4  IREF VSUBS sky130_fd_pr__res_xhigh_po_0p35 l=500000u
X2 pmirror_pfet_64x_flat_0/G8  IREF VSUBS sky130_fd_pr__res_xhigh_po_0p35 l=500000u
X3 pmirror_pfet_64x_flat_0/G2  IREF VSUBS sky130_fd_pr__res_xhigh_po_0p35 l=500000u
X5 pmirror_pfet_64x_flat_0/G16 IREF VSUBS sky130_fd_pr__res_xhigh_po_0p35 l=500000u

X7 VHI pmirror_pfet_64x_flat_0/G32 IOUT VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u
+ l=300000u
X8 IOUT pmirror_pfet_64x_flat_0/G32 VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u
+ l=300000u
X11 IOUT pmirror_pfet_64x_flat_0/G32 VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u
+ w=1e+06u l=300000u
X16 VHI pmirror_pfet_64x_flat_0/G32 IOUT VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u
+ w=1e+06u l=300000u
X17 VHI pmirror_pfet_64x_flat_0/G32 IOUT VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u
+ w=1e+06u l=300000u
X18 VHI pmirror_pfet_64x_flat_0/G32 IOUT VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u
+ w=1e+06u l=300000u
X21 IOUT pmirror_pfet_64x_flat_0/G32 VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u
+ w=1e+06u l=300000u
X22 IOUT pmirror_pfet_64x_flat_0/G32 VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u
+ w=1e+06u l=300000u
X27 IOUT pmirror_pfet_64x_flat_0/G32 VHI VHI sky130_fd_pr__pfet_01v8 ad=1p pd=0u as=0p ps=0u
+ w=1e+06u l=300000u
X28 IOUT pmirror_pfet_64x_flat_0/G32 VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u
+ w=1e+06u l=300000u
X29 VHI pmirror_pfet_64x_flat_0/G32 IOUT VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u
+ w=1e+06u l=300000u
X25 VHI pmirror_pfet_64x_flat_0/G32 IOUT VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u
+ w=1e+06u l=300000u
X35 VHI pmirror_pfet_64x_flat_0/G32 IOUT VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u
+ w=1e+06u l=300000u
X38 VHI pmirror_pfet_64x_flat_0/G32 IOUT VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u
+ w=1e+06u l=300000u
X41 VHI pmirror_pfet_64x_flat_0/G32 IOUT VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u
+ w=1e+06u l=300000u
X43 IOUT pmirror_pfet_64x_flat_0/G32 VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u
+ w=1e+06u l=300000u
X44 IOUT pmirror_pfet_64x_flat_0/G32 VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u
+ w=1e+06u l=300000u
X46 VHI pmirror_pfet_64x_flat_0/G32 IOUT VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u
+ w=1e+06u l=300000u
X54 VHI pmirror_pfet_64x_flat_0/G32 IOUT VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u
+ w=1e+06u l=300000u
X55 IOUT pmirror_pfet_64x_flat_0/G32 VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u
+ w=1e+06u l=300000u
X56 IOUT pmirror_pfet_64x_flat_0/G32 VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u
+ w=1e+06u l=300000u
X60 IOUT pmirror_pfet_64x_flat_0/G32 VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u
+ w=1e+06u l=300000u
X61 IOUT pmirror_pfet_64x_flat_0/G32 VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u
+ w=1e+06u l=300000u
X62 VHI pmirror_pfet_64x_flat_0/G32 IOUT VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u
+ w=1e+06u l=300000u
X67 IOUT pmirror_pfet_64x_flat_0/G32 VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u
+ w=1e+06u l=300000u
X68 IOUT pmirror_pfet_64x_flat_0/G32 VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u
+ w=1e+06u l=300000u
X50 VHI pmirror_pfet_64x_flat_0/G32 IOUT VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u
+ w=1e+06u l=300000u
X73 VHI pmirror_pfet_64x_flat_0/G32 IOUT VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u
+ w=1e+06u l=300000u
X74 IOUT pmirror_pfet_64x_flat_0/G32 VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u
+ w=1e+06u l=300000u
X75 IOUT pmirror_pfet_64x_flat_0/G32 VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u
+ w=1e+06u l=300000u
X69 VHI pmirror_pfet_64x_flat_0/G32 IOUT VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u
+ w=1e+06u l=300000u
X81 VHI pmirror_pfet_64x_flat_0/G32 IOUT VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u
+ w=1e+06u l=300000u

X49 VHI VHI IOUT VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X79 IREF IREF VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u

X6 IOUT pmirror_pfet_64x_flat_0/G16 VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u
+ l=300000u
X9 VHI pmirror_pfet_64x_flat_0/G16 IOUT VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u
+ l=300000u
X10 IOUT pmirror_pfet_64x_flat_0/G16 VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u
+ w=1e+06u l=300000u
X19 IOUT pmirror_pfet_64x_flat_0/G16 VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u
+ w=1e+06u l=300000u
X20 IOUT pmirror_pfet_64x_flat_0/G16 VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u
+ w=1e+06u l=300000u
X26 VHI pmirror_pfet_64x_flat_0/G16 IOUT VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u
+ w=1e+06u l=300000u
X30 IOUT pmirror_pfet_64x_flat_0/G16 VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u
+ w=1e+06u l=300000u
X33 IOUT pmirror_pfet_64x_flat_0/G16 VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u
+ w=1e+06u l=300000u
X36 VHI pmirror_pfet_64x_flat_0/G16 IOUT VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u
+ w=1e+06u l=300000u
X45 VHI pmirror_pfet_64x_flat_0/G16 IOUT VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u
+ w=1e+06u l=300000u
X53 VHI pmirror_pfet_64x_flat_0/G16 IOUT VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u
+ w=1e+06u l=300000u
X57 VHI pmirror_pfet_64x_flat_0/G16 IOUT VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u
+ w=1e+06u l=300000u
X58 VHI pmirror_pfet_64x_flat_0/G16 IOUT VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u
+ w=1e+06u l=300000u
X65 VHI pmirror_pfet_64x_flat_0/G16 IOUT VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u
+ w=1e+06u l=300000u
X82 IOUT pmirror_pfet_64x_flat_0/G16 VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u
+ w=1e+06u l=300000u
X83 IOUT pmirror_pfet_64x_flat_0/G16 VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u
+ w=1e+06u l=300000u

X14 IOUT pmirror_pfet_64x_flat_0/G8 VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u
+ l=300000u
X23 VHI pmirror_pfet_64x_flat_0/G8 IOUT VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u
+ l=300000u
X31 VHI pmirror_pfet_64x_flat_0/G8 IOUT VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u
+ l=300000u
X32 VHI pmirror_pfet_64x_flat_0/G8 IOUT VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u
+ l=300000u
X42 VHI pmirror_pfet_64x_flat_0/G8 IOUT VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u
+ l=300000u
X72 IOUT pmirror_pfet_64x_flat_0/G8 VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u
+ l=300000u
X80 IOUT pmirror_pfet_64x_flat_0/G8 VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u
+ l=300000u
X84 IOUT pmirror_pfet_64x_flat_0/G8 VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u
+ l=300000u

X85 IOUT pmirror_pfet_64x_flat_0/G4 VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u
+ l=300000u
X39 VHI pmirror_pfet_64x_flat_0/G4 IOUT VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u
+ l=300000u
X40 VHI pmirror_pfet_64x_flat_0/G4 IOUT VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u
+ l=300000u
X70 IOUT pmirror_pfet_64x_flat_0/G4 VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u
+ l=300000u

X48 VHI pmirror_pfet_64x_flat_0/G2 IOUT VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u
+ l=300000u
X15 IOUT pmirror_pfet_64x_flat_0/G2 VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u
+ l=300000u

X86 VHI G32 pmirror_pfet_64x_flat_0/G32 VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u
+ w=30e+06u l=150000u
X87 VHI G16 pmirror_pfet_64x_flat_0/G16 VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u
+ w=30e+06u l=150000u
X88 VHI G2 pmirror_pfet_64x_flat_0/G2 VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=30e+06u
+ l=150000u
X89 VHI G4 pmirror_pfet_64x_flat_0/G4 VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=30e+06u
+ l=150000u
X90 VHI G8 pmirror_pfet_64x_flat_0/G8 VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=30e+06u
+ l=150000u

C0 VHI pmirror_pfet_64x_flat_0/G8 10.15fF
C1 pmirror_pfet_64x_flat_0/G16 IOUT 2.36fF
C2 pmirror_pfet_64x_flat_0/G4 VHI 4.30fF
C3 pmirror_pfet_64x_flat_0/G2 IREF 2.13fF
C4 pmirror_pfet_64x_flat_0/G16 pmirror_pfet_64x_flat_0/G8 4.66fF
C5 pmirror_pfet_64x_flat_0/G4 pmirror_pfet_64x_flat_0/G8 3.24fF
C6 pmirror_pfet_64x_flat_0/G2 VHI 4.48fF
C7 pmirror_pfet_64x_flat_0/G4 pmirror_pfet_64x_flat_0/G2 2.55fF
C8 VHI IREF 4.53fF
C9 VHI pmirror_pfet_64x_flat_0/G32 15.40fF
C10 IOUT pmirror_pfet_64x_flat_0/G32 5.39fF
C11 pmirror_pfet_64x_flat_0/G16 pmirror_pfet_64x_flat_0/G32 3.74fF
C12 VHI IOUT 24.04fF
C13 pmirror_pfet_64x_flat_0/G16 VHI 4.93fF
C14 VHI VSUBS 46.10fF


**** end user architecture code
.ends

.GLOBAL GND
.end
