magic
tech sky130B
magscale 1 2
timestamp 1668465492
<< error_p >>
rect -1037 272 -979 278
rect -845 272 -787 278
rect -653 272 -595 278
rect -461 272 -403 278
rect -269 272 -211 278
rect -77 272 -19 278
rect 115 272 173 278
rect 307 272 365 278
rect 499 272 557 278
rect 691 272 749 278
rect 883 272 941 278
rect 1075 272 1133 278
rect -1037 238 -1025 272
rect -845 238 -833 272
rect -653 238 -641 272
rect -461 238 -449 272
rect -269 238 -257 272
rect -77 238 -65 272
rect 115 238 127 272
rect 307 238 319 272
rect 499 238 511 272
rect 691 238 703 272
rect 883 238 895 272
rect 1075 238 1087 272
rect -1037 232 -979 238
rect -845 232 -787 238
rect -653 232 -595 238
rect -461 232 -403 238
rect -269 232 -211 238
rect -77 232 -19 238
rect 115 232 173 238
rect 307 232 365 238
rect 499 232 557 238
rect 691 232 749 238
rect 883 232 941 238
rect 1075 232 1133 238
rect -1133 -238 -1075 -232
rect -941 -238 -883 -232
rect -749 -238 -691 -232
rect -557 -238 -499 -232
rect -365 -238 -307 -232
rect -173 -238 -115 -232
rect 19 -238 77 -232
rect 211 -238 269 -232
rect 403 -238 461 -232
rect 595 -238 653 -232
rect 787 -238 845 -232
rect 979 -238 1037 -232
rect -1133 -272 -1121 -238
rect -941 -272 -929 -238
rect -749 -272 -737 -238
rect -557 -272 -545 -238
rect -365 -272 -353 -238
rect -173 -272 -161 -238
rect 19 -272 31 -238
rect 211 -272 223 -238
rect 403 -272 415 -238
rect 595 -272 607 -238
rect 787 -272 799 -238
rect 979 -272 991 -238
rect -1133 -278 -1075 -272
rect -941 -278 -883 -272
rect -749 -278 -691 -272
rect -557 -278 -499 -272
rect -365 -278 -307 -272
rect -173 -278 -115 -272
rect 19 -278 77 -272
rect 211 -278 269 -272
rect 403 -278 461 -272
rect 595 -278 653 -272
rect 787 -278 845 -272
rect 979 -278 1037 -272
<< pwell >>
rect -1319 -410 1319 410
<< nmos >>
rect -1119 -200 -1089 200
rect -1023 -200 -993 200
rect -927 -200 -897 200
rect -831 -200 -801 200
rect -735 -200 -705 200
rect -639 -200 -609 200
rect -543 -200 -513 200
rect -447 -200 -417 200
rect -351 -200 -321 200
rect -255 -200 -225 200
rect -159 -200 -129 200
rect -63 -200 -33 200
rect 33 -200 63 200
rect 129 -200 159 200
rect 225 -200 255 200
rect 321 -200 351 200
rect 417 -200 447 200
rect 513 -200 543 200
rect 609 -200 639 200
rect 705 -200 735 200
rect 801 -200 831 200
rect 897 -200 927 200
rect 993 -200 1023 200
rect 1089 -200 1119 200
<< ndiff >>
rect -1181 188 -1119 200
rect -1181 -188 -1169 188
rect -1135 -188 -1119 188
rect -1181 -200 -1119 -188
rect -1089 188 -1023 200
rect -1089 -188 -1073 188
rect -1039 -188 -1023 188
rect -1089 -200 -1023 -188
rect -993 188 -927 200
rect -993 -188 -977 188
rect -943 -188 -927 188
rect -993 -200 -927 -188
rect -897 188 -831 200
rect -897 -188 -881 188
rect -847 -188 -831 188
rect -897 -200 -831 -188
rect -801 188 -735 200
rect -801 -188 -785 188
rect -751 -188 -735 188
rect -801 -200 -735 -188
rect -705 188 -639 200
rect -705 -188 -689 188
rect -655 -188 -639 188
rect -705 -200 -639 -188
rect -609 188 -543 200
rect -609 -188 -593 188
rect -559 -188 -543 188
rect -609 -200 -543 -188
rect -513 188 -447 200
rect -513 -188 -497 188
rect -463 -188 -447 188
rect -513 -200 -447 -188
rect -417 188 -351 200
rect -417 -188 -401 188
rect -367 -188 -351 188
rect -417 -200 -351 -188
rect -321 188 -255 200
rect -321 -188 -305 188
rect -271 -188 -255 188
rect -321 -200 -255 -188
rect -225 188 -159 200
rect -225 -188 -209 188
rect -175 -188 -159 188
rect -225 -200 -159 -188
rect -129 188 -63 200
rect -129 -188 -113 188
rect -79 -188 -63 188
rect -129 -200 -63 -188
rect -33 188 33 200
rect -33 -188 -17 188
rect 17 -188 33 188
rect -33 -200 33 -188
rect 63 188 129 200
rect 63 -188 79 188
rect 113 -188 129 188
rect 63 -200 129 -188
rect 159 188 225 200
rect 159 -188 175 188
rect 209 -188 225 188
rect 159 -200 225 -188
rect 255 188 321 200
rect 255 -188 271 188
rect 305 -188 321 188
rect 255 -200 321 -188
rect 351 188 417 200
rect 351 -188 367 188
rect 401 -188 417 188
rect 351 -200 417 -188
rect 447 188 513 200
rect 447 -188 463 188
rect 497 -188 513 188
rect 447 -200 513 -188
rect 543 188 609 200
rect 543 -188 559 188
rect 593 -188 609 188
rect 543 -200 609 -188
rect 639 188 705 200
rect 639 -188 655 188
rect 689 -188 705 188
rect 639 -200 705 -188
rect 735 188 801 200
rect 735 -188 751 188
rect 785 -188 801 188
rect 735 -200 801 -188
rect 831 188 897 200
rect 831 -188 847 188
rect 881 -188 897 188
rect 831 -200 897 -188
rect 927 188 993 200
rect 927 -188 943 188
rect 977 -188 993 188
rect 927 -200 993 -188
rect 1023 188 1089 200
rect 1023 -188 1039 188
rect 1073 -188 1089 188
rect 1023 -200 1089 -188
rect 1119 188 1181 200
rect 1119 -188 1135 188
rect 1169 -188 1181 188
rect 1119 -200 1181 -188
<< ndiffc >>
rect -1169 -188 -1135 188
rect -1073 -188 -1039 188
rect -977 -188 -943 188
rect -881 -188 -847 188
rect -785 -188 -751 188
rect -689 -188 -655 188
rect -593 -188 -559 188
rect -497 -188 -463 188
rect -401 -188 -367 188
rect -305 -188 -271 188
rect -209 -188 -175 188
rect -113 -188 -79 188
rect -17 -188 17 188
rect 79 -188 113 188
rect 175 -188 209 188
rect 271 -188 305 188
rect 367 -188 401 188
rect 463 -188 497 188
rect 559 -188 593 188
rect 655 -188 689 188
rect 751 -188 785 188
rect 847 -188 881 188
rect 943 -188 977 188
rect 1039 -188 1073 188
rect 1135 -188 1169 188
<< psubdiff >>
rect -1283 340 -1187 374
rect 1187 340 1283 374
rect -1283 278 -1249 340
rect 1249 278 1283 340
rect -1283 -340 -1249 -278
rect 1249 -340 1283 -278
rect -1283 -374 -1187 -340
rect 1187 -374 1283 -340
<< psubdiffcont >>
rect -1187 340 1187 374
rect -1283 -278 -1249 278
rect 1249 -278 1283 278
rect -1187 -374 1187 -340
<< poly >>
rect -1041 272 -975 288
rect -1041 238 -1025 272
rect -991 238 -975 272
rect -1119 200 -1089 226
rect -1041 222 -975 238
rect -849 272 -783 288
rect -849 238 -833 272
rect -799 238 -783 272
rect -1023 200 -993 222
rect -927 200 -897 226
rect -849 222 -783 238
rect -657 272 -591 288
rect -657 238 -641 272
rect -607 238 -591 272
rect -831 200 -801 222
rect -735 200 -705 226
rect -657 222 -591 238
rect -465 272 -399 288
rect -465 238 -449 272
rect -415 238 -399 272
rect -639 200 -609 222
rect -543 200 -513 226
rect -465 222 -399 238
rect -273 272 -207 288
rect -273 238 -257 272
rect -223 238 -207 272
rect -447 200 -417 222
rect -351 200 -321 226
rect -273 222 -207 238
rect -81 272 -15 288
rect -81 238 -65 272
rect -31 238 -15 272
rect -255 200 -225 222
rect -159 200 -129 226
rect -81 222 -15 238
rect 111 272 177 288
rect 111 238 127 272
rect 161 238 177 272
rect -63 200 -33 222
rect 33 200 63 226
rect 111 222 177 238
rect 303 272 369 288
rect 303 238 319 272
rect 353 238 369 272
rect 129 200 159 222
rect 225 200 255 226
rect 303 222 369 238
rect 495 272 561 288
rect 495 238 511 272
rect 545 238 561 272
rect 321 200 351 222
rect 417 200 447 226
rect 495 222 561 238
rect 687 272 753 288
rect 687 238 703 272
rect 737 238 753 272
rect 513 200 543 222
rect 609 200 639 226
rect 687 222 753 238
rect 879 272 945 288
rect 879 238 895 272
rect 929 238 945 272
rect 705 200 735 222
rect 801 200 831 226
rect 879 222 945 238
rect 1071 272 1137 288
rect 1071 238 1087 272
rect 1121 238 1137 272
rect 897 200 927 222
rect 993 200 1023 226
rect 1071 222 1137 238
rect 1089 200 1119 222
rect -1119 -222 -1089 -200
rect -1137 -238 -1071 -222
rect -1023 -226 -993 -200
rect -927 -222 -897 -200
rect -1137 -272 -1121 -238
rect -1087 -272 -1071 -238
rect -1137 -288 -1071 -272
rect -945 -238 -879 -222
rect -831 -226 -801 -200
rect -735 -222 -705 -200
rect -945 -272 -929 -238
rect -895 -272 -879 -238
rect -945 -288 -879 -272
rect -753 -238 -687 -222
rect -639 -226 -609 -200
rect -543 -222 -513 -200
rect -753 -272 -737 -238
rect -703 -272 -687 -238
rect -753 -288 -687 -272
rect -561 -238 -495 -222
rect -447 -226 -417 -200
rect -351 -222 -321 -200
rect -561 -272 -545 -238
rect -511 -272 -495 -238
rect -561 -288 -495 -272
rect -369 -238 -303 -222
rect -255 -226 -225 -200
rect -159 -222 -129 -200
rect -369 -272 -353 -238
rect -319 -272 -303 -238
rect -369 -288 -303 -272
rect -177 -238 -111 -222
rect -63 -226 -33 -200
rect 33 -222 63 -200
rect -177 -272 -161 -238
rect -127 -272 -111 -238
rect -177 -288 -111 -272
rect 15 -238 81 -222
rect 129 -226 159 -200
rect 225 -222 255 -200
rect 15 -272 31 -238
rect 65 -272 81 -238
rect 15 -288 81 -272
rect 207 -238 273 -222
rect 321 -226 351 -200
rect 417 -222 447 -200
rect 207 -272 223 -238
rect 257 -272 273 -238
rect 207 -288 273 -272
rect 399 -238 465 -222
rect 513 -226 543 -200
rect 609 -222 639 -200
rect 399 -272 415 -238
rect 449 -272 465 -238
rect 399 -288 465 -272
rect 591 -238 657 -222
rect 705 -226 735 -200
rect 801 -222 831 -200
rect 591 -272 607 -238
rect 641 -272 657 -238
rect 591 -288 657 -272
rect 783 -238 849 -222
rect 897 -226 927 -200
rect 993 -222 1023 -200
rect 783 -272 799 -238
rect 833 -272 849 -238
rect 783 -288 849 -272
rect 975 -238 1041 -222
rect 1089 -226 1119 -200
rect 975 -272 991 -238
rect 1025 -272 1041 -238
rect 975 -288 1041 -272
<< polycont >>
rect -1025 238 -991 272
rect -833 238 -799 272
rect -641 238 -607 272
rect -449 238 -415 272
rect -257 238 -223 272
rect -65 238 -31 272
rect 127 238 161 272
rect 319 238 353 272
rect 511 238 545 272
rect 703 238 737 272
rect 895 238 929 272
rect 1087 238 1121 272
rect -1121 -272 -1087 -238
rect -929 -272 -895 -238
rect -737 -272 -703 -238
rect -545 -272 -511 -238
rect -353 -272 -319 -238
rect -161 -272 -127 -238
rect 31 -272 65 -238
rect 223 -272 257 -238
rect 415 -272 449 -238
rect 607 -272 641 -238
rect 799 -272 833 -238
rect 991 -272 1025 -238
<< locali >>
rect -1283 340 -1187 374
rect 1187 340 1283 374
rect -1283 278 -1249 340
rect 1249 278 1283 340
rect -1041 238 -1025 272
rect -991 238 -975 272
rect -849 238 -833 272
rect -799 238 -783 272
rect -657 238 -641 272
rect -607 238 -591 272
rect -465 238 -449 272
rect -415 238 -399 272
rect -273 238 -257 272
rect -223 238 -207 272
rect -81 238 -65 272
rect -31 238 -15 272
rect 111 238 127 272
rect 161 238 177 272
rect 303 238 319 272
rect 353 238 369 272
rect 495 238 511 272
rect 545 238 561 272
rect 687 238 703 272
rect 737 238 753 272
rect 879 238 895 272
rect 929 238 945 272
rect 1071 238 1087 272
rect 1121 238 1137 272
rect -1169 188 -1135 204
rect -1169 -204 -1135 -188
rect -1073 188 -1039 204
rect -1073 -204 -1039 -188
rect -977 188 -943 204
rect -977 -204 -943 -188
rect -881 188 -847 204
rect -881 -204 -847 -188
rect -785 188 -751 204
rect -785 -204 -751 -188
rect -689 188 -655 204
rect -689 -204 -655 -188
rect -593 188 -559 204
rect -593 -204 -559 -188
rect -497 188 -463 204
rect -497 -204 -463 -188
rect -401 188 -367 204
rect -401 -204 -367 -188
rect -305 188 -271 204
rect -305 -204 -271 -188
rect -209 188 -175 204
rect -209 -204 -175 -188
rect -113 188 -79 204
rect -113 -204 -79 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 79 188 113 204
rect 79 -204 113 -188
rect 175 188 209 204
rect 175 -204 209 -188
rect 271 188 305 204
rect 271 -204 305 -188
rect 367 188 401 204
rect 367 -204 401 -188
rect 463 188 497 204
rect 463 -204 497 -188
rect 559 188 593 204
rect 559 -204 593 -188
rect 655 188 689 204
rect 655 -204 689 -188
rect 751 188 785 204
rect 751 -204 785 -188
rect 847 188 881 204
rect 847 -204 881 -188
rect 943 188 977 204
rect 943 -204 977 -188
rect 1039 188 1073 204
rect 1039 -204 1073 -188
rect 1135 188 1169 204
rect 1135 -204 1169 -188
rect -1137 -272 -1121 -238
rect -1087 -272 -1071 -238
rect -945 -272 -929 -238
rect -895 -272 -879 -238
rect -753 -272 -737 -238
rect -703 -272 -687 -238
rect -561 -272 -545 -238
rect -511 -272 -495 -238
rect -369 -272 -353 -238
rect -319 -272 -303 -238
rect -177 -272 -161 -238
rect -127 -272 -111 -238
rect 15 -272 31 -238
rect 65 -272 81 -238
rect 207 -272 223 -238
rect 257 -272 273 -238
rect 399 -272 415 -238
rect 449 -272 465 -238
rect 591 -272 607 -238
rect 641 -272 657 -238
rect 783 -272 799 -238
rect 833 -272 849 -238
rect 975 -272 991 -238
rect 1025 -272 1041 -238
rect -1283 -340 -1249 -278
rect 1249 -340 1283 -278
rect -1283 -374 -1187 -340
rect 1187 -374 1283 -340
<< viali >>
rect -1025 238 -991 272
rect -833 238 -799 272
rect -641 238 -607 272
rect -449 238 -415 272
rect -257 238 -223 272
rect -65 238 -31 272
rect 127 238 161 272
rect 319 238 353 272
rect 511 238 545 272
rect 703 238 737 272
rect 895 238 929 272
rect 1087 238 1121 272
rect -1169 -188 -1135 188
rect -1073 -188 -1039 188
rect -977 -188 -943 188
rect -881 -188 -847 188
rect -785 -188 -751 188
rect -689 -188 -655 188
rect -593 -188 -559 188
rect -497 -188 -463 188
rect -401 -188 -367 188
rect -305 -188 -271 188
rect -209 -188 -175 188
rect -113 -188 -79 188
rect -17 -188 17 188
rect 79 -188 113 188
rect 175 -188 209 188
rect 271 -188 305 188
rect 367 -188 401 188
rect 463 -188 497 188
rect 559 -188 593 188
rect 655 -188 689 188
rect 751 -188 785 188
rect 847 -188 881 188
rect 943 -188 977 188
rect 1039 -188 1073 188
rect 1135 -188 1169 188
rect -1121 -272 -1087 -238
rect -929 -272 -895 -238
rect -737 -272 -703 -238
rect -545 -272 -511 -238
rect -353 -272 -319 -238
rect -161 -272 -127 -238
rect 31 -272 65 -238
rect 223 -272 257 -238
rect 415 -272 449 -238
rect 607 -272 641 -238
rect 799 -272 833 -238
rect 991 -272 1025 -238
<< metal1 >>
rect -1037 272 -979 278
rect -1037 238 -1025 272
rect -991 238 -979 272
rect -1037 232 -979 238
rect -845 272 -787 278
rect -845 238 -833 272
rect -799 238 -787 272
rect -845 232 -787 238
rect -653 272 -595 278
rect -653 238 -641 272
rect -607 238 -595 272
rect -653 232 -595 238
rect -461 272 -403 278
rect -461 238 -449 272
rect -415 238 -403 272
rect -461 232 -403 238
rect -269 272 -211 278
rect -269 238 -257 272
rect -223 238 -211 272
rect -269 232 -211 238
rect -77 272 -19 278
rect -77 238 -65 272
rect -31 238 -19 272
rect -77 232 -19 238
rect 115 272 173 278
rect 115 238 127 272
rect 161 238 173 272
rect 115 232 173 238
rect 307 272 365 278
rect 307 238 319 272
rect 353 238 365 272
rect 307 232 365 238
rect 499 272 557 278
rect 499 238 511 272
rect 545 238 557 272
rect 499 232 557 238
rect 691 272 749 278
rect 691 238 703 272
rect 737 238 749 272
rect 691 232 749 238
rect 883 272 941 278
rect 883 238 895 272
rect 929 238 941 272
rect 883 232 941 238
rect 1075 272 1133 278
rect 1075 238 1087 272
rect 1121 238 1133 272
rect 1075 232 1133 238
rect -1175 188 -1129 200
rect -1175 -188 -1169 188
rect -1135 -188 -1129 188
rect -1175 -200 -1129 -188
rect -1079 188 -1033 200
rect -1079 -188 -1073 188
rect -1039 -188 -1033 188
rect -1079 -200 -1033 -188
rect -983 188 -937 200
rect -983 -188 -977 188
rect -943 -188 -937 188
rect -983 -200 -937 -188
rect -887 188 -841 200
rect -887 -188 -881 188
rect -847 -188 -841 188
rect -887 -200 -841 -188
rect -791 188 -745 200
rect -791 -188 -785 188
rect -751 -188 -745 188
rect -791 -200 -745 -188
rect -695 188 -649 200
rect -695 -188 -689 188
rect -655 -188 -649 188
rect -695 -200 -649 -188
rect -599 188 -553 200
rect -599 -188 -593 188
rect -559 -188 -553 188
rect -599 -200 -553 -188
rect -503 188 -457 200
rect -503 -188 -497 188
rect -463 -188 -457 188
rect -503 -200 -457 -188
rect -407 188 -361 200
rect -407 -188 -401 188
rect -367 -188 -361 188
rect -407 -200 -361 -188
rect -311 188 -265 200
rect -311 -188 -305 188
rect -271 -188 -265 188
rect -311 -200 -265 -188
rect -215 188 -169 200
rect -215 -188 -209 188
rect -175 -188 -169 188
rect -215 -200 -169 -188
rect -119 188 -73 200
rect -119 -188 -113 188
rect -79 -188 -73 188
rect -119 -200 -73 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 73 188 119 200
rect 73 -188 79 188
rect 113 -188 119 188
rect 73 -200 119 -188
rect 169 188 215 200
rect 169 -188 175 188
rect 209 -188 215 188
rect 169 -200 215 -188
rect 265 188 311 200
rect 265 -188 271 188
rect 305 -188 311 188
rect 265 -200 311 -188
rect 361 188 407 200
rect 361 -188 367 188
rect 401 -188 407 188
rect 361 -200 407 -188
rect 457 188 503 200
rect 457 -188 463 188
rect 497 -188 503 188
rect 457 -200 503 -188
rect 553 188 599 200
rect 553 -188 559 188
rect 593 -188 599 188
rect 553 -200 599 -188
rect 649 188 695 200
rect 649 -188 655 188
rect 689 -188 695 188
rect 649 -200 695 -188
rect 745 188 791 200
rect 745 -188 751 188
rect 785 -188 791 188
rect 745 -200 791 -188
rect 841 188 887 200
rect 841 -188 847 188
rect 881 -188 887 188
rect 841 -200 887 -188
rect 937 188 983 200
rect 937 -188 943 188
rect 977 -188 983 188
rect 937 -200 983 -188
rect 1033 188 1079 200
rect 1033 -188 1039 188
rect 1073 -188 1079 188
rect 1033 -200 1079 -188
rect 1129 188 1175 200
rect 1129 -188 1135 188
rect 1169 -188 1175 188
rect 1129 -200 1175 -188
rect -1133 -238 -1075 -232
rect -1133 -272 -1121 -238
rect -1087 -272 -1075 -238
rect -1133 -278 -1075 -272
rect -941 -238 -883 -232
rect -941 -272 -929 -238
rect -895 -272 -883 -238
rect -941 -278 -883 -272
rect -749 -238 -691 -232
rect -749 -272 -737 -238
rect -703 -272 -691 -238
rect -749 -278 -691 -272
rect -557 -238 -499 -232
rect -557 -272 -545 -238
rect -511 -272 -499 -238
rect -557 -278 -499 -272
rect -365 -238 -307 -232
rect -365 -272 -353 -238
rect -319 -272 -307 -238
rect -365 -278 -307 -272
rect -173 -238 -115 -232
rect -173 -272 -161 -238
rect -127 -272 -115 -238
rect -173 -278 -115 -272
rect 19 -238 77 -232
rect 19 -272 31 -238
rect 65 -272 77 -238
rect 19 -278 77 -272
rect 211 -238 269 -232
rect 211 -272 223 -238
rect 257 -272 269 -238
rect 211 -278 269 -272
rect 403 -238 461 -232
rect 403 -272 415 -238
rect 449 -272 461 -238
rect 403 -278 461 -272
rect 595 -238 653 -232
rect 595 -272 607 -238
rect 641 -272 653 -238
rect 595 -278 653 -272
rect 787 -238 845 -232
rect 787 -272 799 -238
rect 833 -272 845 -238
rect 787 -278 845 -272
rect 979 -238 1037 -232
rect 979 -272 991 -238
rect 1025 -272 1037 -238
rect 979 -278 1037 -272
<< properties >>
string FIXED_BBOX -1266 -357 1266 357
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 0.150 m 1 nf 24 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
