magic
tech sky130A
magscale 1 2
timestamp 1672168347
<< nwell >>
rect 3898 1418 6064 3856
<< pwell >>
rect 3897 -3 6063 1417
<< nmos >>
rect 4093 207 4493 1207
rect 4551 207 4951 1207
rect 5009 207 5409 1207
rect 5467 207 5867 1207
<< pmos >>
rect 4094 1637 4494 3637
rect 4552 1637 4952 3637
rect 5010 1637 5410 3637
rect 5468 1637 5868 3637
<< ndiff >>
rect 4035 1195 4093 1207
rect 4035 219 4047 1195
rect 4081 219 4093 1195
rect 4035 207 4093 219
rect 4493 1195 4551 1207
rect 4493 219 4505 1195
rect 4539 219 4551 1195
rect 4493 207 4551 219
rect 4951 1195 5009 1207
rect 4951 219 4963 1195
rect 4997 219 5009 1195
rect 4951 207 5009 219
rect 5409 1195 5467 1207
rect 5409 219 5421 1195
rect 5455 219 5467 1195
rect 5409 207 5467 219
rect 5867 1195 5925 1207
rect 5867 219 5879 1195
rect 5913 219 5925 1195
rect 5867 207 5925 219
<< pdiff >>
rect 4036 3625 4094 3637
rect 4036 1649 4048 3625
rect 4082 1649 4094 3625
rect 4036 1637 4094 1649
rect 4494 3625 4552 3637
rect 4494 1649 4506 3625
rect 4540 1649 4552 3625
rect 4494 1637 4552 1649
rect 4952 3625 5010 3637
rect 4952 1649 4964 3625
rect 4998 1649 5010 3625
rect 4952 1637 5010 1649
rect 5410 3625 5468 3637
rect 5410 1649 5422 3625
rect 5456 1649 5468 3625
rect 5410 1637 5468 1649
rect 5868 3625 5926 3637
rect 5868 1649 5880 3625
rect 5914 1649 5926 3625
rect 5868 1637 5926 1649
<< ndiffc >>
rect 4047 219 4081 1195
rect 4505 219 4539 1195
rect 4963 219 4997 1195
rect 5421 219 5455 1195
rect 5879 219 5913 1195
<< pdiffc >>
rect 4048 1649 4082 3625
rect 4506 1649 4540 3625
rect 4964 1649 4998 3625
rect 5422 1649 5456 3625
rect 5880 1649 5914 3625
<< psubdiff >>
rect 3933 1347 4029 1381
rect 5931 1347 6027 1381
rect 3933 1285 3967 1347
rect 5993 1285 6027 1347
rect 3933 67 3967 129
rect 5993 67 6027 129
rect 3933 33 4029 67
rect 5931 33 6027 67
<< nsubdiff >>
rect 3934 3786 4030 3820
rect 5932 3786 6028 3820
rect 3934 3724 3968 3786
rect 5994 3724 6028 3786
rect 3934 1488 3968 1550
rect 5994 1488 6028 1550
rect 3934 1454 4030 1488
rect 5932 1454 6028 1488
<< psubdiffcont >>
rect 4029 1347 5931 1381
rect 3933 129 3967 1285
rect 5993 129 6027 1285
rect 4029 33 5931 67
<< nsubdiffcont >>
rect 4030 3786 5932 3820
rect 3934 1550 3968 3724
rect 5994 1550 6028 3724
rect 4030 1454 5932 1488
<< poly >>
rect 4094 3718 4494 3734
rect 4094 3684 4110 3718
rect 4478 3684 4494 3718
rect 4094 3637 4494 3684
rect 4552 3718 4952 3734
rect 4552 3684 4568 3718
rect 4936 3684 4952 3718
rect 4552 3637 4952 3684
rect 5010 3718 5410 3734
rect 5010 3684 5026 3718
rect 5394 3684 5410 3718
rect 5010 3637 5410 3684
rect 5468 3718 5868 3734
rect 5468 3684 5484 3718
rect 5852 3684 5868 3718
rect 5468 3637 5868 3684
rect 4094 1590 4494 1637
rect 4094 1556 4110 1590
rect 4478 1556 4494 1590
rect 4094 1540 4494 1556
rect 4552 1590 4952 1637
rect 4552 1556 4568 1590
rect 4936 1556 4952 1590
rect 4552 1540 4952 1556
rect 5010 1590 5410 1637
rect 5010 1556 5026 1590
rect 5394 1556 5410 1590
rect 5010 1540 5410 1556
rect 5468 1590 5868 1637
rect 5468 1556 5484 1590
rect 5852 1556 5868 1590
rect 5468 1540 5868 1556
rect 4093 1279 4493 1295
rect 4093 1245 4109 1279
rect 4477 1245 4493 1279
rect 4093 1207 4493 1245
rect 4551 1279 4951 1295
rect 4551 1245 4567 1279
rect 4935 1245 4951 1279
rect 4551 1207 4951 1245
rect 5009 1279 5409 1295
rect 5009 1245 5025 1279
rect 5393 1245 5409 1279
rect 5009 1207 5409 1245
rect 5467 1279 5867 1295
rect 5467 1245 5483 1279
rect 5851 1245 5867 1279
rect 5467 1207 5867 1245
rect 4093 169 4493 207
rect 4093 135 4109 169
rect 4477 135 4493 169
rect 4093 119 4493 135
rect 4551 169 4951 207
rect 4551 135 4567 169
rect 4835 135 4951 169
rect 4551 119 4951 135
rect 5009 169 5409 207
rect 5009 135 5125 169
rect 5393 135 5409 169
rect 5009 119 5409 135
rect 5467 169 5867 207
rect 5467 135 5483 169
rect 5851 135 5867 169
rect 5467 119 5867 135
<< polycont >>
rect 4110 3684 4478 3718
rect 4568 3684 4936 3718
rect 5026 3684 5394 3718
rect 5484 3684 5852 3718
rect 4110 1556 4478 1590
rect 4568 1556 4936 1590
rect 5026 1556 5394 1590
rect 5484 1556 5852 1590
rect 4109 1245 4477 1279
rect 4567 1245 4935 1279
rect 5025 1245 5393 1279
rect 5483 1245 5851 1279
rect 4109 135 4477 169
rect 4567 135 4835 169
rect 5125 135 5393 169
rect 5483 135 5851 169
<< locali >>
rect 3960 3860 6020 3880
rect 3960 3820 4000 3860
rect 5980 3820 6020 3860
rect 3934 3786 4030 3820
rect 5932 3786 6028 3820
rect 3934 3724 3968 3786
rect 5994 3724 6028 3786
rect 4094 3684 4110 3718
rect 4478 3684 4494 3718
rect 4552 3684 4568 3718
rect 4936 3684 4952 3718
rect 5010 3684 5026 3718
rect 5394 3684 5410 3718
rect 5468 3684 5484 3718
rect 5852 3684 5868 3718
rect 4048 3625 4082 3641
rect 4048 1633 4082 1649
rect 4506 3625 4540 3641
rect 4506 1633 4540 1649
rect 4964 3625 4998 3641
rect 4964 1633 4998 1649
rect 5422 3625 5456 3641
rect 5422 1633 5456 1649
rect 5880 3625 5914 3641
rect 5880 1633 5914 1649
rect 4094 1556 4110 1590
rect 4478 1556 4494 1590
rect 4552 1556 4568 1590
rect 4936 1556 4952 1590
rect 5010 1556 5026 1590
rect 5394 1556 5410 1590
rect 5468 1556 5484 1590
rect 5852 1556 5868 1590
rect 3934 1488 3968 1550
rect 5994 1488 6028 1550
rect 3934 1454 4030 1488
rect 5932 1454 6028 1488
rect 3933 1347 4029 1381
rect 5931 1347 6027 1381
rect 3933 1285 3967 1347
rect 3933 67 3967 129
rect 4047 1279 4081 1347
rect 5879 1279 5913 1347
rect 4047 1245 4109 1279
rect 4477 1245 4493 1279
rect 4551 1245 4567 1279
rect 4935 1245 4951 1279
rect 5009 1245 5025 1279
rect 5393 1245 5409 1279
rect 5467 1245 5483 1279
rect 5851 1245 5913 1279
rect 4047 1195 4081 1245
rect 4047 169 4081 219
rect 4505 1195 4539 1211
rect 4505 203 4539 219
rect 4963 1195 4997 1211
rect 4047 135 4109 169
rect 4477 135 4493 169
rect 4551 135 4567 169
rect 4835 135 4851 169
rect 4047 67 4081 135
rect 4963 67 4997 219
rect 5421 1195 5455 1211
rect 5421 203 5455 219
rect 5879 1195 5913 1245
rect 5879 169 5913 219
rect 5109 135 5125 169
rect 5393 135 5409 169
rect 5467 135 5483 169
rect 5851 135 5913 169
rect 5879 67 5913 135
rect 5993 1285 6027 1347
rect 5993 67 6027 129
rect 3933 40 4029 67
rect 5931 40 6027 67
rect 3933 33 4000 40
rect 5960 33 6027 40
rect 3960 0 4000 33
rect 5960 0 6000 33
rect 3960 -20 6000 0
<< viali >>
rect 4000 3820 5980 3860
rect 4110 3684 4478 3718
rect 4568 3684 4936 3718
rect 5026 3684 5394 3718
rect 5484 3684 5852 3718
rect 4048 1649 4082 3625
rect 4506 1649 4540 3625
rect 4964 1649 4998 3625
rect 5422 1649 5456 3625
rect 5880 1649 5914 3625
rect 4110 1556 4478 1590
rect 4568 1556 4936 1590
rect 5026 1556 5394 1590
rect 5484 1556 5852 1590
rect 4109 1245 4477 1279
rect 4567 1245 4935 1279
rect 5025 1245 5393 1279
rect 5483 1245 5851 1279
rect 4047 219 4081 1195
rect 4505 219 4539 1195
rect 4963 219 4997 1195
rect 4109 135 4477 169
rect 4567 135 4835 169
rect 5421 219 5455 1195
rect 5879 219 5913 1195
rect 5125 135 5393 169
rect 5483 135 5851 169
rect 4000 33 4029 40
rect 4029 33 5931 40
rect 5931 33 5960 40
rect 4000 0 5960 33
<< metal1 >>
rect 3960 3800 4000 3880
rect 5980 3800 6020 3880
rect 4098 3718 4490 3724
rect 4098 3684 4110 3718
rect 4478 3684 4490 3718
rect 4098 3678 4490 3684
rect 4556 3718 4948 3724
rect 4556 3684 4568 3718
rect 4936 3684 4948 3718
rect 4556 3678 4948 3684
rect 5014 3718 5406 3724
rect 5014 3684 5026 3718
rect 5394 3684 5406 3718
rect 5014 3678 5406 3684
rect 5472 3718 5864 3724
rect 5472 3684 5484 3718
rect 5852 3684 5864 3718
rect 5472 3678 5864 3684
rect 4042 3625 4088 3637
rect 4042 1649 4048 3625
rect 4082 1649 4088 3625
rect 4042 1637 4088 1649
rect 4497 3625 4549 3637
rect 4955 3625 5007 3637
rect 4549 1649 4607 1695
rect 4497 1637 4607 1649
rect 4955 1637 5007 1649
rect 5413 3625 5465 3637
rect 5413 1637 5465 1649
rect 5874 3625 5920 3637
rect 5874 1649 5880 3625
rect 5914 1649 5920 3625
rect 5874 1637 5920 1649
rect 4552 1596 4607 1637
rect 4098 1590 4490 1596
rect 4098 1556 4110 1590
rect 4478 1556 4490 1590
rect 4552 1590 5406 1596
rect 4552 1556 4568 1590
rect 4936 1556 5026 1590
rect 5394 1556 5406 1590
rect 4098 1550 4490 1556
rect 4556 1550 5406 1556
rect 5472 1590 5864 1596
rect 5472 1556 5484 1590
rect 5852 1556 5864 1590
rect 5472 1550 5864 1556
rect 3940 1440 4260 1460
rect 3940 1360 3960 1440
rect 4240 1420 4260 1440
rect 4240 1360 4920 1420
rect 5520 1406 5540 1440
rect 3940 1332 4920 1360
rect 5349 1345 5540 1406
rect 3940 1320 4946 1332
rect 4555 1285 4946 1320
rect 5349 1285 5410 1345
rect 5520 1340 5540 1345
rect 5920 1340 5940 1440
rect 4097 1279 4489 1285
rect 4097 1245 4109 1279
rect 4477 1245 4489 1279
rect 4097 1239 4489 1245
rect 4555 1279 4947 1285
rect 4555 1245 4567 1279
rect 4935 1245 4947 1279
rect 4555 1239 4947 1245
rect 5013 1279 5410 1285
rect 5013 1245 5025 1279
rect 5393 1245 5410 1279
rect 5013 1239 5410 1245
rect 5471 1279 5863 1285
rect 5471 1245 5483 1279
rect 5851 1245 5863 1279
rect 5471 1239 5863 1245
rect 5349 1207 5410 1239
rect 4041 1195 4087 1207
rect 4041 219 4047 1195
rect 4081 219 4087 1195
rect 4041 207 4087 219
rect 4496 1195 4548 1207
rect 4496 207 4548 219
rect 4954 1195 5006 1207
rect 5349 1195 5464 1207
rect 5349 1146 5412 1195
rect 4954 207 5006 219
rect 5412 207 5464 219
rect 5873 1195 5919 1207
rect 5873 219 5879 1195
rect 5913 219 5919 1195
rect 5873 207 5919 219
rect 4097 169 4489 175
rect 4097 135 4109 169
rect 4477 135 4489 169
rect 4097 129 4489 135
rect 4555 169 4847 175
rect 4555 135 4567 169
rect 4835 135 4847 169
rect 4555 129 4847 135
rect 5113 169 5405 175
rect 5113 135 5125 169
rect 5393 135 5405 169
rect 5113 129 5405 135
rect 5471 169 5863 175
rect 5471 135 5483 169
rect 5851 135 5863 169
rect 5471 129 5863 135
rect 3960 -20 4000 60
rect 5960 -20 6000 60
<< via1 >>
rect 4000 3860 5980 3880
rect 4000 3820 5980 3860
rect 4000 3800 5980 3820
rect 4497 1649 4506 3625
rect 4506 1649 4540 3625
rect 4540 1649 4549 3625
rect 4955 1649 4964 3625
rect 4964 1649 4998 3625
rect 4998 1649 5007 3625
rect 5413 1649 5422 3625
rect 5422 1649 5456 3625
rect 5456 1649 5465 3625
rect 3960 1360 4240 1440
rect 5540 1340 5920 1440
rect 4496 219 4505 1195
rect 4505 219 4539 1195
rect 4539 219 4548 1195
rect 4954 219 4963 1195
rect 4963 219 4997 1195
rect 4997 219 5006 1195
rect 5412 219 5421 1195
rect 5421 219 5455 1195
rect 5455 219 5464 1195
rect 4000 40 5960 60
rect 4000 0 5960 40
rect 4000 -20 5960 0
<< metal2 >>
rect 3960 3800 4000 3880
rect 5980 3800 6020 3880
rect 4497 3625 4549 3637
rect 4496 1649 4497 3188
rect 4496 1637 4549 1649
rect 4955 3625 5007 3800
rect 5413 3625 5465 3637
rect 4955 1637 5007 1649
rect 5412 1649 5413 1659
rect 5412 1637 5465 1649
rect 3900 1440 4260 1460
rect 3900 1360 3960 1440
rect 4240 1360 4260 1440
rect 3900 1340 4260 1360
rect 3900 1320 3960 1340
rect 4496 1195 4548 1637
rect 4496 207 4548 219
rect 4954 1195 5006 1207
rect 4954 60 5006 219
rect 5412 1195 5464 1637
rect 5520 1340 5540 1440
rect 5920 1340 5940 1440
rect 5412 207 5464 219
rect 3960 -20 4000 60
rect 5960 -20 6000 60
<< labels >>
rlabel metal2 5920 1340 5940 1440 1 OUT
port 2 n
rlabel metal2 3960 3800 4000 3880 1 VHI
port 3 n
rlabel metal2 3960 -20 4000 60 1 VLO
port 4 n
rlabel metal2 3900 1320 3960 1460 1 IN
<< end >>
