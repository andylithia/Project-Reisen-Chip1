magic
tech sky130A
magscale 1 2
timestamp 1672465491
<< nwell >>
rect 4180 -758 4706 609
<< pwell >>
rect 4180 609 4706 2657
<< nmos >>
rect 4380 819 4410 1319
rect 4476 819 4506 1319
<< pmos >>
rect 4380 -610 4410 390
rect 4476 -610 4506 390
<< ndiff >>
rect 4318 1307 4380 1319
rect 4318 831 4330 1307
rect 4364 831 4380 1307
rect 4318 819 4380 831
rect 4410 1307 4476 1319
rect 4410 831 4426 1307
rect 4460 831 4476 1307
rect 4410 819 4476 831
rect 4506 1307 4568 1319
rect 4506 831 4522 1307
rect 4556 831 4568 1307
rect 4506 819 4568 831
<< pdiff >>
rect 4318 378 4380 390
rect 4318 -598 4330 378
rect 4364 -598 4380 378
rect 4318 -610 4380 -598
rect 4410 378 4476 390
rect 4410 -598 4426 378
rect 4460 -598 4476 378
rect 4410 -610 4476 -598
rect 4506 378 4568 390
rect 4506 -598 4522 378
rect 4556 -598 4568 378
rect 4506 -610 4568 -598
<< ndiffc >>
rect 4330 831 4364 1307
rect 4426 831 4460 1307
rect 4522 831 4556 1307
<< pdiffc >>
rect 4330 -598 4364 378
rect 4426 -598 4460 378
rect 4522 -598 4556 378
<< psubdiff >>
rect 4216 2587 4312 2621
rect 4518 2587 4670 2621
rect 4216 2525 4250 2587
rect 4580 1431 4670 2587
rect 4250 1397 4670 1431
rect 4216 679 4250 741
rect 4636 679 4670 1397
rect 4216 645 4312 679
rect 4574 645 4670 679
<< nsubdiff >>
rect 4216 539 4312 573
rect 4574 539 4670 573
rect 4216 477 4250 539
rect 4216 -688 4250 -626
rect 4636 -688 4670 539
rect 4216 -722 4312 -688
rect 4515 -722 4670 -688
<< psubdiffcont >>
rect 4312 2587 4518 2621
rect 4216 741 4250 2525
rect 4312 645 4574 679
<< nsubdiffcont >>
rect 4312 539 4574 573
rect 4216 -626 4250 477
rect 4312 -722 4515 -688
<< poly >>
rect 4380 1319 4410 1345
rect 4476 1319 4506 1345
rect 4380 797 4410 819
rect 4476 797 4506 819
rect 4362 781 4524 797
rect 4362 747 4378 781
rect 4508 747 4524 781
rect 4362 731 4524 747
rect 4362 471 4524 487
rect 4362 437 4378 471
rect 4508 437 4524 471
rect 4362 421 4524 437
rect 4380 390 4410 421
rect 4476 390 4506 421
rect 4380 -636 4410 -610
rect 4476 -636 4506 -610
<< polycont >>
rect 4378 747 4508 781
rect 4378 437 4508 471
<< xpolycontact >>
rect 4346 2059 4484 2491
rect 4346 1527 4484 1959
<< ppolyres >>
rect 4346 1959 4484 2059
<< locali >>
rect 4216 2621 4287 2658
rect 4216 2587 4312 2621
rect 4518 2587 4580 2621
rect 4216 2574 4287 2587
rect 4216 2525 4229 2574
rect 4274 1319 4287 2574
rect 4330 1319 4364 1323
rect 4274 1313 4364 1319
rect 4292 1307 4364 1313
rect 4292 1224 4330 1307
rect 4274 1217 4330 1224
rect 4274 991 4287 1217
rect 4250 944 4287 991
rect 4330 815 4364 831
rect 4426 1307 4460 1323
rect 4426 815 4460 831
rect 4522 1307 4556 1323
rect 4522 815 4556 831
rect 4362 747 4378 781
rect 4508 747 4524 781
rect 4216 679 4250 741
rect 4216 645 4312 679
rect 4574 645 4670 679
rect 4216 539 4312 573
rect 4574 539 4670 573
rect 4216 477 4250 539
rect 4362 437 4378 471
rect 4508 437 4524 471
rect 4330 378 4364 394
rect 4330 -614 4364 -598
rect 4426 378 4460 394
rect 4426 -614 4460 -598
rect 4522 378 4556 394
rect 4522 -614 4556 -598
rect 4216 -688 4250 -626
rect 4216 -722 4312 -688
rect 4515 -722 4670 -688
rect 4337 -736 4547 -722
rect 4337 -776 4357 -736
rect 4527 -776 4547 -736
rect 4337 -796 4547 -776
<< viali >>
rect 4229 2525 4274 2574
rect 4229 991 4250 2525
rect 4250 1313 4274 2525
rect 4362 2076 4468 2473
rect 4362 1545 4468 1942
rect 4250 1224 4292 1313
rect 4250 991 4274 1224
rect 4330 831 4364 1307
rect 4426 831 4460 1307
rect 4522 831 4556 1307
rect 4378 747 4508 781
rect 4378 437 4508 471
rect 4330 -598 4364 378
rect 4426 -598 4460 378
rect 4522 -598 4556 378
rect 4357 -776 4527 -736
<< metal1 >>
rect 4216 2574 4287 2658
rect 4216 991 4225 2574
rect 4277 1319 4287 2574
rect 4356 2473 4474 2485
rect 4356 2076 4362 2473
rect 4468 2076 4474 2473
rect 4356 2064 4474 2076
rect 4346 1942 4484 1959
rect 4346 1545 4362 1942
rect 4468 1545 4484 1942
rect 4346 1527 4484 1545
rect 4277 1313 4373 1319
rect 4292 1307 4373 1313
rect 4292 1224 4321 1307
rect 4277 1217 4321 1224
rect 4277 991 4287 1217
rect 4216 944 4287 991
rect 4321 819 4373 831
rect 4417 1307 4469 1319
rect 4417 819 4469 831
rect 4513 1307 4565 1319
rect 4513 819 4565 831
rect 4173 781 4520 787
rect 4173 747 4378 781
rect 4508 747 4520 781
rect 4173 741 4520 747
rect 4173 -920 4219 741
rect 4247 471 4520 477
rect 4247 437 4378 471
rect 4508 437 4520 471
rect 4247 431 4520 437
rect 4247 -850 4293 431
rect 4321 378 4373 390
rect 4321 -610 4373 -598
rect 4417 378 4469 390
rect 4417 -610 4469 -598
rect 4513 378 4565 390
rect 4513 -610 4565 -598
rect 4337 -726 4547 -716
rect 4337 -786 4347 -726
rect 4537 -786 4547 -726
rect 4337 -796 4547 -786
rect 4247 -870 4610 -850
rect 4247 -890 4540 -870
rect 4173 -930 4380 -920
rect 4173 -960 4310 -930
rect 4540 -960 4610 -950
rect 4310 -1020 4380 -1010
<< via1 >>
rect 4225 991 4229 2574
rect 4229 1313 4274 2574
rect 4274 1313 4277 2574
rect 4362 2076 4468 2473
rect 4362 1545 4468 1942
rect 4229 1224 4292 1313
rect 4229 991 4274 1224
rect 4274 991 4277 1224
rect 4321 831 4330 1307
rect 4330 831 4364 1307
rect 4364 831 4373 1307
rect 4417 831 4426 1307
rect 4426 831 4460 1307
rect 4460 831 4469 1307
rect 4513 831 4522 1307
rect 4522 831 4556 1307
rect 4556 831 4565 1307
rect 4321 -598 4330 378
rect 4330 -598 4364 378
rect 4364 -598 4373 378
rect 4417 -598 4426 378
rect 4426 -598 4460 378
rect 4460 -598 4469 378
rect 4513 -598 4522 378
rect 4522 -598 4556 378
rect 4556 -598 4565 378
rect 4347 -736 4537 -726
rect 4347 -776 4357 -736
rect 4357 -776 4527 -736
rect 4527 -776 4537 -736
rect 4347 -786 4537 -776
rect 4310 -1010 4380 -930
rect 4540 -950 4610 -870
<< metal2 >>
rect 4250 2658 4280 2670
rect 4216 2574 4287 2658
rect 4216 991 4225 2574
rect 4277 1319 4287 2574
rect 4346 2473 4484 2491
rect 4346 2076 4362 2473
rect 4468 2076 4484 2473
rect 4346 2059 4484 2076
rect 4346 1942 4484 1959
rect 4346 1545 4362 1942
rect 4468 1545 4484 1942
rect 4346 1527 4484 1545
rect 4277 1313 4373 1319
rect 4364 1307 4373 1313
rect 4277 1217 4321 1223
rect 4277 991 4287 1217
rect 4216 944 4287 991
rect 4321 378 4373 831
rect 4321 -638 4373 -598
rect 4417 1307 4469 1527
rect 4417 378 4469 831
rect 4417 -610 4469 -598
rect 4513 1313 4670 1319
rect 4513 1307 4522 1313
rect 4586 1223 4670 1313
rect 4565 1217 4670 1223
rect 4513 378 4565 831
rect 4513 -638 4565 -598
rect 4321 -690 4565 -638
rect 4337 -786 4347 -726
rect 4537 -786 4547 -726
rect 4337 -796 4547 -786
rect 4540 -870 4610 -860
rect 4310 -930 4380 -920
rect 4310 -1030 4380 -1010
rect 4540 -1030 4610 -950
<< via2 >>
rect 4362 2076 4468 2473
rect 4250 1224 4292 1313
rect 4292 1307 4364 1313
rect 4292 1224 4321 1307
rect 4250 1223 4277 1224
rect 4277 1223 4321 1224
rect 4321 1223 4364 1307
rect 4522 1307 4586 1313
rect 4522 1223 4565 1307
rect 4565 1223 4586 1307
rect 4347 -786 4537 -726
<< metal3 >>
rect 4346 2473 4484 2491
rect 4346 2440 4362 2473
rect 4190 2380 4362 2440
rect 4330 2340 4362 2380
rect 4346 2076 4362 2340
rect 4468 2440 4484 2473
rect 4468 2340 4670 2440
rect 4468 2076 4484 2340
rect 4346 2059 4484 2076
rect 4216 1313 4670 1319
rect 4216 1223 4250 1313
rect 4364 1223 4522 1313
rect 4586 1223 4670 1313
rect 4216 1217 4670 1223
rect 4337 -786 4347 -716
rect 4537 -786 4547 -716
rect 4337 -796 4547 -786
<< via3 >>
rect 4347 -726 4537 -716
rect 4347 -786 4537 -726
<< metal4 >>
rect 4216 2650 4287 2658
rect 4200 2580 4287 2650
rect 4216 -656 4287 2580
rect 4216 -702 4297 -656
rect 4216 -706 4308 -702
rect 4216 -716 4567 -706
rect 4216 -722 4347 -716
rect 4227 -786 4347 -722
rect 4537 -786 4567 -716
rect 4227 -796 4567 -786
<< labels >>
rlabel metal2 4310 -1030 4380 -1020 1 S
port 4 n
rlabel metal2 4540 -1030 4610 -1020 1 SBAR
port 5 n
rlabel metal4 4200 2580 4210 2650 1 VHI
port 3 n
rlabel metal2 4250 2660 4280 2670 5 VLO
port 2 s
rlabel metal3 4650 2340 4670 2440 1 IO
port 1 n
rlabel metal2 4430 1360 4460 1420 1 SWNODE
<< end >>
