magic
tech sky130A
magscale 1 2
timestamp 1672475742
<< pwell >>
rect 1063 558 1589 3120
<< nmos >>
rect 1263 868 1293 1868
rect 1359 868 1389 1868
<< ndiff >>
rect 1201 1856 1263 1868
rect 1201 880 1213 1856
rect 1247 880 1263 1856
rect 1201 868 1263 880
rect 1293 1856 1359 1868
rect 1293 880 1309 1856
rect 1343 880 1359 1856
rect 1293 868 1359 880
rect 1389 1856 1451 1868
rect 1389 880 1405 1856
rect 1439 880 1451 1856
rect 1389 868 1451 880
<< ndiffc >>
rect 1213 880 1247 1856
rect 1309 880 1343 1856
rect 1405 880 1439 1856
<< psubdiff >>
rect 1099 3050 1223 3084
rect 1429 3050 1553 3084
rect 1099 2960 1133 3050
rect 1099 628 1133 718
rect 1519 628 1553 3050
rect 1099 594 1195 628
rect 1457 594 1553 628
<< psubdiffcont >>
rect 1223 3050 1429 3084
rect 1099 718 1133 2960
rect 1195 594 1457 628
<< poly >>
rect 1263 1868 1293 1894
rect 1359 1868 1389 1894
rect 1263 846 1293 868
rect 1227 830 1293 846
rect 1227 675 1243 830
rect 1277 675 1293 830
rect 1227 648 1293 675
rect 1359 846 1389 868
rect 1359 830 1425 846
rect 1359 675 1375 830
rect 1409 675 1425 830
rect 1359 648 1425 675
<< polycont >>
rect 1243 675 1277 830
rect 1375 675 1409 830
<< xpolycontact >>
rect 1257 2522 1395 2954
rect 1257 1990 1395 2422
<< ppolyres >>
rect 1257 2422 1395 2522
<< locali >>
rect 1099 3050 1223 3084
rect 1429 3050 1445 3084
rect 1099 2960 1133 3050
rect 1133 2954 1167 2960
rect 1155 724 1167 2954
rect 1213 1856 1247 1872
rect 1213 864 1247 880
rect 1309 1856 1343 1872
rect 1309 864 1343 880
rect 1405 1856 1439 1872
rect 1405 864 1439 880
rect 1133 718 1167 724
rect 1099 628 1133 718
rect 1227 675 1243 830
rect 1277 675 1293 830
rect 1227 668 1293 675
rect 1359 675 1375 830
rect 1409 675 1425 830
rect 1359 668 1425 675
rect 1231 662 1289 668
rect 1363 662 1421 668
rect 1099 594 1195 628
rect 1457 594 1473 628
<< viali >>
rect 1111 724 1133 2954
rect 1133 724 1155 2954
rect 1273 2539 1379 2936
rect 1273 2008 1379 2405
rect 1213 880 1247 1856
rect 1309 880 1343 1856
rect 1405 880 1439 1856
rect 1243 675 1277 830
rect 1375 675 1409 830
<< metal1 >>
rect 1099 2954 1220 2960
rect 1099 724 1111 2954
rect 1155 2950 1220 2954
rect 1155 2810 1160 2950
rect 1155 2800 1220 2810
rect 1257 2936 1395 2954
rect 1155 724 1167 2800
rect 1257 2539 1273 2936
rect 1379 2539 1395 2936
rect 1257 2527 1395 2539
rect 1267 2405 1385 2417
rect 1267 2008 1273 2405
rect 1379 2008 1385 2405
rect 1267 1996 1385 2008
rect 1203 1856 1257 1868
rect 1203 868 1257 880
rect 1303 1856 1349 1996
rect 1303 880 1309 1856
rect 1343 880 1349 1856
rect 1303 868 1349 880
rect 1395 1856 1449 1868
rect 1395 868 1449 880
rect 1099 718 1167 724
rect 1231 830 1289 836
rect 1231 675 1243 830
rect 1277 675 1289 830
rect 1231 662 1289 675
rect 1363 830 1421 836
rect 1363 675 1375 830
rect 1409 675 1421 830
rect 1363 662 1421 675
rect 1240 570 1280 662
rect 1200 510 1210 570
rect 1270 510 1280 570
rect 1370 570 1410 662
rect 1370 510 1380 570
rect 1440 510 1450 570
<< via1 >>
rect 1160 2810 1220 2950
rect 1273 2539 1379 2936
rect 1203 880 1213 1856
rect 1213 880 1247 1856
rect 1247 880 1257 1856
rect 1395 880 1405 1856
rect 1405 880 1439 1856
rect 1439 880 1449 1856
rect 1210 510 1270 570
rect 1380 510 1440 570
<< metal2 >>
rect 1420 3360 1500 3370
rect 1420 3300 1430 3360
rect 1490 3300 1500 3360
rect 1420 3290 1500 3300
rect 1150 3190 1230 3200
rect 1150 3130 1160 3190
rect 1220 3130 1230 3190
rect 1150 3120 1230 3130
rect 1160 2950 1220 3120
rect 1160 2800 1220 2810
rect 1257 2936 1395 2954
rect 1257 2610 1273 2936
rect 1379 2610 1395 2936
rect 1257 2550 1270 2610
rect 1380 2550 1395 2610
rect 1257 2539 1273 2550
rect 1379 2539 1395 2550
rect 1257 2527 1395 2539
rect 1428 1896 1482 3290
rect 1395 1868 1482 1896
rect 1203 1860 1257 1868
rect 1180 1856 1257 1860
rect 1180 1850 1203 1856
rect 1180 1790 1190 1850
rect 1180 1780 1203 1790
rect 1203 868 1257 880
rect 1395 1856 1449 1868
rect 1395 868 1449 880
rect 1200 500 1210 570
rect 1270 500 1280 570
rect 1200 490 1280 500
rect 1370 500 1380 570
rect 1440 500 1450 570
rect 1370 490 1450 500
<< via2 >>
rect 1430 3300 1490 3360
rect 1160 3130 1220 3190
rect 1270 2550 1273 2610
rect 1273 2550 1379 2610
rect 1379 2550 1380 2610
rect 1190 1790 1203 1850
rect 1203 1790 1250 1850
rect 1210 510 1270 560
rect 1210 500 1270 510
rect 1380 510 1440 560
rect 1380 500 1440 510
<< metal3 >>
rect 1060 3360 1590 3370
rect 1060 3300 1430 3360
rect 1490 3300 1590 3360
rect 1060 3290 1590 3300
rect 1060 3190 1590 3200
rect 1060 3130 1160 3190
rect 1220 3130 1590 3190
rect 1060 3120 1590 3130
rect 1060 2610 1590 2620
rect 1060 2550 1270 2610
rect 1380 2550 1590 2610
rect 1060 2540 1590 2550
rect 1060 1850 1590 1860
rect 1060 1790 1190 1850
rect 1250 1790 1590 1850
rect 1060 1780 1590 1790
rect 1200 560 1280 570
rect 1200 500 1210 560
rect 1270 500 1280 560
rect 1200 450 1280 500
rect 1370 560 1450 570
rect 1370 500 1380 560
rect 1440 500 1450 560
rect 1370 450 1450 500
<< comment >>
rect 1099 2960 1133 3084
rect 1099 594 1133 718
<< labels >>
rlabel metal3 1060 3290 1130 3370 1 BUS_OUT
port 1 n
rlabel metal3 1520 3120 1560 3200 1 VSUB
port 4 n
rlabel metal3 1570 2540 1590 2620 1 IN
port 5 n
rlabel metal3 1370 450 1450 470 1 SOUT
port 2 n
rlabel metal3 1200 450 1280 470 1 SGND
port 3 n
rlabel metal3 1060 1780 1100 1860 1 VMID
port 6 n
rlabel metal1 1310 1900 1330 1940 1 SWNODE
<< end >>
