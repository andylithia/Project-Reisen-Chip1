VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cfgsr
  CLASS BLOCK ;
  FOREIGN cfgsr ;
  ORIGIN 0.000 0.000 ;
  SIZE 800.000 BY 80.000 ;
  PIN dq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.930 76.000 48.210 80.000 ;
    END
  END dq[0]
  PIN dq[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.930 76.000 324.210 80.000 ;
    END
  END dq[100]
  PIN dq[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.690 76.000 326.970 80.000 ;
    END
  END dq[101]
  PIN dq[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.450 76.000 329.730 80.000 ;
    END
  END dq[102]
  PIN dq[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.210 76.000 332.490 80.000 ;
    END
  END dq[103]
  PIN dq[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 76.000 335.250 80.000 ;
    END
  END dq[104]
  PIN dq[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.730 76.000 338.010 80.000 ;
    END
  END dq[105]
  PIN dq[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.490 76.000 340.770 80.000 ;
    END
  END dq[106]
  PIN dq[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.250 76.000 343.530 80.000 ;
    END
  END dq[107]
  PIN dq[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.010 76.000 346.290 80.000 ;
    END
  END dq[108]
  PIN dq[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.770 76.000 349.050 80.000 ;
    END
  END dq[109]
  PIN dq[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.530 76.000 75.810 80.000 ;
    END
  END dq[10]
  PIN dq[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.530 76.000 351.810 80.000 ;
    END
  END dq[110]
  PIN dq[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 76.000 354.570 80.000 ;
    END
  END dq[111]
  PIN dq[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.050 76.000 357.330 80.000 ;
    END
  END dq[112]
  PIN dq[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.810 76.000 360.090 80.000 ;
    END
  END dq[113]
  PIN dq[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.570 76.000 362.850 80.000 ;
    END
  END dq[114]
  PIN dq[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.330 76.000 365.610 80.000 ;
    END
  END dq[115]
  PIN dq[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.090 76.000 368.370 80.000 ;
    END
  END dq[116]
  PIN dq[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.850 76.000 371.130 80.000 ;
    END
  END dq[117]
  PIN dq[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.610 76.000 373.890 80.000 ;
    END
  END dq[118]
  PIN dq[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.370 76.000 376.650 80.000 ;
    END
  END dq[119]
  PIN dq[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 76.000 78.570 80.000 ;
    END
  END dq[11]
  PIN dq[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.130 76.000 379.410 80.000 ;
    END
  END dq[120]
  PIN dq[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.890 76.000 382.170 80.000 ;
    END
  END dq[121]
  PIN dq[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.650 76.000 384.930 80.000 ;
    END
  END dq[122]
  PIN dq[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.410 76.000 387.690 80.000 ;
    END
  END dq[123]
  PIN dq[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.170 76.000 390.450 80.000 ;
    END
  END dq[124]
  PIN dq[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 76.000 393.210 80.000 ;
    END
  END dq[125]
  PIN dq[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.690 76.000 395.970 80.000 ;
    END
  END dq[126]
  PIN dq[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.450 76.000 398.730 80.000 ;
    END
  END dq[127]
  PIN dq[128]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.210 76.000 401.490 80.000 ;
    END
  END dq[128]
  PIN dq[129]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.970 76.000 404.250 80.000 ;
    END
  END dq[129]
  PIN dq[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 76.000 81.330 80.000 ;
    END
  END dq[12]
  PIN dq[130]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.730 76.000 407.010 80.000 ;
    END
  END dq[130]
  PIN dq[131]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.490 76.000 409.770 80.000 ;
    END
  END dq[131]
  PIN dq[132]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 76.000 412.530 80.000 ;
    END
  END dq[132]
  PIN dq[133]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.010 76.000 415.290 80.000 ;
    END
  END dq[133]
  PIN dq[134]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.770 76.000 418.050 80.000 ;
    END
  END dq[134]
  PIN dq[135]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.530 76.000 420.810 80.000 ;
    END
  END dq[135]
  PIN dq[136]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.290 76.000 423.570 80.000 ;
    END
  END dq[136]
  PIN dq[137]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.050 76.000 426.330 80.000 ;
    END
  END dq[137]
  PIN dq[138]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.810 76.000 429.090 80.000 ;
    END
  END dq[138]
  PIN dq[139]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.570 76.000 431.850 80.000 ;
    END
  END dq[139]
  PIN dq[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 76.000 84.090 80.000 ;
    END
  END dq[13]
  PIN dq[140]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.330 76.000 434.610 80.000 ;
    END
  END dq[140]
  PIN dq[141]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.090 76.000 437.370 80.000 ;
    END
  END dq[141]
  PIN dq[142]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.850 76.000 440.130 80.000 ;
    END
  END dq[142]
  PIN dq[143]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.610 76.000 442.890 80.000 ;
    END
  END dq[143]
  PIN dq[144]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.370 76.000 445.650 80.000 ;
    END
  END dq[144]
  PIN dq[145]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.130 76.000 448.410 80.000 ;
    END
  END dq[145]
  PIN dq[146]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 76.000 451.170 80.000 ;
    END
  END dq[146]
  PIN dq[147]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.650 76.000 453.930 80.000 ;
    END
  END dq[147]
  PIN dq[148]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.410 76.000 456.690 80.000 ;
    END
  END dq[148]
  PIN dq[149]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 459.170 76.000 459.450 80.000 ;
    END
  END dq[149]
  PIN dq[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.570 76.000 86.850 80.000 ;
    END
  END dq[14]
  PIN dq[150]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.930 76.000 462.210 80.000 ;
    END
  END dq[150]
  PIN dq[151]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.690 76.000 464.970 80.000 ;
    END
  END dq[151]
  PIN dq[152]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.450 76.000 467.730 80.000 ;
    END
  END dq[152]
  PIN dq[153]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.210 76.000 470.490 80.000 ;
    END
  END dq[153]
  PIN dq[154]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.970 76.000 473.250 80.000 ;
    END
  END dq[154]
  PIN dq[155]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.730 76.000 476.010 80.000 ;
    END
  END dq[155]
  PIN dq[156]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.490 76.000 478.770 80.000 ;
    END
  END dq[156]
  PIN dq[157]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.250 76.000 481.530 80.000 ;
    END
  END dq[157]
  PIN dq[158]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.010 76.000 484.290 80.000 ;
    END
  END dq[158]
  PIN dq[159]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.770 76.000 487.050 80.000 ;
    END
  END dq[159]
  PIN dq[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 76.000 89.610 80.000 ;
    END
  END dq[15]
  PIN dq[160]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.530 76.000 489.810 80.000 ;
    END
  END dq[160]
  PIN dq[161]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.290 76.000 492.570 80.000 ;
    END
  END dq[161]
  PIN dq[162]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.050 76.000 495.330 80.000 ;
    END
  END dq[162]
  PIN dq[163]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 497.810 76.000 498.090 80.000 ;
    END
  END dq[163]
  PIN dq[164]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 500.570 76.000 500.850 80.000 ;
    END
  END dq[164]
  PIN dq[165]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 503.330 76.000 503.610 80.000 ;
    END
  END dq[165]
  PIN dq[166]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.090 76.000 506.370 80.000 ;
    END
  END dq[166]
  PIN dq[167]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.850 76.000 509.130 80.000 ;
    END
  END dq[167]
  PIN dq[168]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.610 76.000 511.890 80.000 ;
    END
  END dq[168]
  PIN dq[169]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.370 76.000 514.650 80.000 ;
    END
  END dq[169]
  PIN dq[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 76.000 92.370 80.000 ;
    END
  END dq[16]
  PIN dq[170]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.130 76.000 517.410 80.000 ;
    END
  END dq[170]
  PIN dq[171]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.890 76.000 520.170 80.000 ;
    END
  END dq[171]
  PIN dq[172]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.650 76.000 522.930 80.000 ;
    END
  END dq[172]
  PIN dq[173]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 525.410 76.000 525.690 80.000 ;
    END
  END dq[173]
  PIN dq[174]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 76.000 528.450 80.000 ;
    END
  END dq[174]
  PIN dq[175]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.930 76.000 531.210 80.000 ;
    END
  END dq[175]
  PIN dq[176]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 533.690 76.000 533.970 80.000 ;
    END
  END dq[176]
  PIN dq[177]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 536.450 76.000 536.730 80.000 ;
    END
  END dq[177]
  PIN dq[178]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 539.210 76.000 539.490 80.000 ;
    END
  END dq[178]
  PIN dq[179]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.970 76.000 542.250 80.000 ;
    END
  END dq[179]
  PIN dq[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 76.000 95.130 80.000 ;
    END
  END dq[17]
  PIN dq[180]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.730 76.000 545.010 80.000 ;
    END
  END dq[180]
  PIN dq[181]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.490 76.000 547.770 80.000 ;
    END
  END dq[181]
  PIN dq[182]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.250 76.000 550.530 80.000 ;
    END
  END dq[182]
  PIN dq[183]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.010 76.000 553.290 80.000 ;
    END
  END dq[183]
  PIN dq[184]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 555.770 76.000 556.050 80.000 ;
    END
  END dq[184]
  PIN dq[185]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.530 76.000 558.810 80.000 ;
    END
  END dq[185]
  PIN dq[186]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.290 76.000 561.570 80.000 ;
    END
  END dq[186]
  PIN dq[187]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.050 76.000 564.330 80.000 ;
    END
  END dq[187]
  PIN dq[188]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.810 76.000 567.090 80.000 ;
    END
  END dq[188]
  PIN dq[189]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.570 76.000 569.850 80.000 ;
    END
  END dq[189]
  PIN dq[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.610 76.000 97.890 80.000 ;
    END
  END dq[18]
  PIN dq[190]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.330 76.000 572.610 80.000 ;
    END
  END dq[190]
  PIN dq[191]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.090 76.000 575.370 80.000 ;
    END
  END dq[191]
  PIN dq[192]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.850 76.000 578.130 80.000 ;
    END
  END dq[192]
  PIN dq[193]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 580.610 76.000 580.890 80.000 ;
    END
  END dq[193]
  PIN dq[194]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 583.370 76.000 583.650 80.000 ;
    END
  END dq[194]
  PIN dq[195]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.130 76.000 586.410 80.000 ;
    END
  END dq[195]
  PIN dq[196]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 588.890 76.000 589.170 80.000 ;
    END
  END dq[196]
  PIN dq[197]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.650 76.000 591.930 80.000 ;
    END
  END dq[197]
  PIN dq[198]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 594.410 76.000 594.690 80.000 ;
    END
  END dq[198]
  PIN dq[199]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.170 76.000 597.450 80.000 ;
    END
  END dq[199]
  PIN dq[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.370 76.000 100.650 80.000 ;
    END
  END dq[19]
  PIN dq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 76.000 50.970 80.000 ;
    END
  END dq[1]
  PIN dq[200]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.930 76.000 600.210 80.000 ;
    END
  END dq[200]
  PIN dq[201]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.690 76.000 602.970 80.000 ;
    END
  END dq[201]
  PIN dq[202]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.450 76.000 605.730 80.000 ;
    END
  END dq[202]
  PIN dq[203]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.210 76.000 608.490 80.000 ;
    END
  END dq[203]
  PIN dq[204]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.970 76.000 611.250 80.000 ;
    END
  END dq[204]
  PIN dq[205]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 613.730 76.000 614.010 80.000 ;
    END
  END dq[205]
  PIN dq[206]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.490 76.000 616.770 80.000 ;
    END
  END dq[206]
  PIN dq[207]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 619.250 76.000 619.530 80.000 ;
    END
  END dq[207]
  PIN dq[208]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.010 76.000 622.290 80.000 ;
    END
  END dq[208]
  PIN dq[209]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.770 76.000 625.050 80.000 ;
    END
  END dq[209]
  PIN dq[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 76.000 103.410 80.000 ;
    END
  END dq[20]
  PIN dq[210]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.530 76.000 627.810 80.000 ;
    END
  END dq[210]
  PIN dq[211]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 630.290 76.000 630.570 80.000 ;
    END
  END dq[211]
  PIN dq[212]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.050 76.000 633.330 80.000 ;
    END
  END dq[212]
  PIN dq[213]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 635.810 76.000 636.090 80.000 ;
    END
  END dq[213]
  PIN dq[214]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 638.570 76.000 638.850 80.000 ;
    END
  END dq[214]
  PIN dq[215]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 641.330 76.000 641.610 80.000 ;
    END
  END dq[215]
  PIN dq[216]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.090 76.000 644.370 80.000 ;
    END
  END dq[216]
  PIN dq[217]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.850 76.000 647.130 80.000 ;
    END
  END dq[217]
  PIN dq[218]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 649.610 76.000 649.890 80.000 ;
    END
  END dq[218]
  PIN dq[219]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.370 76.000 652.650 80.000 ;
    END
  END dq[219]
  PIN dq[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 76.000 106.170 80.000 ;
    END
  END dq[21]
  PIN dq[220]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 655.130 76.000 655.410 80.000 ;
    END
  END dq[220]
  PIN dq[221]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.890 76.000 658.170 80.000 ;
    END
  END dq[221]
  PIN dq[222]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.650 76.000 660.930 80.000 ;
    END
  END dq[222]
  PIN dq[223]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.410 76.000 663.690 80.000 ;
    END
  END dq[223]
  PIN dq[224]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.170 76.000 666.450 80.000 ;
    END
  END dq[224]
  PIN dq[225]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.930 76.000 669.210 80.000 ;
    END
  END dq[225]
  PIN dq[226]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 671.690 76.000 671.970 80.000 ;
    END
  END dq[226]
  PIN dq[227]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.450 76.000 674.730 80.000 ;
    END
  END dq[227]
  PIN dq[228]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 677.210 76.000 677.490 80.000 ;
    END
  END dq[228]
  PIN dq[229]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.970 76.000 680.250 80.000 ;
    END
  END dq[229]
  PIN dq[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.650 76.000 108.930 80.000 ;
    END
  END dq[22]
  PIN dq[230]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.730 76.000 683.010 80.000 ;
    END
  END dq[230]
  PIN dq[231]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.490 76.000 685.770 80.000 ;
    END
  END dq[231]
  PIN dq[232]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.250 76.000 688.530 80.000 ;
    END
  END dq[232]
  PIN dq[233]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 691.010 76.000 691.290 80.000 ;
    END
  END dq[233]
  PIN dq[234]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 693.770 76.000 694.050 80.000 ;
    END
  END dq[234]
  PIN dq[235]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.530 76.000 696.810 80.000 ;
    END
  END dq[235]
  PIN dq[236]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.290 76.000 699.570 80.000 ;
    END
  END dq[236]
  PIN dq[237]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.050 76.000 702.330 80.000 ;
    END
  END dq[237]
  PIN dq[238]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 704.810 76.000 705.090 80.000 ;
    END
  END dq[238]
  PIN dq[239]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 707.570 76.000 707.850 80.000 ;
    END
  END dq[239]
  PIN dq[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.410 76.000 111.690 80.000 ;
    END
  END dq[23]
  PIN dq[240]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 710.330 76.000 710.610 80.000 ;
    END
  END dq[240]
  PIN dq[241]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 713.090 76.000 713.370 80.000 ;
    END
  END dq[241]
  PIN dq[242]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.850 76.000 716.130 80.000 ;
    END
  END dq[242]
  PIN dq[243]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.610 76.000 718.890 80.000 ;
    END
  END dq[243]
  PIN dq[244]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.370 76.000 721.650 80.000 ;
    END
  END dq[244]
  PIN dq[245]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.130 76.000 724.410 80.000 ;
    END
  END dq[245]
  PIN dq[246]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 726.890 76.000 727.170 80.000 ;
    END
  END dq[246]
  PIN dq[247]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.650 76.000 729.930 80.000 ;
    END
  END dq[247]
  PIN dq[248]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 732.410 76.000 732.690 80.000 ;
    END
  END dq[248]
  PIN dq[249]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.170 76.000 735.450 80.000 ;
    END
  END dq[249]
  PIN dq[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 76.000 114.450 80.000 ;
    END
  END dq[24]
  PIN dq[250]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.930 76.000 738.210 80.000 ;
    END
  END dq[250]
  PIN dq[251]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.690 76.000 740.970 80.000 ;
    END
  END dq[251]
  PIN dq[252]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.450 76.000 743.730 80.000 ;
    END
  END dq[252]
  PIN dq[253]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 746.210 76.000 746.490 80.000 ;
    END
  END dq[253]
  PIN dq[254]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.970 76.000 749.250 80.000 ;
    END
  END dq[254]
  PIN dq[255]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 751.730 76.000 752.010 80.000 ;
    END
  END dq[255]
  PIN dq[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.930 76.000 117.210 80.000 ;
    END
  END dq[25]
  PIN dq[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 76.000 119.970 80.000 ;
    END
  END dq[26]
  PIN dq[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 76.000 122.730 80.000 ;
    END
  END dq[27]
  PIN dq[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.210 76.000 125.490 80.000 ;
    END
  END dq[28]
  PIN dq[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.970 76.000 128.250 80.000 ;
    END
  END dq[29]
  PIN dq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.450 76.000 53.730 80.000 ;
    END
  END dq[2]
  PIN dq[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.730 76.000 131.010 80.000 ;
    END
  END dq[30]
  PIN dq[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.490 76.000 133.770 80.000 ;
    END
  END dq[31]
  PIN dq[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.250 76.000 136.530 80.000 ;
    END
  END dq[32]
  PIN dq[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.010 76.000 139.290 80.000 ;
    END
  END dq[33]
  PIN dq[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 76.000 142.050 80.000 ;
    END
  END dq[34]
  PIN dq[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 76.000 144.810 80.000 ;
    END
  END dq[35]
  PIN dq[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 76.000 147.570 80.000 ;
    END
  END dq[36]
  PIN dq[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.050 76.000 150.330 80.000 ;
    END
  END dq[37]
  PIN dq[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.810 76.000 153.090 80.000 ;
    END
  END dq[38]
  PIN dq[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.570 76.000 155.850 80.000 ;
    END
  END dq[39]
  PIN dq[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 76.000 56.490 80.000 ;
    END
  END dq[3]
  PIN dq[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.330 76.000 158.610 80.000 ;
    END
  END dq[40]
  PIN dq[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 76.000 161.370 80.000 ;
    END
  END dq[41]
  PIN dq[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.850 76.000 164.130 80.000 ;
    END
  END dq[42]
  PIN dq[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.610 76.000 166.890 80.000 ;
    END
  END dq[43]
  PIN dq[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.370 76.000 169.650 80.000 ;
    END
  END dq[44]
  PIN dq[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.130 76.000 172.410 80.000 ;
    END
  END dq[45]
  PIN dq[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 76.000 175.170 80.000 ;
    END
  END dq[46]
  PIN dq[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.650 76.000 177.930 80.000 ;
    END
  END dq[47]
  PIN dq[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 76.000 180.690 80.000 ;
    END
  END dq[48]
  PIN dq[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.170 76.000 183.450 80.000 ;
    END
  END dq[49]
  PIN dq[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 76.000 59.250 80.000 ;
    END
  END dq[4]
  PIN dq[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.930 76.000 186.210 80.000 ;
    END
  END dq[50]
  PIN dq[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.690 76.000 188.970 80.000 ;
    END
  END dq[51]
  PIN dq[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.450 76.000 191.730 80.000 ;
    END
  END dq[52]
  PIN dq[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.210 76.000 194.490 80.000 ;
    END
  END dq[53]
  PIN dq[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.970 76.000 197.250 80.000 ;
    END
  END dq[54]
  PIN dq[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 76.000 200.010 80.000 ;
    END
  END dq[55]
  PIN dq[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.490 76.000 202.770 80.000 ;
    END
  END dq[56]
  PIN dq[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.250 76.000 205.530 80.000 ;
    END
  END dq[57]
  PIN dq[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.010 76.000 208.290 80.000 ;
    END
  END dq[58]
  PIN dq[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.770 76.000 211.050 80.000 ;
    END
  END dq[59]
  PIN dq[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 76.000 62.010 80.000 ;
    END
  END dq[5]
  PIN dq[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.530 76.000 213.810 80.000 ;
    END
  END dq[60]
  PIN dq[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.290 76.000 216.570 80.000 ;
    END
  END dq[61]
  PIN dq[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 76.000 219.330 80.000 ;
    END
  END dq[62]
  PIN dq[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.810 76.000 222.090 80.000 ;
    END
  END dq[63]
  PIN dq[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.570 76.000 224.850 80.000 ;
    END
  END dq[64]
  PIN dq[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.330 76.000 227.610 80.000 ;
    END
  END dq[65]
  PIN dq[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.090 76.000 230.370 80.000 ;
    END
  END dq[66]
  PIN dq[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.850 76.000 233.130 80.000 ;
    END
  END dq[67]
  PIN dq[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.610 76.000 235.890 80.000 ;
    END
  END dq[68]
  PIN dq[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 76.000 238.650 80.000 ;
    END
  END dq[69]
  PIN dq[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 76.000 64.770 80.000 ;
    END
  END dq[6]
  PIN dq[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.130 76.000 241.410 80.000 ;
    END
  END dq[70]
  PIN dq[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.890 76.000 244.170 80.000 ;
    END
  END dq[71]
  PIN dq[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.650 76.000 246.930 80.000 ;
    END
  END dq[72]
  PIN dq[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.410 76.000 249.690 80.000 ;
    END
  END dq[73]
  PIN dq[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.170 76.000 252.450 80.000 ;
    END
  END dq[74]
  PIN dq[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.930 76.000 255.210 80.000 ;
    END
  END dq[75]
  PIN dq[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 76.000 257.970 80.000 ;
    END
  END dq[76]
  PIN dq[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.450 76.000 260.730 80.000 ;
    END
  END dq[77]
  PIN dq[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.210 76.000 263.490 80.000 ;
    END
  END dq[78]
  PIN dq[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.970 76.000 266.250 80.000 ;
    END
  END dq[79]
  PIN dq[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.250 76.000 67.530 80.000 ;
    END
  END dq[7]
  PIN dq[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.730 76.000 269.010 80.000 ;
    END
  END dq[80]
  PIN dq[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.490 76.000 271.770 80.000 ;
    END
  END dq[81]
  PIN dq[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.250 76.000 274.530 80.000 ;
    END
  END dq[82]
  PIN dq[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 76.000 277.290 80.000 ;
    END
  END dq[83]
  PIN dq[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.770 76.000 280.050 80.000 ;
    END
  END dq[84]
  PIN dq[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.530 76.000 282.810 80.000 ;
    END
  END dq[85]
  PIN dq[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.290 76.000 285.570 80.000 ;
    END
  END dq[86]
  PIN dq[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.050 76.000 288.330 80.000 ;
    END
  END dq[87]
  PIN dq[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.810 76.000 291.090 80.000 ;
    END
  END dq[88]
  PIN dq[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.570 76.000 293.850 80.000 ;
    END
  END dq[89]
  PIN dq[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.010 76.000 70.290 80.000 ;
    END
  END dq[8]
  PIN dq[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 76.000 296.610 80.000 ;
    END
  END dq[90]
  PIN dq[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.090 76.000 299.370 80.000 ;
    END
  END dq[91]
  PIN dq[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.850 76.000 302.130 80.000 ;
    END
  END dq[92]
  PIN dq[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.610 76.000 304.890 80.000 ;
    END
  END dq[93]
  PIN dq[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.370 76.000 307.650 80.000 ;
    END
  END dq[94]
  PIN dq[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.130 76.000 310.410 80.000 ;
    END
  END dq[95]
  PIN dq[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.890 76.000 313.170 80.000 ;
    END
  END dq[96]
  PIN dq[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 76.000 315.930 80.000 ;
    END
  END dq[97]
  PIN dq[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.410 76.000 318.690 80.000 ;
    END
  END dq[98]
  PIN dq[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.170 76.000 321.450 80.000 ;
    END
  END dq[99]
  PIN dq[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 76.000 73.050 80.000 ;
    END
  END dq[9]
  PIN latch
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 4.000 49.600 ;
    END
  END latch
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 9.560 4.000 10.160 ;
    END
  END rst_n
  PIN sclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.720 4.000 69.320 ;
    END
  END sclk
  PIN sdi
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.280 4.000 29.880 ;
    END
  END sdi
  PIN sdo
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 39.480 800.000 40.080 ;
    END
  END sdo
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 103.330 10.640 104.930 68.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 300.555 10.640 302.155 68.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 497.780 10.640 499.380 68.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 695.005 10.640 696.605 68.240 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 201.940 10.640 203.540 68.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 399.165 10.640 400.765 68.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 596.390 10.640 597.990 68.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 793.615 10.640 795.215 68.240 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 794.420 68.085 ;
      LAYER met1 ;
        RECT 5.520 4.800 797.570 75.440 ;
      LAYER met2 ;
        RECT 7.910 75.720 47.650 76.570 ;
        RECT 48.490 75.720 50.410 76.570 ;
        RECT 51.250 75.720 53.170 76.570 ;
        RECT 54.010 75.720 55.930 76.570 ;
        RECT 56.770 75.720 58.690 76.570 ;
        RECT 59.530 75.720 61.450 76.570 ;
        RECT 62.290 75.720 64.210 76.570 ;
        RECT 65.050 75.720 66.970 76.570 ;
        RECT 67.810 75.720 69.730 76.570 ;
        RECT 70.570 75.720 72.490 76.570 ;
        RECT 73.330 75.720 75.250 76.570 ;
        RECT 76.090 75.720 78.010 76.570 ;
        RECT 78.850 75.720 80.770 76.570 ;
        RECT 81.610 75.720 83.530 76.570 ;
        RECT 84.370 75.720 86.290 76.570 ;
        RECT 87.130 75.720 89.050 76.570 ;
        RECT 89.890 75.720 91.810 76.570 ;
        RECT 92.650 75.720 94.570 76.570 ;
        RECT 95.410 75.720 97.330 76.570 ;
        RECT 98.170 75.720 100.090 76.570 ;
        RECT 100.930 75.720 102.850 76.570 ;
        RECT 103.690 75.720 105.610 76.570 ;
        RECT 106.450 75.720 108.370 76.570 ;
        RECT 109.210 75.720 111.130 76.570 ;
        RECT 111.970 75.720 113.890 76.570 ;
        RECT 114.730 75.720 116.650 76.570 ;
        RECT 117.490 75.720 119.410 76.570 ;
        RECT 120.250 75.720 122.170 76.570 ;
        RECT 123.010 75.720 124.930 76.570 ;
        RECT 125.770 75.720 127.690 76.570 ;
        RECT 128.530 75.720 130.450 76.570 ;
        RECT 131.290 75.720 133.210 76.570 ;
        RECT 134.050 75.720 135.970 76.570 ;
        RECT 136.810 75.720 138.730 76.570 ;
        RECT 139.570 75.720 141.490 76.570 ;
        RECT 142.330 75.720 144.250 76.570 ;
        RECT 145.090 75.720 147.010 76.570 ;
        RECT 147.850 75.720 149.770 76.570 ;
        RECT 150.610 75.720 152.530 76.570 ;
        RECT 153.370 75.720 155.290 76.570 ;
        RECT 156.130 75.720 158.050 76.570 ;
        RECT 158.890 75.720 160.810 76.570 ;
        RECT 161.650 75.720 163.570 76.570 ;
        RECT 164.410 75.720 166.330 76.570 ;
        RECT 167.170 75.720 169.090 76.570 ;
        RECT 169.930 75.720 171.850 76.570 ;
        RECT 172.690 75.720 174.610 76.570 ;
        RECT 175.450 75.720 177.370 76.570 ;
        RECT 178.210 75.720 180.130 76.570 ;
        RECT 180.970 75.720 182.890 76.570 ;
        RECT 183.730 75.720 185.650 76.570 ;
        RECT 186.490 75.720 188.410 76.570 ;
        RECT 189.250 75.720 191.170 76.570 ;
        RECT 192.010 75.720 193.930 76.570 ;
        RECT 194.770 75.720 196.690 76.570 ;
        RECT 197.530 75.720 199.450 76.570 ;
        RECT 200.290 75.720 202.210 76.570 ;
        RECT 203.050 75.720 204.970 76.570 ;
        RECT 205.810 75.720 207.730 76.570 ;
        RECT 208.570 75.720 210.490 76.570 ;
        RECT 211.330 75.720 213.250 76.570 ;
        RECT 214.090 75.720 216.010 76.570 ;
        RECT 216.850 75.720 218.770 76.570 ;
        RECT 219.610 75.720 221.530 76.570 ;
        RECT 222.370 75.720 224.290 76.570 ;
        RECT 225.130 75.720 227.050 76.570 ;
        RECT 227.890 75.720 229.810 76.570 ;
        RECT 230.650 75.720 232.570 76.570 ;
        RECT 233.410 75.720 235.330 76.570 ;
        RECT 236.170 75.720 238.090 76.570 ;
        RECT 238.930 75.720 240.850 76.570 ;
        RECT 241.690 75.720 243.610 76.570 ;
        RECT 244.450 75.720 246.370 76.570 ;
        RECT 247.210 75.720 249.130 76.570 ;
        RECT 249.970 75.720 251.890 76.570 ;
        RECT 252.730 75.720 254.650 76.570 ;
        RECT 255.490 75.720 257.410 76.570 ;
        RECT 258.250 75.720 260.170 76.570 ;
        RECT 261.010 75.720 262.930 76.570 ;
        RECT 263.770 75.720 265.690 76.570 ;
        RECT 266.530 75.720 268.450 76.570 ;
        RECT 269.290 75.720 271.210 76.570 ;
        RECT 272.050 75.720 273.970 76.570 ;
        RECT 274.810 75.720 276.730 76.570 ;
        RECT 277.570 75.720 279.490 76.570 ;
        RECT 280.330 75.720 282.250 76.570 ;
        RECT 283.090 75.720 285.010 76.570 ;
        RECT 285.850 75.720 287.770 76.570 ;
        RECT 288.610 75.720 290.530 76.570 ;
        RECT 291.370 75.720 293.290 76.570 ;
        RECT 294.130 75.720 296.050 76.570 ;
        RECT 296.890 75.720 298.810 76.570 ;
        RECT 299.650 75.720 301.570 76.570 ;
        RECT 302.410 75.720 304.330 76.570 ;
        RECT 305.170 75.720 307.090 76.570 ;
        RECT 307.930 75.720 309.850 76.570 ;
        RECT 310.690 75.720 312.610 76.570 ;
        RECT 313.450 75.720 315.370 76.570 ;
        RECT 316.210 75.720 318.130 76.570 ;
        RECT 318.970 75.720 320.890 76.570 ;
        RECT 321.730 75.720 323.650 76.570 ;
        RECT 324.490 75.720 326.410 76.570 ;
        RECT 327.250 75.720 329.170 76.570 ;
        RECT 330.010 75.720 331.930 76.570 ;
        RECT 332.770 75.720 334.690 76.570 ;
        RECT 335.530 75.720 337.450 76.570 ;
        RECT 338.290 75.720 340.210 76.570 ;
        RECT 341.050 75.720 342.970 76.570 ;
        RECT 343.810 75.720 345.730 76.570 ;
        RECT 346.570 75.720 348.490 76.570 ;
        RECT 349.330 75.720 351.250 76.570 ;
        RECT 352.090 75.720 354.010 76.570 ;
        RECT 354.850 75.720 356.770 76.570 ;
        RECT 357.610 75.720 359.530 76.570 ;
        RECT 360.370 75.720 362.290 76.570 ;
        RECT 363.130 75.720 365.050 76.570 ;
        RECT 365.890 75.720 367.810 76.570 ;
        RECT 368.650 75.720 370.570 76.570 ;
        RECT 371.410 75.720 373.330 76.570 ;
        RECT 374.170 75.720 376.090 76.570 ;
        RECT 376.930 75.720 378.850 76.570 ;
        RECT 379.690 75.720 381.610 76.570 ;
        RECT 382.450 75.720 384.370 76.570 ;
        RECT 385.210 75.720 387.130 76.570 ;
        RECT 387.970 75.720 389.890 76.570 ;
        RECT 390.730 75.720 392.650 76.570 ;
        RECT 393.490 75.720 395.410 76.570 ;
        RECT 396.250 75.720 398.170 76.570 ;
        RECT 399.010 75.720 400.930 76.570 ;
        RECT 401.770 75.720 403.690 76.570 ;
        RECT 404.530 75.720 406.450 76.570 ;
        RECT 407.290 75.720 409.210 76.570 ;
        RECT 410.050 75.720 411.970 76.570 ;
        RECT 412.810 75.720 414.730 76.570 ;
        RECT 415.570 75.720 417.490 76.570 ;
        RECT 418.330 75.720 420.250 76.570 ;
        RECT 421.090 75.720 423.010 76.570 ;
        RECT 423.850 75.720 425.770 76.570 ;
        RECT 426.610 75.720 428.530 76.570 ;
        RECT 429.370 75.720 431.290 76.570 ;
        RECT 432.130 75.720 434.050 76.570 ;
        RECT 434.890 75.720 436.810 76.570 ;
        RECT 437.650 75.720 439.570 76.570 ;
        RECT 440.410 75.720 442.330 76.570 ;
        RECT 443.170 75.720 445.090 76.570 ;
        RECT 445.930 75.720 447.850 76.570 ;
        RECT 448.690 75.720 450.610 76.570 ;
        RECT 451.450 75.720 453.370 76.570 ;
        RECT 454.210 75.720 456.130 76.570 ;
        RECT 456.970 75.720 458.890 76.570 ;
        RECT 459.730 75.720 461.650 76.570 ;
        RECT 462.490 75.720 464.410 76.570 ;
        RECT 465.250 75.720 467.170 76.570 ;
        RECT 468.010 75.720 469.930 76.570 ;
        RECT 470.770 75.720 472.690 76.570 ;
        RECT 473.530 75.720 475.450 76.570 ;
        RECT 476.290 75.720 478.210 76.570 ;
        RECT 479.050 75.720 480.970 76.570 ;
        RECT 481.810 75.720 483.730 76.570 ;
        RECT 484.570 75.720 486.490 76.570 ;
        RECT 487.330 75.720 489.250 76.570 ;
        RECT 490.090 75.720 492.010 76.570 ;
        RECT 492.850 75.720 494.770 76.570 ;
        RECT 495.610 75.720 497.530 76.570 ;
        RECT 498.370 75.720 500.290 76.570 ;
        RECT 501.130 75.720 503.050 76.570 ;
        RECT 503.890 75.720 505.810 76.570 ;
        RECT 506.650 75.720 508.570 76.570 ;
        RECT 509.410 75.720 511.330 76.570 ;
        RECT 512.170 75.720 514.090 76.570 ;
        RECT 514.930 75.720 516.850 76.570 ;
        RECT 517.690 75.720 519.610 76.570 ;
        RECT 520.450 75.720 522.370 76.570 ;
        RECT 523.210 75.720 525.130 76.570 ;
        RECT 525.970 75.720 527.890 76.570 ;
        RECT 528.730 75.720 530.650 76.570 ;
        RECT 531.490 75.720 533.410 76.570 ;
        RECT 534.250 75.720 536.170 76.570 ;
        RECT 537.010 75.720 538.930 76.570 ;
        RECT 539.770 75.720 541.690 76.570 ;
        RECT 542.530 75.720 544.450 76.570 ;
        RECT 545.290 75.720 547.210 76.570 ;
        RECT 548.050 75.720 549.970 76.570 ;
        RECT 550.810 75.720 552.730 76.570 ;
        RECT 553.570 75.720 555.490 76.570 ;
        RECT 556.330 75.720 558.250 76.570 ;
        RECT 559.090 75.720 561.010 76.570 ;
        RECT 561.850 75.720 563.770 76.570 ;
        RECT 564.610 75.720 566.530 76.570 ;
        RECT 567.370 75.720 569.290 76.570 ;
        RECT 570.130 75.720 572.050 76.570 ;
        RECT 572.890 75.720 574.810 76.570 ;
        RECT 575.650 75.720 577.570 76.570 ;
        RECT 578.410 75.720 580.330 76.570 ;
        RECT 581.170 75.720 583.090 76.570 ;
        RECT 583.930 75.720 585.850 76.570 ;
        RECT 586.690 75.720 588.610 76.570 ;
        RECT 589.450 75.720 591.370 76.570 ;
        RECT 592.210 75.720 594.130 76.570 ;
        RECT 594.970 75.720 596.890 76.570 ;
        RECT 597.730 75.720 599.650 76.570 ;
        RECT 600.490 75.720 602.410 76.570 ;
        RECT 603.250 75.720 605.170 76.570 ;
        RECT 606.010 75.720 607.930 76.570 ;
        RECT 608.770 75.720 610.690 76.570 ;
        RECT 611.530 75.720 613.450 76.570 ;
        RECT 614.290 75.720 616.210 76.570 ;
        RECT 617.050 75.720 618.970 76.570 ;
        RECT 619.810 75.720 621.730 76.570 ;
        RECT 622.570 75.720 624.490 76.570 ;
        RECT 625.330 75.720 627.250 76.570 ;
        RECT 628.090 75.720 630.010 76.570 ;
        RECT 630.850 75.720 632.770 76.570 ;
        RECT 633.610 75.720 635.530 76.570 ;
        RECT 636.370 75.720 638.290 76.570 ;
        RECT 639.130 75.720 641.050 76.570 ;
        RECT 641.890 75.720 643.810 76.570 ;
        RECT 644.650 75.720 646.570 76.570 ;
        RECT 647.410 75.720 649.330 76.570 ;
        RECT 650.170 75.720 652.090 76.570 ;
        RECT 652.930 75.720 654.850 76.570 ;
        RECT 655.690 75.720 657.610 76.570 ;
        RECT 658.450 75.720 660.370 76.570 ;
        RECT 661.210 75.720 663.130 76.570 ;
        RECT 663.970 75.720 665.890 76.570 ;
        RECT 666.730 75.720 668.650 76.570 ;
        RECT 669.490 75.720 671.410 76.570 ;
        RECT 672.250 75.720 674.170 76.570 ;
        RECT 675.010 75.720 676.930 76.570 ;
        RECT 677.770 75.720 679.690 76.570 ;
        RECT 680.530 75.720 682.450 76.570 ;
        RECT 683.290 75.720 685.210 76.570 ;
        RECT 686.050 75.720 687.970 76.570 ;
        RECT 688.810 75.720 690.730 76.570 ;
        RECT 691.570 75.720 693.490 76.570 ;
        RECT 694.330 75.720 696.250 76.570 ;
        RECT 697.090 75.720 699.010 76.570 ;
        RECT 699.850 75.720 701.770 76.570 ;
        RECT 702.610 75.720 704.530 76.570 ;
        RECT 705.370 75.720 707.290 76.570 ;
        RECT 708.130 75.720 710.050 76.570 ;
        RECT 710.890 75.720 712.810 76.570 ;
        RECT 713.650 75.720 715.570 76.570 ;
        RECT 716.410 75.720 718.330 76.570 ;
        RECT 719.170 75.720 721.090 76.570 ;
        RECT 721.930 75.720 723.850 76.570 ;
        RECT 724.690 75.720 726.610 76.570 ;
        RECT 727.450 75.720 729.370 76.570 ;
        RECT 730.210 75.720 732.130 76.570 ;
        RECT 732.970 75.720 734.890 76.570 ;
        RECT 735.730 75.720 737.650 76.570 ;
        RECT 738.490 75.720 740.410 76.570 ;
        RECT 741.250 75.720 743.170 76.570 ;
        RECT 744.010 75.720 745.930 76.570 ;
        RECT 746.770 75.720 748.690 76.570 ;
        RECT 749.530 75.720 751.450 76.570 ;
        RECT 752.290 75.720 797.540 76.570 ;
        RECT 7.910 4.770 797.540 75.720 ;
      LAYER met3 ;
        RECT 4.000 69.720 796.655 72.585 ;
        RECT 4.400 68.320 796.655 69.720 ;
        RECT 4.000 50.000 796.655 68.320 ;
        RECT 4.400 48.600 796.655 50.000 ;
        RECT 4.000 40.480 796.655 48.600 ;
        RECT 4.000 39.080 795.600 40.480 ;
        RECT 4.000 30.280 796.655 39.080 ;
        RECT 4.400 28.880 796.655 30.280 ;
        RECT 4.000 10.560 796.655 28.880 ;
        RECT 4.400 9.160 796.655 10.560 ;
        RECT 4.000 4.935 796.655 9.160 ;
      LAYER met4 ;
        RECT 621.295 68.640 784.465 72.585 ;
        RECT 621.295 10.240 694.605 68.640 ;
        RECT 697.005 10.240 784.465 68.640 ;
        RECT 621.295 5.615 784.465 10.240 ;
  END
END cfgsr
END LIBRARY

