magic
tech sky130A
magscale 1 2
timestamp 1671334348
<< pwell >>
rect -361 -933 361 933
<< psubdiff >>
rect -325 863 -229 897
rect 229 863 325 897
rect -325 801 -291 863
rect 291 801 325 863
rect -325 -863 -291 -801
rect 291 -863 325 -801
rect -325 -897 -229 -863
rect 229 -897 325 -863
<< psubdiffcont >>
rect -229 863 229 897
rect -325 -801 -291 801
rect 291 -801 325 801
rect -229 -897 229 -863
<< poly >>
rect -195 -717 -129 -337
rect -195 -751 -179 -717
rect -145 -751 -129 -717
rect -195 -767 -129 -751
rect 129 -717 195 -337
rect 129 -751 145 -717
rect 179 -751 195 -717
rect 129 -767 195 -751
<< polycont >>
rect -179 -751 -145 -717
rect 145 -751 179 -717
<< npolyres >>
rect -195 701 -21 767
rect -195 -337 -129 701
rect -87 -167 -21 701
rect 21 701 195 767
rect 21 -167 87 701
rect -87 -233 87 -167
rect 129 -337 195 701
<< locali >>
rect -325 863 -229 897
rect 229 863 325 897
rect -325 801 -291 863
rect 291 801 325 863
rect -195 -751 -179 -717
rect -145 -751 -129 -717
rect 129 -751 145 -717
rect 179 -751 195 -717
rect -325 -863 -291 -801
rect 291 -863 325 -801
rect -325 -897 -229 -863
rect 229 -897 325 -863
<< properties >>
string FIXED_BBOX -308 -880 308 880
string gencell sky130_fd_pr__res_generic_po
string library sky130
string parameters w 0.33 l 5.0 m 1 nx 4 wmin 0.330 lmin 1.650 rho 48.2 val 3.241k dummy 0 dw 0.0 term 0.0 sterm 0.0 caplen 0.4 snake 1 guard 1 glc 1 grc 1 gtc 1 gbc 1 roverlap 0 endcov 100 full_metal 1 hv_guard 0 n_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
