magic
tech sky130A
magscale 1 2
timestamp 1671850507
<< nwell >>
rect 222 249 666 570
<< pwell >>
rect 263 26 349 183
rect 357 1 535 191
rect 539 26 625 183
rect 381 -29 415 1
<< psubdiff >>
rect 289 133 323 157
rect 289 52 323 99
rect 565 133 599 157
rect 565 52 599 99
<< nsubdiff >>
rect 289 444 323 468
rect 289 351 323 410
rect 289 293 323 317
rect 565 444 599 468
rect 565 351 599 410
rect 565 293 599 317
<< psubdiffcont >>
rect 289 99 323 133
rect 565 99 599 133
<< nsubdiffcont >>
rect 289 410 323 444
rect 289 317 323 351
rect 565 410 599 444
rect 565 317 599 351
<< pdiode >>
rect 383 475 509 493
rect 383 305 392 475
rect 500 305 509 475
rect 383 285 509 305
<< ndiode >>
rect 383 147 509 165
rect 383 45 392 147
rect 501 45 509 147
rect 383 27 509 45
<< pdiodec >>
rect 392 305 500 475
<< ndiodec >>
rect 392 45 501 147
<< locali >>
rect 260 515 289 549
rect 323 515 381 549
rect 415 515 473 549
rect 507 515 565 549
rect 599 515 628 549
rect 277 444 335 515
rect 277 410 289 444
rect 323 410 335 444
rect 277 351 335 410
rect 277 317 289 351
rect 323 317 335 351
rect 277 282 335 317
rect 369 475 519 481
rect 369 305 392 475
rect 500 305 519 475
rect 369 240 519 305
rect 553 444 611 515
rect 553 410 565 444
rect 599 410 611 444
rect 553 351 611 410
rect 553 317 565 351
rect 599 317 611 351
rect 553 282 611 317
rect 369 200 384 240
rect 504 200 519 240
rect 277 133 335 150
rect 277 99 289 133
rect 323 99 335 133
rect 277 5 335 99
rect 369 147 519 200
rect 369 45 392 147
rect 501 45 519 147
rect 369 39 519 45
rect 553 133 611 150
rect 553 99 565 133
rect 599 99 611 133
rect 553 5 611 99
rect 260 -29 289 5
rect 323 -29 381 5
rect 415 -29 473 5
rect 507 -29 565 5
rect 599 -29 628 5
<< viali >>
rect 289 515 323 549
rect 381 515 415 549
rect 473 515 507 549
rect 565 515 599 549
rect 384 200 504 240
rect 289 -29 323 5
rect 381 -29 415 5
rect 473 -29 507 5
rect 565 -29 599 5
<< metal1 >>
rect 260 549 628 580
rect 260 515 289 549
rect 323 515 381 549
rect 415 515 473 549
rect 507 515 565 549
rect 599 515 628 549
rect 260 484 628 515
rect 369 240 519 249
rect 369 200 384 240
rect 504 200 519 240
rect 369 191 519 200
rect 260 5 628 36
rect 260 -29 289 5
rect 323 -29 381 5
rect 415 -29 473 5
rect 507 -29 565 5
rect 599 -29 628 5
rect 260 -60 628 -29
<< labels >>
rlabel metal1 370 192 518 248 1 DIODE
rlabel metal1 262 486 626 578 1 VPWR
rlabel metal1 262 -58 626 34 1 VGND
<< end >>
