magic
tech sky130A
magscale 1 2
timestamp 1671154011
<< error_p >>
rect -845 572 -787 578
rect -653 572 -595 578
rect -461 572 -403 578
rect -269 572 -211 578
rect -77 572 -19 578
rect 115 572 173 578
rect 307 572 365 578
rect 499 572 557 578
rect 691 572 749 578
rect 883 572 941 578
rect -845 538 -833 572
rect -653 538 -641 572
rect -461 538 -449 572
rect -269 538 -257 572
rect -77 538 -65 572
rect 115 538 127 572
rect 307 538 319 572
rect 499 538 511 572
rect 691 538 703 572
rect 883 538 895 572
rect -845 532 -787 538
rect -653 532 -595 538
rect -461 532 -403 538
rect -269 532 -211 538
rect -77 532 -19 538
rect 115 532 173 538
rect 307 532 365 538
rect 499 532 557 538
rect 691 532 749 538
rect 883 532 941 538
rect -941 -538 -883 -532
rect -749 -538 -691 -532
rect -557 -538 -499 -532
rect -365 -538 -307 -532
rect -173 -538 -115 -532
rect 19 -538 77 -532
rect 211 -538 269 -532
rect 403 -538 461 -532
rect 595 -538 653 -532
rect 787 -538 845 -532
rect -941 -572 -929 -538
rect -749 -572 -737 -538
rect -557 -572 -545 -538
rect -365 -572 -353 -538
rect -173 -572 -161 -538
rect 19 -572 31 -538
rect 211 -572 223 -538
rect 403 -572 415 -538
rect 595 -572 607 -538
rect 787 -572 799 -538
rect -941 -578 -883 -572
rect -749 -578 -691 -572
rect -557 -578 -499 -572
rect -365 -578 -307 -572
rect -173 -578 -115 -572
rect 19 -578 77 -572
rect 211 -578 269 -572
rect 403 -578 461 -572
rect 595 -578 653 -572
rect 787 -578 845 -572
<< pwell >>
rect -1127 -710 1127 710
<< nmos >>
rect -927 -500 -897 500
rect -831 -500 -801 500
rect -735 -500 -705 500
rect -639 -500 -609 500
rect -543 -500 -513 500
rect -447 -500 -417 500
rect -351 -500 -321 500
rect -255 -500 -225 500
rect -159 -500 -129 500
rect -63 -500 -33 500
rect 33 -500 63 500
rect 129 -500 159 500
rect 225 -500 255 500
rect 321 -500 351 500
rect 417 -500 447 500
rect 513 -500 543 500
rect 609 -500 639 500
rect 705 -500 735 500
rect 801 -500 831 500
rect 897 -500 927 500
<< ndiff >>
rect -989 488 -927 500
rect -989 -488 -977 488
rect -943 -488 -927 488
rect -989 -500 -927 -488
rect -897 488 -831 500
rect -897 -488 -881 488
rect -847 -488 -831 488
rect -897 -500 -831 -488
rect -801 488 -735 500
rect -801 -488 -785 488
rect -751 -488 -735 488
rect -801 -500 -735 -488
rect -705 488 -639 500
rect -705 -488 -689 488
rect -655 -488 -639 488
rect -705 -500 -639 -488
rect -609 488 -543 500
rect -609 -488 -593 488
rect -559 -488 -543 488
rect -609 -500 -543 -488
rect -513 488 -447 500
rect -513 -488 -497 488
rect -463 -488 -447 488
rect -513 -500 -447 -488
rect -417 488 -351 500
rect -417 -488 -401 488
rect -367 -488 -351 488
rect -417 -500 -351 -488
rect -321 488 -255 500
rect -321 -488 -305 488
rect -271 -488 -255 488
rect -321 -500 -255 -488
rect -225 488 -159 500
rect -225 -488 -209 488
rect -175 -488 -159 488
rect -225 -500 -159 -488
rect -129 488 -63 500
rect -129 -488 -113 488
rect -79 -488 -63 488
rect -129 -500 -63 -488
rect -33 488 33 500
rect -33 -488 -17 488
rect 17 -488 33 488
rect -33 -500 33 -488
rect 63 488 129 500
rect 63 -488 79 488
rect 113 -488 129 488
rect 63 -500 129 -488
rect 159 488 225 500
rect 159 -488 175 488
rect 209 -488 225 488
rect 159 -500 225 -488
rect 255 488 321 500
rect 255 -488 271 488
rect 305 -488 321 488
rect 255 -500 321 -488
rect 351 488 417 500
rect 351 -488 367 488
rect 401 -488 417 488
rect 351 -500 417 -488
rect 447 488 513 500
rect 447 -488 463 488
rect 497 -488 513 488
rect 447 -500 513 -488
rect 543 488 609 500
rect 543 -488 559 488
rect 593 -488 609 488
rect 543 -500 609 -488
rect 639 488 705 500
rect 639 -488 655 488
rect 689 -488 705 488
rect 639 -500 705 -488
rect 735 488 801 500
rect 735 -488 751 488
rect 785 -488 801 488
rect 735 -500 801 -488
rect 831 488 897 500
rect 831 -488 847 488
rect 881 -488 897 488
rect 831 -500 897 -488
rect 927 488 989 500
rect 927 -488 943 488
rect 977 -488 989 488
rect 927 -500 989 -488
<< ndiffc >>
rect -977 -488 -943 488
rect -881 -488 -847 488
rect -785 -488 -751 488
rect -689 -488 -655 488
rect -593 -488 -559 488
rect -497 -488 -463 488
rect -401 -488 -367 488
rect -305 -488 -271 488
rect -209 -488 -175 488
rect -113 -488 -79 488
rect -17 -488 17 488
rect 79 -488 113 488
rect 175 -488 209 488
rect 271 -488 305 488
rect 367 -488 401 488
rect 463 -488 497 488
rect 559 -488 593 488
rect 655 -488 689 488
rect 751 -488 785 488
rect 847 -488 881 488
rect 943 -488 977 488
<< psubdiff >>
rect -1091 640 -995 674
rect 995 640 1091 674
rect -1091 578 -1057 640
rect 1057 578 1091 640
rect -1091 -640 -1057 -578
rect 1057 -640 1091 -578
rect -1091 -674 -995 -640
rect 995 -674 1091 -640
<< psubdiffcont >>
rect -995 640 995 674
rect -1091 -578 -1057 578
rect 1057 -578 1091 578
rect -995 -674 995 -640
<< poly >>
rect -849 572 -783 588
rect -849 538 -833 572
rect -799 538 -783 572
rect -927 500 -897 526
rect -849 522 -783 538
rect -657 572 -591 588
rect -657 538 -641 572
rect -607 538 -591 572
rect -831 500 -801 522
rect -735 500 -705 526
rect -657 522 -591 538
rect -465 572 -399 588
rect -465 538 -449 572
rect -415 538 -399 572
rect -639 500 -609 522
rect -543 500 -513 526
rect -465 522 -399 538
rect -273 572 -207 588
rect -273 538 -257 572
rect -223 538 -207 572
rect -447 500 -417 522
rect -351 500 -321 526
rect -273 522 -207 538
rect -81 572 -15 588
rect -81 538 -65 572
rect -31 538 -15 572
rect -255 500 -225 522
rect -159 500 -129 526
rect -81 522 -15 538
rect 111 572 177 588
rect 111 538 127 572
rect 161 538 177 572
rect -63 500 -33 522
rect 33 500 63 526
rect 111 522 177 538
rect 303 572 369 588
rect 303 538 319 572
rect 353 538 369 572
rect 129 500 159 522
rect 225 500 255 526
rect 303 522 369 538
rect 495 572 561 588
rect 495 538 511 572
rect 545 538 561 572
rect 321 500 351 522
rect 417 500 447 526
rect 495 522 561 538
rect 687 572 753 588
rect 687 538 703 572
rect 737 538 753 572
rect 513 500 543 522
rect 609 500 639 526
rect 687 522 753 538
rect 879 572 945 588
rect 879 538 895 572
rect 929 538 945 572
rect 705 500 735 522
rect 801 500 831 526
rect 879 522 945 538
rect 897 500 927 522
rect -927 -522 -897 -500
rect -945 -538 -879 -522
rect -831 -526 -801 -500
rect -735 -522 -705 -500
rect -945 -572 -929 -538
rect -895 -572 -879 -538
rect -945 -588 -879 -572
rect -753 -538 -687 -522
rect -639 -526 -609 -500
rect -543 -522 -513 -500
rect -753 -572 -737 -538
rect -703 -572 -687 -538
rect -753 -588 -687 -572
rect -561 -538 -495 -522
rect -447 -526 -417 -500
rect -351 -522 -321 -500
rect -561 -572 -545 -538
rect -511 -572 -495 -538
rect -561 -588 -495 -572
rect -369 -538 -303 -522
rect -255 -526 -225 -500
rect -159 -522 -129 -500
rect -369 -572 -353 -538
rect -319 -572 -303 -538
rect -369 -588 -303 -572
rect -177 -538 -111 -522
rect -63 -526 -33 -500
rect 33 -522 63 -500
rect -177 -572 -161 -538
rect -127 -572 -111 -538
rect -177 -588 -111 -572
rect 15 -538 81 -522
rect 129 -526 159 -500
rect 225 -522 255 -500
rect 15 -572 31 -538
rect 65 -572 81 -538
rect 15 -588 81 -572
rect 207 -538 273 -522
rect 321 -526 351 -500
rect 417 -522 447 -500
rect 207 -572 223 -538
rect 257 -572 273 -538
rect 207 -588 273 -572
rect 399 -538 465 -522
rect 513 -526 543 -500
rect 609 -522 639 -500
rect 399 -572 415 -538
rect 449 -572 465 -538
rect 399 -588 465 -572
rect 591 -538 657 -522
rect 705 -526 735 -500
rect 801 -522 831 -500
rect 591 -572 607 -538
rect 641 -572 657 -538
rect 591 -588 657 -572
rect 783 -538 849 -522
rect 897 -526 927 -500
rect 783 -572 799 -538
rect 833 -572 849 -538
rect 783 -588 849 -572
<< polycont >>
rect -833 538 -799 572
rect -641 538 -607 572
rect -449 538 -415 572
rect -257 538 -223 572
rect -65 538 -31 572
rect 127 538 161 572
rect 319 538 353 572
rect 511 538 545 572
rect 703 538 737 572
rect 895 538 929 572
rect -929 -572 -895 -538
rect -737 -572 -703 -538
rect -545 -572 -511 -538
rect -353 -572 -319 -538
rect -161 -572 -127 -538
rect 31 -572 65 -538
rect 223 -572 257 -538
rect 415 -572 449 -538
rect 607 -572 641 -538
rect 799 -572 833 -538
<< locali >>
rect -1091 640 -995 674
rect 995 640 1091 674
rect -1091 578 -1057 640
rect 1057 578 1091 640
rect -849 538 -833 572
rect -799 538 -783 572
rect -657 538 -641 572
rect -607 538 -591 572
rect -465 538 -449 572
rect -415 538 -399 572
rect -273 538 -257 572
rect -223 538 -207 572
rect -81 538 -65 572
rect -31 538 -15 572
rect 111 538 127 572
rect 161 538 177 572
rect 303 538 319 572
rect 353 538 369 572
rect 495 538 511 572
rect 545 538 561 572
rect 687 538 703 572
rect 737 538 753 572
rect 879 538 895 572
rect 929 538 945 572
rect -977 488 -943 504
rect -977 -504 -943 -488
rect -881 488 -847 504
rect -881 -504 -847 -488
rect -785 488 -751 504
rect -785 -504 -751 -488
rect -689 488 -655 504
rect -689 -504 -655 -488
rect -593 488 -559 504
rect -593 -504 -559 -488
rect -497 488 -463 504
rect -497 -504 -463 -488
rect -401 488 -367 504
rect -401 -504 -367 -488
rect -305 488 -271 504
rect -305 -504 -271 -488
rect -209 488 -175 504
rect -209 -504 -175 -488
rect -113 488 -79 504
rect -113 -504 -79 -488
rect -17 488 17 504
rect -17 -504 17 -488
rect 79 488 113 504
rect 79 -504 113 -488
rect 175 488 209 504
rect 175 -504 209 -488
rect 271 488 305 504
rect 271 -504 305 -488
rect 367 488 401 504
rect 367 -504 401 -488
rect 463 488 497 504
rect 463 -504 497 -488
rect 559 488 593 504
rect 559 -504 593 -488
rect 655 488 689 504
rect 655 -504 689 -488
rect 751 488 785 504
rect 751 -504 785 -488
rect 847 488 881 504
rect 847 -504 881 -488
rect 943 488 977 504
rect 943 -504 977 -488
rect -945 -572 -929 -538
rect -895 -572 -879 -538
rect -753 -572 -737 -538
rect -703 -572 -687 -538
rect -561 -572 -545 -538
rect -511 -572 -495 -538
rect -369 -572 -353 -538
rect -319 -572 -303 -538
rect -177 -572 -161 -538
rect -127 -572 -111 -538
rect 15 -572 31 -538
rect 65 -572 81 -538
rect 207 -572 223 -538
rect 257 -572 273 -538
rect 399 -572 415 -538
rect 449 -572 465 -538
rect 591 -572 607 -538
rect 641 -572 657 -538
rect 783 -572 799 -538
rect 833 -572 849 -538
rect -1091 -640 -1057 -578
rect 1057 -640 1091 -578
rect -1091 -674 -995 -640
rect 995 -674 1091 -640
<< viali >>
rect -833 538 -799 572
rect -641 538 -607 572
rect -449 538 -415 572
rect -257 538 -223 572
rect -65 538 -31 572
rect 127 538 161 572
rect 319 538 353 572
rect 511 538 545 572
rect 703 538 737 572
rect 895 538 929 572
rect -977 -488 -943 488
rect -881 -488 -847 488
rect -785 -488 -751 488
rect -689 -488 -655 488
rect -593 -488 -559 488
rect -497 -488 -463 488
rect -401 -488 -367 488
rect -305 -488 -271 488
rect -209 -488 -175 488
rect -113 -488 -79 488
rect -17 -488 17 488
rect 79 -488 113 488
rect 175 -488 209 488
rect 271 -488 305 488
rect 367 -488 401 488
rect 463 -488 497 488
rect 559 -488 593 488
rect 655 -488 689 488
rect 751 -488 785 488
rect 847 -488 881 488
rect 943 -488 977 488
rect -929 -572 -895 -538
rect -737 -572 -703 -538
rect -545 -572 -511 -538
rect -353 -572 -319 -538
rect -161 -572 -127 -538
rect 31 -572 65 -538
rect 223 -572 257 -538
rect 415 -572 449 -538
rect 607 -572 641 -538
rect 799 -572 833 -538
<< metal1 >>
rect -845 572 -787 578
rect -845 538 -833 572
rect -799 538 -787 572
rect -845 532 -787 538
rect -653 572 -595 578
rect -653 538 -641 572
rect -607 538 -595 572
rect -653 532 -595 538
rect -461 572 -403 578
rect -461 538 -449 572
rect -415 538 -403 572
rect -461 532 -403 538
rect -269 572 -211 578
rect -269 538 -257 572
rect -223 538 -211 572
rect -269 532 -211 538
rect -77 572 -19 578
rect -77 538 -65 572
rect -31 538 -19 572
rect -77 532 -19 538
rect 115 572 173 578
rect 115 538 127 572
rect 161 538 173 572
rect 115 532 173 538
rect 307 572 365 578
rect 307 538 319 572
rect 353 538 365 572
rect 307 532 365 538
rect 499 572 557 578
rect 499 538 511 572
rect 545 538 557 572
rect 499 532 557 538
rect 691 572 749 578
rect 691 538 703 572
rect 737 538 749 572
rect 691 532 749 538
rect 883 572 941 578
rect 883 538 895 572
rect 929 538 941 572
rect 883 532 941 538
rect -983 488 -937 500
rect -983 -488 -977 488
rect -943 -488 -937 488
rect -983 -500 -937 -488
rect -887 488 -841 500
rect -887 -488 -881 488
rect -847 -488 -841 488
rect -887 -500 -841 -488
rect -791 488 -745 500
rect -791 -488 -785 488
rect -751 -488 -745 488
rect -791 -500 -745 -488
rect -695 488 -649 500
rect -695 -488 -689 488
rect -655 -488 -649 488
rect -695 -500 -649 -488
rect -599 488 -553 500
rect -599 -488 -593 488
rect -559 -488 -553 488
rect -599 -500 -553 -488
rect -503 488 -457 500
rect -503 -488 -497 488
rect -463 -488 -457 488
rect -503 -500 -457 -488
rect -407 488 -361 500
rect -407 -488 -401 488
rect -367 -488 -361 488
rect -407 -500 -361 -488
rect -311 488 -265 500
rect -311 -488 -305 488
rect -271 -488 -265 488
rect -311 -500 -265 -488
rect -215 488 -169 500
rect -215 -488 -209 488
rect -175 -488 -169 488
rect -215 -500 -169 -488
rect -119 488 -73 500
rect -119 -488 -113 488
rect -79 -488 -73 488
rect -119 -500 -73 -488
rect -23 488 23 500
rect -23 -488 -17 488
rect 17 -488 23 488
rect -23 -500 23 -488
rect 73 488 119 500
rect 73 -488 79 488
rect 113 -488 119 488
rect 73 -500 119 -488
rect 169 488 215 500
rect 169 -488 175 488
rect 209 -488 215 488
rect 169 -500 215 -488
rect 265 488 311 500
rect 265 -488 271 488
rect 305 -488 311 488
rect 265 -500 311 -488
rect 361 488 407 500
rect 361 -488 367 488
rect 401 -488 407 488
rect 361 -500 407 -488
rect 457 488 503 500
rect 457 -488 463 488
rect 497 -488 503 488
rect 457 -500 503 -488
rect 553 488 599 500
rect 553 -488 559 488
rect 593 -488 599 488
rect 553 -500 599 -488
rect 649 488 695 500
rect 649 -488 655 488
rect 689 -488 695 488
rect 649 -500 695 -488
rect 745 488 791 500
rect 745 -488 751 488
rect 785 -488 791 488
rect 745 -500 791 -488
rect 841 488 887 500
rect 841 -488 847 488
rect 881 -488 887 488
rect 841 -500 887 -488
rect 937 488 983 500
rect 937 -488 943 488
rect 977 -488 983 488
rect 937 -500 983 -488
rect -941 -538 -883 -532
rect -941 -572 -929 -538
rect -895 -572 -883 -538
rect -941 -578 -883 -572
rect -749 -538 -691 -532
rect -749 -572 -737 -538
rect -703 -572 -691 -538
rect -749 -578 -691 -572
rect -557 -538 -499 -532
rect -557 -572 -545 -538
rect -511 -572 -499 -538
rect -557 -578 -499 -572
rect -365 -538 -307 -532
rect -365 -572 -353 -538
rect -319 -572 -307 -538
rect -365 -578 -307 -572
rect -173 -538 -115 -532
rect -173 -572 -161 -538
rect -127 -572 -115 -538
rect -173 -578 -115 -572
rect 19 -538 77 -532
rect 19 -572 31 -538
rect 65 -572 77 -538
rect 19 -578 77 -572
rect 211 -538 269 -532
rect 211 -572 223 -538
rect 257 -572 269 -538
rect 211 -578 269 -572
rect 403 -538 461 -532
rect 403 -572 415 -538
rect 449 -572 461 -538
rect 403 -578 461 -572
rect 595 -538 653 -532
rect 595 -572 607 -538
rect 641 -572 653 -538
rect 595 -578 653 -572
rect 787 -538 845 -532
rect 787 -572 799 -538
rect 833 -572 845 -538
rect 787 -578 845 -572
<< properties >>
string FIXED_BBOX -1074 -657 1074 657
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 5 l 0.150 m 1 nf 20 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
