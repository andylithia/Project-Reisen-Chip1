magic
tech sky130A
timestamp 1671647065
<< metal1 >>
rect -6003 1876 -2003 2000
rect -6003 1850 -5696 1876
rect -5670 1850 -5536 1876
rect -5510 1850 -5376 1876
rect -5350 1850 -5216 1876
rect -5190 1850 -5056 1876
rect -5030 1850 -4896 1876
rect -4870 1850 -4736 1876
rect -4710 1850 -4576 1876
rect -4550 1850 -4416 1876
rect -4390 1850 -4256 1876
rect -4230 1850 -4096 1876
rect -4070 1850 -3936 1876
rect -3910 1850 -3776 1876
rect -3750 1850 -3616 1876
rect -3590 1850 -3456 1876
rect -3430 1850 -3296 1876
rect -3270 1850 -3136 1876
rect -3110 1850 -2976 1876
rect -2950 1850 -2816 1876
rect -2790 1850 -2656 1876
rect -2630 1850 -2496 1876
rect -2470 1850 -2336 1876
rect -2310 1850 -2003 1876
rect -6003 1773 -2003 1850
rect -6003 1747 -5881 1773
rect -5855 1747 -2148 1773
rect -2122 1747 -2003 1773
rect -6003 1730 -2003 1747
rect -6003 1613 -5733 1730
rect -6003 1587 -5881 1613
rect -5855 1587 -5733 1613
rect -6003 1453 -5733 1587
rect -6003 1427 -5881 1453
rect -5855 1427 -5733 1453
rect -6003 1293 -5733 1427
rect -6003 1267 -5881 1293
rect -5855 1267 -5733 1293
rect -6003 1133 -5733 1267
rect -6003 1107 -5881 1133
rect -5855 1107 -5733 1133
rect -6003 973 -5733 1107
rect -6003 947 -5881 973
rect -5855 947 -5733 973
rect -6003 813 -5733 947
rect -6003 787 -5881 813
rect -5855 787 -5733 813
rect -6003 653 -5733 787
rect -6003 627 -5881 653
rect -5855 627 -5733 653
rect -6003 493 -5733 627
rect -6003 467 -5881 493
rect -5855 467 -5733 493
rect -6003 333 -5733 467
rect -6003 307 -5881 333
rect -5855 307 -5733 333
rect -6003 173 -5733 307
rect -6003 147 -5881 173
rect -5855 147 -5733 173
rect -6003 13 -5733 147
rect -6003 -13 -5881 13
rect -5855 -13 -5733 13
rect -6003 -147 -5733 -13
rect -6003 -173 -5881 -147
rect -5855 -173 -5733 -147
rect -6003 -307 -5733 -173
rect -6003 -333 -5881 -307
rect -5855 -333 -5733 -307
rect -6003 -467 -5733 -333
rect -6003 -493 -5881 -467
rect -5855 -493 -5733 -467
rect -6003 -627 -5733 -493
rect -6003 -653 -5881 -627
rect -5855 -653 -5733 -627
rect -6003 -787 -5733 -653
rect -6003 -813 -5881 -787
rect -5855 -813 -5733 -787
rect -6003 -947 -5733 -813
rect -6003 -973 -5881 -947
rect -5855 -973 -5733 -947
rect -6003 -1107 -5733 -973
rect -6003 -1133 -5881 -1107
rect -5855 -1133 -5733 -1107
rect -6003 -1267 -5733 -1133
rect -6003 -1293 -5881 -1267
rect -5855 -1293 -5733 -1267
rect -6003 -1427 -5733 -1293
rect -6003 -1453 -5881 -1427
rect -5855 -1453 -5733 -1427
rect -6003 -1587 -5733 -1453
rect -6003 -1613 -5881 -1587
rect -5855 -1613 -5733 -1587
rect -6003 -1730 -5733 -1613
rect -2273 1613 -2003 1730
rect -2273 1587 -2148 1613
rect -2122 1587 -2003 1613
rect -2273 1453 -2003 1587
rect -2273 1427 -2148 1453
rect -2122 1427 -2003 1453
rect -2273 1293 -2003 1427
rect -2273 1267 -2148 1293
rect -2122 1267 -2003 1293
rect -2273 1133 -2003 1267
rect -2273 1107 -2148 1133
rect -2122 1107 -2003 1133
rect -2273 973 -2003 1107
rect -2273 947 -2148 973
rect -2122 947 -2003 973
rect -2273 813 -2003 947
rect -2273 787 -2148 813
rect -2122 787 -2003 813
rect -2273 653 -2003 787
rect -2273 627 -2148 653
rect -2122 627 -2003 653
rect -2273 493 -2003 627
rect -2273 467 -2148 493
rect -2122 467 -2003 493
rect -2273 333 -2003 467
rect -2273 307 -2148 333
rect -2122 307 -2003 333
rect -2273 173 -2003 307
rect -2273 147 -2148 173
rect -2122 147 -2003 173
rect -2273 13 -2003 147
rect -2273 -13 -2148 13
rect -2122 -13 -2003 13
rect -2273 -147 -2003 -13
rect -2273 -173 -2148 -147
rect -2122 -173 -2003 -147
rect -2273 -307 -2003 -173
rect -2273 -333 -2148 -307
rect -2122 -333 -2003 -307
rect -2273 -467 -2003 -333
rect -2273 -493 -2148 -467
rect -2122 -493 -2003 -467
rect -2273 -627 -2003 -493
rect -2273 -653 -2148 -627
rect -2122 -653 -2003 -627
rect -2273 -787 -2003 -653
rect -2273 -813 -2148 -787
rect -2122 -813 -2003 -787
rect -2273 -947 -2003 -813
rect -2273 -973 -2148 -947
rect -2122 -973 -2003 -947
rect -2273 -1107 -2003 -973
rect -2273 -1133 -2148 -1107
rect -2122 -1133 -2003 -1107
rect -2273 -1267 -2003 -1133
rect -2273 -1293 -2148 -1267
rect -2122 -1293 -2003 -1267
rect -2273 -1427 -2003 -1293
rect -2273 -1453 -2148 -1427
rect -2122 -1453 -2003 -1427
rect -2273 -1587 -2003 -1453
rect -2273 -1613 -2148 -1587
rect -2122 -1613 -2003 -1587
rect -2273 -1730 -2003 -1613
rect -6003 -1747 -2003 -1730
rect -6003 -1773 -5881 -1747
rect -5855 -1773 -2148 -1747
rect -2122 -1773 -2003 -1747
rect -6003 -1852 -2003 -1773
rect -6003 -1878 -5696 -1852
rect -5670 -1878 -5536 -1852
rect -5510 -1878 -5376 -1852
rect -5350 -1878 -5216 -1852
rect -5190 -1878 -5056 -1852
rect -5030 -1878 -4896 -1852
rect -4870 -1878 -4736 -1852
rect -4710 -1878 -4576 -1852
rect -4550 -1878 -4416 -1852
rect -4390 -1878 -4256 -1852
rect -4230 -1878 -4096 -1852
rect -4070 -1878 -3936 -1852
rect -3910 -1878 -3776 -1852
rect -3750 -1878 -3616 -1852
rect -3590 -1878 -3456 -1852
rect -3430 -1878 -3296 -1852
rect -3270 -1878 -3136 -1852
rect -3110 -1878 -2976 -1852
rect -2950 -1878 -2816 -1852
rect -2790 -1878 -2656 -1852
rect -2630 -1878 -2496 -1852
rect -2470 -1878 -2336 -1852
rect -2310 -1878 -2003 -1852
rect -6003 -2000 -2003 -1878
<< via1 >>
rect -5696 1850 -5670 1876
rect -5536 1850 -5510 1876
rect -5376 1850 -5350 1876
rect -5216 1850 -5190 1876
rect -5056 1850 -5030 1876
rect -4896 1850 -4870 1876
rect -4736 1850 -4710 1876
rect -4576 1850 -4550 1876
rect -4416 1850 -4390 1876
rect -4256 1850 -4230 1876
rect -4096 1850 -4070 1876
rect -3936 1850 -3910 1876
rect -3776 1850 -3750 1876
rect -3616 1850 -3590 1876
rect -3456 1850 -3430 1876
rect -3296 1850 -3270 1876
rect -3136 1850 -3110 1876
rect -2976 1850 -2950 1876
rect -2816 1850 -2790 1876
rect -2656 1850 -2630 1876
rect -2496 1850 -2470 1876
rect -2336 1850 -2310 1876
rect -5881 1747 -5855 1773
rect -2148 1747 -2122 1773
rect -5881 1587 -5855 1613
rect -5881 1427 -5855 1453
rect -5881 1267 -5855 1293
rect -5881 1107 -5855 1133
rect -5881 947 -5855 973
rect -5881 787 -5855 813
rect -5881 627 -5855 653
rect -5881 467 -5855 493
rect -5881 307 -5855 333
rect -5881 147 -5855 173
rect -5881 -13 -5855 13
rect -5881 -173 -5855 -147
rect -5881 -333 -5855 -307
rect -5881 -493 -5855 -467
rect -5881 -653 -5855 -627
rect -5881 -813 -5855 -787
rect -5881 -973 -5855 -947
rect -5881 -1133 -5855 -1107
rect -5881 -1293 -5855 -1267
rect -5881 -1453 -5855 -1427
rect -5881 -1613 -5855 -1587
rect -2148 1587 -2122 1613
rect -2148 1427 -2122 1453
rect -2148 1267 -2122 1293
rect -2148 1107 -2122 1133
rect -2148 947 -2122 973
rect -2148 787 -2122 813
rect -2148 627 -2122 653
rect -2148 467 -2122 493
rect -2148 307 -2122 333
rect -2148 147 -2122 173
rect -2148 -13 -2122 13
rect -2148 -173 -2122 -147
rect -2148 -333 -2122 -307
rect -2148 -493 -2122 -467
rect -2148 -653 -2122 -627
rect -2148 -813 -2122 -787
rect -2148 -973 -2122 -947
rect -2148 -1133 -2122 -1107
rect -2148 -1293 -2122 -1267
rect -2148 -1453 -2122 -1427
rect -2148 -1613 -2122 -1587
rect -5881 -1773 -5855 -1747
rect -2148 -1773 -2122 -1747
rect -5696 -1878 -5670 -1852
rect -5536 -1878 -5510 -1852
rect -5376 -1878 -5350 -1852
rect -5216 -1878 -5190 -1852
rect -5056 -1878 -5030 -1852
rect -4896 -1878 -4870 -1852
rect -4736 -1878 -4710 -1852
rect -4576 -1878 -4550 -1852
rect -4416 -1878 -4390 -1852
rect -4256 -1878 -4230 -1852
rect -4096 -1878 -4070 -1852
rect -3936 -1878 -3910 -1852
rect -3776 -1878 -3750 -1852
rect -3616 -1878 -3590 -1852
rect -3456 -1878 -3430 -1852
rect -3296 -1878 -3270 -1852
rect -3136 -1878 -3110 -1852
rect -2976 -1878 -2950 -1852
rect -2816 -1878 -2790 -1852
rect -2656 -1878 -2630 -1852
rect -2496 -1878 -2470 -1852
rect -2336 -1878 -2310 -1852
<< metal2 >>
rect -6003 1877 -2003 2000
rect -6003 1849 -5697 1877
rect -5669 1849 -5537 1877
rect -5509 1849 -5377 1877
rect -5349 1849 -5217 1877
rect -5189 1849 -5057 1877
rect -5029 1849 -4897 1877
rect -4869 1849 -4737 1877
rect -4709 1849 -4577 1877
rect -4549 1849 -4417 1877
rect -4389 1849 -4257 1877
rect -4229 1849 -4097 1877
rect -4069 1849 -3937 1877
rect -3909 1849 -3777 1877
rect -3749 1849 -3617 1877
rect -3589 1849 -3457 1877
rect -3429 1849 -3297 1877
rect -3269 1849 -3137 1877
rect -3109 1849 -2977 1877
rect -2949 1849 -2817 1877
rect -2789 1849 -2657 1877
rect -2629 1849 -2497 1877
rect -2469 1849 -2337 1877
rect -2309 1849 -2003 1877
rect -6003 1774 -2003 1849
rect -6003 1746 -5882 1774
rect -5854 1746 -2149 1774
rect -2121 1746 -2003 1774
rect -6003 1730 -2003 1746
rect -6003 1614 -5733 1730
rect -6003 1586 -5882 1614
rect -5854 1586 -5733 1614
rect -6003 1454 -5733 1586
rect -6003 1426 -5882 1454
rect -5854 1426 -5733 1454
rect -6003 1294 -5733 1426
rect -6003 1266 -5882 1294
rect -5854 1266 -5733 1294
rect -6003 1134 -5733 1266
rect -6003 1106 -5882 1134
rect -5854 1106 -5733 1134
rect -6003 974 -5733 1106
rect -6003 946 -5882 974
rect -5854 946 -5733 974
rect -6003 814 -5733 946
rect -6003 786 -5882 814
rect -5854 786 -5733 814
rect -6003 654 -5733 786
rect -6003 626 -5882 654
rect -5854 626 -5733 654
rect -6003 494 -5733 626
rect -6003 466 -5882 494
rect -5854 466 -5733 494
rect -6003 334 -5733 466
rect -6003 306 -5882 334
rect -5854 306 -5733 334
rect -6003 174 -5733 306
rect -6003 146 -5882 174
rect -5854 146 -5733 174
rect -6003 14 -5733 146
rect -6003 -14 -5882 14
rect -5854 -14 -5733 14
rect -6003 -146 -5733 -14
rect -6003 -174 -5882 -146
rect -5854 -174 -5733 -146
rect -6003 -306 -5733 -174
rect -6003 -334 -5882 -306
rect -5854 -334 -5733 -306
rect -6003 -466 -5733 -334
rect -6003 -494 -5882 -466
rect -5854 -494 -5733 -466
rect -6003 -626 -5733 -494
rect -6003 -654 -5882 -626
rect -5854 -654 -5733 -626
rect -6003 -786 -5733 -654
rect -6003 -814 -5882 -786
rect -5854 -814 -5733 -786
rect -6003 -946 -5733 -814
rect -6003 -974 -5882 -946
rect -5854 -974 -5733 -946
rect -6003 -1106 -5733 -974
rect -6003 -1134 -5882 -1106
rect -5854 -1134 -5733 -1106
rect -6003 -1266 -5733 -1134
rect -6003 -1294 -5882 -1266
rect -5854 -1294 -5733 -1266
rect -6003 -1426 -5733 -1294
rect -6003 -1454 -5882 -1426
rect -5854 -1454 -5733 -1426
rect -6003 -1586 -5733 -1454
rect -6003 -1614 -5882 -1586
rect -5854 -1614 -5733 -1586
rect -6003 -1730 -5733 -1614
rect -2273 1614 -2003 1730
rect -2273 1586 -2149 1614
rect -2121 1586 -2003 1614
rect -2273 1454 -2003 1586
rect -2273 1426 -2149 1454
rect -2121 1426 -2003 1454
rect -2273 1294 -2003 1426
rect -2273 1266 -2149 1294
rect -2121 1266 -2003 1294
rect -2273 1134 -2003 1266
rect -2273 1106 -2149 1134
rect -2121 1106 -2003 1134
rect -2273 974 -2003 1106
rect -2273 946 -2149 974
rect -2121 946 -2003 974
rect -2273 814 -2003 946
rect -2273 786 -2149 814
rect -2121 786 -2003 814
rect -2273 654 -2003 786
rect -2273 626 -2149 654
rect -2121 626 -2003 654
rect -2273 494 -2003 626
rect -2273 466 -2149 494
rect -2121 466 -2003 494
rect -2273 334 -2003 466
rect -2273 306 -2149 334
rect -2121 306 -2003 334
rect -2273 174 -2003 306
rect -2273 146 -2149 174
rect -2121 146 -2003 174
rect -2273 14 -2003 146
rect -2273 -14 -2149 14
rect -2121 -14 -2003 14
rect -2273 -146 -2003 -14
rect -2273 -174 -2149 -146
rect -2121 -174 -2003 -146
rect -2273 -306 -2003 -174
rect -2273 -334 -2149 -306
rect -2121 -334 -2003 -306
rect -2273 -466 -2003 -334
rect -2273 -494 -2149 -466
rect -2121 -494 -2003 -466
rect -2273 -626 -2003 -494
rect -2273 -654 -2149 -626
rect -2121 -654 -2003 -626
rect -2273 -786 -2003 -654
rect -2273 -814 -2149 -786
rect -2121 -814 -2003 -786
rect -2273 -946 -2003 -814
rect -2273 -974 -2149 -946
rect -2121 -974 -2003 -946
rect -2273 -1106 -2003 -974
rect -2273 -1134 -2149 -1106
rect -2121 -1134 -2003 -1106
rect -2273 -1266 -2003 -1134
rect -2273 -1294 -2149 -1266
rect -2121 -1294 -2003 -1266
rect -2273 -1426 -2003 -1294
rect -2273 -1454 -2149 -1426
rect -2121 -1454 -2003 -1426
rect -2273 -1586 -2003 -1454
rect -2273 -1614 -2149 -1586
rect -2121 -1614 -2003 -1586
rect -2273 -1730 -2003 -1614
rect -6003 -1746 -2003 -1730
rect -6003 -1774 -5882 -1746
rect -5854 -1774 -2149 -1746
rect -2121 -1774 -2003 -1746
rect -6003 -1851 -2003 -1774
rect -6003 -1879 -5697 -1851
rect -5669 -1879 -5537 -1851
rect -5509 -1879 -5377 -1851
rect -5349 -1879 -5217 -1851
rect -5189 -1879 -5057 -1851
rect -5029 -1879 -4897 -1851
rect -4869 -1879 -4737 -1851
rect -4709 -1879 -4577 -1851
rect -4549 -1879 -4417 -1851
rect -4389 -1879 -4257 -1851
rect -4229 -1879 -4097 -1851
rect -4069 -1879 -3937 -1851
rect -3909 -1879 -3777 -1851
rect -3749 -1879 -3617 -1851
rect -3589 -1879 -3457 -1851
rect -3429 -1879 -3297 -1851
rect -3269 -1879 -3137 -1851
rect -3109 -1879 -2977 -1851
rect -2949 -1879 -2817 -1851
rect -2789 -1879 -2657 -1851
rect -2629 -1879 -2497 -1851
rect -2469 -1879 -2337 -1851
rect -2309 -1879 -2003 -1851
rect -6003 -2000 -2003 -1879
<< via2 >>
rect -5697 1876 -5669 1877
rect -5697 1850 -5696 1876
rect -5696 1850 -5670 1876
rect -5670 1850 -5669 1876
rect -5697 1849 -5669 1850
rect -5537 1876 -5509 1877
rect -5537 1850 -5536 1876
rect -5536 1850 -5510 1876
rect -5510 1850 -5509 1876
rect -5537 1849 -5509 1850
rect -5377 1876 -5349 1877
rect -5377 1850 -5376 1876
rect -5376 1850 -5350 1876
rect -5350 1850 -5349 1876
rect -5377 1849 -5349 1850
rect -5217 1876 -5189 1877
rect -5217 1850 -5216 1876
rect -5216 1850 -5190 1876
rect -5190 1850 -5189 1876
rect -5217 1849 -5189 1850
rect -5057 1876 -5029 1877
rect -5057 1850 -5056 1876
rect -5056 1850 -5030 1876
rect -5030 1850 -5029 1876
rect -5057 1849 -5029 1850
rect -4897 1876 -4869 1877
rect -4897 1850 -4896 1876
rect -4896 1850 -4870 1876
rect -4870 1850 -4869 1876
rect -4897 1849 -4869 1850
rect -4737 1876 -4709 1877
rect -4737 1850 -4736 1876
rect -4736 1850 -4710 1876
rect -4710 1850 -4709 1876
rect -4737 1849 -4709 1850
rect -4577 1876 -4549 1877
rect -4577 1850 -4576 1876
rect -4576 1850 -4550 1876
rect -4550 1850 -4549 1876
rect -4577 1849 -4549 1850
rect -4417 1876 -4389 1877
rect -4417 1850 -4416 1876
rect -4416 1850 -4390 1876
rect -4390 1850 -4389 1876
rect -4417 1849 -4389 1850
rect -4257 1876 -4229 1877
rect -4257 1850 -4256 1876
rect -4256 1850 -4230 1876
rect -4230 1850 -4229 1876
rect -4257 1849 -4229 1850
rect -4097 1876 -4069 1877
rect -4097 1850 -4096 1876
rect -4096 1850 -4070 1876
rect -4070 1850 -4069 1876
rect -4097 1849 -4069 1850
rect -3937 1876 -3909 1877
rect -3937 1850 -3936 1876
rect -3936 1850 -3910 1876
rect -3910 1850 -3909 1876
rect -3937 1849 -3909 1850
rect -3777 1876 -3749 1877
rect -3777 1850 -3776 1876
rect -3776 1850 -3750 1876
rect -3750 1850 -3749 1876
rect -3777 1849 -3749 1850
rect -3617 1876 -3589 1877
rect -3617 1850 -3616 1876
rect -3616 1850 -3590 1876
rect -3590 1850 -3589 1876
rect -3617 1849 -3589 1850
rect -3457 1876 -3429 1877
rect -3457 1850 -3456 1876
rect -3456 1850 -3430 1876
rect -3430 1850 -3429 1876
rect -3457 1849 -3429 1850
rect -3297 1876 -3269 1877
rect -3297 1850 -3296 1876
rect -3296 1850 -3270 1876
rect -3270 1850 -3269 1876
rect -3297 1849 -3269 1850
rect -3137 1876 -3109 1877
rect -3137 1850 -3136 1876
rect -3136 1850 -3110 1876
rect -3110 1850 -3109 1876
rect -3137 1849 -3109 1850
rect -2977 1876 -2949 1877
rect -2977 1850 -2976 1876
rect -2976 1850 -2950 1876
rect -2950 1850 -2949 1876
rect -2977 1849 -2949 1850
rect -2817 1876 -2789 1877
rect -2817 1850 -2816 1876
rect -2816 1850 -2790 1876
rect -2790 1850 -2789 1876
rect -2817 1849 -2789 1850
rect -2657 1876 -2629 1877
rect -2657 1850 -2656 1876
rect -2656 1850 -2630 1876
rect -2630 1850 -2629 1876
rect -2657 1849 -2629 1850
rect -2497 1876 -2469 1877
rect -2497 1850 -2496 1876
rect -2496 1850 -2470 1876
rect -2470 1850 -2469 1876
rect -2497 1849 -2469 1850
rect -2337 1876 -2309 1877
rect -2337 1850 -2336 1876
rect -2336 1850 -2310 1876
rect -2310 1850 -2309 1876
rect -2337 1849 -2309 1850
rect -5882 1773 -5854 1774
rect -5882 1747 -5881 1773
rect -5881 1747 -5855 1773
rect -5855 1747 -5854 1773
rect -5882 1746 -5854 1747
rect -2149 1773 -2121 1774
rect -2149 1747 -2148 1773
rect -2148 1747 -2122 1773
rect -2122 1747 -2121 1773
rect -2149 1746 -2121 1747
rect -5882 1613 -5854 1614
rect -5882 1587 -5881 1613
rect -5881 1587 -5855 1613
rect -5855 1587 -5854 1613
rect -5882 1586 -5854 1587
rect -5882 1453 -5854 1454
rect -5882 1427 -5881 1453
rect -5881 1427 -5855 1453
rect -5855 1427 -5854 1453
rect -5882 1426 -5854 1427
rect -5882 1293 -5854 1294
rect -5882 1267 -5881 1293
rect -5881 1267 -5855 1293
rect -5855 1267 -5854 1293
rect -5882 1266 -5854 1267
rect -5882 1133 -5854 1134
rect -5882 1107 -5881 1133
rect -5881 1107 -5855 1133
rect -5855 1107 -5854 1133
rect -5882 1106 -5854 1107
rect -5882 973 -5854 974
rect -5882 947 -5881 973
rect -5881 947 -5855 973
rect -5855 947 -5854 973
rect -5882 946 -5854 947
rect -5882 813 -5854 814
rect -5882 787 -5881 813
rect -5881 787 -5855 813
rect -5855 787 -5854 813
rect -5882 786 -5854 787
rect -5882 653 -5854 654
rect -5882 627 -5881 653
rect -5881 627 -5855 653
rect -5855 627 -5854 653
rect -5882 626 -5854 627
rect -5882 493 -5854 494
rect -5882 467 -5881 493
rect -5881 467 -5855 493
rect -5855 467 -5854 493
rect -5882 466 -5854 467
rect -5882 333 -5854 334
rect -5882 307 -5881 333
rect -5881 307 -5855 333
rect -5855 307 -5854 333
rect -5882 306 -5854 307
rect -5882 173 -5854 174
rect -5882 147 -5881 173
rect -5881 147 -5855 173
rect -5855 147 -5854 173
rect -5882 146 -5854 147
rect -5882 13 -5854 14
rect -5882 -13 -5881 13
rect -5881 -13 -5855 13
rect -5855 -13 -5854 13
rect -5882 -14 -5854 -13
rect -5882 -147 -5854 -146
rect -5882 -173 -5881 -147
rect -5881 -173 -5855 -147
rect -5855 -173 -5854 -147
rect -5882 -174 -5854 -173
rect -5882 -307 -5854 -306
rect -5882 -333 -5881 -307
rect -5881 -333 -5855 -307
rect -5855 -333 -5854 -307
rect -5882 -334 -5854 -333
rect -5882 -467 -5854 -466
rect -5882 -493 -5881 -467
rect -5881 -493 -5855 -467
rect -5855 -493 -5854 -467
rect -5882 -494 -5854 -493
rect -5882 -627 -5854 -626
rect -5882 -653 -5881 -627
rect -5881 -653 -5855 -627
rect -5855 -653 -5854 -627
rect -5882 -654 -5854 -653
rect -5882 -787 -5854 -786
rect -5882 -813 -5881 -787
rect -5881 -813 -5855 -787
rect -5855 -813 -5854 -787
rect -5882 -814 -5854 -813
rect -5882 -947 -5854 -946
rect -5882 -973 -5881 -947
rect -5881 -973 -5855 -947
rect -5855 -973 -5854 -947
rect -5882 -974 -5854 -973
rect -5882 -1107 -5854 -1106
rect -5882 -1133 -5881 -1107
rect -5881 -1133 -5855 -1107
rect -5855 -1133 -5854 -1107
rect -5882 -1134 -5854 -1133
rect -5882 -1267 -5854 -1266
rect -5882 -1293 -5881 -1267
rect -5881 -1293 -5855 -1267
rect -5855 -1293 -5854 -1267
rect -5882 -1294 -5854 -1293
rect -5882 -1427 -5854 -1426
rect -5882 -1453 -5881 -1427
rect -5881 -1453 -5855 -1427
rect -5855 -1453 -5854 -1427
rect -5882 -1454 -5854 -1453
rect -5882 -1587 -5854 -1586
rect -5882 -1613 -5881 -1587
rect -5881 -1613 -5855 -1587
rect -5855 -1613 -5854 -1587
rect -5882 -1614 -5854 -1613
rect -2149 1613 -2121 1614
rect -2149 1587 -2148 1613
rect -2148 1587 -2122 1613
rect -2122 1587 -2121 1613
rect -2149 1586 -2121 1587
rect -2149 1453 -2121 1454
rect -2149 1427 -2148 1453
rect -2148 1427 -2122 1453
rect -2122 1427 -2121 1453
rect -2149 1426 -2121 1427
rect -2149 1293 -2121 1294
rect -2149 1267 -2148 1293
rect -2148 1267 -2122 1293
rect -2122 1267 -2121 1293
rect -2149 1266 -2121 1267
rect -2149 1133 -2121 1134
rect -2149 1107 -2148 1133
rect -2148 1107 -2122 1133
rect -2122 1107 -2121 1133
rect -2149 1106 -2121 1107
rect -2149 973 -2121 974
rect -2149 947 -2148 973
rect -2148 947 -2122 973
rect -2122 947 -2121 973
rect -2149 946 -2121 947
rect -2149 813 -2121 814
rect -2149 787 -2148 813
rect -2148 787 -2122 813
rect -2122 787 -2121 813
rect -2149 786 -2121 787
rect -2149 653 -2121 654
rect -2149 627 -2148 653
rect -2148 627 -2122 653
rect -2122 627 -2121 653
rect -2149 626 -2121 627
rect -2149 493 -2121 494
rect -2149 467 -2148 493
rect -2148 467 -2122 493
rect -2122 467 -2121 493
rect -2149 466 -2121 467
rect -2149 333 -2121 334
rect -2149 307 -2148 333
rect -2148 307 -2122 333
rect -2122 307 -2121 333
rect -2149 306 -2121 307
rect -2149 173 -2121 174
rect -2149 147 -2148 173
rect -2148 147 -2122 173
rect -2122 147 -2121 173
rect -2149 146 -2121 147
rect -2149 13 -2121 14
rect -2149 -13 -2148 13
rect -2148 -13 -2122 13
rect -2122 -13 -2121 13
rect -2149 -14 -2121 -13
rect -2149 -147 -2121 -146
rect -2149 -173 -2148 -147
rect -2148 -173 -2122 -147
rect -2122 -173 -2121 -147
rect -2149 -174 -2121 -173
rect -2149 -307 -2121 -306
rect -2149 -333 -2148 -307
rect -2148 -333 -2122 -307
rect -2122 -333 -2121 -307
rect -2149 -334 -2121 -333
rect -2149 -467 -2121 -466
rect -2149 -493 -2148 -467
rect -2148 -493 -2122 -467
rect -2122 -493 -2121 -467
rect -2149 -494 -2121 -493
rect -2149 -627 -2121 -626
rect -2149 -653 -2148 -627
rect -2148 -653 -2122 -627
rect -2122 -653 -2121 -627
rect -2149 -654 -2121 -653
rect -2149 -787 -2121 -786
rect -2149 -813 -2148 -787
rect -2148 -813 -2122 -787
rect -2122 -813 -2121 -787
rect -2149 -814 -2121 -813
rect -2149 -947 -2121 -946
rect -2149 -973 -2148 -947
rect -2148 -973 -2122 -947
rect -2122 -973 -2121 -947
rect -2149 -974 -2121 -973
rect -2149 -1107 -2121 -1106
rect -2149 -1133 -2148 -1107
rect -2148 -1133 -2122 -1107
rect -2122 -1133 -2121 -1107
rect -2149 -1134 -2121 -1133
rect -2149 -1267 -2121 -1266
rect -2149 -1293 -2148 -1267
rect -2148 -1293 -2122 -1267
rect -2122 -1293 -2121 -1267
rect -2149 -1294 -2121 -1293
rect -2149 -1427 -2121 -1426
rect -2149 -1453 -2148 -1427
rect -2148 -1453 -2122 -1427
rect -2122 -1453 -2121 -1427
rect -2149 -1454 -2121 -1453
rect -2149 -1587 -2121 -1586
rect -2149 -1613 -2148 -1587
rect -2148 -1613 -2122 -1587
rect -2122 -1613 -2121 -1587
rect -2149 -1614 -2121 -1613
rect -5882 -1747 -5854 -1746
rect -5882 -1773 -5881 -1747
rect -5881 -1773 -5855 -1747
rect -5855 -1773 -5854 -1747
rect -5882 -1774 -5854 -1773
rect -2149 -1747 -2121 -1746
rect -2149 -1773 -2148 -1747
rect -2148 -1773 -2122 -1747
rect -2122 -1773 -2121 -1747
rect -2149 -1774 -2121 -1773
rect -5697 -1852 -5669 -1851
rect -5697 -1878 -5696 -1852
rect -5696 -1878 -5670 -1852
rect -5670 -1878 -5669 -1852
rect -5697 -1879 -5669 -1878
rect -5537 -1852 -5509 -1851
rect -5537 -1878 -5536 -1852
rect -5536 -1878 -5510 -1852
rect -5510 -1878 -5509 -1852
rect -5537 -1879 -5509 -1878
rect -5377 -1852 -5349 -1851
rect -5377 -1878 -5376 -1852
rect -5376 -1878 -5350 -1852
rect -5350 -1878 -5349 -1852
rect -5377 -1879 -5349 -1878
rect -5217 -1852 -5189 -1851
rect -5217 -1878 -5216 -1852
rect -5216 -1878 -5190 -1852
rect -5190 -1878 -5189 -1852
rect -5217 -1879 -5189 -1878
rect -5057 -1852 -5029 -1851
rect -5057 -1878 -5056 -1852
rect -5056 -1878 -5030 -1852
rect -5030 -1878 -5029 -1852
rect -5057 -1879 -5029 -1878
rect -4897 -1852 -4869 -1851
rect -4897 -1878 -4896 -1852
rect -4896 -1878 -4870 -1852
rect -4870 -1878 -4869 -1852
rect -4897 -1879 -4869 -1878
rect -4737 -1852 -4709 -1851
rect -4737 -1878 -4736 -1852
rect -4736 -1878 -4710 -1852
rect -4710 -1878 -4709 -1852
rect -4737 -1879 -4709 -1878
rect -4577 -1852 -4549 -1851
rect -4577 -1878 -4576 -1852
rect -4576 -1878 -4550 -1852
rect -4550 -1878 -4549 -1852
rect -4577 -1879 -4549 -1878
rect -4417 -1852 -4389 -1851
rect -4417 -1878 -4416 -1852
rect -4416 -1878 -4390 -1852
rect -4390 -1878 -4389 -1852
rect -4417 -1879 -4389 -1878
rect -4257 -1852 -4229 -1851
rect -4257 -1878 -4256 -1852
rect -4256 -1878 -4230 -1852
rect -4230 -1878 -4229 -1852
rect -4257 -1879 -4229 -1878
rect -4097 -1852 -4069 -1851
rect -4097 -1878 -4096 -1852
rect -4096 -1878 -4070 -1852
rect -4070 -1878 -4069 -1852
rect -4097 -1879 -4069 -1878
rect -3937 -1852 -3909 -1851
rect -3937 -1878 -3936 -1852
rect -3936 -1878 -3910 -1852
rect -3910 -1878 -3909 -1852
rect -3937 -1879 -3909 -1878
rect -3777 -1852 -3749 -1851
rect -3777 -1878 -3776 -1852
rect -3776 -1878 -3750 -1852
rect -3750 -1878 -3749 -1852
rect -3777 -1879 -3749 -1878
rect -3617 -1852 -3589 -1851
rect -3617 -1878 -3616 -1852
rect -3616 -1878 -3590 -1852
rect -3590 -1878 -3589 -1852
rect -3617 -1879 -3589 -1878
rect -3457 -1852 -3429 -1851
rect -3457 -1878 -3456 -1852
rect -3456 -1878 -3430 -1852
rect -3430 -1878 -3429 -1852
rect -3457 -1879 -3429 -1878
rect -3297 -1852 -3269 -1851
rect -3297 -1878 -3296 -1852
rect -3296 -1878 -3270 -1852
rect -3270 -1878 -3269 -1852
rect -3297 -1879 -3269 -1878
rect -3137 -1852 -3109 -1851
rect -3137 -1878 -3136 -1852
rect -3136 -1878 -3110 -1852
rect -3110 -1878 -3109 -1852
rect -3137 -1879 -3109 -1878
rect -2977 -1852 -2949 -1851
rect -2977 -1878 -2976 -1852
rect -2976 -1878 -2950 -1852
rect -2950 -1878 -2949 -1852
rect -2977 -1879 -2949 -1878
rect -2817 -1852 -2789 -1851
rect -2817 -1878 -2816 -1852
rect -2816 -1878 -2790 -1852
rect -2790 -1878 -2789 -1852
rect -2817 -1879 -2789 -1878
rect -2657 -1852 -2629 -1851
rect -2657 -1878 -2656 -1852
rect -2656 -1878 -2630 -1852
rect -2630 -1878 -2629 -1852
rect -2657 -1879 -2629 -1878
rect -2497 -1852 -2469 -1851
rect -2497 -1878 -2496 -1852
rect -2496 -1878 -2470 -1852
rect -2470 -1878 -2469 -1852
rect -2497 -1879 -2469 -1878
rect -2337 -1852 -2309 -1851
rect -2337 -1878 -2336 -1852
rect -2336 -1878 -2310 -1852
rect -2310 -1878 -2309 -1852
rect -2337 -1879 -2309 -1878
<< metal3 >>
rect -6003 1879 -2003 2000
rect -6003 1847 -5699 1879
rect -5667 1847 -5539 1879
rect -5507 1847 -5379 1879
rect -5347 1847 -5219 1879
rect -5187 1847 -5059 1879
rect -5027 1847 -4899 1879
rect -4867 1847 -4739 1879
rect -4707 1847 -4579 1879
rect -4547 1847 -4419 1879
rect -4387 1847 -4259 1879
rect -4227 1847 -4099 1879
rect -4067 1847 -3939 1879
rect -3907 1847 -3779 1879
rect -3747 1847 -3619 1879
rect -3587 1847 -3459 1879
rect -3427 1847 -3299 1879
rect -3267 1847 -3139 1879
rect -3107 1847 -2979 1879
rect -2947 1847 -2819 1879
rect -2787 1847 -2659 1879
rect -2627 1847 -2499 1879
rect -2467 1847 -2339 1879
rect -2307 1847 -2003 1879
rect -6003 1776 -2003 1847
rect -6003 1744 -5884 1776
rect -5852 1744 -2151 1776
rect -2119 1744 -2003 1776
rect -6003 1730 -2003 1744
rect -6003 1616 -5733 1730
rect -6003 1584 -5884 1616
rect -5852 1584 -5733 1616
rect -6003 1456 -5733 1584
rect -6003 1424 -5884 1456
rect -5852 1424 -5733 1456
rect -6003 1296 -5733 1424
rect -6003 1264 -5884 1296
rect -5852 1264 -5733 1296
rect -6003 1136 -5733 1264
rect -6003 1104 -5884 1136
rect -5852 1104 -5733 1136
rect -6003 976 -5733 1104
rect -6003 944 -5884 976
rect -5852 944 -5733 976
rect -6003 816 -5733 944
rect -6003 784 -5884 816
rect -5852 784 -5733 816
rect -6003 656 -5733 784
rect -6003 624 -5884 656
rect -5852 624 -5733 656
rect -6003 496 -5733 624
rect -6003 464 -5884 496
rect -5852 464 -5733 496
rect -6003 336 -5733 464
rect -6003 304 -5884 336
rect -5852 304 -5733 336
rect -6003 176 -5733 304
rect -6003 144 -5884 176
rect -5852 144 -5733 176
rect -6003 16 -5733 144
rect -6003 -16 -5884 16
rect -5852 -16 -5733 16
rect -6003 -144 -5733 -16
rect -6003 -176 -5884 -144
rect -5852 -176 -5733 -144
rect -6003 -304 -5733 -176
rect -6003 -336 -5884 -304
rect -5852 -336 -5733 -304
rect -6003 -464 -5733 -336
rect -6003 -496 -5884 -464
rect -5852 -496 -5733 -464
rect -6003 -624 -5733 -496
rect -6003 -656 -5884 -624
rect -5852 -656 -5733 -624
rect -6003 -784 -5733 -656
rect -6003 -816 -5884 -784
rect -5852 -816 -5733 -784
rect -6003 -944 -5733 -816
rect -6003 -976 -5884 -944
rect -5852 -976 -5733 -944
rect -6003 -1104 -5733 -976
rect -6003 -1136 -5884 -1104
rect -5852 -1136 -5733 -1104
rect -6003 -1264 -5733 -1136
rect -6003 -1296 -5884 -1264
rect -5852 -1296 -5733 -1264
rect -6003 -1424 -5733 -1296
rect -6003 -1456 -5884 -1424
rect -5852 -1456 -5733 -1424
rect -6003 -1584 -5733 -1456
rect -6003 -1616 -5884 -1584
rect -5852 -1616 -5733 -1584
rect -6003 -1730 -5733 -1616
rect -2273 1616 -2003 1730
rect -2273 1584 -2151 1616
rect -2119 1584 -2003 1616
rect -2273 1456 -2003 1584
rect -2273 1424 -2151 1456
rect -2119 1424 -2003 1456
rect -2273 1296 -2003 1424
rect -2273 1264 -2151 1296
rect -2119 1264 -2003 1296
rect -2273 1136 -2003 1264
rect -2273 1104 -2151 1136
rect -2119 1104 -2003 1136
rect -2273 976 -2003 1104
rect -2273 944 -2151 976
rect -2119 944 -2003 976
rect -2273 816 -2003 944
rect -2273 784 -2151 816
rect -2119 784 -2003 816
rect -2273 656 -2003 784
rect -2273 624 -2151 656
rect -2119 624 -2003 656
rect -2273 496 -2003 624
rect -2273 464 -2151 496
rect -2119 464 -2003 496
rect -2273 336 -2003 464
rect -2273 304 -2151 336
rect -2119 304 -2003 336
rect -2273 176 -2003 304
rect -2273 144 -2151 176
rect -2119 144 -2003 176
rect -2273 16 -2003 144
rect -2273 -16 -2151 16
rect -2119 -16 -2003 16
rect -2273 -144 -2003 -16
rect -2273 -176 -2151 -144
rect -2119 -176 -2003 -144
rect -2273 -304 -2003 -176
rect -2273 -336 -2151 -304
rect -2119 -336 -2003 -304
rect -2273 -464 -2003 -336
rect -2273 -496 -2151 -464
rect -2119 -496 -2003 -464
rect -2273 -624 -2003 -496
rect -2273 -656 -2151 -624
rect -2119 -656 -2003 -624
rect -2273 -784 -2003 -656
rect -2273 -816 -2151 -784
rect -2119 -816 -2003 -784
rect -2273 -944 -2003 -816
rect -2273 -976 -2151 -944
rect -2119 -976 -2003 -944
rect -2273 -1104 -2003 -976
rect -2273 -1136 -2151 -1104
rect -2119 -1136 -2003 -1104
rect -2273 -1264 -2003 -1136
rect -2273 -1296 -2151 -1264
rect -2119 -1296 -2003 -1264
rect -2273 -1424 -2003 -1296
rect -2273 -1456 -2151 -1424
rect -2119 -1456 -2003 -1424
rect -2273 -1584 -2003 -1456
rect -2273 -1616 -2151 -1584
rect -2119 -1616 -2003 -1584
rect -2273 -1730 -2003 -1616
rect -6003 -1744 -2003 -1730
rect -6003 -1776 -5884 -1744
rect -5852 -1776 -2151 -1744
rect -2119 -1776 -2003 -1744
rect -6003 -1849 -2003 -1776
rect -6003 -1881 -5699 -1849
rect -5667 -1881 -5539 -1849
rect -5507 -1881 -5379 -1849
rect -5347 -1881 -5219 -1849
rect -5187 -1881 -5059 -1849
rect -5027 -1881 -4899 -1849
rect -4867 -1881 -4739 -1849
rect -4707 -1881 -4579 -1849
rect -4547 -1881 -4419 -1849
rect -4387 -1881 -4259 -1849
rect -4227 -1881 -4099 -1849
rect -4067 -1881 -3939 -1849
rect -3907 -1881 -3779 -1849
rect -3747 -1881 -3619 -1849
rect -3587 -1881 -3459 -1849
rect -3427 -1881 -3299 -1849
rect -3267 -1881 -3139 -1849
rect -3107 -1881 -2979 -1849
rect -2947 -1881 -2819 -1849
rect -2787 -1881 -2659 -1849
rect -2627 -1881 -2499 -1849
rect -2467 -1881 -2339 -1849
rect -2307 -1881 -2003 -1849
rect -6003 -2000 -2003 -1881
<< via3 >>
rect -5699 1877 -5667 1879
rect -5699 1849 -5697 1877
rect -5697 1849 -5669 1877
rect -5669 1849 -5667 1877
rect -5699 1847 -5667 1849
rect -5539 1877 -5507 1879
rect -5539 1849 -5537 1877
rect -5537 1849 -5509 1877
rect -5509 1849 -5507 1877
rect -5539 1847 -5507 1849
rect -5379 1877 -5347 1879
rect -5379 1849 -5377 1877
rect -5377 1849 -5349 1877
rect -5349 1849 -5347 1877
rect -5379 1847 -5347 1849
rect -5219 1877 -5187 1879
rect -5219 1849 -5217 1877
rect -5217 1849 -5189 1877
rect -5189 1849 -5187 1877
rect -5219 1847 -5187 1849
rect -5059 1877 -5027 1879
rect -5059 1849 -5057 1877
rect -5057 1849 -5029 1877
rect -5029 1849 -5027 1877
rect -5059 1847 -5027 1849
rect -4899 1877 -4867 1879
rect -4899 1849 -4897 1877
rect -4897 1849 -4869 1877
rect -4869 1849 -4867 1877
rect -4899 1847 -4867 1849
rect -4739 1877 -4707 1879
rect -4739 1849 -4737 1877
rect -4737 1849 -4709 1877
rect -4709 1849 -4707 1877
rect -4739 1847 -4707 1849
rect -4579 1877 -4547 1879
rect -4579 1849 -4577 1877
rect -4577 1849 -4549 1877
rect -4549 1849 -4547 1877
rect -4579 1847 -4547 1849
rect -4419 1877 -4387 1879
rect -4419 1849 -4417 1877
rect -4417 1849 -4389 1877
rect -4389 1849 -4387 1877
rect -4419 1847 -4387 1849
rect -4259 1877 -4227 1879
rect -4259 1849 -4257 1877
rect -4257 1849 -4229 1877
rect -4229 1849 -4227 1877
rect -4259 1847 -4227 1849
rect -4099 1877 -4067 1879
rect -4099 1849 -4097 1877
rect -4097 1849 -4069 1877
rect -4069 1849 -4067 1877
rect -4099 1847 -4067 1849
rect -3939 1877 -3907 1879
rect -3939 1849 -3937 1877
rect -3937 1849 -3909 1877
rect -3909 1849 -3907 1877
rect -3939 1847 -3907 1849
rect -3779 1877 -3747 1879
rect -3779 1849 -3777 1877
rect -3777 1849 -3749 1877
rect -3749 1849 -3747 1877
rect -3779 1847 -3747 1849
rect -3619 1877 -3587 1879
rect -3619 1849 -3617 1877
rect -3617 1849 -3589 1877
rect -3589 1849 -3587 1877
rect -3619 1847 -3587 1849
rect -3459 1877 -3427 1879
rect -3459 1849 -3457 1877
rect -3457 1849 -3429 1877
rect -3429 1849 -3427 1877
rect -3459 1847 -3427 1849
rect -3299 1877 -3267 1879
rect -3299 1849 -3297 1877
rect -3297 1849 -3269 1877
rect -3269 1849 -3267 1877
rect -3299 1847 -3267 1849
rect -3139 1877 -3107 1879
rect -3139 1849 -3137 1877
rect -3137 1849 -3109 1877
rect -3109 1849 -3107 1877
rect -3139 1847 -3107 1849
rect -2979 1877 -2947 1879
rect -2979 1849 -2977 1877
rect -2977 1849 -2949 1877
rect -2949 1849 -2947 1877
rect -2979 1847 -2947 1849
rect -2819 1877 -2787 1879
rect -2819 1849 -2817 1877
rect -2817 1849 -2789 1877
rect -2789 1849 -2787 1877
rect -2819 1847 -2787 1849
rect -2659 1877 -2627 1879
rect -2659 1849 -2657 1877
rect -2657 1849 -2629 1877
rect -2629 1849 -2627 1877
rect -2659 1847 -2627 1849
rect -2499 1877 -2467 1879
rect -2499 1849 -2497 1877
rect -2497 1849 -2469 1877
rect -2469 1849 -2467 1877
rect -2499 1847 -2467 1849
rect -2339 1877 -2307 1879
rect -2339 1849 -2337 1877
rect -2337 1849 -2309 1877
rect -2309 1849 -2307 1877
rect -2339 1847 -2307 1849
rect -5884 1774 -5852 1776
rect -5884 1746 -5882 1774
rect -5882 1746 -5854 1774
rect -5854 1746 -5852 1774
rect -5884 1744 -5852 1746
rect -2151 1774 -2119 1776
rect -2151 1746 -2149 1774
rect -2149 1746 -2121 1774
rect -2121 1746 -2119 1774
rect -2151 1744 -2119 1746
rect -5884 1614 -5852 1616
rect -5884 1586 -5882 1614
rect -5882 1586 -5854 1614
rect -5854 1586 -5852 1614
rect -5884 1584 -5852 1586
rect -5884 1454 -5852 1456
rect -5884 1426 -5882 1454
rect -5882 1426 -5854 1454
rect -5854 1426 -5852 1454
rect -5884 1424 -5852 1426
rect -5884 1294 -5852 1296
rect -5884 1266 -5882 1294
rect -5882 1266 -5854 1294
rect -5854 1266 -5852 1294
rect -5884 1264 -5852 1266
rect -5884 1134 -5852 1136
rect -5884 1106 -5882 1134
rect -5882 1106 -5854 1134
rect -5854 1106 -5852 1134
rect -5884 1104 -5852 1106
rect -5884 974 -5852 976
rect -5884 946 -5882 974
rect -5882 946 -5854 974
rect -5854 946 -5852 974
rect -5884 944 -5852 946
rect -5884 814 -5852 816
rect -5884 786 -5882 814
rect -5882 786 -5854 814
rect -5854 786 -5852 814
rect -5884 784 -5852 786
rect -5884 654 -5852 656
rect -5884 626 -5882 654
rect -5882 626 -5854 654
rect -5854 626 -5852 654
rect -5884 624 -5852 626
rect -5884 494 -5852 496
rect -5884 466 -5882 494
rect -5882 466 -5854 494
rect -5854 466 -5852 494
rect -5884 464 -5852 466
rect -5884 334 -5852 336
rect -5884 306 -5882 334
rect -5882 306 -5854 334
rect -5854 306 -5852 334
rect -5884 304 -5852 306
rect -5884 174 -5852 176
rect -5884 146 -5882 174
rect -5882 146 -5854 174
rect -5854 146 -5852 174
rect -5884 144 -5852 146
rect -5884 14 -5852 16
rect -5884 -14 -5882 14
rect -5882 -14 -5854 14
rect -5854 -14 -5852 14
rect -5884 -16 -5852 -14
rect -5884 -146 -5852 -144
rect -5884 -174 -5882 -146
rect -5882 -174 -5854 -146
rect -5854 -174 -5852 -146
rect -5884 -176 -5852 -174
rect -5884 -306 -5852 -304
rect -5884 -334 -5882 -306
rect -5882 -334 -5854 -306
rect -5854 -334 -5852 -306
rect -5884 -336 -5852 -334
rect -5884 -466 -5852 -464
rect -5884 -494 -5882 -466
rect -5882 -494 -5854 -466
rect -5854 -494 -5852 -466
rect -5884 -496 -5852 -494
rect -5884 -626 -5852 -624
rect -5884 -654 -5882 -626
rect -5882 -654 -5854 -626
rect -5854 -654 -5852 -626
rect -5884 -656 -5852 -654
rect -5884 -786 -5852 -784
rect -5884 -814 -5882 -786
rect -5882 -814 -5854 -786
rect -5854 -814 -5852 -786
rect -5884 -816 -5852 -814
rect -5884 -946 -5852 -944
rect -5884 -974 -5882 -946
rect -5882 -974 -5854 -946
rect -5854 -974 -5852 -946
rect -5884 -976 -5852 -974
rect -5884 -1106 -5852 -1104
rect -5884 -1134 -5882 -1106
rect -5882 -1134 -5854 -1106
rect -5854 -1134 -5852 -1106
rect -5884 -1136 -5852 -1134
rect -5884 -1266 -5852 -1264
rect -5884 -1294 -5882 -1266
rect -5882 -1294 -5854 -1266
rect -5854 -1294 -5852 -1266
rect -5884 -1296 -5852 -1294
rect -5884 -1426 -5852 -1424
rect -5884 -1454 -5882 -1426
rect -5882 -1454 -5854 -1426
rect -5854 -1454 -5852 -1426
rect -5884 -1456 -5852 -1454
rect -5884 -1586 -5852 -1584
rect -5884 -1614 -5882 -1586
rect -5882 -1614 -5854 -1586
rect -5854 -1614 -5852 -1586
rect -5884 -1616 -5852 -1614
rect -2151 1614 -2119 1616
rect -2151 1586 -2149 1614
rect -2149 1586 -2121 1614
rect -2121 1586 -2119 1614
rect -2151 1584 -2119 1586
rect -2151 1454 -2119 1456
rect -2151 1426 -2149 1454
rect -2149 1426 -2121 1454
rect -2121 1426 -2119 1454
rect -2151 1424 -2119 1426
rect -2151 1294 -2119 1296
rect -2151 1266 -2149 1294
rect -2149 1266 -2121 1294
rect -2121 1266 -2119 1294
rect -2151 1264 -2119 1266
rect -2151 1134 -2119 1136
rect -2151 1106 -2149 1134
rect -2149 1106 -2121 1134
rect -2121 1106 -2119 1134
rect -2151 1104 -2119 1106
rect -2151 974 -2119 976
rect -2151 946 -2149 974
rect -2149 946 -2121 974
rect -2121 946 -2119 974
rect -2151 944 -2119 946
rect -2151 814 -2119 816
rect -2151 786 -2149 814
rect -2149 786 -2121 814
rect -2121 786 -2119 814
rect -2151 784 -2119 786
rect -2151 654 -2119 656
rect -2151 626 -2149 654
rect -2149 626 -2121 654
rect -2121 626 -2119 654
rect -2151 624 -2119 626
rect -2151 494 -2119 496
rect -2151 466 -2149 494
rect -2149 466 -2121 494
rect -2121 466 -2119 494
rect -2151 464 -2119 466
rect -2151 334 -2119 336
rect -2151 306 -2149 334
rect -2149 306 -2121 334
rect -2121 306 -2119 334
rect -2151 304 -2119 306
rect -2151 174 -2119 176
rect -2151 146 -2149 174
rect -2149 146 -2121 174
rect -2121 146 -2119 174
rect -2151 144 -2119 146
rect -2151 14 -2119 16
rect -2151 -14 -2149 14
rect -2149 -14 -2121 14
rect -2121 -14 -2119 14
rect -2151 -16 -2119 -14
rect -2151 -146 -2119 -144
rect -2151 -174 -2149 -146
rect -2149 -174 -2121 -146
rect -2121 -174 -2119 -146
rect -2151 -176 -2119 -174
rect -2151 -306 -2119 -304
rect -2151 -334 -2149 -306
rect -2149 -334 -2121 -306
rect -2121 -334 -2119 -306
rect -2151 -336 -2119 -334
rect -2151 -466 -2119 -464
rect -2151 -494 -2149 -466
rect -2149 -494 -2121 -466
rect -2121 -494 -2119 -466
rect -2151 -496 -2119 -494
rect -2151 -626 -2119 -624
rect -2151 -654 -2149 -626
rect -2149 -654 -2121 -626
rect -2121 -654 -2119 -626
rect -2151 -656 -2119 -654
rect -2151 -786 -2119 -784
rect -2151 -814 -2149 -786
rect -2149 -814 -2121 -786
rect -2121 -814 -2119 -786
rect -2151 -816 -2119 -814
rect -2151 -946 -2119 -944
rect -2151 -974 -2149 -946
rect -2149 -974 -2121 -946
rect -2121 -974 -2119 -946
rect -2151 -976 -2119 -974
rect -2151 -1106 -2119 -1104
rect -2151 -1134 -2149 -1106
rect -2149 -1134 -2121 -1106
rect -2121 -1134 -2119 -1106
rect -2151 -1136 -2119 -1134
rect -2151 -1266 -2119 -1264
rect -2151 -1294 -2149 -1266
rect -2149 -1294 -2121 -1266
rect -2121 -1294 -2119 -1266
rect -2151 -1296 -2119 -1294
rect -2151 -1426 -2119 -1424
rect -2151 -1454 -2149 -1426
rect -2149 -1454 -2121 -1426
rect -2121 -1454 -2119 -1426
rect -2151 -1456 -2119 -1454
rect -2151 -1586 -2119 -1584
rect -2151 -1614 -2149 -1586
rect -2149 -1614 -2121 -1586
rect -2121 -1614 -2119 -1586
rect -2151 -1616 -2119 -1614
rect -5884 -1746 -5852 -1744
rect -5884 -1774 -5882 -1746
rect -5882 -1774 -5854 -1746
rect -5854 -1774 -5852 -1746
rect -5884 -1776 -5852 -1774
rect -2151 -1746 -2119 -1744
rect -2151 -1774 -2149 -1746
rect -2149 -1774 -2121 -1746
rect -2121 -1774 -2119 -1746
rect -2151 -1776 -2119 -1774
rect -5699 -1851 -5667 -1849
rect -5699 -1879 -5697 -1851
rect -5697 -1879 -5669 -1851
rect -5669 -1879 -5667 -1851
rect -5699 -1881 -5667 -1879
rect -5539 -1851 -5507 -1849
rect -5539 -1879 -5537 -1851
rect -5537 -1879 -5509 -1851
rect -5509 -1879 -5507 -1851
rect -5539 -1881 -5507 -1879
rect -5379 -1851 -5347 -1849
rect -5379 -1879 -5377 -1851
rect -5377 -1879 -5349 -1851
rect -5349 -1879 -5347 -1851
rect -5379 -1881 -5347 -1879
rect -5219 -1851 -5187 -1849
rect -5219 -1879 -5217 -1851
rect -5217 -1879 -5189 -1851
rect -5189 -1879 -5187 -1851
rect -5219 -1881 -5187 -1879
rect -5059 -1851 -5027 -1849
rect -5059 -1879 -5057 -1851
rect -5057 -1879 -5029 -1851
rect -5029 -1879 -5027 -1851
rect -5059 -1881 -5027 -1879
rect -4899 -1851 -4867 -1849
rect -4899 -1879 -4897 -1851
rect -4897 -1879 -4869 -1851
rect -4869 -1879 -4867 -1851
rect -4899 -1881 -4867 -1879
rect -4739 -1851 -4707 -1849
rect -4739 -1879 -4737 -1851
rect -4737 -1879 -4709 -1851
rect -4709 -1879 -4707 -1851
rect -4739 -1881 -4707 -1879
rect -4579 -1851 -4547 -1849
rect -4579 -1879 -4577 -1851
rect -4577 -1879 -4549 -1851
rect -4549 -1879 -4547 -1851
rect -4579 -1881 -4547 -1879
rect -4419 -1851 -4387 -1849
rect -4419 -1879 -4417 -1851
rect -4417 -1879 -4389 -1851
rect -4389 -1879 -4387 -1851
rect -4419 -1881 -4387 -1879
rect -4259 -1851 -4227 -1849
rect -4259 -1879 -4257 -1851
rect -4257 -1879 -4229 -1851
rect -4229 -1879 -4227 -1851
rect -4259 -1881 -4227 -1879
rect -4099 -1851 -4067 -1849
rect -4099 -1879 -4097 -1851
rect -4097 -1879 -4069 -1851
rect -4069 -1879 -4067 -1851
rect -4099 -1881 -4067 -1879
rect -3939 -1851 -3907 -1849
rect -3939 -1879 -3937 -1851
rect -3937 -1879 -3909 -1851
rect -3909 -1879 -3907 -1851
rect -3939 -1881 -3907 -1879
rect -3779 -1851 -3747 -1849
rect -3779 -1879 -3777 -1851
rect -3777 -1879 -3749 -1851
rect -3749 -1879 -3747 -1851
rect -3779 -1881 -3747 -1879
rect -3619 -1851 -3587 -1849
rect -3619 -1879 -3617 -1851
rect -3617 -1879 -3589 -1851
rect -3589 -1879 -3587 -1851
rect -3619 -1881 -3587 -1879
rect -3459 -1851 -3427 -1849
rect -3459 -1879 -3457 -1851
rect -3457 -1879 -3429 -1851
rect -3429 -1879 -3427 -1851
rect -3459 -1881 -3427 -1879
rect -3299 -1851 -3267 -1849
rect -3299 -1879 -3297 -1851
rect -3297 -1879 -3269 -1851
rect -3269 -1879 -3267 -1851
rect -3299 -1881 -3267 -1879
rect -3139 -1851 -3107 -1849
rect -3139 -1879 -3137 -1851
rect -3137 -1879 -3109 -1851
rect -3109 -1879 -3107 -1851
rect -3139 -1881 -3107 -1879
rect -2979 -1851 -2947 -1849
rect -2979 -1879 -2977 -1851
rect -2977 -1879 -2949 -1851
rect -2949 -1879 -2947 -1851
rect -2979 -1881 -2947 -1879
rect -2819 -1851 -2787 -1849
rect -2819 -1879 -2817 -1851
rect -2817 -1879 -2789 -1851
rect -2789 -1879 -2787 -1851
rect -2819 -1881 -2787 -1879
rect -2659 -1851 -2627 -1849
rect -2659 -1879 -2657 -1851
rect -2657 -1879 -2629 -1851
rect -2629 -1879 -2627 -1851
rect -2659 -1881 -2627 -1879
rect -2499 -1851 -2467 -1849
rect -2499 -1879 -2497 -1851
rect -2497 -1879 -2469 -1851
rect -2469 -1879 -2467 -1851
rect -2499 -1881 -2467 -1879
rect -2339 -1851 -2307 -1849
rect -2339 -1879 -2337 -1851
rect -2337 -1879 -2309 -1851
rect -2309 -1879 -2307 -1851
rect -2339 -1881 -2307 -1879
<< metal4 >>
rect -6003 1922 -2003 2000
rect -6003 1819 -5742 1922
rect -6003 1701 -5927 1819
rect -5809 1804 -5742 1819
rect -5624 1804 -5582 1922
rect -5464 1804 -5422 1922
rect -5304 1804 -5262 1922
rect -5144 1804 -5102 1922
rect -4984 1804 -4942 1922
rect -4824 1804 -4782 1922
rect -4664 1804 -4622 1922
rect -4504 1804 -4462 1922
rect -4344 1804 -4302 1922
rect -4184 1804 -4142 1922
rect -4024 1804 -3982 1922
rect -3864 1804 -3822 1922
rect -3704 1804 -3662 1922
rect -3544 1804 -3502 1922
rect -3384 1804 -3342 1922
rect -3224 1804 -3182 1922
rect -3064 1804 -3022 1922
rect -2904 1804 -2862 1922
rect -2744 1804 -2702 1922
rect -2584 1804 -2542 1922
rect -2424 1804 -2382 1922
rect -2264 1819 -2003 1922
rect -2264 1804 -2194 1819
rect -5809 1730 -2194 1804
rect -5809 1701 -5733 1730
rect -6003 1659 -5733 1701
rect -6003 1541 -5927 1659
rect -5809 1541 -5733 1659
rect -6003 1499 -5733 1541
rect -6003 1381 -5927 1499
rect -5809 1381 -5733 1499
rect -6003 1339 -5733 1381
rect -6003 1221 -5927 1339
rect -5809 1221 -5733 1339
rect -6003 1179 -5733 1221
rect -6003 1061 -5927 1179
rect -5809 1061 -5733 1179
rect -6003 1019 -5733 1061
rect -6003 901 -5927 1019
rect -5809 901 -5733 1019
rect -6003 859 -5733 901
rect -6003 741 -5927 859
rect -5809 741 -5733 859
rect -6003 699 -5733 741
rect -6003 581 -5927 699
rect -5809 581 -5733 699
rect -6003 539 -5733 581
rect -6003 421 -5927 539
rect -5809 421 -5733 539
rect -6003 379 -5733 421
rect -6003 261 -5927 379
rect -5809 261 -5733 379
rect -6003 219 -5733 261
rect -6003 101 -5927 219
rect -5809 101 -5733 219
rect -6003 59 -5733 101
rect -6003 -59 -5927 59
rect -5809 -59 -5733 59
rect -6003 -101 -5733 -59
rect -6003 -219 -5927 -101
rect -5809 -219 -5733 -101
rect -6003 -261 -5733 -219
rect -6003 -379 -5927 -261
rect -5809 -379 -5733 -261
rect -6003 -421 -5733 -379
rect -6003 -539 -5927 -421
rect -5809 -539 -5733 -421
rect -6003 -581 -5733 -539
rect -6003 -699 -5927 -581
rect -5809 -699 -5733 -581
rect -6003 -741 -5733 -699
rect -6003 -859 -5927 -741
rect -5809 -859 -5733 -741
rect -6003 -901 -5733 -859
rect -6003 -1019 -5927 -901
rect -5809 -1019 -5733 -901
rect -6003 -1061 -5733 -1019
rect -6003 -1179 -5927 -1061
rect -5809 -1179 -5733 -1061
rect -6003 -1221 -5733 -1179
rect -6003 -1339 -5927 -1221
rect -5809 -1339 -5733 -1221
rect -6003 -1381 -5733 -1339
rect -6003 -1499 -5927 -1381
rect -5809 -1499 -5733 -1381
rect -6003 -1541 -5733 -1499
rect -6003 -1659 -5927 -1541
rect -5809 -1659 -5733 -1541
rect -6003 -1701 -5733 -1659
rect -6003 -1819 -5927 -1701
rect -5809 -1730 -5733 -1701
rect -2273 1701 -2194 1730
rect -2076 1701 -2003 1819
rect -2273 1659 -2003 1701
rect -2273 1541 -2194 1659
rect -2076 1541 -2003 1659
rect -2273 1499 -2003 1541
rect -2273 1381 -2194 1499
rect -2076 1381 -2003 1499
rect -2273 1339 -2003 1381
rect -2273 1221 -2194 1339
rect -2076 1221 -2003 1339
rect -2273 1179 -2003 1221
rect -2273 1061 -2194 1179
rect -2076 1061 -2003 1179
rect -2273 1019 -2003 1061
rect -2273 901 -2194 1019
rect -2076 901 -2003 1019
rect -2273 859 -2003 901
rect -2273 741 -2194 859
rect -2076 741 -2003 859
rect -2273 699 -2003 741
rect -2273 581 -2194 699
rect -2076 581 -2003 699
rect -2273 539 -2003 581
rect -2273 421 -2194 539
rect -2076 421 -2003 539
rect -2273 379 -2003 421
rect -2273 261 -2194 379
rect -2076 261 -2003 379
rect -2273 219 -2003 261
rect -2273 101 -2194 219
rect -2076 101 -2003 219
rect -2273 59 -2003 101
rect -2273 -59 -2194 59
rect -2076 -59 -2003 59
rect -2273 -101 -2003 -59
rect -2273 -219 -2194 -101
rect -2076 -219 -2003 -101
rect -2273 -261 -2003 -219
rect -2273 -379 -2194 -261
rect -2076 -379 -2003 -261
rect -2273 -421 -2003 -379
rect -2273 -539 -2194 -421
rect -2076 -539 -2003 -421
rect -2273 -581 -2003 -539
rect -2273 -699 -2194 -581
rect -2076 -699 -2003 -581
rect -2273 -741 -2003 -699
rect -2273 -859 -2194 -741
rect -2076 -859 -2003 -741
rect -2273 -901 -2003 -859
rect -2273 -1019 -2194 -901
rect -2076 -1019 -2003 -901
rect -2273 -1061 -2003 -1019
rect -2273 -1179 -2194 -1061
rect -2076 -1179 -2003 -1061
rect -2273 -1221 -2003 -1179
rect -2273 -1339 -2194 -1221
rect -2076 -1339 -2003 -1221
rect -2273 -1381 -2003 -1339
rect -2273 -1499 -2194 -1381
rect -2076 -1499 -2003 -1381
rect -2273 -1541 -2003 -1499
rect -2273 -1659 -2194 -1541
rect -2076 -1659 -2003 -1541
rect -2273 -1701 -2003 -1659
rect -2273 -1730 -2194 -1701
rect -5809 -1806 -2194 -1730
rect -5809 -1819 -5742 -1806
rect -6003 -1924 -5742 -1819
rect -5624 -1924 -5582 -1806
rect -5464 -1924 -5422 -1806
rect -5304 -1924 -5262 -1806
rect -5144 -1924 -5102 -1806
rect -4984 -1924 -4942 -1806
rect -4824 -1924 -4782 -1806
rect -4664 -1924 -4622 -1806
rect -4504 -1924 -4462 -1806
rect -4344 -1924 -4302 -1806
rect -4184 -1924 -4142 -1806
rect -4024 -1924 -3982 -1806
rect -3864 -1924 -3822 -1806
rect -3704 -1924 -3662 -1806
rect -3544 -1924 -3502 -1806
rect -3384 -1924 -3342 -1806
rect -3224 -1924 -3182 -1806
rect -3064 -1924 -3022 -1806
rect -2904 -1924 -2862 -1806
rect -2744 -1924 -2702 -1806
rect -2584 -1924 -2542 -1806
rect -2424 -1924 -2382 -1806
rect -2264 -1819 -2194 -1806
rect -2076 -1819 -2003 -1701
rect -2264 -1924 -2003 -1819
rect -6003 -2000 -2003 -1924
<< via4 >>
rect -5742 1879 -5624 1922
rect -5742 1847 -5699 1879
rect -5699 1847 -5667 1879
rect -5667 1847 -5624 1879
rect -5927 1776 -5809 1819
rect -5742 1804 -5624 1847
rect -5582 1879 -5464 1922
rect -5582 1847 -5539 1879
rect -5539 1847 -5507 1879
rect -5507 1847 -5464 1879
rect -5582 1804 -5464 1847
rect -5422 1879 -5304 1922
rect -5422 1847 -5379 1879
rect -5379 1847 -5347 1879
rect -5347 1847 -5304 1879
rect -5422 1804 -5304 1847
rect -5262 1879 -5144 1922
rect -5262 1847 -5219 1879
rect -5219 1847 -5187 1879
rect -5187 1847 -5144 1879
rect -5262 1804 -5144 1847
rect -5102 1879 -4984 1922
rect -5102 1847 -5059 1879
rect -5059 1847 -5027 1879
rect -5027 1847 -4984 1879
rect -5102 1804 -4984 1847
rect -4942 1879 -4824 1922
rect -4942 1847 -4899 1879
rect -4899 1847 -4867 1879
rect -4867 1847 -4824 1879
rect -4942 1804 -4824 1847
rect -4782 1879 -4664 1922
rect -4782 1847 -4739 1879
rect -4739 1847 -4707 1879
rect -4707 1847 -4664 1879
rect -4782 1804 -4664 1847
rect -4622 1879 -4504 1922
rect -4622 1847 -4579 1879
rect -4579 1847 -4547 1879
rect -4547 1847 -4504 1879
rect -4622 1804 -4504 1847
rect -4462 1879 -4344 1922
rect -4462 1847 -4419 1879
rect -4419 1847 -4387 1879
rect -4387 1847 -4344 1879
rect -4462 1804 -4344 1847
rect -4302 1879 -4184 1922
rect -4302 1847 -4259 1879
rect -4259 1847 -4227 1879
rect -4227 1847 -4184 1879
rect -4302 1804 -4184 1847
rect -4142 1879 -4024 1922
rect -4142 1847 -4099 1879
rect -4099 1847 -4067 1879
rect -4067 1847 -4024 1879
rect -4142 1804 -4024 1847
rect -3982 1879 -3864 1922
rect -3982 1847 -3939 1879
rect -3939 1847 -3907 1879
rect -3907 1847 -3864 1879
rect -3982 1804 -3864 1847
rect -3822 1879 -3704 1922
rect -3822 1847 -3779 1879
rect -3779 1847 -3747 1879
rect -3747 1847 -3704 1879
rect -3822 1804 -3704 1847
rect -3662 1879 -3544 1922
rect -3662 1847 -3619 1879
rect -3619 1847 -3587 1879
rect -3587 1847 -3544 1879
rect -3662 1804 -3544 1847
rect -3502 1879 -3384 1922
rect -3502 1847 -3459 1879
rect -3459 1847 -3427 1879
rect -3427 1847 -3384 1879
rect -3502 1804 -3384 1847
rect -3342 1879 -3224 1922
rect -3342 1847 -3299 1879
rect -3299 1847 -3267 1879
rect -3267 1847 -3224 1879
rect -3342 1804 -3224 1847
rect -3182 1879 -3064 1922
rect -3182 1847 -3139 1879
rect -3139 1847 -3107 1879
rect -3107 1847 -3064 1879
rect -3182 1804 -3064 1847
rect -3022 1879 -2904 1922
rect -3022 1847 -2979 1879
rect -2979 1847 -2947 1879
rect -2947 1847 -2904 1879
rect -3022 1804 -2904 1847
rect -2862 1879 -2744 1922
rect -2862 1847 -2819 1879
rect -2819 1847 -2787 1879
rect -2787 1847 -2744 1879
rect -2862 1804 -2744 1847
rect -2702 1879 -2584 1922
rect -2702 1847 -2659 1879
rect -2659 1847 -2627 1879
rect -2627 1847 -2584 1879
rect -2702 1804 -2584 1847
rect -2542 1879 -2424 1922
rect -2542 1847 -2499 1879
rect -2499 1847 -2467 1879
rect -2467 1847 -2424 1879
rect -2542 1804 -2424 1847
rect -2382 1879 -2264 1922
rect -2382 1847 -2339 1879
rect -2339 1847 -2307 1879
rect -2307 1847 -2264 1879
rect -2382 1804 -2264 1847
rect -5927 1744 -5884 1776
rect -5884 1744 -5852 1776
rect -5852 1744 -5809 1776
rect -5927 1701 -5809 1744
rect -2194 1776 -2076 1819
rect -2194 1744 -2151 1776
rect -2151 1744 -2119 1776
rect -2119 1744 -2076 1776
rect -5927 1616 -5809 1659
rect -5927 1584 -5884 1616
rect -5884 1584 -5852 1616
rect -5852 1584 -5809 1616
rect -5927 1541 -5809 1584
rect -5927 1456 -5809 1499
rect -5927 1424 -5884 1456
rect -5884 1424 -5852 1456
rect -5852 1424 -5809 1456
rect -5927 1381 -5809 1424
rect -5927 1296 -5809 1339
rect -5927 1264 -5884 1296
rect -5884 1264 -5852 1296
rect -5852 1264 -5809 1296
rect -5927 1221 -5809 1264
rect -5927 1136 -5809 1179
rect -5927 1104 -5884 1136
rect -5884 1104 -5852 1136
rect -5852 1104 -5809 1136
rect -5927 1061 -5809 1104
rect -5927 976 -5809 1019
rect -5927 944 -5884 976
rect -5884 944 -5852 976
rect -5852 944 -5809 976
rect -5927 901 -5809 944
rect -5927 816 -5809 859
rect -5927 784 -5884 816
rect -5884 784 -5852 816
rect -5852 784 -5809 816
rect -5927 741 -5809 784
rect -5927 656 -5809 699
rect -5927 624 -5884 656
rect -5884 624 -5852 656
rect -5852 624 -5809 656
rect -5927 581 -5809 624
rect -5927 496 -5809 539
rect -5927 464 -5884 496
rect -5884 464 -5852 496
rect -5852 464 -5809 496
rect -5927 421 -5809 464
rect -5927 336 -5809 379
rect -5927 304 -5884 336
rect -5884 304 -5852 336
rect -5852 304 -5809 336
rect -5927 261 -5809 304
rect -5927 176 -5809 219
rect -5927 144 -5884 176
rect -5884 144 -5852 176
rect -5852 144 -5809 176
rect -5927 101 -5809 144
rect -5927 16 -5809 59
rect -5927 -16 -5884 16
rect -5884 -16 -5852 16
rect -5852 -16 -5809 16
rect -5927 -59 -5809 -16
rect -5927 -144 -5809 -101
rect -5927 -176 -5884 -144
rect -5884 -176 -5852 -144
rect -5852 -176 -5809 -144
rect -5927 -219 -5809 -176
rect -5927 -304 -5809 -261
rect -5927 -336 -5884 -304
rect -5884 -336 -5852 -304
rect -5852 -336 -5809 -304
rect -5927 -379 -5809 -336
rect -5927 -464 -5809 -421
rect -5927 -496 -5884 -464
rect -5884 -496 -5852 -464
rect -5852 -496 -5809 -464
rect -5927 -539 -5809 -496
rect -5927 -624 -5809 -581
rect -5927 -656 -5884 -624
rect -5884 -656 -5852 -624
rect -5852 -656 -5809 -624
rect -5927 -699 -5809 -656
rect -5927 -784 -5809 -741
rect -5927 -816 -5884 -784
rect -5884 -816 -5852 -784
rect -5852 -816 -5809 -784
rect -5927 -859 -5809 -816
rect -5927 -944 -5809 -901
rect -5927 -976 -5884 -944
rect -5884 -976 -5852 -944
rect -5852 -976 -5809 -944
rect -5927 -1019 -5809 -976
rect -5927 -1104 -5809 -1061
rect -5927 -1136 -5884 -1104
rect -5884 -1136 -5852 -1104
rect -5852 -1136 -5809 -1104
rect -5927 -1179 -5809 -1136
rect -5927 -1264 -5809 -1221
rect -5927 -1296 -5884 -1264
rect -5884 -1296 -5852 -1264
rect -5852 -1296 -5809 -1264
rect -5927 -1339 -5809 -1296
rect -5927 -1424 -5809 -1381
rect -5927 -1456 -5884 -1424
rect -5884 -1456 -5852 -1424
rect -5852 -1456 -5809 -1424
rect -5927 -1499 -5809 -1456
rect -5927 -1584 -5809 -1541
rect -5927 -1616 -5884 -1584
rect -5884 -1616 -5852 -1584
rect -5852 -1616 -5809 -1584
rect -5927 -1659 -5809 -1616
rect -5927 -1744 -5809 -1701
rect -2194 1701 -2076 1744
rect -2194 1616 -2076 1659
rect -2194 1584 -2151 1616
rect -2151 1584 -2119 1616
rect -2119 1584 -2076 1616
rect -2194 1541 -2076 1584
rect -2194 1456 -2076 1499
rect -2194 1424 -2151 1456
rect -2151 1424 -2119 1456
rect -2119 1424 -2076 1456
rect -2194 1381 -2076 1424
rect -2194 1296 -2076 1339
rect -2194 1264 -2151 1296
rect -2151 1264 -2119 1296
rect -2119 1264 -2076 1296
rect -2194 1221 -2076 1264
rect -2194 1136 -2076 1179
rect -2194 1104 -2151 1136
rect -2151 1104 -2119 1136
rect -2119 1104 -2076 1136
rect -2194 1061 -2076 1104
rect -2194 976 -2076 1019
rect -2194 944 -2151 976
rect -2151 944 -2119 976
rect -2119 944 -2076 976
rect -2194 901 -2076 944
rect -2194 816 -2076 859
rect -2194 784 -2151 816
rect -2151 784 -2119 816
rect -2119 784 -2076 816
rect -2194 741 -2076 784
rect -2194 656 -2076 699
rect -2194 624 -2151 656
rect -2151 624 -2119 656
rect -2119 624 -2076 656
rect -2194 581 -2076 624
rect -2194 496 -2076 539
rect -2194 464 -2151 496
rect -2151 464 -2119 496
rect -2119 464 -2076 496
rect -2194 421 -2076 464
rect -2194 336 -2076 379
rect -2194 304 -2151 336
rect -2151 304 -2119 336
rect -2119 304 -2076 336
rect -2194 261 -2076 304
rect -2194 176 -2076 219
rect -2194 144 -2151 176
rect -2151 144 -2119 176
rect -2119 144 -2076 176
rect -2194 101 -2076 144
rect -2194 16 -2076 59
rect -2194 -16 -2151 16
rect -2151 -16 -2119 16
rect -2119 -16 -2076 16
rect -2194 -59 -2076 -16
rect -2194 -144 -2076 -101
rect -2194 -176 -2151 -144
rect -2151 -176 -2119 -144
rect -2119 -176 -2076 -144
rect -2194 -219 -2076 -176
rect -2194 -304 -2076 -261
rect -2194 -336 -2151 -304
rect -2151 -336 -2119 -304
rect -2119 -336 -2076 -304
rect -2194 -379 -2076 -336
rect -2194 -464 -2076 -421
rect -2194 -496 -2151 -464
rect -2151 -496 -2119 -464
rect -2119 -496 -2076 -464
rect -2194 -539 -2076 -496
rect -2194 -624 -2076 -581
rect -2194 -656 -2151 -624
rect -2151 -656 -2119 -624
rect -2119 -656 -2076 -624
rect -2194 -699 -2076 -656
rect -2194 -784 -2076 -741
rect -2194 -816 -2151 -784
rect -2151 -816 -2119 -784
rect -2119 -816 -2076 -784
rect -2194 -859 -2076 -816
rect -2194 -944 -2076 -901
rect -2194 -976 -2151 -944
rect -2151 -976 -2119 -944
rect -2119 -976 -2076 -944
rect -2194 -1019 -2076 -976
rect -2194 -1104 -2076 -1061
rect -2194 -1136 -2151 -1104
rect -2151 -1136 -2119 -1104
rect -2119 -1136 -2076 -1104
rect -2194 -1179 -2076 -1136
rect -2194 -1264 -2076 -1221
rect -2194 -1296 -2151 -1264
rect -2151 -1296 -2119 -1264
rect -2119 -1296 -2076 -1264
rect -2194 -1339 -2076 -1296
rect -2194 -1424 -2076 -1381
rect -2194 -1456 -2151 -1424
rect -2151 -1456 -2119 -1424
rect -2119 -1456 -2076 -1424
rect -2194 -1499 -2076 -1456
rect -2194 -1584 -2076 -1541
rect -2194 -1616 -2151 -1584
rect -2151 -1616 -2119 -1584
rect -2119 -1616 -2076 -1584
rect -2194 -1659 -2076 -1616
rect -5927 -1776 -5884 -1744
rect -5884 -1776 -5852 -1744
rect -5852 -1776 -5809 -1744
rect -5927 -1819 -5809 -1776
rect -2194 -1744 -2076 -1701
rect -2194 -1776 -2151 -1744
rect -2151 -1776 -2119 -1744
rect -2119 -1776 -2076 -1744
rect -5742 -1849 -5624 -1806
rect -5742 -1881 -5699 -1849
rect -5699 -1881 -5667 -1849
rect -5667 -1881 -5624 -1849
rect -5742 -1924 -5624 -1881
rect -5582 -1849 -5464 -1806
rect -5582 -1881 -5539 -1849
rect -5539 -1881 -5507 -1849
rect -5507 -1881 -5464 -1849
rect -5582 -1924 -5464 -1881
rect -5422 -1849 -5304 -1806
rect -5422 -1881 -5379 -1849
rect -5379 -1881 -5347 -1849
rect -5347 -1881 -5304 -1849
rect -5422 -1924 -5304 -1881
rect -5262 -1849 -5144 -1806
rect -5262 -1881 -5219 -1849
rect -5219 -1881 -5187 -1849
rect -5187 -1881 -5144 -1849
rect -5262 -1924 -5144 -1881
rect -5102 -1849 -4984 -1806
rect -5102 -1881 -5059 -1849
rect -5059 -1881 -5027 -1849
rect -5027 -1881 -4984 -1849
rect -5102 -1924 -4984 -1881
rect -4942 -1849 -4824 -1806
rect -4942 -1881 -4899 -1849
rect -4899 -1881 -4867 -1849
rect -4867 -1881 -4824 -1849
rect -4942 -1924 -4824 -1881
rect -4782 -1849 -4664 -1806
rect -4782 -1881 -4739 -1849
rect -4739 -1881 -4707 -1849
rect -4707 -1881 -4664 -1849
rect -4782 -1924 -4664 -1881
rect -4622 -1849 -4504 -1806
rect -4622 -1881 -4579 -1849
rect -4579 -1881 -4547 -1849
rect -4547 -1881 -4504 -1849
rect -4622 -1924 -4504 -1881
rect -4462 -1849 -4344 -1806
rect -4462 -1881 -4419 -1849
rect -4419 -1881 -4387 -1849
rect -4387 -1881 -4344 -1849
rect -4462 -1924 -4344 -1881
rect -4302 -1849 -4184 -1806
rect -4302 -1881 -4259 -1849
rect -4259 -1881 -4227 -1849
rect -4227 -1881 -4184 -1849
rect -4302 -1924 -4184 -1881
rect -4142 -1849 -4024 -1806
rect -4142 -1881 -4099 -1849
rect -4099 -1881 -4067 -1849
rect -4067 -1881 -4024 -1849
rect -4142 -1924 -4024 -1881
rect -3982 -1849 -3864 -1806
rect -3982 -1881 -3939 -1849
rect -3939 -1881 -3907 -1849
rect -3907 -1881 -3864 -1849
rect -3982 -1924 -3864 -1881
rect -3822 -1849 -3704 -1806
rect -3822 -1881 -3779 -1849
rect -3779 -1881 -3747 -1849
rect -3747 -1881 -3704 -1849
rect -3822 -1924 -3704 -1881
rect -3662 -1849 -3544 -1806
rect -3662 -1881 -3619 -1849
rect -3619 -1881 -3587 -1849
rect -3587 -1881 -3544 -1849
rect -3662 -1924 -3544 -1881
rect -3502 -1849 -3384 -1806
rect -3502 -1881 -3459 -1849
rect -3459 -1881 -3427 -1849
rect -3427 -1881 -3384 -1849
rect -3502 -1924 -3384 -1881
rect -3342 -1849 -3224 -1806
rect -3342 -1881 -3299 -1849
rect -3299 -1881 -3267 -1849
rect -3267 -1881 -3224 -1849
rect -3342 -1924 -3224 -1881
rect -3182 -1849 -3064 -1806
rect -3182 -1881 -3139 -1849
rect -3139 -1881 -3107 -1849
rect -3107 -1881 -3064 -1849
rect -3182 -1924 -3064 -1881
rect -3022 -1849 -2904 -1806
rect -3022 -1881 -2979 -1849
rect -2979 -1881 -2947 -1849
rect -2947 -1881 -2904 -1849
rect -3022 -1924 -2904 -1881
rect -2862 -1849 -2744 -1806
rect -2862 -1881 -2819 -1849
rect -2819 -1881 -2787 -1849
rect -2787 -1881 -2744 -1849
rect -2862 -1924 -2744 -1881
rect -2702 -1849 -2584 -1806
rect -2702 -1881 -2659 -1849
rect -2659 -1881 -2627 -1849
rect -2627 -1881 -2584 -1849
rect -2702 -1924 -2584 -1881
rect -2542 -1849 -2424 -1806
rect -2542 -1881 -2499 -1849
rect -2499 -1881 -2467 -1849
rect -2467 -1881 -2424 -1849
rect -2542 -1924 -2424 -1881
rect -2382 -1849 -2264 -1806
rect -2194 -1819 -2076 -1776
rect -2382 -1881 -2339 -1849
rect -2339 -1881 -2307 -1849
rect -2307 -1881 -2264 -1849
rect -2382 -1924 -2264 -1881
<< metal5 >>
rect -6003 1922 -2003 2000
rect -6003 1819 -5742 1922
rect -6003 1701 -5927 1819
rect -5809 1804 -5742 1819
rect -5624 1804 -5582 1922
rect -5464 1804 -5422 1922
rect -5304 1804 -5262 1922
rect -5144 1804 -5102 1922
rect -4984 1804 -4942 1922
rect -4824 1804 -4782 1922
rect -4664 1804 -4622 1922
rect -4504 1804 -4462 1922
rect -4344 1804 -4302 1922
rect -4184 1804 -4142 1922
rect -4024 1804 -3982 1922
rect -3864 1804 -3822 1922
rect -3704 1804 -3662 1922
rect -3544 1804 -3502 1922
rect -3384 1804 -3342 1922
rect -3224 1804 -3182 1922
rect -3064 1804 -3022 1922
rect -2904 1804 -2862 1922
rect -2744 1804 -2702 1922
rect -2584 1804 -2542 1922
rect -2424 1804 -2382 1922
rect -2264 1819 -2003 1922
rect -2264 1804 -2194 1819
rect -5809 1701 -2194 1804
rect -2076 1701 -2003 1819
rect -6003 1659 -2003 1701
rect -6003 1541 -5927 1659
rect -5809 1541 -2194 1659
rect -2076 1541 -2003 1659
rect -6003 1499 -2003 1541
rect -6003 1381 -5927 1499
rect -5809 1381 -2194 1499
rect -2076 1381 -2003 1499
rect -6003 1339 -2003 1381
rect -6003 1221 -5927 1339
rect -5809 1221 -2194 1339
rect -2076 1221 -2003 1339
rect -6003 1179 -2003 1221
rect -6003 1061 -5927 1179
rect -5809 1061 -2194 1179
rect -2076 1061 -2003 1179
rect -6003 1019 -2003 1061
rect -6003 901 -5927 1019
rect -5809 901 -2194 1019
rect -2076 901 -2003 1019
rect -6003 859 -2003 901
rect -6003 741 -5927 859
rect -5809 741 -2194 859
rect -2076 741 -2003 859
rect -6003 699 -2003 741
rect -6003 581 -5927 699
rect -5809 581 -2194 699
rect -2076 581 -2003 699
rect -6003 539 -2003 581
rect -6003 421 -5927 539
rect -5809 421 -2194 539
rect -2076 421 -2003 539
rect -6003 379 -2003 421
rect -6003 261 -5927 379
rect -5809 261 -2194 379
rect -2076 261 -2003 379
rect -6003 219 -2003 261
rect -6003 101 -5927 219
rect -5809 101 -2194 219
rect -2076 101 -2003 219
rect -6003 59 -2003 101
rect -6003 -59 -5927 59
rect -5809 -59 -2194 59
rect -2076 -59 -2003 59
rect -6003 -101 -2003 -59
rect -6003 -219 -5927 -101
rect -5809 -219 -2194 -101
rect -2076 -219 -2003 -101
rect -6003 -261 -2003 -219
rect -6003 -379 -5927 -261
rect -5809 -379 -2194 -261
rect -2076 -379 -2003 -261
rect -6003 -421 -2003 -379
rect -6003 -539 -5927 -421
rect -5809 -539 -2194 -421
rect -2076 -539 -2003 -421
rect -6003 -581 -2003 -539
rect -6003 -699 -5927 -581
rect -5809 -699 -2194 -581
rect -2076 -699 -2003 -581
rect -6003 -741 -2003 -699
rect -6003 -859 -5927 -741
rect -5809 -859 -2194 -741
rect -2076 -859 -2003 -741
rect -6003 -901 -2003 -859
rect -6003 -1019 -5927 -901
rect -5809 -1019 -2194 -901
rect -2076 -1019 -2003 -901
rect -6003 -1061 -2003 -1019
rect -6003 -1179 -5927 -1061
rect -5809 -1179 -2194 -1061
rect -2076 -1179 -2003 -1061
rect -6003 -1221 -2003 -1179
rect -6003 -1339 -5927 -1221
rect -5809 -1339 -2194 -1221
rect -2076 -1339 -2003 -1221
rect -6003 -1381 -2003 -1339
rect -6003 -1499 -5927 -1381
rect -5809 -1499 -2194 -1381
rect -2076 -1499 -2003 -1381
rect -6003 -1541 -2003 -1499
rect -6003 -1659 -5927 -1541
rect -5809 -1659 -2194 -1541
rect -2076 -1659 -2003 -1541
rect -6003 -1701 -2003 -1659
rect -6003 -1819 -5927 -1701
rect -5809 -1806 -2194 -1701
rect -5809 -1819 -5742 -1806
rect -6003 -1924 -5742 -1819
rect -5624 -1924 -5582 -1806
rect -5464 -1924 -5422 -1806
rect -5304 -1924 -5262 -1806
rect -5144 -1924 -5102 -1806
rect -4984 -1924 -4942 -1806
rect -4824 -1924 -4782 -1806
rect -4664 -1924 -4622 -1806
rect -4504 -1924 -4462 -1806
rect -4344 -1924 -4302 -1806
rect -4184 -1924 -4142 -1806
rect -4024 -1924 -3982 -1806
rect -3864 -1924 -3822 -1806
rect -3704 -1924 -3662 -1806
rect -3544 -1924 -3502 -1806
rect -3384 -1924 -3342 -1806
rect -3224 -1924 -3182 -1806
rect -3064 -1924 -3022 -1806
rect -2904 -1924 -2862 -1806
rect -2744 -1924 -2702 -1806
rect -2584 -1924 -2542 -1806
rect -2424 -1924 -2382 -1806
rect -2264 -1819 -2194 -1806
rect -2076 -1819 -2003 -1701
rect -2264 -1924 -2003 -1819
rect -6003 -2000 -2003 -1924
<< glass >>
rect -5888 -1880 -2118 1880
<< labels >>
<< end >>
