magic
tech sky130B
timestamp 1668125262
<< metal4 >>
rect 1580 4420 2420 4520
rect 1580 -160 1640 4420
rect 1670 -160 1770 4390
rect 1800 -160 1920 4420
rect 1950 -160 2050 4390
rect 2080 -160 2200 4420
rect 2230 -160 2330 4390
rect 2360 -160 2420 4420
<< fillblock >>
rect 1860 -160 2140 4520
<< labels >>
rlabel metal4 1950 -160 2050 -100 1 TOP
rlabel metal4 1920 4420 2080 4520 1 BOT
rlabel metal4 1640 4420 1800 4520 1 BOT
rlabel metal4 2230 -160 2330 -100 1 TOPR
rlabel metal4 1670 -160 1770 -100 1 TOPL
<< end >>
