magic
tech sky130A
magscale 1 2
timestamp 1671334348
<< pwell >>
rect -201 -648 201 648
<< psubdiff >>
rect -165 578 -69 612
rect 69 578 165 612
rect -165 516 -131 578
rect 131 516 165 578
rect -165 -578 -131 -516
rect 131 -578 165 -516
rect -165 -612 -69 -578
rect 69 -612 165 -578
<< psubdiffcont >>
rect -69 578 69 612
rect -165 -516 -131 516
rect 131 -516 165 516
rect -69 -612 69 -578
<< xpolycontact >>
rect -35 50 35 482
rect -35 -482 35 -50
<< xpolyres >>
rect -35 -50 35 50
<< locali >>
rect -165 578 -69 612
rect 69 578 165 612
rect -165 516 -131 578
rect 131 516 165 578
rect -165 -578 -131 -516
rect 131 -578 165 -516
rect -165 -612 -69 -578
rect 69 -612 165 -578
<< viali >>
rect -19 67 19 464
rect -19 -464 19 -67
<< metal1 >>
rect -25 464 25 476
rect -25 67 -19 464
rect 19 67 25 464
rect -25 55 25 67
rect -25 -67 25 -55
rect -25 -464 -19 -67
rect 19 -464 25 -67
rect -25 -476 25 -464
<< res0p35 >>
rect -37 -52 37 52
<< properties >>
string FIXED_BBOX -148 -595 148 595
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.35 l 0.5 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 3.932k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 1 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
