magic
tech sky130A
magscale 1 2
timestamp 1671169241
<< nwell >>
rect -1438 4672 4088 7110
<< pmos >>
rect -1242 4891 -1182 6891
rect -1124 4891 -1064 6891
rect -1006 4891 -946 6891
rect -888 4891 -828 6891
rect -770 4891 -710 6891
rect -652 4891 -592 6891
rect -534 4891 -474 6891
rect -416 4891 -356 6891
rect -298 4891 -238 6891
rect -180 4891 -120 6891
rect -62 4891 -2 6891
rect 56 4891 116 6891
rect 174 4891 234 6891
rect 292 4891 352 6891
rect 410 4891 470 6891
rect 528 4891 588 6891
rect 646 4891 706 6891
rect 764 4891 824 6891
rect 882 4891 942 6891
rect 1000 4891 1060 6891
rect 1118 4891 1178 6891
rect 1236 4891 1296 6891
rect 1354 4891 1414 6891
rect 1472 4891 1532 6891
rect 1590 4891 1650 6891
rect 1708 4891 1768 6891
rect 1826 4891 1886 6891
rect 1944 4891 2004 6891
rect 2062 4891 2122 6891
rect 2180 4891 2240 6891
rect 2298 4891 2358 6891
rect 2416 4891 2476 6891
rect 2534 4891 2594 6891
rect 2652 4891 2712 6891
rect 2770 4891 2830 6891
rect 2888 4891 2948 6891
rect 3006 4891 3066 6891
rect 3124 4891 3184 6891
rect 3242 4891 3302 6891
rect 3360 4891 3420 6891
rect 3478 4891 3538 6891
rect 3596 4891 3656 6891
rect 3714 4891 3774 6891
rect 3832 4891 3892 6891
<< pdiff >>
rect -1300 6879 -1242 6891
rect -1300 4903 -1288 6879
rect -1254 4903 -1242 6879
rect -1300 4891 -1242 4903
rect -1182 6879 -1124 6891
rect -1182 4903 -1170 6879
rect -1136 4903 -1124 6879
rect -1182 4891 -1124 4903
rect -1064 6879 -1006 6891
rect -1064 4903 -1052 6879
rect -1018 4903 -1006 6879
rect -1064 4891 -1006 4903
rect -946 6879 -888 6891
rect -946 4903 -934 6879
rect -900 4903 -888 6879
rect -946 4891 -888 4903
rect -828 6879 -770 6891
rect -828 4903 -816 6879
rect -782 4903 -770 6879
rect -828 4891 -770 4903
rect -710 6879 -652 6891
rect -710 4903 -698 6879
rect -664 4903 -652 6879
rect -710 4891 -652 4903
rect -592 6879 -534 6891
rect -592 4903 -580 6879
rect -546 4903 -534 6879
rect -592 4891 -534 4903
rect -474 6879 -416 6891
rect -474 4903 -462 6879
rect -428 4903 -416 6879
rect -474 4891 -416 4903
rect -356 6879 -298 6891
rect -356 4903 -344 6879
rect -310 4903 -298 6879
rect -356 4891 -298 4903
rect -238 6879 -180 6891
rect -238 4903 -226 6879
rect -192 4903 -180 6879
rect -238 4891 -180 4903
rect -120 6879 -62 6891
rect -120 4903 -108 6879
rect -74 4903 -62 6879
rect -120 4891 -62 4903
rect -2 6879 56 6891
rect -2 4903 10 6879
rect 44 4903 56 6879
rect -2 4891 56 4903
rect 116 6879 174 6891
rect 116 4903 128 6879
rect 162 4903 174 6879
rect 116 4891 174 4903
rect 234 6879 292 6891
rect 234 4903 246 6879
rect 280 4903 292 6879
rect 234 4891 292 4903
rect 352 6879 410 6891
rect 352 4903 364 6879
rect 398 4903 410 6879
rect 352 4891 410 4903
rect 470 6879 528 6891
rect 470 4903 482 6879
rect 516 4903 528 6879
rect 470 4891 528 4903
rect 588 6879 646 6891
rect 588 4903 600 6879
rect 634 4903 646 6879
rect 588 4891 646 4903
rect 706 6879 764 6891
rect 706 4903 718 6879
rect 752 4903 764 6879
rect 706 4891 764 4903
rect 824 6879 882 6891
rect 824 4903 836 6879
rect 870 4903 882 6879
rect 824 4891 882 4903
rect 942 6879 1000 6891
rect 942 4903 954 6879
rect 988 4903 1000 6879
rect 942 4891 1000 4903
rect 1060 6879 1118 6891
rect 1060 4903 1072 6879
rect 1106 4903 1118 6879
rect 1060 4891 1118 4903
rect 1178 6879 1236 6891
rect 1178 4903 1190 6879
rect 1224 4903 1236 6879
rect 1178 4891 1236 4903
rect 1296 6879 1354 6891
rect 1296 4903 1308 6879
rect 1342 4903 1354 6879
rect 1296 4891 1354 4903
rect 1414 6879 1472 6891
rect 1414 4903 1426 6879
rect 1460 4903 1472 6879
rect 1414 4891 1472 4903
rect 1532 6879 1590 6891
rect 1532 4903 1544 6879
rect 1578 4903 1590 6879
rect 1532 4891 1590 4903
rect 1650 6879 1708 6891
rect 1650 4903 1662 6879
rect 1696 4903 1708 6879
rect 1650 4891 1708 4903
rect 1768 6879 1826 6891
rect 1768 4903 1780 6879
rect 1814 4903 1826 6879
rect 1768 4891 1826 4903
rect 1886 6879 1944 6891
rect 1886 4903 1898 6879
rect 1932 4903 1944 6879
rect 1886 4891 1944 4903
rect 2004 6879 2062 6891
rect 2004 4903 2016 6879
rect 2050 4903 2062 6879
rect 2004 4891 2062 4903
rect 2122 6879 2180 6891
rect 2122 4903 2134 6879
rect 2168 4903 2180 6879
rect 2122 4891 2180 4903
rect 2240 6879 2298 6891
rect 2240 4903 2252 6879
rect 2286 4903 2298 6879
rect 2240 4891 2298 4903
rect 2358 6879 2416 6891
rect 2358 4903 2370 6879
rect 2404 4903 2416 6879
rect 2358 4891 2416 4903
rect 2476 6879 2534 6891
rect 2476 4903 2488 6879
rect 2522 4903 2534 6879
rect 2476 4891 2534 4903
rect 2594 6879 2652 6891
rect 2594 4903 2606 6879
rect 2640 4903 2652 6879
rect 2594 4891 2652 4903
rect 2712 6879 2770 6891
rect 2712 4903 2724 6879
rect 2758 4903 2770 6879
rect 2712 4891 2770 4903
rect 2830 6879 2888 6891
rect 2830 4903 2842 6879
rect 2876 4903 2888 6879
rect 2830 4891 2888 4903
rect 2948 6879 3006 6891
rect 2948 4903 2960 6879
rect 2994 4903 3006 6879
rect 2948 4891 3006 4903
rect 3066 6879 3124 6891
rect 3066 4903 3078 6879
rect 3112 4903 3124 6879
rect 3066 4891 3124 4903
rect 3184 6879 3242 6891
rect 3184 4903 3196 6879
rect 3230 4903 3242 6879
rect 3184 4891 3242 4903
rect 3302 6879 3360 6891
rect 3302 4903 3314 6879
rect 3348 4903 3360 6879
rect 3302 4891 3360 4903
rect 3420 6879 3478 6891
rect 3420 4903 3432 6879
rect 3466 4903 3478 6879
rect 3420 4891 3478 4903
rect 3538 6879 3596 6891
rect 3538 4903 3550 6879
rect 3584 4903 3596 6879
rect 3538 4891 3596 4903
rect 3656 6879 3714 6891
rect 3656 4903 3668 6879
rect 3702 4903 3714 6879
rect 3656 4891 3714 4903
rect 3774 6879 3832 6891
rect 3774 4903 3786 6879
rect 3820 4903 3832 6879
rect 3774 4891 3832 4903
rect 3892 6879 3950 6891
rect 3892 4903 3904 6879
rect 3938 4903 3950 6879
rect 3892 4891 3950 4903
<< pdiffc >>
rect -1288 4903 -1254 6879
rect -1170 4903 -1136 6879
rect -1052 4903 -1018 6879
rect -934 4903 -900 6879
rect -816 4903 -782 6879
rect -698 4903 -664 6879
rect -580 4903 -546 6879
rect -462 4903 -428 6879
rect -344 4903 -310 6879
rect -226 4903 -192 6879
rect -108 4903 -74 6879
rect 10 4903 44 6879
rect 128 4903 162 6879
rect 246 4903 280 6879
rect 364 4903 398 6879
rect 482 4903 516 6879
rect 600 4903 634 6879
rect 718 4903 752 6879
rect 836 4903 870 6879
rect 954 4903 988 6879
rect 1072 4903 1106 6879
rect 1190 4903 1224 6879
rect 1308 4903 1342 6879
rect 1426 4903 1460 6879
rect 1544 4903 1578 6879
rect 1662 4903 1696 6879
rect 1780 4903 1814 6879
rect 1898 4903 1932 6879
rect 2016 4903 2050 6879
rect 2134 4903 2168 6879
rect 2252 4903 2286 6879
rect 2370 4903 2404 6879
rect 2488 4903 2522 6879
rect 2606 4903 2640 6879
rect 2724 4903 2758 6879
rect 2842 4903 2876 6879
rect 2960 4903 2994 6879
rect 3078 4903 3112 6879
rect 3196 4903 3230 6879
rect 3314 4903 3348 6879
rect 3432 4903 3466 6879
rect 3550 4903 3584 6879
rect 3668 4903 3702 6879
rect 3786 4903 3820 6879
rect 3904 4903 3938 6879
<< nsubdiff >>
rect -1402 7040 -1306 7074
rect 3956 7040 4052 7074
rect -1402 6978 -1368 7040
rect 4018 6978 4052 7040
rect -1402 4742 -1368 4804
rect 4018 4742 4052 4804
rect -1402 4708 -1306 4742
rect 3956 4708 4052 4742
<< nsubdiffcont >>
rect -1306 7040 3956 7074
rect -1402 4804 -1368 6978
rect 4018 4804 4052 6978
rect -1306 4708 3956 4742
<< poly >>
rect -1245 6972 -1179 6988
rect -1245 6938 -1229 6972
rect -1195 6938 -1179 6972
rect -1245 6922 -1179 6938
rect -1127 6972 -1061 6988
rect -1127 6938 -1111 6972
rect -1077 6938 -1061 6972
rect -1127 6922 -1061 6938
rect -1009 6972 -943 6988
rect -1009 6938 -993 6972
rect -959 6938 -943 6972
rect -1009 6922 -943 6938
rect -891 6972 -825 6988
rect -891 6938 -875 6972
rect -841 6938 -825 6972
rect -891 6922 -825 6938
rect -773 6972 -707 6988
rect -773 6938 -757 6972
rect -723 6938 -707 6972
rect -773 6922 -707 6938
rect -655 6972 -589 6988
rect -655 6938 -639 6972
rect -605 6938 -589 6972
rect -655 6922 -589 6938
rect -537 6972 -471 6988
rect -537 6938 -521 6972
rect -487 6938 -471 6972
rect -537 6922 -471 6938
rect -419 6972 -353 6988
rect -419 6938 -403 6972
rect -369 6938 -353 6972
rect -419 6922 -353 6938
rect -301 6972 -235 6988
rect -301 6938 -285 6972
rect -251 6938 -235 6972
rect -301 6922 -235 6938
rect -183 6972 -117 6988
rect -183 6938 -167 6972
rect -133 6938 -117 6972
rect -183 6922 -117 6938
rect -65 6972 1 6988
rect -65 6938 -49 6972
rect -15 6938 1 6972
rect -65 6922 1 6938
rect 53 6972 119 6988
rect 53 6938 69 6972
rect 103 6938 119 6972
rect 53 6922 119 6938
rect 171 6972 237 6988
rect 171 6938 187 6972
rect 221 6938 237 6972
rect 171 6922 237 6938
rect 289 6972 355 6988
rect 289 6938 305 6972
rect 339 6938 355 6972
rect 289 6922 355 6938
rect 407 6972 473 6988
rect 407 6938 423 6972
rect 457 6938 473 6972
rect 407 6922 473 6938
rect 525 6972 591 6988
rect 525 6938 541 6972
rect 575 6938 591 6972
rect 525 6922 591 6938
rect 643 6972 709 6988
rect 643 6938 659 6972
rect 693 6938 709 6972
rect 643 6922 709 6938
rect 761 6972 827 6988
rect 761 6938 777 6972
rect 811 6938 827 6972
rect 761 6922 827 6938
rect 879 6972 945 6988
rect 879 6938 895 6972
rect 929 6938 945 6972
rect 879 6922 945 6938
rect 997 6972 1063 6988
rect 997 6938 1013 6972
rect 1047 6938 1063 6972
rect 997 6922 1063 6938
rect 1115 6922 1181 6988
rect 1233 6922 1299 6988
rect 1351 6922 1417 6988
rect 1469 6922 1535 6988
rect 1587 6972 1653 6988
rect 1587 6938 1603 6972
rect 1637 6938 1653 6972
rect 1587 6922 1653 6938
rect 1705 6972 1771 6988
rect 1705 6938 1721 6972
rect 1755 6938 1771 6972
rect 1705 6922 1771 6938
rect 1823 6972 1889 6988
rect 1823 6938 1839 6972
rect 1873 6938 1889 6972
rect 1823 6922 1889 6938
rect 1941 6972 2007 6988
rect 1941 6938 1957 6972
rect 1991 6938 2007 6972
rect 1941 6922 2007 6938
rect 2059 6972 2125 6988
rect 2059 6938 2075 6972
rect 2109 6938 2125 6972
rect 2059 6922 2125 6938
rect 2177 6972 2243 6988
rect 2177 6938 2193 6972
rect 2227 6938 2243 6972
rect 2177 6922 2243 6938
rect 2295 6972 2361 6988
rect 2295 6938 2311 6972
rect 2345 6938 2361 6972
rect 2295 6922 2361 6938
rect 2413 6972 2479 6988
rect 2413 6938 2429 6972
rect 2463 6938 2479 6972
rect 2413 6922 2479 6938
rect 2531 6972 2597 6988
rect 2531 6938 2547 6972
rect 2581 6938 2597 6972
rect 2531 6922 2597 6938
rect 2649 6972 2715 6988
rect 2649 6938 2665 6972
rect 2699 6938 2715 6972
rect 2649 6922 2715 6938
rect 2767 6972 2833 6988
rect 2767 6938 2783 6972
rect 2817 6938 2833 6972
rect 2767 6922 2833 6938
rect 2885 6972 2951 6988
rect 2885 6938 2901 6972
rect 2935 6938 2951 6972
rect 2885 6922 2951 6938
rect 3003 6972 3069 6988
rect 3003 6938 3019 6972
rect 3053 6938 3069 6972
rect 3003 6922 3069 6938
rect 3121 6972 3187 6988
rect 3121 6938 3137 6972
rect 3171 6938 3187 6972
rect 3121 6922 3187 6938
rect 3239 6972 3305 6988
rect 3239 6938 3255 6972
rect 3289 6938 3305 6972
rect 3239 6922 3305 6938
rect 3357 6972 3423 6988
rect 3357 6938 3373 6972
rect 3407 6938 3423 6972
rect 3357 6922 3423 6938
rect 3475 6972 3541 6988
rect 3475 6938 3491 6972
rect 3525 6938 3541 6972
rect 3475 6922 3541 6938
rect 3593 6972 3659 6988
rect 3593 6938 3609 6972
rect 3643 6938 3659 6972
rect 3593 6922 3659 6938
rect 3711 6972 3777 6988
rect 3711 6938 3727 6972
rect 3761 6938 3777 6972
rect 3711 6922 3777 6938
rect 3829 6972 3895 6988
rect 3829 6938 3845 6972
rect 3879 6938 3895 6972
rect 3829 6922 3895 6938
rect -1242 6891 -1182 6922
rect -1124 6891 -1064 6922
rect -1006 6891 -946 6922
rect -888 6891 -828 6922
rect -770 6891 -710 6922
rect -652 6891 -592 6922
rect -534 6891 -474 6922
rect -416 6891 -356 6922
rect -298 6891 -238 6922
rect -180 6891 -120 6922
rect -62 6891 -2 6922
rect 56 6891 116 6922
rect 174 6891 234 6922
rect 292 6891 352 6922
rect 410 6891 470 6922
rect 528 6891 588 6922
rect 646 6891 706 6922
rect 764 6891 824 6922
rect 882 6891 942 6922
rect 1000 6891 1060 6922
rect 1118 6891 1178 6922
rect 1236 6891 1296 6922
rect 1354 6891 1414 6922
rect 1472 6891 1532 6922
rect 1590 6891 1650 6922
rect 1708 6891 1768 6922
rect 1826 6891 1886 6922
rect 1944 6891 2004 6922
rect 2062 6891 2122 6922
rect 2180 6891 2240 6922
rect 2298 6891 2358 6922
rect 2416 6891 2476 6922
rect 2534 6891 2594 6922
rect 2652 6891 2712 6922
rect 2770 6891 2830 6922
rect 2888 6891 2948 6922
rect 3006 6891 3066 6922
rect 3124 6891 3184 6922
rect 3242 6891 3302 6922
rect 3360 6891 3420 6922
rect 3478 6891 3538 6922
rect 3596 6891 3656 6922
rect 3714 6891 3774 6922
rect 3832 6891 3892 6922
rect -1242 4860 -1182 4891
rect -1124 4860 -1064 4891
rect -1006 4860 -946 4891
rect -888 4860 -828 4891
rect -770 4860 -710 4891
rect -652 4860 -592 4891
rect -534 4860 -474 4891
rect -416 4860 -356 4891
rect -298 4860 -238 4891
rect -180 4860 -120 4891
rect -62 4860 -2 4891
rect 56 4860 116 4891
rect 174 4860 234 4891
rect 292 4860 352 4891
rect 410 4860 470 4891
rect 528 4860 588 4891
rect 646 4860 706 4891
rect 764 4860 824 4891
rect 882 4860 942 4891
rect 1000 4860 1060 4891
rect 1118 4860 1178 4891
rect 1236 4860 1296 4891
rect 1354 4860 1414 4891
rect 1472 4860 1532 4891
rect 1590 4860 1650 4891
rect 1708 4860 1768 4891
rect 1826 4860 1886 4891
rect 1944 4860 2004 4891
rect 2062 4860 2122 4891
rect 2180 4860 2240 4891
rect 2298 4860 2358 4891
rect 2416 4860 2476 4891
rect 2534 4860 2594 4891
rect 2652 4860 2712 4891
rect 2770 4860 2830 4891
rect 2888 4860 2948 4891
rect 3006 4860 3066 4891
rect 3124 4860 3184 4891
rect 3242 4860 3302 4891
rect 3360 4860 3420 4891
rect 3478 4860 3538 4891
rect 3596 4860 3656 4891
rect 3714 4860 3774 4891
rect 3832 4860 3892 4891
rect -1245 4844 -1179 4860
rect -1245 4810 -1229 4844
rect -1195 4810 -1179 4844
rect -1245 4794 -1179 4810
rect -1127 4844 -1061 4860
rect -1127 4810 -1111 4844
rect -1077 4810 -1061 4844
rect -1127 4794 -1061 4810
rect -1009 4844 -943 4860
rect -1009 4810 -993 4844
rect -959 4810 -943 4844
rect -1009 4794 -943 4810
rect -891 4844 -825 4860
rect -891 4810 -875 4844
rect -841 4810 -825 4844
rect -891 4794 -825 4810
rect -773 4844 -707 4860
rect -773 4810 -757 4844
rect -723 4810 -707 4844
rect -773 4794 -707 4810
rect -655 4844 -589 4860
rect -655 4810 -639 4844
rect -605 4810 -589 4844
rect -655 4794 -589 4810
rect -537 4844 -471 4860
rect -537 4810 -521 4844
rect -487 4810 -471 4844
rect -537 4794 -471 4810
rect -419 4844 -353 4860
rect -419 4810 -403 4844
rect -369 4810 -353 4844
rect -419 4794 -353 4810
rect -301 4844 -235 4860
rect -301 4810 -285 4844
rect -251 4810 -235 4844
rect -301 4794 -235 4810
rect -183 4844 -117 4860
rect -183 4810 -167 4844
rect -133 4810 -117 4844
rect -183 4794 -117 4810
rect -65 4844 1 4860
rect -65 4810 -49 4844
rect -15 4810 1 4844
rect -65 4794 1 4810
rect 53 4844 119 4860
rect 53 4810 69 4844
rect 103 4810 119 4844
rect 53 4794 119 4810
rect 171 4844 237 4860
rect 171 4810 187 4844
rect 221 4810 237 4844
rect 171 4794 237 4810
rect 289 4844 355 4860
rect 289 4810 305 4844
rect 339 4810 355 4844
rect 289 4794 355 4810
rect 407 4844 473 4860
rect 407 4810 423 4844
rect 457 4810 473 4844
rect 407 4794 473 4810
rect 525 4844 591 4860
rect 525 4810 541 4844
rect 575 4810 591 4844
rect 525 4794 591 4810
rect 643 4844 709 4860
rect 643 4810 659 4844
rect 693 4810 709 4844
rect 643 4794 709 4810
rect 761 4844 827 4860
rect 761 4810 777 4844
rect 811 4810 827 4844
rect 761 4794 827 4810
rect 879 4844 945 4860
rect 879 4810 895 4844
rect 929 4810 945 4844
rect 879 4794 945 4810
rect 997 4844 1063 4860
rect 997 4810 1013 4844
rect 1047 4810 1063 4844
rect 997 4794 1063 4810
rect 1115 4844 1181 4860
rect 1115 4810 1131 4844
rect 1165 4810 1181 4844
rect 1115 4794 1181 4810
rect 1233 4844 1299 4860
rect 1233 4810 1249 4844
rect 1283 4810 1299 4844
rect 1233 4794 1299 4810
rect 1351 4844 1417 4860
rect 1351 4810 1367 4844
rect 1401 4810 1417 4844
rect 1351 4794 1417 4810
rect 1469 4844 1535 4860
rect 1469 4810 1485 4844
rect 1519 4810 1535 4844
rect 1469 4794 1535 4810
rect 1587 4844 1653 4860
rect 1587 4810 1603 4844
rect 1637 4810 1653 4844
rect 1587 4794 1653 4810
rect 1705 4844 1771 4860
rect 1705 4810 1721 4844
rect 1755 4810 1771 4844
rect 1705 4794 1771 4810
rect 1823 4844 1889 4860
rect 1823 4810 1839 4844
rect 1873 4810 1889 4844
rect 1823 4794 1889 4810
rect 1941 4844 2007 4860
rect 1941 4810 1957 4844
rect 1991 4810 2007 4844
rect 1941 4794 2007 4810
rect 2059 4844 2125 4860
rect 2059 4810 2075 4844
rect 2109 4810 2125 4844
rect 2059 4794 2125 4810
rect 2177 4844 2243 4860
rect 2177 4810 2193 4844
rect 2227 4810 2243 4844
rect 2177 4794 2243 4810
rect 2295 4844 2361 4860
rect 2295 4810 2311 4844
rect 2345 4810 2361 4844
rect 2295 4794 2361 4810
rect 2413 4844 2479 4860
rect 2413 4810 2429 4844
rect 2463 4810 2479 4844
rect 2413 4794 2479 4810
rect 2531 4844 2597 4860
rect 2531 4810 2547 4844
rect 2581 4810 2597 4844
rect 2531 4794 2597 4810
rect 2649 4844 2715 4860
rect 2649 4810 2665 4844
rect 2699 4810 2715 4844
rect 2649 4794 2715 4810
rect 2767 4844 2833 4860
rect 2767 4810 2783 4844
rect 2817 4810 2833 4844
rect 2767 4794 2833 4810
rect 2885 4844 2951 4860
rect 2885 4810 2901 4844
rect 2935 4810 2951 4844
rect 2885 4794 2951 4810
rect 3003 4844 3069 4860
rect 3003 4810 3019 4844
rect 3053 4810 3069 4844
rect 3003 4794 3069 4810
rect 3121 4844 3187 4860
rect 3121 4810 3137 4844
rect 3171 4810 3187 4844
rect 3121 4794 3187 4810
rect 3239 4844 3305 4860
rect 3239 4810 3255 4844
rect 3289 4810 3305 4844
rect 3239 4794 3305 4810
rect 3357 4844 3423 4860
rect 3357 4810 3373 4844
rect 3407 4810 3423 4844
rect 3357 4794 3423 4810
rect 3475 4844 3541 4860
rect 3475 4810 3491 4844
rect 3525 4810 3541 4844
rect 3475 4794 3541 4810
rect 3593 4844 3659 4860
rect 3593 4810 3609 4844
rect 3643 4810 3659 4844
rect 3593 4794 3659 4810
rect 3711 4844 3777 4860
rect 3711 4810 3727 4844
rect 3761 4810 3777 4844
rect 3711 4794 3777 4810
rect 3829 4844 3895 4860
rect 3829 4810 3845 4844
rect 3879 4810 3895 4844
rect 3829 4794 3895 4810
<< polycont >>
rect -1229 6938 -1195 6972
rect -1111 6938 -1077 6972
rect -993 6938 -959 6972
rect -875 6938 -841 6972
rect -757 6938 -723 6972
rect -639 6938 -605 6972
rect -521 6938 -487 6972
rect -403 6938 -369 6972
rect -285 6938 -251 6972
rect -167 6938 -133 6972
rect -49 6938 -15 6972
rect 69 6938 103 6972
rect 187 6938 221 6972
rect 305 6938 339 6972
rect 423 6938 457 6972
rect 541 6938 575 6972
rect 659 6938 693 6972
rect 777 6938 811 6972
rect 895 6938 929 6972
rect 1013 6938 1047 6972
rect 1603 6938 1637 6972
rect 1721 6938 1755 6972
rect 1839 6938 1873 6972
rect 1957 6938 1991 6972
rect 2075 6938 2109 6972
rect 2193 6938 2227 6972
rect 2311 6938 2345 6972
rect 2429 6938 2463 6972
rect 2547 6938 2581 6972
rect 2665 6938 2699 6972
rect 2783 6938 2817 6972
rect 2901 6938 2935 6972
rect 3019 6938 3053 6972
rect 3137 6938 3171 6972
rect 3255 6938 3289 6972
rect 3373 6938 3407 6972
rect 3491 6938 3525 6972
rect 3609 6938 3643 6972
rect 3727 6938 3761 6972
rect 3845 6938 3879 6972
rect -1229 4810 -1195 4844
rect -1111 4810 -1077 4844
rect -993 4810 -959 4844
rect -875 4810 -841 4844
rect -757 4810 -723 4844
rect -639 4810 -605 4844
rect -521 4810 -487 4844
rect -403 4810 -369 4844
rect -285 4810 -251 4844
rect -167 4810 -133 4844
rect -49 4810 -15 4844
rect 69 4810 103 4844
rect 187 4810 221 4844
rect 305 4810 339 4844
rect 423 4810 457 4844
rect 541 4810 575 4844
rect 659 4810 693 4844
rect 777 4810 811 4844
rect 895 4810 929 4844
rect 1013 4810 1047 4844
rect 1131 4810 1165 4844
rect 1249 4810 1283 4844
rect 1367 4810 1401 4844
rect 1485 4810 1519 4844
rect 1603 4810 1637 4844
rect 1721 4810 1755 4844
rect 1839 4810 1873 4844
rect 1957 4810 1991 4844
rect 2075 4810 2109 4844
rect 2193 4810 2227 4844
rect 2311 4810 2345 4844
rect 2429 4810 2463 4844
rect 2547 4810 2581 4844
rect 2665 4810 2699 4844
rect 2783 4810 2817 4844
rect 2901 4810 2935 4844
rect 3019 4810 3053 4844
rect 3137 4810 3171 4844
rect 3255 4810 3289 4844
rect 3373 4810 3407 4844
rect 3491 4810 3525 4844
rect 3609 4810 3643 4844
rect 3727 4810 3761 4844
rect 3845 4810 3879 4844
<< locali >>
rect -1402 7040 -1306 7074
rect 3956 7040 4052 7074
rect -1402 6978 -1368 7040
rect 4018 6978 4052 7040
rect -1245 6938 -1229 6972
rect -1195 6938 -1179 6972
rect -1127 6938 -1111 6972
rect -1077 6938 -1061 6972
rect -1009 6938 -993 6972
rect -959 6938 -943 6972
rect -891 6938 -875 6972
rect -841 6938 -825 6972
rect -773 6938 -757 6972
rect -723 6938 -707 6972
rect -655 6938 -639 6972
rect -605 6938 -589 6972
rect -537 6938 -521 6972
rect -487 6938 -471 6972
rect -419 6938 -403 6972
rect -369 6938 -353 6972
rect -301 6938 -285 6972
rect -251 6938 -235 6972
rect -183 6938 -167 6972
rect -133 6938 -117 6972
rect -65 6938 -49 6972
rect -15 6938 1 6972
rect 53 6938 69 6972
rect 103 6938 119 6972
rect 171 6938 187 6972
rect 221 6938 237 6972
rect 289 6938 305 6972
rect 339 6938 355 6972
rect 407 6938 423 6972
rect 457 6938 473 6972
rect 525 6938 541 6972
rect 575 6938 591 6972
rect 643 6938 659 6972
rect 693 6938 709 6972
rect 761 6938 777 6972
rect 811 6938 827 6972
rect 879 6938 895 6972
rect 929 6938 945 6972
rect 997 6938 1013 6972
rect 1047 6938 1063 6972
rect 1587 6938 1603 6972
rect 1637 6938 1653 6972
rect 1705 6938 1721 6972
rect 1755 6938 1771 6972
rect 1823 6938 1839 6972
rect 1873 6938 1889 6972
rect 1941 6938 1957 6972
rect 1991 6938 2007 6972
rect 2059 6938 2075 6972
rect 2109 6938 2125 6972
rect 2177 6938 2193 6972
rect 2227 6938 2243 6972
rect 2295 6938 2311 6972
rect 2345 6938 2361 6972
rect 2413 6938 2429 6972
rect 2463 6938 2479 6972
rect 2531 6938 2547 6972
rect 2581 6938 2597 6972
rect 2649 6938 2665 6972
rect 2699 6938 2715 6972
rect 2767 6938 2783 6972
rect 2817 6938 2833 6972
rect 2885 6938 2901 6972
rect 2935 6938 2951 6972
rect 3003 6938 3019 6972
rect 3053 6938 3069 6972
rect 3121 6938 3137 6972
rect 3171 6938 3187 6972
rect 3239 6938 3255 6972
rect 3289 6938 3305 6972
rect 3357 6938 3373 6972
rect 3407 6938 3423 6972
rect 3475 6938 3491 6972
rect 3525 6938 3541 6972
rect 3593 6938 3609 6972
rect 3643 6938 3659 6972
rect 3711 6938 3727 6972
rect 3761 6938 3777 6972
rect 3829 6938 3845 6972
rect 3879 6938 3895 6972
rect -1288 6879 -1254 6895
rect -1288 4887 -1254 4903
rect -1170 6879 -1136 6895
rect -1170 4887 -1136 4903
rect -1052 6879 -1018 6895
rect -1052 4887 -1018 4903
rect -934 6879 -900 6895
rect -934 4887 -900 4903
rect -816 6879 -782 6895
rect -816 4887 -782 4903
rect -698 6879 -664 6895
rect -698 4887 -664 4903
rect -580 6879 -546 6895
rect -580 4887 -546 4903
rect -462 6879 -428 6895
rect -462 4887 -428 4903
rect -344 6879 -310 6895
rect -344 4887 -310 4903
rect -226 6879 -192 6895
rect -226 4887 -192 4903
rect -108 6879 -74 6895
rect -108 4887 -74 4903
rect 10 6879 44 6895
rect 10 4887 44 4903
rect 128 6879 162 6895
rect 128 4887 162 4903
rect 246 6879 280 6895
rect 246 4887 280 4903
rect 364 6879 398 6895
rect 364 4887 398 4903
rect 482 6879 516 6895
rect 482 4887 516 4903
rect 600 6879 634 6895
rect 600 4887 634 4903
rect 718 6879 752 6895
rect 718 4887 752 4903
rect 836 6879 870 6895
rect 836 4887 870 4903
rect 954 6879 988 6895
rect 954 4887 988 4903
rect 1072 6879 1106 6895
rect 1072 4887 1106 4903
rect 1190 6879 1224 6895
rect 1190 4887 1224 4903
rect 1308 6879 1342 6895
rect 1308 4887 1342 4903
rect 1426 6879 1460 6895
rect 1426 4887 1460 4903
rect 1544 6879 1578 6895
rect 1544 4887 1578 4903
rect 1662 6879 1696 6895
rect 1662 4887 1696 4903
rect 1780 6879 1814 6895
rect 1780 4887 1814 4903
rect 1898 6879 1932 6895
rect 1898 4887 1932 4903
rect 2016 6879 2050 6895
rect 2016 4887 2050 4903
rect 2134 6879 2168 6895
rect 2134 4887 2168 4903
rect 2252 6879 2286 6895
rect 2252 4887 2286 4903
rect 2370 6879 2404 6895
rect 2370 4887 2404 4903
rect 2488 6879 2522 6895
rect 2488 4887 2522 4903
rect 2606 6879 2640 6895
rect 2606 4887 2640 4903
rect 2724 6879 2758 6895
rect 2724 4887 2758 4903
rect 2842 6879 2876 6895
rect 2842 4887 2876 4903
rect 2960 6879 2994 6895
rect 2960 4887 2994 4903
rect 3078 6879 3112 6895
rect 3078 4887 3112 4903
rect 3196 6879 3230 6895
rect 3196 4887 3230 4903
rect 3314 6879 3348 6895
rect 3314 4887 3348 4903
rect 3432 6879 3466 6895
rect 3432 4887 3466 4903
rect 3550 6879 3584 6895
rect 3550 4887 3584 4903
rect 3668 6879 3702 6895
rect 3668 4887 3702 4903
rect 3786 6879 3820 6895
rect 3786 4887 3820 4903
rect 3904 6879 3938 6895
rect 3904 4887 3938 4903
rect -1245 4810 -1229 4844
rect -1195 4810 -1179 4844
rect -1127 4810 -1111 4844
rect -1077 4810 -1061 4844
rect -1009 4810 -993 4844
rect -959 4810 -943 4844
rect -891 4810 -875 4844
rect -841 4810 -825 4844
rect -773 4810 -757 4844
rect -723 4810 -707 4844
rect -655 4810 -639 4844
rect -605 4810 -589 4844
rect -537 4810 -521 4844
rect -487 4810 -471 4844
rect -419 4810 -403 4844
rect -369 4810 -353 4844
rect -301 4810 -285 4844
rect -251 4810 -235 4844
rect -183 4810 -167 4844
rect -133 4810 -117 4844
rect -65 4810 -49 4844
rect -15 4810 1 4844
rect 53 4810 69 4844
rect 103 4810 119 4844
rect 171 4810 187 4844
rect 221 4810 237 4844
rect 289 4810 305 4844
rect 339 4810 355 4844
rect 407 4810 423 4844
rect 457 4810 473 4844
rect 525 4810 541 4844
rect 575 4810 591 4844
rect 643 4810 659 4844
rect 693 4810 709 4844
rect 761 4810 777 4844
rect 811 4810 827 4844
rect 879 4810 895 4844
rect 929 4810 945 4844
rect 997 4810 1013 4844
rect 1047 4810 1063 4844
rect 1115 4810 1131 4844
rect 1165 4810 1181 4844
rect 1233 4810 1249 4844
rect 1283 4810 1299 4844
rect 1351 4810 1367 4844
rect 1401 4810 1417 4844
rect 1469 4810 1485 4844
rect 1519 4810 1535 4844
rect 1587 4810 1603 4844
rect 1637 4810 1653 4844
rect 1705 4810 1721 4844
rect 1755 4810 1771 4844
rect 1823 4810 1839 4844
rect 1873 4810 1889 4844
rect 1941 4810 1957 4844
rect 1991 4810 2007 4844
rect 2059 4810 2075 4844
rect 2109 4810 2125 4844
rect 2177 4810 2193 4844
rect 2227 4810 2243 4844
rect 2295 4810 2311 4844
rect 2345 4810 2361 4844
rect 2413 4810 2429 4844
rect 2463 4810 2479 4844
rect 2531 4810 2547 4844
rect 2581 4810 2597 4844
rect 2649 4810 2665 4844
rect 2699 4810 2715 4844
rect 2767 4810 2783 4844
rect 2817 4810 2833 4844
rect 2885 4810 2901 4844
rect 2935 4810 2951 4844
rect 3003 4810 3019 4844
rect 3053 4810 3069 4844
rect 3121 4810 3137 4844
rect 3171 4810 3187 4844
rect 3239 4810 3255 4844
rect 3289 4810 3305 4844
rect 3357 4810 3373 4844
rect 3407 4810 3423 4844
rect 3475 4810 3491 4844
rect 3525 4810 3541 4844
rect 3593 4810 3609 4844
rect 3643 4810 3659 4844
rect 3711 4810 3727 4844
rect 3761 4810 3777 4844
rect 3829 4810 3845 4844
rect 3879 4810 3895 4844
rect -1402 4742 -1368 4804
rect 4018 4742 4052 4804
rect -1402 4708 -1306 4742
rect 3956 4708 4052 4742
<< viali >>
rect -1229 6938 -1195 6972
rect -1111 6938 -1077 6972
rect -993 6938 -959 6972
rect -875 6938 -841 6972
rect -757 6938 -723 6972
rect -639 6938 -605 6972
rect -521 6938 -487 6972
rect -403 6938 -369 6972
rect -285 6938 -251 6972
rect -167 6938 -133 6972
rect -49 6938 -15 6972
rect 69 6938 103 6972
rect 187 6938 221 6972
rect 305 6938 339 6972
rect 423 6938 457 6972
rect 541 6938 575 6972
rect 659 6938 693 6972
rect 777 6938 811 6972
rect 895 6938 929 6972
rect 1013 6938 1047 6972
rect 1603 6938 1637 6972
rect 1721 6938 1755 6972
rect 1839 6938 1873 6972
rect 1957 6938 1991 6972
rect 2075 6938 2109 6972
rect 2193 6938 2227 6972
rect 2311 6938 2345 6972
rect 2429 6938 2463 6972
rect 2547 6938 2581 6972
rect 2665 6938 2699 6972
rect 2783 6938 2817 6972
rect 2901 6938 2935 6972
rect 3019 6938 3053 6972
rect 3137 6938 3171 6972
rect 3255 6938 3289 6972
rect 3373 6938 3407 6972
rect 3491 6938 3525 6972
rect 3609 6938 3643 6972
rect 3727 6938 3761 6972
rect 3845 6938 3879 6972
rect -1402 6491 -1368 6891
rect -1402 4891 -1368 5291
rect -1288 4903 -1254 6879
rect -1170 4903 -1136 6879
rect -1052 4903 -1018 6879
rect -934 4903 -900 6879
rect -816 4903 -782 6879
rect -698 4903 -664 6879
rect -580 4903 -546 6879
rect -462 4903 -428 6879
rect -344 4903 -310 6879
rect -226 4903 -192 6879
rect -108 4903 -74 6879
rect 10 4903 44 6879
rect 128 4903 162 6879
rect 246 4903 280 6879
rect 364 4903 398 6879
rect 482 4903 516 6879
rect 600 4903 634 6879
rect 718 4903 752 6879
rect 836 4903 870 6879
rect 954 4903 988 6879
rect 1072 4903 1106 6879
rect 1190 4903 1224 6879
rect 1308 4903 1342 6879
rect 1426 4903 1460 6879
rect 1544 4903 1578 6879
rect 1662 4903 1696 6879
rect 1780 4903 1814 6879
rect 1898 4903 1932 6879
rect 2016 4903 2050 6879
rect 2134 4903 2168 6879
rect 2252 4903 2286 6879
rect 2370 4903 2404 6879
rect 2488 4903 2522 6879
rect 2606 4903 2640 6879
rect 2724 4903 2758 6879
rect 2842 4903 2876 6879
rect 2960 4903 2994 6879
rect 3078 4903 3112 6879
rect 3196 4903 3230 6879
rect 3314 4903 3348 6879
rect 3432 4903 3466 6879
rect 3550 4903 3584 6879
rect 3668 4903 3702 6879
rect 3786 4903 3820 6879
rect 3904 4903 3938 6879
rect 4018 6491 4052 6891
rect 4018 4891 4052 5291
rect -1229 4810 -1195 4844
rect -1111 4810 -1077 4844
rect -993 4810 -959 4844
rect -875 4810 -841 4844
rect -757 4810 -723 4844
rect -639 4810 -605 4844
rect -521 4810 -487 4844
rect -403 4810 -369 4844
rect -285 4810 -251 4844
rect -167 4810 -133 4844
rect -49 4810 -15 4844
rect 69 4810 103 4844
rect 187 4810 221 4844
rect 305 4810 339 4844
rect 423 4810 457 4844
rect 541 4810 575 4844
rect 659 4810 693 4844
rect 777 4810 811 4844
rect 895 4810 929 4844
rect 1013 4810 1047 4844
rect 1131 4810 1165 4844
rect 1249 4810 1283 4844
rect 1367 4810 1401 4844
rect 1485 4810 1519 4844
rect 1603 4810 1637 4844
rect 1721 4810 1755 4844
rect 1839 4810 1873 4844
rect 1957 4810 1991 4844
rect 2075 4810 2109 4844
rect 2193 4810 2227 4844
rect 2311 4810 2345 4844
rect 2429 4810 2463 4844
rect 2547 4810 2581 4844
rect 2665 4810 2699 4844
rect 2783 4810 2817 4844
rect 2901 4810 2935 4844
rect 3019 4810 3053 4844
rect 3137 4810 3171 4844
rect 3255 4810 3289 4844
rect 3373 4810 3407 4844
rect 3491 4810 3525 4844
rect 3609 4810 3643 4844
rect 3727 4810 3761 4844
rect 3845 4810 3879 4844
<< metal1 >>
rect -1297 6972 -1065 6978
rect -1297 6938 -1229 6972
rect -1195 6938 -1111 6972
rect -1077 6938 -1065 6972
rect -1297 6932 -1065 6938
rect -1005 6972 1059 6978
rect -1005 6938 -993 6972
rect -959 6938 -875 6972
rect -841 6938 -757 6972
rect -723 6938 -639 6972
rect -605 6938 -521 6972
rect -487 6938 -403 6972
rect -369 6938 -285 6972
rect -251 6938 -167 6972
rect -133 6938 -49 6972
rect -15 6938 69 6972
rect 103 6938 187 6972
rect 221 6938 305 6972
rect 339 6938 423 6972
rect 457 6938 541 6972
rect 575 6938 659 6972
rect 693 6938 777 6972
rect 811 6938 895 6972
rect 929 6938 1013 6972
rect 1047 6938 1059 6972
rect -1005 6932 1059 6938
rect 1591 6972 3655 6978
rect 1591 6938 1603 6972
rect 1637 6938 1721 6972
rect 1755 6938 1839 6972
rect 1873 6938 1957 6972
rect 1991 6938 2075 6972
rect 2109 6938 2193 6972
rect 2227 6938 2311 6972
rect 2345 6938 2429 6972
rect 2463 6938 2547 6972
rect 2581 6938 2665 6972
rect 2699 6938 2783 6972
rect 2817 6938 2901 6972
rect 2935 6938 3019 6972
rect 3053 6938 3137 6972
rect 3171 6938 3255 6972
rect 3289 6938 3373 6972
rect 3407 6938 3491 6972
rect 3525 6938 3609 6972
rect 3643 6938 3655 6972
rect 1591 6932 3655 6938
rect 3715 6972 3947 6978
rect 3715 6938 3727 6972
rect 3761 6938 3845 6972
rect 3879 6938 3947 6972
rect 3715 6932 3947 6938
rect -1408 6891 -1362 6903
rect -1297 6891 -1245 6932
rect -1408 6491 -1402 6891
rect -1368 6879 -1245 6891
rect -1368 6491 -1297 6879
rect -1408 6479 -1362 6491
rect -1408 5291 -1362 5303
rect -1408 4891 -1402 5291
rect -1368 4903 -1297 5291
rect -1368 4891 -1245 4903
rect -1408 4879 -1362 4891
rect -1297 4850 -1245 4891
rect -1179 6879 -1127 6932
rect -1179 4850 -1127 4903
rect -1061 6879 -1009 6891
rect -1061 4891 -1009 4903
rect -943 6879 -891 6891
rect -943 4891 -891 4903
rect -825 6879 -773 6891
rect -825 4891 -773 4903
rect -707 6879 -655 6891
rect -707 4891 -655 4903
rect -589 6879 -537 6891
rect -589 4891 -537 4903
rect -471 6879 -419 6891
rect -471 4891 -419 4903
rect -353 6879 -301 6891
rect -353 4891 -301 4903
rect -235 6879 -183 6891
rect -235 4891 -183 4903
rect -117 6879 -65 6891
rect -117 4891 -65 4903
rect 1 6879 53 6891
rect 1 4891 53 4903
rect 119 6879 171 6891
rect 119 4891 171 4903
rect 237 6879 289 6891
rect 237 4891 289 4903
rect 355 6879 407 6891
rect 355 4891 407 4903
rect 473 6879 525 6891
rect 473 4891 525 4903
rect 591 6879 643 6891
rect 591 4891 643 4903
rect 709 6879 761 6891
rect 709 4891 761 4903
rect 827 6879 879 6891
rect 827 4891 879 4903
rect 945 6879 997 6932
rect 945 4850 997 4903
rect 1063 6879 1115 6891
rect 1063 4891 1115 4903
rect 1181 6879 1233 6891
rect 1181 4891 1233 4903
rect 1299 6879 1351 6891
rect 1299 4891 1351 4903
rect 1417 6879 1469 6891
rect 1417 4891 1469 4903
rect 1535 6879 1587 6891
rect 1535 4891 1587 4903
rect 1653 6879 1705 6932
rect 1233 4850 1299 4856
rect 1653 4850 1705 4903
rect 1771 6879 1823 6891
rect 1771 4891 1823 4903
rect 1889 6879 1941 6891
rect 1889 4891 1941 4903
rect 2007 6879 2059 6891
rect 2007 4891 2059 4903
rect 2125 6879 2177 6891
rect 2125 4891 2177 4903
rect 2243 6879 2295 6891
rect 2243 4891 2295 4903
rect 2361 6879 2413 6891
rect 2361 4891 2413 4903
rect 2479 6879 2531 6891
rect 2479 4891 2531 4903
rect 2597 6879 2649 6891
rect 2597 4891 2649 4903
rect 2715 6879 2767 6891
rect 2715 4891 2767 4903
rect 2833 6879 2885 6891
rect 2833 4891 2885 4903
rect 2951 6879 3003 6891
rect 2951 4891 3003 4903
rect 3069 6879 3121 6891
rect 3069 4891 3121 4903
rect 3187 6879 3239 6891
rect 3187 4891 3239 4903
rect 3305 6879 3357 6891
rect 3305 4891 3357 4903
rect 3423 6879 3475 6891
rect 3423 4891 3475 4903
rect 3541 6879 3593 6891
rect 3541 4891 3593 4903
rect 3659 6879 3711 6891
rect 3659 4891 3711 4903
rect 3777 6879 3829 6932
rect 3777 4850 3829 4903
rect 3895 6891 3947 6932
rect 4012 6891 4058 6903
rect 3895 6879 4018 6891
rect 3947 6491 4018 6879
rect 4052 6491 4058 6891
rect 4012 6479 4058 6491
rect 4012 5291 4058 5303
rect 3947 4903 4018 5291
rect 3895 4891 4018 4903
rect 4052 4891 4058 5291
rect 3895 4850 3947 4891
rect 4012 4879 4058 4891
rect -1297 4844 -1065 4850
rect -1297 4810 -1229 4844
rect -1195 4810 -1111 4844
rect -1077 4810 -1065 4844
rect -1297 4804 -1065 4810
rect -1005 4844 1237 4850
rect -1005 4810 -993 4844
rect -959 4810 -875 4844
rect -841 4810 -757 4844
rect -723 4810 -639 4844
rect -605 4810 -521 4844
rect -487 4810 -403 4844
rect -369 4810 -285 4844
rect -251 4810 -167 4844
rect -133 4810 -49 4844
rect -15 4810 69 4844
rect 103 4810 187 4844
rect 221 4810 305 4844
rect 339 4810 423 4844
rect 457 4810 541 4844
rect 575 4810 659 4844
rect 693 4810 777 4844
rect 811 4810 895 4844
rect 929 4810 1013 4844
rect 1047 4810 1131 4844
rect 1165 4810 1237 4844
rect -1005 4804 1237 4810
rect 1233 4793 1237 4804
rect 1296 4793 1299 4850
rect 1233 4787 1299 4793
rect 1355 4844 3655 4850
rect 1355 4810 1367 4844
rect 1401 4810 1485 4844
rect 1519 4810 1603 4844
rect 1637 4810 1721 4844
rect 1755 4810 1839 4844
rect 1873 4810 1957 4844
rect 1991 4810 2075 4844
rect 2109 4810 2193 4844
rect 2227 4810 2311 4844
rect 2345 4810 2429 4844
rect 2463 4810 2547 4844
rect 2581 4810 2665 4844
rect 2699 4810 2783 4844
rect 2817 4810 2901 4844
rect 2935 4810 3019 4844
rect 3053 4810 3137 4844
rect 3171 4810 3255 4844
rect 3289 4810 3373 4844
rect 3407 4810 3491 4844
rect 3525 4810 3609 4844
rect 3643 4810 3655 4844
rect 1355 4804 3655 4810
rect 3715 4844 3947 4850
rect 3715 4810 3727 4844
rect 3761 4810 3845 4844
rect 3879 4810 3947 4844
rect 3715 4804 3947 4810
rect 1355 4793 1414 4804
rect 1355 4730 1414 4736
<< via1 >>
rect -1297 4903 -1288 6879
rect -1288 4903 -1254 6879
rect -1254 4903 -1245 6879
rect -1179 4903 -1170 6879
rect -1170 4903 -1136 6879
rect -1136 4903 -1127 6879
rect -1061 4903 -1052 6879
rect -1052 4903 -1018 6879
rect -1018 4903 -1009 6879
rect -943 4903 -934 6879
rect -934 4903 -900 6879
rect -900 4903 -891 6879
rect -825 4903 -816 6879
rect -816 4903 -782 6879
rect -782 4903 -773 6879
rect -707 4903 -698 6879
rect -698 4903 -664 6879
rect -664 4903 -655 6879
rect -589 4903 -580 6879
rect -580 4903 -546 6879
rect -546 4903 -537 6879
rect -471 4903 -462 6879
rect -462 4903 -428 6879
rect -428 4903 -419 6879
rect -353 4903 -344 6879
rect -344 4903 -310 6879
rect -310 4903 -301 6879
rect -235 4903 -226 6879
rect -226 4903 -192 6879
rect -192 4903 -183 6879
rect -117 4903 -108 6879
rect -108 4903 -74 6879
rect -74 4903 -65 6879
rect 1 4903 10 6879
rect 10 4903 44 6879
rect 44 4903 53 6879
rect 119 4903 128 6879
rect 128 4903 162 6879
rect 162 4903 171 6879
rect 237 4903 246 6879
rect 246 4903 280 6879
rect 280 4903 289 6879
rect 355 4903 364 6879
rect 364 4903 398 6879
rect 398 4903 407 6879
rect 473 4903 482 6879
rect 482 4903 516 6879
rect 516 4903 525 6879
rect 591 4903 600 6879
rect 600 4903 634 6879
rect 634 4903 643 6879
rect 709 4903 718 6879
rect 718 4903 752 6879
rect 752 4903 761 6879
rect 827 4903 836 6879
rect 836 4903 870 6879
rect 870 4903 879 6879
rect 945 4903 954 6879
rect 954 4903 988 6879
rect 988 4903 997 6879
rect 1063 4903 1072 6879
rect 1072 4903 1106 6879
rect 1106 4903 1115 6879
rect 1181 4903 1190 6879
rect 1190 4903 1224 6879
rect 1224 4903 1233 6879
rect 1299 4903 1308 6879
rect 1308 4903 1342 6879
rect 1342 4903 1351 6879
rect 1417 4903 1426 6879
rect 1426 4903 1460 6879
rect 1460 4903 1469 6879
rect 1535 4903 1544 6879
rect 1544 4903 1578 6879
rect 1578 4903 1587 6879
rect 1653 4903 1662 6879
rect 1662 4903 1696 6879
rect 1696 4903 1705 6879
rect 1771 4903 1780 6879
rect 1780 4903 1814 6879
rect 1814 4903 1823 6879
rect 1889 4903 1898 6879
rect 1898 4903 1932 6879
rect 1932 4903 1941 6879
rect 2007 4903 2016 6879
rect 2016 4903 2050 6879
rect 2050 4903 2059 6879
rect 2125 4903 2134 6879
rect 2134 4903 2168 6879
rect 2168 4903 2177 6879
rect 2243 4903 2252 6879
rect 2252 4903 2286 6879
rect 2286 4903 2295 6879
rect 2361 4903 2370 6879
rect 2370 4903 2404 6879
rect 2404 4903 2413 6879
rect 2479 4903 2488 6879
rect 2488 4903 2522 6879
rect 2522 4903 2531 6879
rect 2597 4903 2606 6879
rect 2606 4903 2640 6879
rect 2640 4903 2649 6879
rect 2715 4903 2724 6879
rect 2724 4903 2758 6879
rect 2758 4903 2767 6879
rect 2833 4903 2842 6879
rect 2842 4903 2876 6879
rect 2876 4903 2885 6879
rect 2951 4903 2960 6879
rect 2960 4903 2994 6879
rect 2994 4903 3003 6879
rect 3069 4903 3078 6879
rect 3078 4903 3112 6879
rect 3112 4903 3121 6879
rect 3187 4903 3196 6879
rect 3196 4903 3230 6879
rect 3230 4903 3239 6879
rect 3305 4903 3314 6879
rect 3314 4903 3348 6879
rect 3348 4903 3357 6879
rect 3423 4903 3432 6879
rect 3432 4903 3466 6879
rect 3466 4903 3475 6879
rect 3541 4903 3550 6879
rect 3550 4903 3584 6879
rect 3584 4903 3593 6879
rect 3659 4903 3668 6879
rect 3668 4903 3702 6879
rect 3702 4903 3711 6879
rect 3777 4903 3786 6879
rect 3786 4903 3820 6879
rect 3820 4903 3829 6879
rect 3895 4903 3904 6879
rect 3904 4903 3938 6879
rect 3938 4903 3947 6879
rect 1237 4844 1296 4850
rect 1237 4810 1249 4844
rect 1249 4810 1283 4844
rect 1283 4810 1296 4844
rect 1237 4793 1296 4810
rect 1355 4736 1414 4793
<< metal2 >>
rect -1297 7040 3947 7142
rect -1297 6879 -1245 7040
rect -1297 4891 -1245 4903
rect -1179 6879 -1127 7040
rect -1179 4891 -1127 4903
rect -1061 6879 -1009 7040
rect -1061 4891 -1009 4903
rect -943 6879 -891 6891
rect -943 4742 -891 4903
rect -825 6879 -773 7040
rect -825 4891 -773 4903
rect -707 6879 -655 6891
rect -707 4742 -655 4903
rect -589 6879 -537 7040
rect -589 4891 -537 4903
rect -471 6879 -419 6891
rect -471 4742 -419 4903
rect -353 6879 -301 7040
rect -353 4891 -301 4903
rect -235 6879 -183 6891
rect -235 4742 -183 4903
rect -117 6879 -65 7040
rect -117 4891 -65 4903
rect 1 6879 53 6891
rect 1 4742 53 4903
rect 119 6879 171 7040
rect 119 4891 171 4903
rect 237 6879 289 6891
rect 237 4742 289 4903
rect 355 6879 407 7040
rect 355 4891 407 4903
rect 473 6879 525 6891
rect 473 4742 525 4903
rect 591 6879 643 7040
rect 591 4891 643 4903
rect 709 6879 761 6891
rect 709 4742 761 4903
rect 827 6879 879 7040
rect 827 4891 879 4903
rect 945 6879 997 6891
rect -943 4640 761 4742
rect 945 4708 997 4903
rect 1063 6879 1115 7040
rect 1063 4891 1115 4903
rect 1181 6879 1233 6891
rect 1181 4887 1233 4903
rect 1299 6879 1351 7040
rect 1299 4891 1351 4903
rect 1417 6879 1469 6891
rect 1417 4891 1469 4903
rect 1535 6879 1587 7040
rect 1535 4891 1587 4903
rect 1653 6879 1705 6891
rect 1181 4758 1209 4887
rect 1440 4856 1468 4891
rect 1237 4850 1468 4856
rect 1296 4828 1468 4850
rect 1296 4793 1299 4828
rect 1237 4787 1299 4793
rect 1355 4793 1414 4799
rect 1181 4736 1355 4758
rect 1181 4730 1414 4736
rect 1653 4707 1705 4903
rect 1771 6879 1823 7040
rect 1889 6879 1941 6891
rect 1771 4891 1823 4903
rect 1888 4903 1889 4971
rect 1888 4891 1941 4903
rect 2007 6879 2059 7040
rect 2125 6879 2177 6891
rect 2007 4891 2059 4903
rect 2124 4903 2125 4971
rect 2124 4891 2177 4903
rect 2243 6879 2295 7040
rect 2361 6879 2413 6891
rect 2243 4891 2295 4903
rect 2360 4903 2361 4971
rect 2360 4891 2413 4903
rect 2479 6879 2531 7040
rect 2597 6879 2649 6891
rect 2479 4891 2531 4903
rect 2596 4903 2597 4971
rect 2596 4891 2649 4903
rect 2715 6879 2767 7040
rect 2833 6879 2885 6891
rect 2715 4891 2767 4903
rect 2832 4903 2833 4971
rect 2832 4891 2885 4903
rect 2951 6879 3003 7040
rect 3069 6879 3121 6891
rect 2951 4891 3003 4903
rect 3068 4903 3069 4971
rect 3068 4891 3121 4903
rect 3187 6879 3239 7040
rect 3305 6879 3357 6891
rect 3187 4891 3239 4903
rect 3304 4903 3305 4971
rect 3304 4891 3357 4903
rect 3423 6879 3475 7040
rect 3541 6879 3593 6891
rect 3423 4891 3475 4903
rect 3540 4903 3541 4971
rect 3540 4891 3593 4903
rect 3659 6879 3711 7040
rect 3777 6879 3829 7040
rect 3659 4891 3711 4903
rect 3776 4903 3777 4971
rect 3776 4891 3829 4903
rect 3895 6879 3947 7040
rect 3895 4891 3947 4903
rect 1888 4742 1940 4891
rect 2124 4742 2176 4891
rect 2360 4742 2412 4891
rect 2596 4742 2648 4891
rect 2832 4742 2884 4891
rect 3068 4742 3120 4891
rect 3304 4742 3356 4891
rect 3540 4742 3592 4891
rect 1888 4640 3592 4742
<< labels >>
rlabel metal2 -1297 7098 -1233 7142 1 VDD
rlabel metal2 -943 4640 -872 4693 1 IOUT1
rlabel metal2 945 4708 997 4742 1 IIN1
rlabel metal2 1653 4707 1705 4741 1 IIN2
rlabel metal2 3540 4640 3592 4674 1 IOUT2
<< end >>
