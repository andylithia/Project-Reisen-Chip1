magic
tech sky130B
timestamp 1668465492
<< error_p >>
rect -1117 136 -1088 139
rect -907 136 -878 139
rect -697 136 -668 139
rect -487 136 -458 139
rect -277 136 -248 139
rect -67 136 -38 139
rect 143 136 172 139
rect 353 136 382 139
rect 563 136 592 139
rect 773 136 802 139
rect 983 136 1012 139
rect 1193 136 1222 139
rect -1117 119 -1111 136
rect -907 119 -901 136
rect -697 119 -691 136
rect -487 119 -481 136
rect -277 119 -271 136
rect -67 119 -61 136
rect 143 119 149 136
rect 353 119 359 136
rect 563 119 569 136
rect 773 119 779 136
rect 983 119 989 136
rect 1193 119 1199 136
rect -1117 116 -1088 119
rect -907 116 -878 119
rect -697 116 -668 119
rect -487 116 -458 119
rect -277 116 -248 119
rect -67 116 -38 119
rect 143 116 172 119
rect 353 116 382 119
rect 563 116 592 119
rect 773 116 802 119
rect 983 116 1012 119
rect 1193 116 1222 119
rect -1222 -119 -1193 -116
rect -1012 -119 -983 -116
rect -802 -119 -773 -116
rect -592 -119 -563 -116
rect -382 -119 -353 -116
rect -172 -119 -143 -116
rect 38 -119 67 -116
rect 248 -119 277 -116
rect 458 -119 487 -116
rect 668 -119 697 -116
rect 878 -119 907 -116
rect 1088 -119 1117 -116
rect -1222 -136 -1216 -119
rect -1012 -136 -1006 -119
rect -802 -136 -796 -119
rect -592 -136 -586 -119
rect -382 -136 -376 -119
rect -172 -136 -166 -119
rect 38 -136 44 -119
rect 248 -136 254 -119
rect 458 -136 464 -119
rect 668 -136 674 -119
rect 878 -136 884 -119
rect 1088 -136 1094 -119
rect -1222 -139 -1193 -136
rect -1012 -139 -983 -136
rect -802 -139 -773 -136
rect -592 -139 -563 -136
rect -382 -139 -353 -136
rect -172 -139 -143 -136
rect 38 -139 67 -136
rect 248 -139 277 -136
rect 458 -139 487 -136
rect 668 -139 697 -136
rect 878 -139 907 -136
rect 1088 -139 1117 -136
<< pwell >>
rect -1315 -205 1315 205
<< nmos >>
rect -1215 -100 -1200 100
rect -1110 -100 -1095 100
rect -1005 -100 -990 100
rect -900 -100 -885 100
rect -795 -100 -780 100
rect -690 -100 -675 100
rect -585 -100 -570 100
rect -480 -100 -465 100
rect -375 -100 -360 100
rect -270 -100 -255 100
rect -165 -100 -150 100
rect -60 -100 -45 100
rect 45 -100 60 100
rect 150 -100 165 100
rect 255 -100 270 100
rect 360 -100 375 100
rect 465 -100 480 100
rect 570 -100 585 100
rect 675 -100 690 100
rect 780 -100 795 100
rect 885 -100 900 100
rect 990 -100 1005 100
rect 1095 -100 1110 100
rect 1200 -100 1215 100
<< ndiff >>
rect -1246 94 -1215 100
rect -1246 -94 -1240 94
rect -1223 -94 -1215 94
rect -1246 -100 -1215 -94
rect -1200 94 -1169 100
rect -1200 -94 -1192 94
rect -1175 -94 -1169 94
rect -1200 -100 -1169 -94
rect -1141 94 -1110 100
rect -1141 -94 -1135 94
rect -1118 -94 -1110 94
rect -1141 -100 -1110 -94
rect -1095 94 -1064 100
rect -1095 -94 -1087 94
rect -1070 -94 -1064 94
rect -1095 -100 -1064 -94
rect -1036 94 -1005 100
rect -1036 -94 -1030 94
rect -1013 -94 -1005 94
rect -1036 -100 -1005 -94
rect -990 94 -959 100
rect -990 -94 -982 94
rect -965 -94 -959 94
rect -990 -100 -959 -94
rect -931 94 -900 100
rect -931 -94 -925 94
rect -908 -94 -900 94
rect -931 -100 -900 -94
rect -885 94 -854 100
rect -885 -94 -877 94
rect -860 -94 -854 94
rect -885 -100 -854 -94
rect -826 94 -795 100
rect -826 -94 -820 94
rect -803 -94 -795 94
rect -826 -100 -795 -94
rect -780 94 -749 100
rect -780 -94 -772 94
rect -755 -94 -749 94
rect -780 -100 -749 -94
rect -721 94 -690 100
rect -721 -94 -715 94
rect -698 -94 -690 94
rect -721 -100 -690 -94
rect -675 94 -644 100
rect -675 -94 -667 94
rect -650 -94 -644 94
rect -675 -100 -644 -94
rect -616 94 -585 100
rect -616 -94 -610 94
rect -593 -94 -585 94
rect -616 -100 -585 -94
rect -570 94 -539 100
rect -570 -94 -562 94
rect -545 -94 -539 94
rect -570 -100 -539 -94
rect -511 94 -480 100
rect -511 -94 -505 94
rect -488 -94 -480 94
rect -511 -100 -480 -94
rect -465 94 -434 100
rect -465 -94 -457 94
rect -440 -94 -434 94
rect -465 -100 -434 -94
rect -406 94 -375 100
rect -406 -94 -400 94
rect -383 -94 -375 94
rect -406 -100 -375 -94
rect -360 94 -329 100
rect -360 -94 -352 94
rect -335 -94 -329 94
rect -360 -100 -329 -94
rect -301 94 -270 100
rect -301 -94 -295 94
rect -278 -94 -270 94
rect -301 -100 -270 -94
rect -255 94 -224 100
rect -255 -94 -247 94
rect -230 -94 -224 94
rect -255 -100 -224 -94
rect -196 94 -165 100
rect -196 -94 -190 94
rect -173 -94 -165 94
rect -196 -100 -165 -94
rect -150 94 -119 100
rect -150 -94 -142 94
rect -125 -94 -119 94
rect -150 -100 -119 -94
rect -91 94 -60 100
rect -91 -94 -85 94
rect -68 -94 -60 94
rect -91 -100 -60 -94
rect -45 94 -14 100
rect -45 -94 -37 94
rect -20 -94 -14 94
rect -45 -100 -14 -94
rect 14 94 45 100
rect 14 -94 20 94
rect 37 -94 45 94
rect 14 -100 45 -94
rect 60 94 91 100
rect 60 -94 68 94
rect 85 -94 91 94
rect 60 -100 91 -94
rect 119 94 150 100
rect 119 -94 125 94
rect 142 -94 150 94
rect 119 -100 150 -94
rect 165 94 196 100
rect 165 -94 173 94
rect 190 -94 196 94
rect 165 -100 196 -94
rect 224 94 255 100
rect 224 -94 230 94
rect 247 -94 255 94
rect 224 -100 255 -94
rect 270 94 301 100
rect 270 -94 278 94
rect 295 -94 301 94
rect 270 -100 301 -94
rect 329 94 360 100
rect 329 -94 335 94
rect 352 -94 360 94
rect 329 -100 360 -94
rect 375 94 406 100
rect 375 -94 383 94
rect 400 -94 406 94
rect 375 -100 406 -94
rect 434 94 465 100
rect 434 -94 440 94
rect 457 -94 465 94
rect 434 -100 465 -94
rect 480 94 511 100
rect 480 -94 488 94
rect 505 -94 511 94
rect 480 -100 511 -94
rect 539 94 570 100
rect 539 -94 545 94
rect 562 -94 570 94
rect 539 -100 570 -94
rect 585 94 616 100
rect 585 -94 593 94
rect 610 -94 616 94
rect 585 -100 616 -94
rect 644 94 675 100
rect 644 -94 650 94
rect 667 -94 675 94
rect 644 -100 675 -94
rect 690 94 721 100
rect 690 -94 698 94
rect 715 -94 721 94
rect 690 -100 721 -94
rect 749 94 780 100
rect 749 -94 755 94
rect 772 -94 780 94
rect 749 -100 780 -94
rect 795 94 826 100
rect 795 -94 803 94
rect 820 -94 826 94
rect 795 -100 826 -94
rect 854 94 885 100
rect 854 -94 860 94
rect 877 -94 885 94
rect 854 -100 885 -94
rect 900 94 931 100
rect 900 -94 908 94
rect 925 -94 931 94
rect 900 -100 931 -94
rect 959 94 990 100
rect 959 -94 965 94
rect 982 -94 990 94
rect 959 -100 990 -94
rect 1005 94 1036 100
rect 1005 -94 1013 94
rect 1030 -94 1036 94
rect 1005 -100 1036 -94
rect 1064 94 1095 100
rect 1064 -94 1070 94
rect 1087 -94 1095 94
rect 1064 -100 1095 -94
rect 1110 94 1141 100
rect 1110 -94 1118 94
rect 1135 -94 1141 94
rect 1110 -100 1141 -94
rect 1169 94 1200 100
rect 1169 -94 1175 94
rect 1192 -94 1200 94
rect 1169 -100 1200 -94
rect 1215 94 1246 100
rect 1215 -94 1223 94
rect 1240 -94 1246 94
rect 1215 -100 1246 -94
<< ndiffc >>
rect -1240 -94 -1223 94
rect -1192 -94 -1175 94
rect -1135 -94 -1118 94
rect -1087 -94 -1070 94
rect -1030 -94 -1013 94
rect -982 -94 -965 94
rect -925 -94 -908 94
rect -877 -94 -860 94
rect -820 -94 -803 94
rect -772 -94 -755 94
rect -715 -94 -698 94
rect -667 -94 -650 94
rect -610 -94 -593 94
rect -562 -94 -545 94
rect -505 -94 -488 94
rect -457 -94 -440 94
rect -400 -94 -383 94
rect -352 -94 -335 94
rect -295 -94 -278 94
rect -247 -94 -230 94
rect -190 -94 -173 94
rect -142 -94 -125 94
rect -85 -94 -68 94
rect -37 -94 -20 94
rect 20 -94 37 94
rect 68 -94 85 94
rect 125 -94 142 94
rect 173 -94 190 94
rect 230 -94 247 94
rect 278 -94 295 94
rect 335 -94 352 94
rect 383 -94 400 94
rect 440 -94 457 94
rect 488 -94 505 94
rect 545 -94 562 94
rect 593 -94 610 94
rect 650 -94 667 94
rect 698 -94 715 94
rect 755 -94 772 94
rect 803 -94 820 94
rect 860 -94 877 94
rect 908 -94 925 94
rect 965 -94 982 94
rect 1013 -94 1030 94
rect 1070 -94 1087 94
rect 1118 -94 1135 94
rect 1175 -94 1192 94
rect 1223 -94 1240 94
<< psubdiff >>
rect -1297 170 -1249 187
rect 1249 170 1297 187
rect -1297 139 -1280 170
rect 1280 139 1297 170
rect -1297 -170 -1280 -139
rect 1280 -170 1297 -139
rect -1297 -187 -1249 -170
rect 1249 -187 1297 -170
<< psubdiffcont >>
rect -1249 170 1249 187
rect -1297 -139 -1280 139
rect 1280 -139 1297 139
rect -1249 -187 1249 -170
<< poly >>
rect -1119 136 -1086 144
rect -1119 119 -1111 136
rect -1094 119 -1086 136
rect -1215 100 -1200 113
rect -1119 111 -1086 119
rect -909 136 -876 144
rect -909 119 -901 136
rect -884 119 -876 136
rect -1110 100 -1095 111
rect -1005 100 -990 113
rect -909 111 -876 119
rect -699 136 -666 144
rect -699 119 -691 136
rect -674 119 -666 136
rect -900 100 -885 111
rect -795 100 -780 113
rect -699 111 -666 119
rect -489 136 -456 144
rect -489 119 -481 136
rect -464 119 -456 136
rect -690 100 -675 111
rect -585 100 -570 113
rect -489 111 -456 119
rect -279 136 -246 144
rect -279 119 -271 136
rect -254 119 -246 136
rect -480 100 -465 111
rect -375 100 -360 113
rect -279 111 -246 119
rect -69 136 -36 144
rect -69 119 -61 136
rect -44 119 -36 136
rect -270 100 -255 111
rect -165 100 -150 113
rect -69 111 -36 119
rect 141 136 174 144
rect 141 119 149 136
rect 166 119 174 136
rect -60 100 -45 111
rect 45 100 60 113
rect 141 111 174 119
rect 351 136 384 144
rect 351 119 359 136
rect 376 119 384 136
rect 150 100 165 111
rect 255 100 270 113
rect 351 111 384 119
rect 561 136 594 144
rect 561 119 569 136
rect 586 119 594 136
rect 360 100 375 111
rect 465 100 480 113
rect 561 111 594 119
rect 771 136 804 144
rect 771 119 779 136
rect 796 119 804 136
rect 570 100 585 111
rect 675 100 690 113
rect 771 111 804 119
rect 981 136 1014 144
rect 981 119 989 136
rect 1006 119 1014 136
rect 780 100 795 111
rect 885 100 900 113
rect 981 111 1014 119
rect 1191 136 1224 144
rect 1191 119 1199 136
rect 1216 119 1224 136
rect 990 100 1005 111
rect 1095 100 1110 113
rect 1191 111 1224 119
rect 1200 100 1215 111
rect -1215 -111 -1200 -100
rect -1224 -119 -1191 -111
rect -1110 -113 -1095 -100
rect -1005 -111 -990 -100
rect -1224 -136 -1216 -119
rect -1199 -136 -1191 -119
rect -1224 -144 -1191 -136
rect -1014 -119 -981 -111
rect -900 -113 -885 -100
rect -795 -111 -780 -100
rect -1014 -136 -1006 -119
rect -989 -136 -981 -119
rect -1014 -144 -981 -136
rect -804 -119 -771 -111
rect -690 -113 -675 -100
rect -585 -111 -570 -100
rect -804 -136 -796 -119
rect -779 -136 -771 -119
rect -804 -144 -771 -136
rect -594 -119 -561 -111
rect -480 -113 -465 -100
rect -375 -111 -360 -100
rect -594 -136 -586 -119
rect -569 -136 -561 -119
rect -594 -144 -561 -136
rect -384 -119 -351 -111
rect -270 -113 -255 -100
rect -165 -111 -150 -100
rect -384 -136 -376 -119
rect -359 -136 -351 -119
rect -384 -144 -351 -136
rect -174 -119 -141 -111
rect -60 -113 -45 -100
rect 45 -111 60 -100
rect -174 -136 -166 -119
rect -149 -136 -141 -119
rect -174 -144 -141 -136
rect 36 -119 69 -111
rect 150 -113 165 -100
rect 255 -111 270 -100
rect 36 -136 44 -119
rect 61 -136 69 -119
rect 36 -144 69 -136
rect 246 -119 279 -111
rect 360 -113 375 -100
rect 465 -111 480 -100
rect 246 -136 254 -119
rect 271 -136 279 -119
rect 246 -144 279 -136
rect 456 -119 489 -111
rect 570 -113 585 -100
rect 675 -111 690 -100
rect 456 -136 464 -119
rect 481 -136 489 -119
rect 456 -144 489 -136
rect 666 -119 699 -111
rect 780 -113 795 -100
rect 885 -111 900 -100
rect 666 -136 674 -119
rect 691 -136 699 -119
rect 666 -144 699 -136
rect 876 -119 909 -111
rect 990 -113 1005 -100
rect 1095 -111 1110 -100
rect 876 -136 884 -119
rect 901 -136 909 -119
rect 876 -144 909 -136
rect 1086 -119 1119 -111
rect 1200 -113 1215 -100
rect 1086 -136 1094 -119
rect 1111 -136 1119 -119
rect 1086 -144 1119 -136
<< polycont >>
rect -1111 119 -1094 136
rect -901 119 -884 136
rect -691 119 -674 136
rect -481 119 -464 136
rect -271 119 -254 136
rect -61 119 -44 136
rect 149 119 166 136
rect 359 119 376 136
rect 569 119 586 136
rect 779 119 796 136
rect 989 119 1006 136
rect 1199 119 1216 136
rect -1216 -136 -1199 -119
rect -1006 -136 -989 -119
rect -796 -136 -779 -119
rect -586 -136 -569 -119
rect -376 -136 -359 -119
rect -166 -136 -149 -119
rect 44 -136 61 -119
rect 254 -136 271 -119
rect 464 -136 481 -119
rect 674 -136 691 -119
rect 884 -136 901 -119
rect 1094 -136 1111 -119
<< locali >>
rect -1297 170 -1249 187
rect 1249 170 1297 187
rect -1297 139 -1280 170
rect 1280 139 1297 170
rect -1119 119 -1111 136
rect -1094 119 -1086 136
rect -909 119 -901 136
rect -884 119 -876 136
rect -699 119 -691 136
rect -674 119 -666 136
rect -489 119 -481 136
rect -464 119 -456 136
rect -279 119 -271 136
rect -254 119 -246 136
rect -69 119 -61 136
rect -44 119 -36 136
rect 141 119 149 136
rect 166 119 174 136
rect 351 119 359 136
rect 376 119 384 136
rect 561 119 569 136
rect 586 119 594 136
rect 771 119 779 136
rect 796 119 804 136
rect 981 119 989 136
rect 1006 119 1014 136
rect 1191 119 1199 136
rect 1216 119 1224 136
rect -1240 94 -1223 102
rect -1240 -102 -1223 -94
rect -1192 94 -1175 102
rect -1192 -102 -1175 -94
rect -1135 94 -1118 102
rect -1135 -102 -1118 -94
rect -1087 94 -1070 102
rect -1087 -102 -1070 -94
rect -1030 94 -1013 102
rect -1030 -102 -1013 -94
rect -982 94 -965 102
rect -982 -102 -965 -94
rect -925 94 -908 102
rect -925 -102 -908 -94
rect -877 94 -860 102
rect -877 -102 -860 -94
rect -820 94 -803 102
rect -820 -102 -803 -94
rect -772 94 -755 102
rect -772 -102 -755 -94
rect -715 94 -698 102
rect -715 -102 -698 -94
rect -667 94 -650 102
rect -667 -102 -650 -94
rect -610 94 -593 102
rect -610 -102 -593 -94
rect -562 94 -545 102
rect -562 -102 -545 -94
rect -505 94 -488 102
rect -505 -102 -488 -94
rect -457 94 -440 102
rect -457 -102 -440 -94
rect -400 94 -383 102
rect -400 -102 -383 -94
rect -352 94 -335 102
rect -352 -102 -335 -94
rect -295 94 -278 102
rect -295 -102 -278 -94
rect -247 94 -230 102
rect -247 -102 -230 -94
rect -190 94 -173 102
rect -190 -102 -173 -94
rect -142 94 -125 102
rect -142 -102 -125 -94
rect -85 94 -68 102
rect -85 -102 -68 -94
rect -37 94 -20 102
rect -37 -102 -20 -94
rect 20 94 37 102
rect 20 -102 37 -94
rect 68 94 85 102
rect 68 -102 85 -94
rect 125 94 142 102
rect 125 -102 142 -94
rect 173 94 190 102
rect 173 -102 190 -94
rect 230 94 247 102
rect 230 -102 247 -94
rect 278 94 295 102
rect 278 -102 295 -94
rect 335 94 352 102
rect 335 -102 352 -94
rect 383 94 400 102
rect 383 -102 400 -94
rect 440 94 457 102
rect 440 -102 457 -94
rect 488 94 505 102
rect 488 -102 505 -94
rect 545 94 562 102
rect 545 -102 562 -94
rect 593 94 610 102
rect 593 -102 610 -94
rect 650 94 667 102
rect 650 -102 667 -94
rect 698 94 715 102
rect 698 -102 715 -94
rect 755 94 772 102
rect 755 -102 772 -94
rect 803 94 820 102
rect 803 -102 820 -94
rect 860 94 877 102
rect 860 -102 877 -94
rect 908 94 925 102
rect 908 -102 925 -94
rect 965 94 982 102
rect 965 -102 982 -94
rect 1013 94 1030 102
rect 1013 -102 1030 -94
rect 1070 94 1087 102
rect 1070 -102 1087 -94
rect 1118 94 1135 102
rect 1118 -102 1135 -94
rect 1175 94 1192 102
rect 1175 -102 1192 -94
rect 1223 94 1240 102
rect 1223 -102 1240 -94
rect -1224 -136 -1216 -119
rect -1199 -136 -1191 -119
rect -1014 -136 -1006 -119
rect -989 -136 -981 -119
rect -804 -136 -796 -119
rect -779 -136 -771 -119
rect -594 -136 -586 -119
rect -569 -136 -561 -119
rect -384 -136 -376 -119
rect -359 -136 -351 -119
rect -174 -136 -166 -119
rect -149 -136 -141 -119
rect 36 -136 44 -119
rect 61 -136 69 -119
rect 246 -136 254 -119
rect 271 -136 279 -119
rect 456 -136 464 -119
rect 481 -136 489 -119
rect 666 -136 674 -119
rect 691 -136 699 -119
rect 876 -136 884 -119
rect 901 -136 909 -119
rect 1086 -136 1094 -119
rect 1111 -136 1119 -119
rect -1297 -170 -1280 -139
rect 1280 -170 1297 -139
rect -1297 -187 -1249 -170
rect 1249 -187 1297 -170
<< viali >>
rect -1111 119 -1094 136
rect -901 119 -884 136
rect -691 119 -674 136
rect -481 119 -464 136
rect -271 119 -254 136
rect -61 119 -44 136
rect 149 119 166 136
rect 359 119 376 136
rect 569 119 586 136
rect 779 119 796 136
rect 989 119 1006 136
rect 1199 119 1216 136
rect -1240 -94 -1223 94
rect -1192 -94 -1175 94
rect -1135 -94 -1118 94
rect -1087 -94 -1070 94
rect -1030 -94 -1013 94
rect -982 -94 -965 94
rect -925 -94 -908 94
rect -877 -94 -860 94
rect -820 -94 -803 94
rect -772 -94 -755 94
rect -715 -94 -698 94
rect -667 -94 -650 94
rect -610 -94 -593 94
rect -562 -94 -545 94
rect -505 -94 -488 94
rect -457 -94 -440 94
rect -400 -94 -383 94
rect -352 -94 -335 94
rect -295 -94 -278 94
rect -247 -94 -230 94
rect -190 -94 -173 94
rect -142 -94 -125 94
rect -85 -94 -68 94
rect -37 -94 -20 94
rect 20 -94 37 94
rect 68 -94 85 94
rect 125 -94 142 94
rect 173 -94 190 94
rect 230 -94 247 94
rect 278 -94 295 94
rect 335 -94 352 94
rect 383 -94 400 94
rect 440 -94 457 94
rect 488 -94 505 94
rect 545 -94 562 94
rect 593 -94 610 94
rect 650 -94 667 94
rect 698 -94 715 94
rect 755 -94 772 94
rect 803 -94 820 94
rect 860 -94 877 94
rect 908 -94 925 94
rect 965 -94 982 94
rect 1013 -94 1030 94
rect 1070 -94 1087 94
rect 1118 -94 1135 94
rect 1175 -94 1192 94
rect 1223 -94 1240 94
rect -1216 -136 -1199 -119
rect -1006 -136 -989 -119
rect -796 -136 -779 -119
rect -586 -136 -569 -119
rect -376 -136 -359 -119
rect -166 -136 -149 -119
rect 44 -136 61 -119
rect 254 -136 271 -119
rect 464 -136 481 -119
rect 674 -136 691 -119
rect 884 -136 901 -119
rect 1094 -136 1111 -119
<< metal1 >>
rect -1117 136 -1088 139
rect -1117 119 -1111 136
rect -1094 119 -1088 136
rect -1117 116 -1088 119
rect -907 136 -878 139
rect -907 119 -901 136
rect -884 119 -878 136
rect -907 116 -878 119
rect -697 136 -668 139
rect -697 119 -691 136
rect -674 119 -668 136
rect -697 116 -668 119
rect -487 136 -458 139
rect -487 119 -481 136
rect -464 119 -458 136
rect -487 116 -458 119
rect -277 136 -248 139
rect -277 119 -271 136
rect -254 119 -248 136
rect -277 116 -248 119
rect -67 136 -38 139
rect -67 119 -61 136
rect -44 119 -38 136
rect -67 116 -38 119
rect 143 136 172 139
rect 143 119 149 136
rect 166 119 172 136
rect 143 116 172 119
rect 353 136 382 139
rect 353 119 359 136
rect 376 119 382 136
rect 353 116 382 119
rect 563 136 592 139
rect 563 119 569 136
rect 586 119 592 136
rect 563 116 592 119
rect 773 136 802 139
rect 773 119 779 136
rect 796 119 802 136
rect 773 116 802 119
rect 983 136 1012 139
rect 983 119 989 136
rect 1006 119 1012 136
rect 983 116 1012 119
rect 1193 136 1222 139
rect 1193 119 1199 136
rect 1216 119 1222 136
rect 1193 116 1222 119
rect -1243 94 -1220 100
rect -1243 -94 -1240 94
rect -1223 -94 -1220 94
rect -1243 -100 -1220 -94
rect -1195 94 -1172 100
rect -1195 -94 -1192 94
rect -1175 -94 -1172 94
rect -1195 -100 -1172 -94
rect -1138 94 -1115 100
rect -1138 -94 -1135 94
rect -1118 -94 -1115 94
rect -1138 -100 -1115 -94
rect -1090 94 -1067 100
rect -1090 -94 -1087 94
rect -1070 -94 -1067 94
rect -1090 -100 -1067 -94
rect -1033 94 -1010 100
rect -1033 -94 -1030 94
rect -1013 -94 -1010 94
rect -1033 -100 -1010 -94
rect -985 94 -962 100
rect -985 -94 -982 94
rect -965 -94 -962 94
rect -985 -100 -962 -94
rect -928 94 -905 100
rect -928 -94 -925 94
rect -908 -94 -905 94
rect -928 -100 -905 -94
rect -880 94 -857 100
rect -880 -94 -877 94
rect -860 -94 -857 94
rect -880 -100 -857 -94
rect -823 94 -800 100
rect -823 -94 -820 94
rect -803 -94 -800 94
rect -823 -100 -800 -94
rect -775 94 -752 100
rect -775 -94 -772 94
rect -755 -94 -752 94
rect -775 -100 -752 -94
rect -718 94 -695 100
rect -718 -94 -715 94
rect -698 -94 -695 94
rect -718 -100 -695 -94
rect -670 94 -647 100
rect -670 -94 -667 94
rect -650 -94 -647 94
rect -670 -100 -647 -94
rect -613 94 -590 100
rect -613 -94 -610 94
rect -593 -94 -590 94
rect -613 -100 -590 -94
rect -565 94 -542 100
rect -565 -94 -562 94
rect -545 -94 -542 94
rect -565 -100 -542 -94
rect -508 94 -485 100
rect -508 -94 -505 94
rect -488 -94 -485 94
rect -508 -100 -485 -94
rect -460 94 -437 100
rect -460 -94 -457 94
rect -440 -94 -437 94
rect -460 -100 -437 -94
rect -403 94 -380 100
rect -403 -94 -400 94
rect -383 -94 -380 94
rect -403 -100 -380 -94
rect -355 94 -332 100
rect -355 -94 -352 94
rect -335 -94 -332 94
rect -355 -100 -332 -94
rect -298 94 -275 100
rect -298 -94 -295 94
rect -278 -94 -275 94
rect -298 -100 -275 -94
rect -250 94 -227 100
rect -250 -94 -247 94
rect -230 -94 -227 94
rect -250 -100 -227 -94
rect -193 94 -170 100
rect -193 -94 -190 94
rect -173 -94 -170 94
rect -193 -100 -170 -94
rect -145 94 -122 100
rect -145 -94 -142 94
rect -125 -94 -122 94
rect -145 -100 -122 -94
rect -88 94 -65 100
rect -88 -94 -85 94
rect -68 -94 -65 94
rect -88 -100 -65 -94
rect -40 94 -17 100
rect -40 -94 -37 94
rect -20 -94 -17 94
rect -40 -100 -17 -94
rect 17 94 40 100
rect 17 -94 20 94
rect 37 -94 40 94
rect 17 -100 40 -94
rect 65 94 88 100
rect 65 -94 68 94
rect 85 -94 88 94
rect 65 -100 88 -94
rect 122 94 145 100
rect 122 -94 125 94
rect 142 -94 145 94
rect 122 -100 145 -94
rect 170 94 193 100
rect 170 -94 173 94
rect 190 -94 193 94
rect 170 -100 193 -94
rect 227 94 250 100
rect 227 -94 230 94
rect 247 -94 250 94
rect 227 -100 250 -94
rect 275 94 298 100
rect 275 -94 278 94
rect 295 -94 298 94
rect 275 -100 298 -94
rect 332 94 355 100
rect 332 -94 335 94
rect 352 -94 355 94
rect 332 -100 355 -94
rect 380 94 403 100
rect 380 -94 383 94
rect 400 -94 403 94
rect 380 -100 403 -94
rect 437 94 460 100
rect 437 -94 440 94
rect 457 -94 460 94
rect 437 -100 460 -94
rect 485 94 508 100
rect 485 -94 488 94
rect 505 -94 508 94
rect 485 -100 508 -94
rect 542 94 565 100
rect 542 -94 545 94
rect 562 -94 565 94
rect 542 -100 565 -94
rect 590 94 613 100
rect 590 -94 593 94
rect 610 -94 613 94
rect 590 -100 613 -94
rect 647 94 670 100
rect 647 -94 650 94
rect 667 -94 670 94
rect 647 -100 670 -94
rect 695 94 718 100
rect 695 -94 698 94
rect 715 -94 718 94
rect 695 -100 718 -94
rect 752 94 775 100
rect 752 -94 755 94
rect 772 -94 775 94
rect 752 -100 775 -94
rect 800 94 823 100
rect 800 -94 803 94
rect 820 -94 823 94
rect 800 -100 823 -94
rect 857 94 880 100
rect 857 -94 860 94
rect 877 -94 880 94
rect 857 -100 880 -94
rect 905 94 928 100
rect 905 -94 908 94
rect 925 -94 928 94
rect 905 -100 928 -94
rect 962 94 985 100
rect 962 -94 965 94
rect 982 -94 985 94
rect 962 -100 985 -94
rect 1010 94 1033 100
rect 1010 -94 1013 94
rect 1030 -94 1033 94
rect 1010 -100 1033 -94
rect 1067 94 1090 100
rect 1067 -94 1070 94
rect 1087 -94 1090 94
rect 1067 -100 1090 -94
rect 1115 94 1138 100
rect 1115 -94 1118 94
rect 1135 -94 1138 94
rect 1115 -100 1138 -94
rect 1172 94 1195 100
rect 1172 -94 1175 94
rect 1192 -94 1195 94
rect 1172 -100 1195 -94
rect 1220 94 1243 100
rect 1220 -94 1223 94
rect 1240 -94 1243 94
rect 1220 -100 1243 -94
rect -1222 -119 -1193 -116
rect -1222 -136 -1216 -119
rect -1199 -136 -1193 -119
rect -1222 -139 -1193 -136
rect -1012 -119 -983 -116
rect -1012 -136 -1006 -119
rect -989 -136 -983 -119
rect -1012 -139 -983 -136
rect -802 -119 -773 -116
rect -802 -136 -796 -119
rect -779 -136 -773 -119
rect -802 -139 -773 -136
rect -592 -119 -563 -116
rect -592 -136 -586 -119
rect -569 -136 -563 -119
rect -592 -139 -563 -136
rect -382 -119 -353 -116
rect -382 -136 -376 -119
rect -359 -136 -353 -119
rect -382 -139 -353 -136
rect -172 -119 -143 -116
rect -172 -136 -166 -119
rect -149 -136 -143 -119
rect -172 -139 -143 -136
rect 38 -119 67 -116
rect 38 -136 44 -119
rect 61 -136 67 -119
rect 38 -139 67 -136
rect 248 -119 277 -116
rect 248 -136 254 -119
rect 271 -136 277 -119
rect 248 -139 277 -136
rect 458 -119 487 -116
rect 458 -136 464 -119
rect 481 -136 487 -119
rect 458 -139 487 -136
rect 668 -119 697 -116
rect 668 -136 674 -119
rect 691 -136 697 -119
rect 668 -139 697 -136
rect 878 -119 907 -116
rect 878 -136 884 -119
rect 901 -136 907 -119
rect 878 -139 907 -136
rect 1088 -119 1117 -116
rect 1088 -136 1094 -119
rect 1111 -136 1117 -119
rect 1088 -139 1117 -136
<< properties >>
string FIXED_BBOX -1288 -178 1288 178
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 0.150 m 1 nf 24 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
