magic
tech sky130A
magscale 1 2
timestamp 1671207568
<< error_p >>
rect -383 281 -325 287
rect -265 281 -207 287
rect -147 281 -89 287
rect -29 281 29 287
rect 89 281 147 287
rect 207 281 265 287
rect 325 281 383 287
rect -383 247 -371 281
rect -265 247 -253 281
rect -147 247 -135 281
rect -29 247 -17 281
rect 89 247 101 281
rect 207 247 219 281
rect 325 247 337 281
rect -383 241 -325 247
rect -265 241 -207 247
rect -147 241 -89 247
rect -29 241 29 247
rect 89 241 147 247
rect 207 241 265 247
rect 325 241 383 247
rect -383 -247 -325 -241
rect -265 -247 -207 -241
rect -147 -247 -89 -241
rect -29 -247 29 -241
rect 89 -247 147 -241
rect 207 -247 265 -241
rect 325 -247 383 -241
rect -383 -281 -371 -247
rect -265 -281 -253 -247
rect -147 -281 -135 -247
rect -29 -281 -17 -247
rect 89 -281 101 -247
rect 207 -281 219 -247
rect 325 -281 337 -247
rect -383 -287 -325 -281
rect -265 -287 -207 -281
rect -147 -287 -89 -281
rect -29 -287 29 -281
rect 89 -287 147 -281
rect 207 -287 265 -281
rect 325 -287 383 -281
<< nwell >>
rect -580 -419 580 419
<< pmos >>
rect -384 -200 -324 200
rect -266 -200 -206 200
rect -148 -200 -88 200
rect -30 -200 30 200
rect 88 -200 148 200
rect 206 -200 266 200
rect 324 -200 384 200
<< pdiff >>
rect -442 188 -384 200
rect -442 -188 -430 188
rect -396 -188 -384 188
rect -442 -200 -384 -188
rect -324 188 -266 200
rect -324 -188 -312 188
rect -278 -188 -266 188
rect -324 -200 -266 -188
rect -206 188 -148 200
rect -206 -188 -194 188
rect -160 -188 -148 188
rect -206 -200 -148 -188
rect -88 188 -30 200
rect -88 -188 -76 188
rect -42 -188 -30 188
rect -88 -200 -30 -188
rect 30 188 88 200
rect 30 -188 42 188
rect 76 -188 88 188
rect 30 -200 88 -188
rect 148 188 206 200
rect 148 -188 160 188
rect 194 -188 206 188
rect 148 -200 206 -188
rect 266 188 324 200
rect 266 -188 278 188
rect 312 -188 324 188
rect 266 -200 324 -188
rect 384 188 442 200
rect 384 -188 396 188
rect 430 -188 442 188
rect 384 -200 442 -188
<< pdiffc >>
rect -430 -188 -396 188
rect -312 -188 -278 188
rect -194 -188 -160 188
rect -76 -188 -42 188
rect 42 -188 76 188
rect 160 -188 194 188
rect 278 -188 312 188
rect 396 -188 430 188
<< nsubdiff >>
rect -544 349 -448 383
rect 448 349 544 383
rect -544 287 -510 349
rect 510 287 544 349
rect -544 -349 -510 -287
rect 510 -349 544 -287
rect -544 -383 -448 -349
rect 448 -383 544 -349
<< nsubdiffcont >>
rect -448 349 448 383
rect -544 -287 -510 287
rect 510 -287 544 287
rect -448 -383 448 -349
<< poly >>
rect -387 281 -321 297
rect -387 247 -371 281
rect -337 247 -321 281
rect -387 231 -321 247
rect -269 281 -203 297
rect -269 247 -253 281
rect -219 247 -203 281
rect -269 231 -203 247
rect -151 281 -85 297
rect -151 247 -135 281
rect -101 247 -85 281
rect -151 231 -85 247
rect -33 281 33 297
rect -33 247 -17 281
rect 17 247 33 281
rect -33 231 33 247
rect 85 281 151 297
rect 85 247 101 281
rect 135 247 151 281
rect 85 231 151 247
rect 203 281 269 297
rect 203 247 219 281
rect 253 247 269 281
rect 203 231 269 247
rect 321 281 387 297
rect 321 247 337 281
rect 371 247 387 281
rect 321 231 387 247
rect -384 200 -324 231
rect -266 200 -206 231
rect -148 200 -88 231
rect -30 200 30 231
rect 88 200 148 231
rect 206 200 266 231
rect 324 200 384 231
rect -384 -231 -324 -200
rect -266 -231 -206 -200
rect -148 -231 -88 -200
rect -30 -231 30 -200
rect 88 -231 148 -200
rect 206 -231 266 -200
rect 324 -231 384 -200
rect -387 -247 -321 -231
rect -387 -281 -371 -247
rect -337 -281 -321 -247
rect -387 -297 -321 -281
rect -269 -247 -203 -231
rect -269 -281 -253 -247
rect -219 -281 -203 -247
rect -269 -297 -203 -281
rect -151 -247 -85 -231
rect -151 -281 -135 -247
rect -101 -281 -85 -247
rect -151 -297 -85 -281
rect -33 -247 33 -231
rect -33 -281 -17 -247
rect 17 -281 33 -247
rect -33 -297 33 -281
rect 85 -247 151 -231
rect 85 -281 101 -247
rect 135 -281 151 -247
rect 85 -297 151 -281
rect 203 -247 269 -231
rect 203 -281 219 -247
rect 253 -281 269 -247
rect 203 -297 269 -281
rect 321 -247 387 -231
rect 321 -281 337 -247
rect 371 -281 387 -247
rect 321 -297 387 -281
<< polycont >>
rect -371 247 -337 281
rect -253 247 -219 281
rect -135 247 -101 281
rect -17 247 17 281
rect 101 247 135 281
rect 219 247 253 281
rect 337 247 371 281
rect -371 -281 -337 -247
rect -253 -281 -219 -247
rect -135 -281 -101 -247
rect -17 -281 17 -247
rect 101 -281 135 -247
rect 219 -281 253 -247
rect 337 -281 371 -247
<< locali >>
rect -544 349 -448 383
rect 448 349 544 383
rect -544 287 -510 349
rect 510 287 544 349
rect -387 247 -371 281
rect -337 247 -321 281
rect -269 247 -253 281
rect -219 247 -203 281
rect -151 247 -135 281
rect -101 247 -85 281
rect -33 247 -17 281
rect 17 247 33 281
rect 85 247 101 281
rect 135 247 151 281
rect 203 247 219 281
rect 253 247 269 281
rect 321 247 337 281
rect 371 247 387 281
rect -430 188 -396 204
rect -430 -204 -396 -188
rect -312 188 -278 204
rect -312 -204 -278 -188
rect -194 188 -160 204
rect -194 -204 -160 -188
rect -76 188 -42 204
rect -76 -204 -42 -188
rect 42 188 76 204
rect 42 -204 76 -188
rect 160 188 194 204
rect 160 -204 194 -188
rect 278 188 312 204
rect 278 -204 312 -188
rect 396 188 430 204
rect 396 -204 430 -188
rect -387 -281 -371 -247
rect -337 -281 -321 -247
rect -269 -281 -253 -247
rect -219 -281 -203 -247
rect -151 -281 -135 -247
rect -101 -281 -85 -247
rect -33 -281 -17 -247
rect 17 -281 33 -247
rect 85 -281 101 -247
rect 135 -281 151 -247
rect 203 -281 219 -247
rect 253 -281 269 -247
rect 321 -281 337 -247
rect 371 -281 387 -247
rect -544 -349 -510 -287
rect 510 -349 544 -287
rect -544 -383 -448 -349
rect 448 -383 544 -349
<< viali >>
rect -371 247 -337 281
rect -253 247 -219 281
rect -135 247 -101 281
rect -17 247 17 281
rect 101 247 135 281
rect 219 247 253 281
rect 337 247 371 281
rect -430 -188 -396 188
rect -312 -188 -278 188
rect -194 -188 -160 188
rect -76 -188 -42 188
rect 42 -188 76 188
rect 160 -188 194 188
rect 278 -188 312 188
rect 396 -188 430 188
rect -371 -281 -337 -247
rect -253 -281 -219 -247
rect -135 -281 -101 -247
rect -17 -281 17 -247
rect 101 -281 135 -247
rect 219 -281 253 -247
rect 337 -281 371 -247
<< metal1 >>
rect -383 281 -325 287
rect -383 247 -371 281
rect -337 247 -325 281
rect -383 241 -325 247
rect -265 281 -207 287
rect -265 247 -253 281
rect -219 247 -207 281
rect -265 241 -207 247
rect -147 281 -89 287
rect -147 247 -135 281
rect -101 247 -89 281
rect -147 241 -89 247
rect -29 281 29 287
rect -29 247 -17 281
rect 17 247 29 281
rect -29 241 29 247
rect 89 281 147 287
rect 89 247 101 281
rect 135 247 147 281
rect 89 241 147 247
rect 207 281 265 287
rect 207 247 219 281
rect 253 247 265 281
rect 207 241 265 247
rect 325 281 383 287
rect 325 247 337 281
rect 371 247 383 281
rect 325 241 383 247
rect -436 188 -390 200
rect -436 -188 -430 188
rect -396 -188 -390 188
rect -436 -200 -390 -188
rect -318 188 -272 200
rect -318 -188 -312 188
rect -278 -188 -272 188
rect -318 -200 -272 -188
rect -200 188 -154 200
rect -200 -188 -194 188
rect -160 -188 -154 188
rect -200 -200 -154 -188
rect -82 188 -36 200
rect -82 -188 -76 188
rect -42 -188 -36 188
rect -82 -200 -36 -188
rect 36 188 82 200
rect 36 -188 42 188
rect 76 -188 82 188
rect 36 -200 82 -188
rect 154 188 200 200
rect 154 -188 160 188
rect 194 -188 200 188
rect 154 -200 200 -188
rect 272 188 318 200
rect 272 -188 278 188
rect 312 -188 318 188
rect 272 -200 318 -188
rect 390 188 436 200
rect 390 -188 396 188
rect 430 -188 436 188
rect 390 -200 436 -188
rect -383 -247 -325 -241
rect -383 -281 -371 -247
rect -337 -281 -325 -247
rect -383 -287 -325 -281
rect -265 -247 -207 -241
rect -265 -281 -253 -247
rect -219 -281 -207 -247
rect -265 -287 -207 -281
rect -147 -247 -89 -241
rect -147 -281 -135 -247
rect -101 -281 -89 -247
rect -147 -287 -89 -281
rect -29 -247 29 -241
rect -29 -281 -17 -247
rect 17 -281 29 -247
rect -29 -287 29 -281
rect 89 -247 147 -241
rect 89 -281 101 -247
rect 135 -281 147 -247
rect 89 -287 147 -281
rect 207 -247 265 -241
rect 207 -281 219 -247
rect 253 -281 265 -247
rect 207 -287 265 -281
rect 325 -247 383 -241
rect 325 -281 337 -247
rect 371 -281 383 -247
rect 325 -287 383 -281
<< properties >>
string FIXED_BBOX -527 -366 527 366
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2 l 0.3 m 1 nf 7 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
