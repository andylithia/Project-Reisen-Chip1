magic
tech sky130A
magscale 1 2
timestamp 1671297949
<< error_p >>
rect -676 -1906 -666 -1888
rect -676 -1956 -638 -1938
<< error_s >>
rect 3482 1184 3716 1188
rect -2523 396 -954 440
rect 1405 -206 1406 -205
rect 1406 -207 1407 -206
rect 196 -1748 234 -1730
rect 224 -1798 234 -1780
rect -676 -1878 -638 -1860
rect -676 -1928 -666 -1910
<< error_ps >>
rect -1194 -3780 -1136 -3774
rect -1002 -3780 -944 -3774
rect -810 -3780 -752 -3774
rect -618 -3780 -560 -3774
rect -1194 -3814 -1182 -3780
rect -1002 -3814 -990 -3780
rect -810 -3814 -798 -3780
rect -618 -3814 -606 -3780
rect -1194 -3820 -1136 -3814
rect -1002 -3820 -944 -3814
rect -810 -3820 -752 -3814
rect -618 -3820 -560 -3814
rect -1098 -4090 -1040 -4084
rect -906 -4090 -848 -4084
rect -714 -4090 -656 -4084
rect -522 -4090 -464 -4084
rect -1098 -4124 -1086 -4090
rect -906 -4124 -894 -4090
rect -714 -4124 -702 -4090
rect -522 -4124 -510 -4090
rect -1098 -4130 -1040 -4124
rect -906 -4130 -848 -4124
rect -714 -4130 -656 -4124
rect -522 -4130 -464 -4124
rect -1194 -4450 -1136 -4444
rect -1002 -4450 -944 -4444
rect -810 -4450 -752 -4444
rect -618 -4450 -560 -4444
rect -1194 -4484 -1182 -4450
rect -1002 -4484 -990 -4450
rect -810 -4484 -798 -4450
rect -618 -4484 -606 -4450
rect -1194 -4490 -1136 -4484
rect -1002 -4490 -944 -4484
rect -810 -4490 -752 -4484
rect -618 -4490 -560 -4484
rect -1098 -4978 -1040 -4972
rect -906 -4978 -848 -4972
rect -714 -4978 -656 -4972
rect -522 -4978 -464 -4972
rect -1098 -5012 -1086 -4978
rect -906 -5012 -894 -4978
rect -714 -5012 -702 -4978
rect -522 -5012 -510 -4978
rect -1098 -5018 -1040 -5012
rect -906 -5018 -848 -5012
rect -714 -5018 -656 -5012
rect -522 -5018 -464 -5012
<< metal3 >>
rect -464 1584 4234 2492
rect -464 -426 4242 1584
rect 1160 -5880 4242 -426
<< mimcap >>
rect -232 1188 4008 2332
rect -232 1184 3480 1188
rect 3482 1184 4008 1188
rect -232 -206 1546 1184
rect 1406 -5550 1546 -206
rect 3890 -5550 4008 1184
rect 1406 -5656 4008 -5550
<< mimcapcontact >>
rect 3480 1184 3482 1188
rect 1546 -5550 3890 1184
<< metal4 >>
rect -464 1584 4234 2492
rect -464 1188 4242 1584
rect -464 1184 3480 1188
rect 3482 1184 4242 1188
rect -464 -426 1546 1184
rect 1160 -5550 1546 -426
rect 3890 -5550 4242 1184
rect 1160 -5880 4242 -5550
<< mimcap2 >>
rect -232 1188 4008 2332
rect -232 1184 3480 1188
rect 3482 1184 4008 1188
rect -232 -206 1546 1184
rect 1406 -5550 1546 -206
rect 3890 -5550 4008 1184
rect 1406 -5656 4008 -5550
<< mimcap2contact >>
rect 3480 1184 3482 1188
rect 1546 -5550 3890 1184
<< metal5 >>
rect -464 1584 4234 2492
rect -464 1188 4242 1584
rect -464 1184 3480 1188
rect 3482 1184 4242 1188
rect -464 -426 1546 1184
rect 1160 -5550 1546 -426
rect 3890 -5550 4242 1184
rect 1160 -5880 4242 -5550
use QCS_unit1_flat_dnw  QCS_unit1_flat_dnw_0
timestamp 1668748373
transform 1 0 -4554 0 1 996
box 1520 -680 3680 1480
use cmota_1_flat_1  cmota_1_flat_1_0
timestamp 1671204228
transform 1 0 -7488 0 1 6126
box -164 -3800 5363 2800
use cmota_1_flat_1  cmota_1_flat_1_1
timestamp 1671204228
transform 1 0 -1544 0 1 6126
box -164 -3800 5363 2800
use dnw_test  dnw_test_0
timestamp 1671210538
transform 1 0 -4738 0 -1 -138
box -2940 -620 5635 8540
use sky130_fd_pr__res_xhigh_po_0p35_KL8RQM  sky130_fd_pr__res_xhigh_po_0p35_KL8RQM_0
timestamp 1671210538
transform 1 0 1294 0 -1 1370
box -1778 -934 1778 934
<< end >>
