** sch_path: /home/andylithia/openmpw/Project-Reisen-Chip1/xschem/adc_strongarm_tb.sch
**.subckt adc_strongarm_tb
V1 VDD GND 1.8
.save i(v1)
V2 CKIN GND PULSE(0 1.8 0 0.01n 0.01n 0.5n 1n)
.save i(v2)
V3 net1 GND PULSE(0.8 1.0 0 100n 0 1 2)
.save i(v3)
x3 asclk GND GND VDD VDD net12 sky130_fd_sc_hs__clkbuf_4
R2 net9 net1 0.5k m=1
x8 net5 net4 VDD GND net2 net3 adc_strongarm_latch
x9 VDD net2 net3 net9 net8 net12 GND net6 adc_strongarm
V5 net7 GND 0.9
.save i(v5)
R4 net8 net7 0.5k m=1
x1 net2 net3 gnd gnd vdd vdd asclk sky130_fd_sc_hs__xnor2_2
V7 net10 GND PULSE(0.8 1.0 0 100n 0 1 2)
.save i(v7)
x4 asclk1 GND GND VDD VDD net13 sky130_fd_sc_hs__clkbuf_4
R1 VIP net10 0.5k m=1
x5 VONL VOPL VDD GND VOP VON adc_strongarm_latch
x7 VDD VOP VON VIP VIN net13 GND CKBUF adc_strongarm
V8 net11 GND 0.9
.save i(v8)
R3 VIN net11 0.5k m=1
x12 VOP VON gnd gnd vdd vdd asclk1 sky130_fd_sc_hs__and2_2
**** begin user architecture code

.tran 1p 100n
.save all
.control
run
display
plot CKIN CKBUF
plot VIP VIN
plot VOP VON CKBUF VIP VIN
plot VONL VOPL
.endc


.lib /home/andylithia/openmpw/pdk_1/sky130B/libs.tech/ngspice/sky130.lib.spice tt
.include /home/andylithia/openmpw/pdk_1/sky130B/libs.ref/sky130_fd_sc_hs/spice/sky130_fd_sc_hs.spice

**** end user architecture code
**.ends

* expanding   symbol:  adc_strongarm_latch.sym # of pins=6
** sym_path: /home/andylithia/openmpw/Project-Reisen-Chip1/xschem/adc_strongarm_latch.sym
** sch_path: /home/andylithia/openmpw/Project-Reisen-Chip1/xschem/adc_strongarm_latch.sch
.subckt adc_strongarm_latch VONL VOPL vdd gnd VP VN
*.iopin vdd
*.iopin gnd
*.ipin VP
*.ipin VN
*.opin VOPL
*.opin VONL
XM11 VOPL net1 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM12 VONL net2 gnd gnd sky130_fd_pr__nfet_01v8 L=0.15 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
x6 VOPL gnd gnd vdd vdd VONL sky130_fd_sc_hs__inv_1
x7 VONL gnd gnd vdd vdd VOPL sky130_fd_sc_hs__inv_1
x1 VP gnd gnd vdd vdd net1 sky130_fd_sc_hs__inv_1
x2 VN gnd gnd vdd vdd net2 sky130_fd_sc_hs__inv_1
.ends


* expanding   symbol:  adc_strongarm.sym # of pins=8
** sym_path: /home/andylithia/openmpw/Project-Reisen-Chip1/xschem/adc_strongarm.sym
** sch_path: /home/andylithia/openmpw/Project-Reisen-Chip1/xschem/adc_strongarm.sch
.subckt adc_strongarm vdd vop von vip vin ckin_c16 gnd ckbuf
*.ipin vip
*.ipin vin
*.iopin gnd
*.iopin vdd
*.opin vop
*.opin von
*.iopin ckin_c16
*.opin ckbuf
XM1 net3 vip net1 gnd sky130_fd_pr__nfet_01v8 L=0.15 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2
XM2 net2 vin net1 gnd sky130_fd_pr__nfet_01v8 L=0.15 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2
XM3 net1 ckbuf gnd gnd sky130_fd_pr__nfet_01v8 L=0.15 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2
XM4 vop von net3 gnd sky130_fd_pr__nfet_01v8 L=0.15 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2
XM5 von vop net2 gnd sky130_fd_pr__nfet_01v8 L=0.15 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2
XM6 von vop vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2
XM7 vop von vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2
XM8 vop ckbuf vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2
XM9 von ckbuf vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2
x1 ckbuf gnd gnd vdd vdd net4 sky130_fd_sc_hs__inv_4
XM10 net2 net4 net3 gnd sky130_fd_pr__nfet_01v8 L=0.15 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2
x2 ckin_c16 gnd gnd vdd vdd ckbuf sky130_fd_sc_hs__clkbuf_16
.ends

.GLOBAL GND
.end
