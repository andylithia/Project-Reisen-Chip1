magic
tech sky130A
magscale 1 2
timestamp 1671634351
<< pwell >>
rect 1066 781 2200 860
rect 1066 772 1308 781
rect 1414 772 2200 781
rect 1066 744 2200 772
rect 1066 698 1730 744
rect 1734 698 2200 744
rect 1066 -60 2200 698
<< nmos >>
rect 1682 150 1712 650
rect 1778 150 1808 650
rect 1874 150 1904 650
rect 1970 150 2000 650
<< ndiff >>
rect 1620 638 1682 650
rect 1620 162 1632 638
rect 1666 162 1682 638
rect 1620 150 1682 162
rect 1712 638 1778 650
rect 1712 162 1728 638
rect 1762 162 1778 638
rect 1712 150 1778 162
rect 1808 638 1874 650
rect 1808 162 1824 638
rect 1858 162 1874 638
rect 1808 150 1874 162
rect 1904 638 1970 650
rect 1904 162 1920 638
rect 1954 162 1970 638
rect 1904 150 1970 162
rect 2000 638 2062 650
rect 2000 162 2016 638
rect 2050 162 2062 638
rect 2000 150 2062 162
<< ndiffc >>
rect 1632 162 1666 638
rect 1728 162 1762 638
rect 1824 162 1858 638
rect 1920 162 1954 638
rect 2016 162 2050 638
<< psubdiff >>
rect 1102 790 1218 824
rect 2068 790 2164 824
rect 1102 728 1136 790
rect 2130 728 2164 790
rect 1102 10 1136 72
rect 2130 10 2164 72
rect 1102 -24 1218 10
rect 2068 -24 2164 10
<< psubdiffcont >>
rect 1218 790 2068 824
rect 1102 72 1136 728
rect 2130 72 2164 728
rect 1218 -24 2068 10
<< poly >>
rect 1682 650 1712 676
rect 1778 650 1808 676
rect 1874 650 1904 676
rect 1970 650 2000 676
rect 1682 128 1712 150
rect 1778 128 1808 150
rect 1682 112 1808 128
rect 1682 78 1758 112
rect 1792 78 1808 112
rect 1682 62 1808 78
rect 1874 128 1904 150
rect 1970 128 2000 150
rect 1874 112 2000 128
rect 1874 78 1950 112
rect 1984 78 2000 112
rect 1874 62 2000 78
<< polycont >>
rect 1758 78 1792 112
rect 1950 78 1984 112
<< xpolycontact >>
rect 1278 106 1348 538
rect 1444 106 1514 538
<< xpolyres >>
rect 1278 604 1514 674
rect 1278 538 1348 604
rect 1444 538 1514 604
<< locali >>
rect 1068 960 2028 980
rect 1068 900 1088 960
rect 2008 900 2028 960
rect 1068 858 2028 900
rect 1068 824 2198 858
rect 1068 790 1218 824
rect 2068 790 2198 824
rect 1068 728 1136 790
rect 1068 72 1102 728
rect 1632 638 1666 654
rect 1068 10 1136 72
rect 1278 90 1287 106
rect 1340 90 1348 106
rect 1278 67 1348 90
rect 1632 118 1666 162
rect 1728 638 1762 790
rect 2130 728 2198 790
rect 1728 146 1762 162
rect 1824 638 1858 654
rect 1824 146 1858 162
rect 1920 638 1954 654
rect 1920 146 1954 162
rect 2016 638 2050 654
rect 2016 146 2050 162
rect 1514 106 1666 118
rect 1444 67 1666 106
rect 1742 78 1758 112
rect 1792 78 1808 112
rect 1934 78 1950 112
rect 1984 78 2000 112
rect 2164 72 2198 728
rect 2130 10 2198 72
rect 1068 -24 1218 10
rect 2068 -24 2198 10
rect 1068 -58 2198 -24
<< viali >>
rect 1088 900 2008 960
rect 1287 106 1340 522
rect 1287 90 1340 106
rect 1632 162 1666 638
rect 1728 162 1762 638
rect 1824 162 1858 638
rect 1920 162 1954 638
rect 2016 162 2050 638
rect 1758 78 1792 112
rect 1950 78 1984 112
<< metal1 >>
rect 1068 1100 2028 1120
rect 1068 900 1088 1100
rect 2008 900 2028 1100
rect 1068 880 2028 900
rect 1626 718 2056 758
rect 1626 638 1672 718
rect 1278 522 1348 538
rect 1278 519 1287 522
rect 1340 519 1348 522
rect 1626 162 1632 638
rect 1666 162 1672 638
rect 1626 150 1672 162
rect 1722 638 1768 650
rect 1722 162 1728 638
rect 1762 162 1768 638
rect 1722 150 1768 162
rect 1818 638 1864 718
rect 1818 162 1824 638
rect 1858 162 1864 638
rect 1818 150 1864 162
rect 1911 638 1963 650
rect 1911 635 1920 638
rect 1954 635 1963 638
rect 1911 162 1920 166
rect 1954 162 1963 166
rect 1911 149 1963 162
rect 2010 638 2056 718
rect 2010 162 2016 638
rect 2050 162 2056 638
rect 2010 150 2056 162
rect 1278 67 1348 90
rect 1728 112 1808 118
rect 1728 78 1758 112
rect 1792 78 1808 112
rect 1728 72 1808 78
rect 1920 112 2000 118
rect 1920 78 1950 112
rect 1984 78 2000 112
rect 1920 72 2000 78
rect 1728 33 1762 72
rect 1038 -1 1762 33
rect 1920 -29 1954 72
rect 1039 -63 1954 -29
<< via1 >>
rect 1088 960 2008 1100
rect 1088 900 2008 960
rect 1278 90 1287 519
rect 1287 90 1340 519
rect 1340 90 1348 519
rect 1911 166 1920 635
rect 1920 166 1954 635
rect 1954 166 1963 635
<< metal2 >>
rect 1068 1100 2028 1120
rect 1068 900 1088 1100
rect 2008 900 2028 1100
rect 1068 880 2028 900
rect 1911 635 2199 650
rect 1963 630 2199 635
rect 1278 519 1348 538
rect 1100 100 1278 300
rect 2180 420 2199 630
rect 1963 400 2199 420
rect 1911 149 1963 166
rect 1278 67 1348 90
<< via2 >>
rect 1088 900 2008 1100
rect 1960 420 1963 630
rect 1963 420 2180 630
<< metal3 >>
rect 1068 1180 2028 1200
rect 1068 900 1088 1180
rect 2008 900 2028 1180
rect 1068 880 2028 900
rect 2200 800 7800 1200
rect 1200 700 7800 800
rect 1200 0 1300 700
rect 1700 630 7800 700
rect 1700 420 1960 630
rect 2180 420 7800 630
rect 1700 0 7800 420
rect 1200 -100 7800 0
<< via3 >>
rect 1088 1100 2008 1180
rect 1088 980 2008 1100
rect 1300 0 1700 700
<< mimcap >>
rect 2300 1060 7700 1100
rect 2300 40 2340 1060
rect 7660 40 7700 1060
rect 2300 0 7700 40
<< mimcapcontact >>
rect 2340 40 7660 1060
<< metal4 >>
rect 1068 1180 7800 1200
rect 1068 980 1088 1180
rect 2008 1060 7800 1180
rect 2008 980 2340 1060
rect 1068 960 2340 980
rect 1200 700 1800 800
rect 1200 0 1300 700
rect 1700 0 1800 700
rect 1200 -100 1800 0
rect 2200 40 2340 960
rect 7660 40 7800 1060
rect 2200 -100 7800 40
<< via4 >>
rect 1300 0 1700 700
<< mimcap2 >>
rect 2300 1060 7700 1100
rect 2300 40 2340 1060
rect 7660 40 7700 1060
rect 2300 0 7700 40
<< mimcap2contact >>
rect 2340 40 7660 1060
<< metal5 >>
rect 2200 1060 7800 1200
rect 2200 800 2340 1060
rect 1200 700 2340 800
rect 1200 0 1300 700
rect 1700 40 2340 700
rect 7660 40 7800 1060
rect 1700 0 7800 40
rect 1200 -100 7800 0
<< labels >>
rlabel metal2 1100 100 1158 300 1 IN
rlabel locali 1068 862 1324 880 1 VSUB
rlabel metal5 2070 740 2198 798 1 OUT
rlabel metal1 1040 0 1064 32 1 SBAR
rlabel metal1 1040 -62 1064 -30 1 S
<< end >>
