magic
tech sky130A
magscale 1 2
timestamp 1672206111
<< metal1 >>
rect -1142 -4438 -1078 -4430
rect -1142 -4510 -1078 -4502
rect -3769 -7084 -3729 -6884
rect -3701 -7084 -3661 -6884
<< via1 >>
rect -1142 -4502 -1078 -4438
<< metal2 >>
rect -4930 590 -4750 600
rect -4930 120 -4920 590
rect -4760 120 -4750 590
rect -4930 -2810 -4750 120
rect -2000 0 1400 100
rect -2000 -500 -1900 0
rect 1300 -500 1400 0
rect -2000 -600 1400 -500
rect 1682 -3140 1802 -3134
rect 1680 -3180 1802 -3140
rect 1682 -3186 1802 -3180
rect -1400 -4438 -1078 -4430
rect -1400 -4440 -1142 -4438
rect -1400 -4500 -1390 -4440
rect -1230 -4500 -1142 -4440
rect -1400 -4502 -1142 -4500
rect -1400 -4510 -1078 -4502
rect -2440 -6700 -1600 -5800
rect 1600 -6000 2000 -5800
rect -3600 -7040 -3340 -6900
rect -2820 -7000 -1600 -6700
rect 1200 -7000 2000 -6000
rect -3600 -7084 -3520 -7040
rect -2600 -7100 -1200 -7000
rect -2600 -7700 -2500 -7100
rect -1300 -7700 -1200 -7100
rect -2600 -7800 -1200 -7700
rect 600 -7100 2000 -7000
rect 600 -7700 700 -7100
rect 1900 -7700 2000 -7100
rect 600 -7800 2000 -7700
<< via2 >>
rect -4920 120 -4760 590
rect -1900 -500 1300 0
rect -1390 -4500 -1230 -4440
rect -2500 -7700 -1300 -7100
rect 700 -7700 1900 -7100
<< metal3 >>
rect -4930 590 -4750 600
rect -4930 120 -4920 590
rect -4760 120 -4750 590
rect -4930 110 -4750 120
rect -2000 0 1400 100
rect -7000 -7100 -4200 -200
rect -2000 -500 -1900 0
rect 1300 -500 1400 0
rect -2000 -600 1400 -500
rect -660 -4200 -620 -4180
rect 120 -4200 160 -4180
rect -1400 -4440 -1220 -4430
rect -1400 -4500 -1390 -4440
rect -1230 -4500 -1220 -4440
rect -3200 -5800 -3000 -5600
rect -2600 -5700 -2100 -5500
rect -1400 -5700 -1220 -4500
rect -2400 -6000 -1220 -5700
rect -7000 -7700 -6900 -7100
rect -4300 -7700 -4200 -7100
rect -7000 -7800 -4200 -7700
rect -2600 -7100 -1200 -7000
rect -2600 -7700 -2500 -7100
rect -1300 -7700 -1200 -7100
rect -2600 -7800 -1200 -7700
rect 600 -7100 2000 -7000
rect 600 -7700 700 -7100
rect 1900 -7700 2000 -7100
rect 600 -7800 2000 -7700
<< via3 >>
rect -4920 120 -4760 590
rect -1900 -500 1300 0
rect -6900 -7700 -4300 -7100
rect -2500 -7700 -1300 -7100
rect 700 -7700 1900 -7100
<< mimcap >>
rect -6900 -340 -4300 -300
rect -6900 -6460 -6860 -340
rect -4340 -6460 -4300 -340
rect -6900 -6500 -4300 -6460
<< mimcapcontact >>
rect -6860 -6460 -4340 -340
<< metal4 >>
rect -6800 590 1400 600
rect -6800 120 -4920 590
rect -4760 120 1400 590
rect -6800 100 1400 120
rect -6800 -200 -4400 100
rect -2000 0 1400 100
rect -7000 -340 -4200 -200
rect -7000 -6460 -6860 -340
rect -4340 -6460 -4200 -340
rect -2000 -500 -1900 0
rect 1300 -500 1400 0
rect -2000 -600 1400 -500
rect -7000 -6600 -4200 -6460
rect -2740 -7000 -2501 -6832
rect -7000 -7100 -4200 -7000
rect -7000 -7700 -6900 -7100
rect -4300 -7300 -4200 -7100
rect -2740 -7100 2000 -7000
rect -2740 -7300 -2500 -7100
rect -4300 -7700 -2500 -7300
rect -1300 -7700 700 -7100
rect 1900 -7700 2000 -7100
rect -7000 -7800 2000 -7700
<< via4 >>
rect -6900 -7700 -4300 -7100
<< mimcap2 >>
rect -6900 -340 -4300 -300
rect -6900 -6460 -6860 -340
rect -4340 -6460 -4300 -340
rect -6900 -6500 -4300 -6460
<< mimcap2contact >>
rect -6860 -6460 -4340 -340
<< metal5 >>
rect -7000 -340 -4200 -200
rect -7000 -6460 -6860 -340
rect -4340 -6460 -4200 -340
rect -7000 -7100 -4200 -6460
rect -7000 -7700 -6900 -7100
rect -4300 -7700 -4200 -7100
rect -7000 -7800 -4200 -7700
use cmota_gb_rp  cmota_gb_rp_0
timestamp 1671672231
transform 1 0 -2798 0 1 -3200
box 308 -3800 5600 2800
use gated_iref_fix  gated_iref_fix_0
timestamp 1672205966
transform 0 1 -3700 1 0 -7948
box 940 -2420 7820 1220
<< labels >>
rlabel metal3 -660 -4200 -620 -4180 1 VIN
rlabel metal3 120 -4200 160 -4180 1 VIP
rlabel metal4 -3820 320 -3440 600 1 VHI
rlabel metal4 -3440 -7800 -3260 -7300 1 VLO
rlabel metal1 -3701 -7084 -3661 -7044 1 SBAR
rlabel metal1 -3769 -7084 -3729 -7044 1 S
rlabel metal2 -3600 -7084 -3520 -7004 1 VREF
rlabel space 1309 -3186 1682 -3134 1 VOP
rlabel metal3 -2080 -5780 -2020 -5720 1 VREF_GATED
rlabel metal2 1682 -3186 1802 -3134 1 VOP
<< end >>
