magic
tech sky130A
magscale 1 2
timestamp 1671152619
<< error_p >>
rect -1150 2081 -1092 2087
rect -1032 2081 -974 2087
rect -914 2081 -856 2087
rect -796 2081 -738 2087
rect -678 2081 -620 2087
rect -560 2081 -502 2087
rect -442 2081 -384 2087
rect -324 2081 -266 2087
rect -206 2081 -148 2087
rect -88 2081 -30 2087
rect 30 2081 88 2087
rect 148 2081 206 2087
rect 266 2081 324 2087
rect 384 2081 442 2087
rect 502 2081 560 2087
rect 620 2081 678 2087
rect 738 2081 796 2087
rect 856 2081 914 2087
rect 974 2081 1032 2087
rect 1092 2081 1150 2087
rect -1150 2047 -1138 2081
rect -1032 2047 -1020 2081
rect -914 2047 -902 2081
rect -796 2047 -784 2081
rect -678 2047 -666 2081
rect -560 2047 -548 2081
rect -442 2047 -430 2081
rect -324 2047 -312 2081
rect -206 2047 -194 2081
rect -88 2047 -76 2081
rect 30 2047 42 2081
rect 148 2047 160 2081
rect 266 2047 278 2081
rect 384 2047 396 2081
rect 502 2047 514 2081
rect 620 2047 632 2081
rect 738 2047 750 2081
rect 856 2047 868 2081
rect 974 2047 986 2081
rect 1092 2047 1104 2081
rect -1150 2041 -1092 2047
rect -1032 2041 -974 2047
rect -914 2041 -856 2047
rect -796 2041 -738 2047
rect -678 2041 -620 2047
rect -560 2041 -502 2047
rect -442 2041 -384 2047
rect -324 2041 -266 2047
rect -206 2041 -148 2047
rect -88 2041 -30 2047
rect 30 2041 88 2047
rect 148 2041 206 2047
rect 266 2041 324 2047
rect 384 2041 442 2047
rect 502 2041 560 2047
rect 620 2041 678 2047
rect 738 2041 796 2047
rect 856 2041 914 2047
rect 974 2041 1032 2047
rect 1092 2041 1150 2047
rect -1150 -2047 -1092 -2041
rect -1032 -2047 -974 -2041
rect -914 -2047 -856 -2041
rect -796 -2047 -738 -2041
rect -678 -2047 -620 -2041
rect -560 -2047 -502 -2041
rect -442 -2047 -384 -2041
rect -324 -2047 -266 -2041
rect -206 -2047 -148 -2041
rect -88 -2047 -30 -2041
rect 30 -2047 88 -2041
rect 148 -2047 206 -2041
rect 266 -2047 324 -2041
rect 384 -2047 442 -2041
rect 502 -2047 560 -2041
rect 620 -2047 678 -2041
rect 738 -2047 796 -2041
rect 856 -2047 914 -2041
rect 974 -2047 1032 -2041
rect 1092 -2047 1150 -2041
rect -1150 -2081 -1138 -2047
rect -1032 -2081 -1020 -2047
rect -914 -2081 -902 -2047
rect -796 -2081 -784 -2047
rect -678 -2081 -666 -2047
rect -560 -2081 -548 -2047
rect -442 -2081 -430 -2047
rect -324 -2081 -312 -2047
rect -206 -2081 -194 -2047
rect -88 -2081 -76 -2047
rect 30 -2081 42 -2047
rect 148 -2081 160 -2047
rect 266 -2081 278 -2047
rect 384 -2081 396 -2047
rect 502 -2081 514 -2047
rect 620 -2081 632 -2047
rect 738 -2081 750 -2047
rect 856 -2081 868 -2047
rect 974 -2081 986 -2047
rect 1092 -2081 1104 -2047
rect -1150 -2087 -1092 -2081
rect -1032 -2087 -974 -2081
rect -914 -2087 -856 -2081
rect -796 -2087 -738 -2081
rect -678 -2087 -620 -2081
rect -560 -2087 -502 -2081
rect -442 -2087 -384 -2081
rect -324 -2087 -266 -2081
rect -206 -2087 -148 -2081
rect -88 -2087 -30 -2081
rect 30 -2087 88 -2081
rect 148 -2087 206 -2081
rect 266 -2087 324 -2081
rect 384 -2087 442 -2081
rect 502 -2087 560 -2081
rect 620 -2087 678 -2081
rect 738 -2087 796 -2081
rect 856 -2087 914 -2081
rect 974 -2087 1032 -2081
rect 1092 -2087 1150 -2081
<< nwell >>
rect -1347 -2219 1347 2219
<< pmos >>
rect -1151 -2000 -1091 2000
rect -1033 -2000 -973 2000
rect -915 -2000 -855 2000
rect -797 -2000 -737 2000
rect -679 -2000 -619 2000
rect -561 -2000 -501 2000
rect -443 -2000 -383 2000
rect -325 -2000 -265 2000
rect -207 -2000 -147 2000
rect -89 -2000 -29 2000
rect 29 -2000 89 2000
rect 147 -2000 207 2000
rect 265 -2000 325 2000
rect 383 -2000 443 2000
rect 501 -2000 561 2000
rect 619 -2000 679 2000
rect 737 -2000 797 2000
rect 855 -2000 915 2000
rect 973 -2000 1033 2000
rect 1091 -2000 1151 2000
<< pdiff >>
rect -1209 1988 -1151 2000
rect -1209 -1988 -1197 1988
rect -1163 -1988 -1151 1988
rect -1209 -2000 -1151 -1988
rect -1091 1988 -1033 2000
rect -1091 -1988 -1079 1988
rect -1045 -1988 -1033 1988
rect -1091 -2000 -1033 -1988
rect -973 1988 -915 2000
rect -973 -1988 -961 1988
rect -927 -1988 -915 1988
rect -973 -2000 -915 -1988
rect -855 1988 -797 2000
rect -855 -1988 -843 1988
rect -809 -1988 -797 1988
rect -855 -2000 -797 -1988
rect -737 1988 -679 2000
rect -737 -1988 -725 1988
rect -691 -1988 -679 1988
rect -737 -2000 -679 -1988
rect -619 1988 -561 2000
rect -619 -1988 -607 1988
rect -573 -1988 -561 1988
rect -619 -2000 -561 -1988
rect -501 1988 -443 2000
rect -501 -1988 -489 1988
rect -455 -1988 -443 1988
rect -501 -2000 -443 -1988
rect -383 1988 -325 2000
rect -383 -1988 -371 1988
rect -337 -1988 -325 1988
rect -383 -2000 -325 -1988
rect -265 1988 -207 2000
rect -265 -1988 -253 1988
rect -219 -1988 -207 1988
rect -265 -2000 -207 -1988
rect -147 1988 -89 2000
rect -147 -1988 -135 1988
rect -101 -1988 -89 1988
rect -147 -2000 -89 -1988
rect -29 1988 29 2000
rect -29 -1988 -17 1988
rect 17 -1988 29 1988
rect -29 -2000 29 -1988
rect 89 1988 147 2000
rect 89 -1988 101 1988
rect 135 -1988 147 1988
rect 89 -2000 147 -1988
rect 207 1988 265 2000
rect 207 -1988 219 1988
rect 253 -1988 265 1988
rect 207 -2000 265 -1988
rect 325 1988 383 2000
rect 325 -1988 337 1988
rect 371 -1988 383 1988
rect 325 -2000 383 -1988
rect 443 1988 501 2000
rect 443 -1988 455 1988
rect 489 -1988 501 1988
rect 443 -2000 501 -1988
rect 561 1988 619 2000
rect 561 -1988 573 1988
rect 607 -1988 619 1988
rect 561 -2000 619 -1988
rect 679 1988 737 2000
rect 679 -1988 691 1988
rect 725 -1988 737 1988
rect 679 -2000 737 -1988
rect 797 1988 855 2000
rect 797 -1988 809 1988
rect 843 -1988 855 1988
rect 797 -2000 855 -1988
rect 915 1988 973 2000
rect 915 -1988 927 1988
rect 961 -1988 973 1988
rect 915 -2000 973 -1988
rect 1033 1988 1091 2000
rect 1033 -1988 1045 1988
rect 1079 -1988 1091 1988
rect 1033 -2000 1091 -1988
rect 1151 1988 1209 2000
rect 1151 -1988 1163 1988
rect 1197 -1988 1209 1988
rect 1151 -2000 1209 -1988
<< pdiffc >>
rect -1197 -1988 -1163 1988
rect -1079 -1988 -1045 1988
rect -961 -1988 -927 1988
rect -843 -1988 -809 1988
rect -725 -1988 -691 1988
rect -607 -1988 -573 1988
rect -489 -1988 -455 1988
rect -371 -1988 -337 1988
rect -253 -1988 -219 1988
rect -135 -1988 -101 1988
rect -17 -1988 17 1988
rect 101 -1988 135 1988
rect 219 -1988 253 1988
rect 337 -1988 371 1988
rect 455 -1988 489 1988
rect 573 -1988 607 1988
rect 691 -1988 725 1988
rect 809 -1988 843 1988
rect 927 -1988 961 1988
rect 1045 -1988 1079 1988
rect 1163 -1988 1197 1988
<< nsubdiff >>
rect -1311 2149 -1215 2183
rect 1215 2149 1311 2183
rect -1311 2087 -1277 2149
rect 1277 2087 1311 2149
rect -1311 -2149 -1277 -2087
rect 1277 -2149 1311 -2087
rect -1311 -2183 -1215 -2149
rect 1215 -2183 1311 -2149
<< nsubdiffcont >>
rect -1215 2149 1215 2183
rect -1311 -2087 -1277 2087
rect 1277 -2087 1311 2087
rect -1215 -2183 1215 -2149
<< poly >>
rect -1154 2081 -1088 2097
rect -1154 2047 -1138 2081
rect -1104 2047 -1088 2081
rect -1154 2031 -1088 2047
rect -1036 2081 -970 2097
rect -1036 2047 -1020 2081
rect -986 2047 -970 2081
rect -1036 2031 -970 2047
rect -918 2081 -852 2097
rect -918 2047 -902 2081
rect -868 2047 -852 2081
rect -918 2031 -852 2047
rect -800 2081 -734 2097
rect -800 2047 -784 2081
rect -750 2047 -734 2081
rect -800 2031 -734 2047
rect -682 2081 -616 2097
rect -682 2047 -666 2081
rect -632 2047 -616 2081
rect -682 2031 -616 2047
rect -564 2081 -498 2097
rect -564 2047 -548 2081
rect -514 2047 -498 2081
rect -564 2031 -498 2047
rect -446 2081 -380 2097
rect -446 2047 -430 2081
rect -396 2047 -380 2081
rect -446 2031 -380 2047
rect -328 2081 -262 2097
rect -328 2047 -312 2081
rect -278 2047 -262 2081
rect -328 2031 -262 2047
rect -210 2081 -144 2097
rect -210 2047 -194 2081
rect -160 2047 -144 2081
rect -210 2031 -144 2047
rect -92 2081 -26 2097
rect -92 2047 -76 2081
rect -42 2047 -26 2081
rect -92 2031 -26 2047
rect 26 2081 92 2097
rect 26 2047 42 2081
rect 76 2047 92 2081
rect 26 2031 92 2047
rect 144 2081 210 2097
rect 144 2047 160 2081
rect 194 2047 210 2081
rect 144 2031 210 2047
rect 262 2081 328 2097
rect 262 2047 278 2081
rect 312 2047 328 2081
rect 262 2031 328 2047
rect 380 2081 446 2097
rect 380 2047 396 2081
rect 430 2047 446 2081
rect 380 2031 446 2047
rect 498 2081 564 2097
rect 498 2047 514 2081
rect 548 2047 564 2081
rect 498 2031 564 2047
rect 616 2081 682 2097
rect 616 2047 632 2081
rect 666 2047 682 2081
rect 616 2031 682 2047
rect 734 2081 800 2097
rect 734 2047 750 2081
rect 784 2047 800 2081
rect 734 2031 800 2047
rect 852 2081 918 2097
rect 852 2047 868 2081
rect 902 2047 918 2081
rect 852 2031 918 2047
rect 970 2081 1036 2097
rect 970 2047 986 2081
rect 1020 2047 1036 2081
rect 970 2031 1036 2047
rect 1088 2081 1154 2097
rect 1088 2047 1104 2081
rect 1138 2047 1154 2081
rect 1088 2031 1154 2047
rect -1151 2000 -1091 2031
rect -1033 2000 -973 2031
rect -915 2000 -855 2031
rect -797 2000 -737 2031
rect -679 2000 -619 2031
rect -561 2000 -501 2031
rect -443 2000 -383 2031
rect -325 2000 -265 2031
rect -207 2000 -147 2031
rect -89 2000 -29 2031
rect 29 2000 89 2031
rect 147 2000 207 2031
rect 265 2000 325 2031
rect 383 2000 443 2031
rect 501 2000 561 2031
rect 619 2000 679 2031
rect 737 2000 797 2031
rect 855 2000 915 2031
rect 973 2000 1033 2031
rect 1091 2000 1151 2031
rect -1151 -2031 -1091 -2000
rect -1033 -2031 -973 -2000
rect -915 -2031 -855 -2000
rect -797 -2031 -737 -2000
rect -679 -2031 -619 -2000
rect -561 -2031 -501 -2000
rect -443 -2031 -383 -2000
rect -325 -2031 -265 -2000
rect -207 -2031 -147 -2000
rect -89 -2031 -29 -2000
rect 29 -2031 89 -2000
rect 147 -2031 207 -2000
rect 265 -2031 325 -2000
rect 383 -2031 443 -2000
rect 501 -2031 561 -2000
rect 619 -2031 679 -2000
rect 737 -2031 797 -2000
rect 855 -2031 915 -2000
rect 973 -2031 1033 -2000
rect 1091 -2031 1151 -2000
rect -1154 -2047 -1088 -2031
rect -1154 -2081 -1138 -2047
rect -1104 -2081 -1088 -2047
rect -1154 -2097 -1088 -2081
rect -1036 -2047 -970 -2031
rect -1036 -2081 -1020 -2047
rect -986 -2081 -970 -2047
rect -1036 -2097 -970 -2081
rect -918 -2047 -852 -2031
rect -918 -2081 -902 -2047
rect -868 -2081 -852 -2047
rect -918 -2097 -852 -2081
rect -800 -2047 -734 -2031
rect -800 -2081 -784 -2047
rect -750 -2081 -734 -2047
rect -800 -2097 -734 -2081
rect -682 -2047 -616 -2031
rect -682 -2081 -666 -2047
rect -632 -2081 -616 -2047
rect -682 -2097 -616 -2081
rect -564 -2047 -498 -2031
rect -564 -2081 -548 -2047
rect -514 -2081 -498 -2047
rect -564 -2097 -498 -2081
rect -446 -2047 -380 -2031
rect -446 -2081 -430 -2047
rect -396 -2081 -380 -2047
rect -446 -2097 -380 -2081
rect -328 -2047 -262 -2031
rect -328 -2081 -312 -2047
rect -278 -2081 -262 -2047
rect -328 -2097 -262 -2081
rect -210 -2047 -144 -2031
rect -210 -2081 -194 -2047
rect -160 -2081 -144 -2047
rect -210 -2097 -144 -2081
rect -92 -2047 -26 -2031
rect -92 -2081 -76 -2047
rect -42 -2081 -26 -2047
rect -92 -2097 -26 -2081
rect 26 -2047 92 -2031
rect 26 -2081 42 -2047
rect 76 -2081 92 -2047
rect 26 -2097 92 -2081
rect 144 -2047 210 -2031
rect 144 -2081 160 -2047
rect 194 -2081 210 -2047
rect 144 -2097 210 -2081
rect 262 -2047 328 -2031
rect 262 -2081 278 -2047
rect 312 -2081 328 -2047
rect 262 -2097 328 -2081
rect 380 -2047 446 -2031
rect 380 -2081 396 -2047
rect 430 -2081 446 -2047
rect 380 -2097 446 -2081
rect 498 -2047 564 -2031
rect 498 -2081 514 -2047
rect 548 -2081 564 -2047
rect 498 -2097 564 -2081
rect 616 -2047 682 -2031
rect 616 -2081 632 -2047
rect 666 -2081 682 -2047
rect 616 -2097 682 -2081
rect 734 -2047 800 -2031
rect 734 -2081 750 -2047
rect 784 -2081 800 -2047
rect 734 -2097 800 -2081
rect 852 -2047 918 -2031
rect 852 -2081 868 -2047
rect 902 -2081 918 -2047
rect 852 -2097 918 -2081
rect 970 -2047 1036 -2031
rect 970 -2081 986 -2047
rect 1020 -2081 1036 -2047
rect 970 -2097 1036 -2081
rect 1088 -2047 1154 -2031
rect 1088 -2081 1104 -2047
rect 1138 -2081 1154 -2047
rect 1088 -2097 1154 -2081
<< polycont >>
rect -1138 2047 -1104 2081
rect -1020 2047 -986 2081
rect -902 2047 -868 2081
rect -784 2047 -750 2081
rect -666 2047 -632 2081
rect -548 2047 -514 2081
rect -430 2047 -396 2081
rect -312 2047 -278 2081
rect -194 2047 -160 2081
rect -76 2047 -42 2081
rect 42 2047 76 2081
rect 160 2047 194 2081
rect 278 2047 312 2081
rect 396 2047 430 2081
rect 514 2047 548 2081
rect 632 2047 666 2081
rect 750 2047 784 2081
rect 868 2047 902 2081
rect 986 2047 1020 2081
rect 1104 2047 1138 2081
rect -1138 -2081 -1104 -2047
rect -1020 -2081 -986 -2047
rect -902 -2081 -868 -2047
rect -784 -2081 -750 -2047
rect -666 -2081 -632 -2047
rect -548 -2081 -514 -2047
rect -430 -2081 -396 -2047
rect -312 -2081 -278 -2047
rect -194 -2081 -160 -2047
rect -76 -2081 -42 -2047
rect 42 -2081 76 -2047
rect 160 -2081 194 -2047
rect 278 -2081 312 -2047
rect 396 -2081 430 -2047
rect 514 -2081 548 -2047
rect 632 -2081 666 -2047
rect 750 -2081 784 -2047
rect 868 -2081 902 -2047
rect 986 -2081 1020 -2047
rect 1104 -2081 1138 -2047
<< locali >>
rect -1311 2149 -1215 2183
rect 1215 2149 1311 2183
rect -1311 2087 -1277 2149
rect 1277 2087 1311 2149
rect -1154 2047 -1138 2081
rect -1104 2047 -1088 2081
rect -1036 2047 -1020 2081
rect -986 2047 -970 2081
rect -918 2047 -902 2081
rect -868 2047 -852 2081
rect -800 2047 -784 2081
rect -750 2047 -734 2081
rect -682 2047 -666 2081
rect -632 2047 -616 2081
rect -564 2047 -548 2081
rect -514 2047 -498 2081
rect -446 2047 -430 2081
rect -396 2047 -380 2081
rect -328 2047 -312 2081
rect -278 2047 -262 2081
rect -210 2047 -194 2081
rect -160 2047 -144 2081
rect -92 2047 -76 2081
rect -42 2047 -26 2081
rect 26 2047 42 2081
rect 76 2047 92 2081
rect 144 2047 160 2081
rect 194 2047 210 2081
rect 262 2047 278 2081
rect 312 2047 328 2081
rect 380 2047 396 2081
rect 430 2047 446 2081
rect 498 2047 514 2081
rect 548 2047 564 2081
rect 616 2047 632 2081
rect 666 2047 682 2081
rect 734 2047 750 2081
rect 784 2047 800 2081
rect 852 2047 868 2081
rect 902 2047 918 2081
rect 970 2047 986 2081
rect 1020 2047 1036 2081
rect 1088 2047 1104 2081
rect 1138 2047 1154 2081
rect -1197 1988 -1163 2004
rect -1197 -2004 -1163 -1988
rect -1079 1988 -1045 2004
rect -1079 -2004 -1045 -1988
rect -961 1988 -927 2004
rect -961 -2004 -927 -1988
rect -843 1988 -809 2004
rect -843 -2004 -809 -1988
rect -725 1988 -691 2004
rect -725 -2004 -691 -1988
rect -607 1988 -573 2004
rect -607 -2004 -573 -1988
rect -489 1988 -455 2004
rect -489 -2004 -455 -1988
rect -371 1988 -337 2004
rect -371 -2004 -337 -1988
rect -253 1988 -219 2004
rect -253 -2004 -219 -1988
rect -135 1988 -101 2004
rect -135 -2004 -101 -1988
rect -17 1988 17 2004
rect -17 -2004 17 -1988
rect 101 1988 135 2004
rect 101 -2004 135 -1988
rect 219 1988 253 2004
rect 219 -2004 253 -1988
rect 337 1988 371 2004
rect 337 -2004 371 -1988
rect 455 1988 489 2004
rect 455 -2004 489 -1988
rect 573 1988 607 2004
rect 573 -2004 607 -1988
rect 691 1988 725 2004
rect 691 -2004 725 -1988
rect 809 1988 843 2004
rect 809 -2004 843 -1988
rect 927 1988 961 2004
rect 927 -2004 961 -1988
rect 1045 1988 1079 2004
rect 1045 -2004 1079 -1988
rect 1163 1988 1197 2004
rect 1163 -2004 1197 -1988
rect -1154 -2081 -1138 -2047
rect -1104 -2081 -1088 -2047
rect -1036 -2081 -1020 -2047
rect -986 -2081 -970 -2047
rect -918 -2081 -902 -2047
rect -868 -2081 -852 -2047
rect -800 -2081 -784 -2047
rect -750 -2081 -734 -2047
rect -682 -2081 -666 -2047
rect -632 -2081 -616 -2047
rect -564 -2081 -548 -2047
rect -514 -2081 -498 -2047
rect -446 -2081 -430 -2047
rect -396 -2081 -380 -2047
rect -328 -2081 -312 -2047
rect -278 -2081 -262 -2047
rect -210 -2081 -194 -2047
rect -160 -2081 -144 -2047
rect -92 -2081 -76 -2047
rect -42 -2081 -26 -2047
rect 26 -2081 42 -2047
rect 76 -2081 92 -2047
rect 144 -2081 160 -2047
rect 194 -2081 210 -2047
rect 262 -2081 278 -2047
rect 312 -2081 328 -2047
rect 380 -2081 396 -2047
rect 430 -2081 446 -2047
rect 498 -2081 514 -2047
rect 548 -2081 564 -2047
rect 616 -2081 632 -2047
rect 666 -2081 682 -2047
rect 734 -2081 750 -2047
rect 784 -2081 800 -2047
rect 852 -2081 868 -2047
rect 902 -2081 918 -2047
rect 970 -2081 986 -2047
rect 1020 -2081 1036 -2047
rect 1088 -2081 1104 -2047
rect 1138 -2081 1154 -2047
rect -1311 -2149 -1277 -2087
rect 1277 -2149 1311 -2087
rect -1311 -2183 -1215 -2149
rect 1215 -2183 1311 -2149
<< viali >>
rect -1138 2047 -1104 2081
rect -1020 2047 -986 2081
rect -902 2047 -868 2081
rect -784 2047 -750 2081
rect -666 2047 -632 2081
rect -548 2047 -514 2081
rect -430 2047 -396 2081
rect -312 2047 -278 2081
rect -194 2047 -160 2081
rect -76 2047 -42 2081
rect 42 2047 76 2081
rect 160 2047 194 2081
rect 278 2047 312 2081
rect 396 2047 430 2081
rect 514 2047 548 2081
rect 632 2047 666 2081
rect 750 2047 784 2081
rect 868 2047 902 2081
rect 986 2047 1020 2081
rect 1104 2047 1138 2081
rect -1197 -1988 -1163 1988
rect -1079 -1988 -1045 1988
rect -961 -1988 -927 1988
rect -843 -1988 -809 1988
rect -725 -1988 -691 1988
rect -607 -1988 -573 1988
rect -489 -1988 -455 1988
rect -371 -1988 -337 1988
rect -253 -1988 -219 1988
rect -135 -1988 -101 1988
rect -17 -1988 17 1988
rect 101 -1988 135 1988
rect 219 -1988 253 1988
rect 337 -1988 371 1988
rect 455 -1988 489 1988
rect 573 -1988 607 1988
rect 691 -1988 725 1988
rect 809 -1988 843 1988
rect 927 -1988 961 1988
rect 1045 -1988 1079 1988
rect 1163 -1988 1197 1988
rect -1138 -2081 -1104 -2047
rect -1020 -2081 -986 -2047
rect -902 -2081 -868 -2047
rect -784 -2081 -750 -2047
rect -666 -2081 -632 -2047
rect -548 -2081 -514 -2047
rect -430 -2081 -396 -2047
rect -312 -2081 -278 -2047
rect -194 -2081 -160 -2047
rect -76 -2081 -42 -2047
rect 42 -2081 76 -2047
rect 160 -2081 194 -2047
rect 278 -2081 312 -2047
rect 396 -2081 430 -2047
rect 514 -2081 548 -2047
rect 632 -2081 666 -2047
rect 750 -2081 784 -2047
rect 868 -2081 902 -2047
rect 986 -2081 1020 -2047
rect 1104 -2081 1138 -2047
<< metal1 >>
rect -1150 2081 -1092 2087
rect -1150 2047 -1138 2081
rect -1104 2047 -1092 2081
rect -1150 2041 -1092 2047
rect -1032 2081 -974 2087
rect -1032 2047 -1020 2081
rect -986 2047 -974 2081
rect -1032 2041 -974 2047
rect -914 2081 -856 2087
rect -914 2047 -902 2081
rect -868 2047 -856 2081
rect -914 2041 -856 2047
rect -796 2081 -738 2087
rect -796 2047 -784 2081
rect -750 2047 -738 2081
rect -796 2041 -738 2047
rect -678 2081 -620 2087
rect -678 2047 -666 2081
rect -632 2047 -620 2081
rect -678 2041 -620 2047
rect -560 2081 -502 2087
rect -560 2047 -548 2081
rect -514 2047 -502 2081
rect -560 2041 -502 2047
rect -442 2081 -384 2087
rect -442 2047 -430 2081
rect -396 2047 -384 2081
rect -442 2041 -384 2047
rect -324 2081 -266 2087
rect -324 2047 -312 2081
rect -278 2047 -266 2081
rect -324 2041 -266 2047
rect -206 2081 -148 2087
rect -206 2047 -194 2081
rect -160 2047 -148 2081
rect -206 2041 -148 2047
rect -88 2081 -30 2087
rect -88 2047 -76 2081
rect -42 2047 -30 2081
rect -88 2041 -30 2047
rect 30 2081 88 2087
rect 30 2047 42 2081
rect 76 2047 88 2081
rect 30 2041 88 2047
rect 148 2081 206 2087
rect 148 2047 160 2081
rect 194 2047 206 2081
rect 148 2041 206 2047
rect 266 2081 324 2087
rect 266 2047 278 2081
rect 312 2047 324 2081
rect 266 2041 324 2047
rect 384 2081 442 2087
rect 384 2047 396 2081
rect 430 2047 442 2081
rect 384 2041 442 2047
rect 502 2081 560 2087
rect 502 2047 514 2081
rect 548 2047 560 2081
rect 502 2041 560 2047
rect 620 2081 678 2087
rect 620 2047 632 2081
rect 666 2047 678 2081
rect 620 2041 678 2047
rect 738 2081 796 2087
rect 738 2047 750 2081
rect 784 2047 796 2081
rect 738 2041 796 2047
rect 856 2081 914 2087
rect 856 2047 868 2081
rect 902 2047 914 2081
rect 856 2041 914 2047
rect 974 2081 1032 2087
rect 974 2047 986 2081
rect 1020 2047 1032 2081
rect 974 2041 1032 2047
rect 1092 2081 1150 2087
rect 1092 2047 1104 2081
rect 1138 2047 1150 2081
rect 1092 2041 1150 2047
rect -1203 1988 -1157 2000
rect -1203 -1988 -1197 1988
rect -1163 -1988 -1157 1988
rect -1203 -2000 -1157 -1988
rect -1085 1988 -1039 2000
rect -1085 -1988 -1079 1988
rect -1045 -1988 -1039 1988
rect -1085 -2000 -1039 -1988
rect -967 1988 -921 2000
rect -967 -1988 -961 1988
rect -927 -1988 -921 1988
rect -967 -2000 -921 -1988
rect -849 1988 -803 2000
rect -849 -1988 -843 1988
rect -809 -1988 -803 1988
rect -849 -2000 -803 -1988
rect -731 1988 -685 2000
rect -731 -1988 -725 1988
rect -691 -1988 -685 1988
rect -731 -2000 -685 -1988
rect -613 1988 -567 2000
rect -613 -1988 -607 1988
rect -573 -1988 -567 1988
rect -613 -2000 -567 -1988
rect -495 1988 -449 2000
rect -495 -1988 -489 1988
rect -455 -1988 -449 1988
rect -495 -2000 -449 -1988
rect -377 1988 -331 2000
rect -377 -1988 -371 1988
rect -337 -1988 -331 1988
rect -377 -2000 -331 -1988
rect -259 1988 -213 2000
rect -259 -1988 -253 1988
rect -219 -1988 -213 1988
rect -259 -2000 -213 -1988
rect -141 1988 -95 2000
rect -141 -1988 -135 1988
rect -101 -1988 -95 1988
rect -141 -2000 -95 -1988
rect -23 1988 23 2000
rect -23 -1988 -17 1988
rect 17 -1988 23 1988
rect -23 -2000 23 -1988
rect 95 1988 141 2000
rect 95 -1988 101 1988
rect 135 -1988 141 1988
rect 95 -2000 141 -1988
rect 213 1988 259 2000
rect 213 -1988 219 1988
rect 253 -1988 259 1988
rect 213 -2000 259 -1988
rect 331 1988 377 2000
rect 331 -1988 337 1988
rect 371 -1988 377 1988
rect 331 -2000 377 -1988
rect 449 1988 495 2000
rect 449 -1988 455 1988
rect 489 -1988 495 1988
rect 449 -2000 495 -1988
rect 567 1988 613 2000
rect 567 -1988 573 1988
rect 607 -1988 613 1988
rect 567 -2000 613 -1988
rect 685 1988 731 2000
rect 685 -1988 691 1988
rect 725 -1988 731 1988
rect 685 -2000 731 -1988
rect 803 1988 849 2000
rect 803 -1988 809 1988
rect 843 -1988 849 1988
rect 803 -2000 849 -1988
rect 921 1988 967 2000
rect 921 -1988 927 1988
rect 961 -1988 967 1988
rect 921 -2000 967 -1988
rect 1039 1988 1085 2000
rect 1039 -1988 1045 1988
rect 1079 -1988 1085 1988
rect 1039 -2000 1085 -1988
rect 1157 1988 1203 2000
rect 1157 -1988 1163 1988
rect 1197 -1988 1203 1988
rect 1157 -2000 1203 -1988
rect -1150 -2047 -1092 -2041
rect -1150 -2081 -1138 -2047
rect -1104 -2081 -1092 -2047
rect -1150 -2087 -1092 -2081
rect -1032 -2047 -974 -2041
rect -1032 -2081 -1020 -2047
rect -986 -2081 -974 -2047
rect -1032 -2087 -974 -2081
rect -914 -2047 -856 -2041
rect -914 -2081 -902 -2047
rect -868 -2081 -856 -2047
rect -914 -2087 -856 -2081
rect -796 -2047 -738 -2041
rect -796 -2081 -784 -2047
rect -750 -2081 -738 -2047
rect -796 -2087 -738 -2081
rect -678 -2047 -620 -2041
rect -678 -2081 -666 -2047
rect -632 -2081 -620 -2047
rect -678 -2087 -620 -2081
rect -560 -2047 -502 -2041
rect -560 -2081 -548 -2047
rect -514 -2081 -502 -2047
rect -560 -2087 -502 -2081
rect -442 -2047 -384 -2041
rect -442 -2081 -430 -2047
rect -396 -2081 -384 -2047
rect -442 -2087 -384 -2081
rect -324 -2047 -266 -2041
rect -324 -2081 -312 -2047
rect -278 -2081 -266 -2047
rect -324 -2087 -266 -2081
rect -206 -2047 -148 -2041
rect -206 -2081 -194 -2047
rect -160 -2081 -148 -2047
rect -206 -2087 -148 -2081
rect -88 -2047 -30 -2041
rect -88 -2081 -76 -2047
rect -42 -2081 -30 -2047
rect -88 -2087 -30 -2081
rect 30 -2047 88 -2041
rect 30 -2081 42 -2047
rect 76 -2081 88 -2047
rect 30 -2087 88 -2081
rect 148 -2047 206 -2041
rect 148 -2081 160 -2047
rect 194 -2081 206 -2047
rect 148 -2087 206 -2081
rect 266 -2047 324 -2041
rect 266 -2081 278 -2047
rect 312 -2081 324 -2047
rect 266 -2087 324 -2081
rect 384 -2047 442 -2041
rect 384 -2081 396 -2047
rect 430 -2081 442 -2047
rect 384 -2087 442 -2081
rect 502 -2047 560 -2041
rect 502 -2081 514 -2047
rect 548 -2081 560 -2047
rect 502 -2087 560 -2081
rect 620 -2047 678 -2041
rect 620 -2081 632 -2047
rect 666 -2081 678 -2047
rect 620 -2087 678 -2081
rect 738 -2047 796 -2041
rect 738 -2081 750 -2047
rect 784 -2081 796 -2047
rect 738 -2087 796 -2081
rect 856 -2047 914 -2041
rect 856 -2081 868 -2047
rect 902 -2081 914 -2047
rect 856 -2087 914 -2081
rect 974 -2047 1032 -2041
rect 974 -2081 986 -2047
rect 1020 -2081 1032 -2047
rect 974 -2087 1032 -2081
rect 1092 -2047 1150 -2041
rect 1092 -2081 1104 -2047
rect 1138 -2081 1150 -2047
rect 1092 -2087 1150 -2081
<< properties >>
string FIXED_BBOX -1294 -2166 1294 2166
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 20 l 0.3 m 1 nf 20 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
