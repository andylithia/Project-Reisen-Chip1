magic
tech sky130A
timestamp 1672031511
<< metal1 >>
rect -3 62 61 66
rect -3 4 0 62
rect 58 4 61 62
rect -3 0 61 4
<< via1 >>
rect 0 4 58 62
<< metal2 >>
rect -3 62 61 66
rect -3 4 0 62
rect 58 4 61 62
rect -3 0 61 4
<< end >>
