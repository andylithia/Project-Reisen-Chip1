magic
tech sky130A
magscale 1 2
timestamp 1672102789
<< pwell >>
rect 19907 3007 21503 3409
rect 20980 -5420 21600 -3920
<< psubdiff >>
rect 19943 3339 20039 3373
rect 21371 3339 21467 3373
rect 19943 3277 19977 3339
rect 21433 3277 21467 3339
rect 19943 3077 19977 3139
rect 21433 3077 21467 3139
rect 19943 3043 20039 3077
rect 21371 3043 21467 3077
<< psubdiffcont >>
rect 20039 3339 21371 3373
rect 19943 3139 19977 3277
rect 21433 3139 21467 3277
rect 20039 3043 21371 3077
<< xpolycontact >>
rect 20073 3173 20505 3243
rect 20905 3173 21337 3243
<< xpolyres >>
rect 20505 3173 20905 3243
<< locali >>
rect 19943 3339 20039 3373
rect 21371 3339 21467 3373
rect 19943 3277 19977 3339
rect 21433 3277 21467 3339
rect 19943 3077 19977 3139
rect 21433 3077 21467 3139
rect 19943 3043 20039 3077
rect 21371 3043 21467 3077
rect 19980 1760 20300 3043
rect 21100 1800 21420 3043
rect 19980 1460 20020 1760
rect 20260 1460 20300 1760
rect 19980 1420 20300 1460
rect 20340 -1680 20660 -1640
rect 20340 -2200 20380 -1680
rect 20620 -2200 20660 -1680
rect 20340 -2240 20660 -2200
rect 21280 -3060 21560 -3040
rect 21280 -3200 21300 -3060
rect 21540 -3200 21560 -3060
rect 21280 -3220 21560 -3200
rect 20940 -5280 21080 -4120
<< viali >>
rect 20091 3189 20488 3227
rect 20922 3189 21319 3227
rect 20020 1460 20260 1760
rect 20380 -2200 20620 -1680
rect 21300 -3200 21540 -3060
<< metal1 >>
rect 20920 3280 21360 3300
rect 20060 3227 20100 3260
rect 20460 3227 20500 3260
rect 20920 3233 20940 3280
rect 20060 3189 20091 3227
rect 20488 3189 20500 3227
rect 20060 3160 20100 3189
rect 20460 3160 20500 3189
rect 20910 3227 20940 3233
rect 20910 3189 20922 3227
rect 20910 3183 20940 3189
rect 20920 3140 20940 3183
rect 21340 3140 21360 3280
rect 20920 3120 21360 3140
rect 19980 1760 20800 1800
rect 19980 1460 20020 1760
rect 20260 1460 20800 1760
rect 19980 1420 20800 1460
rect 14510 -1100 14560 -1060
rect 14400 -1880 14460 -1860
rect 14400 -1960 14460 -1940
rect 14499 -1960 14539 -1580
rect 20340 -1680 20660 -1640
rect 20340 -2200 20380 -1680
rect 20620 -2200 20660 -1680
rect 20340 -2240 20660 -2200
rect 21280 -3060 21560 -3040
rect 21280 -3200 21300 -3060
rect 21540 -3200 21560 -3060
rect 21280 -3220 21560 -3200
rect 21180 -4100 21420 -4080
rect 21180 -4500 21200 -4100
rect 21400 -4500 21420 -4100
rect 21180 -4520 21420 -4500
rect 21180 -4860 21260 -4820
rect 21180 -5260 21260 -5220
rect 21360 -4860 21440 -4820
rect 21360 -5260 21440 -5220
rect 6000 -11248 14000 -11000
rect 6000 -11300 6614 -11248
rect 6666 -11300 6934 -11248
rect 6986 -11300 7254 -11248
rect 7306 -11300 7574 -11248
rect 7626 -11300 7894 -11248
rect 7946 -11300 8214 -11248
rect 8266 -11300 8534 -11248
rect 8586 -11300 8854 -11248
rect 8906 -11300 9174 -11248
rect 9226 -11300 9494 -11248
rect 9546 -11300 9814 -11248
rect 9866 -11300 10134 -11248
rect 10186 -11300 10454 -11248
rect 10506 -11300 10774 -11248
rect 10826 -11300 11094 -11248
rect 11146 -11300 11414 -11248
rect 11466 -11300 11734 -11248
rect 11786 -11300 12054 -11248
rect 12106 -11300 12374 -11248
rect 12426 -11300 12694 -11248
rect 12746 -11300 13014 -11248
rect 13066 -11300 13334 -11248
rect 13386 -11300 14000 -11248
rect 6000 -11454 14000 -11300
rect 6000 -11506 6244 -11454
rect 6296 -11506 13710 -11454
rect 13762 -11506 14000 -11454
rect 6000 -11540 14000 -11506
rect 6000 -11774 6540 -11540
rect 6000 -11826 6244 -11774
rect 6296 -11826 6540 -11774
rect 6000 -12094 6540 -11826
rect 6000 -12146 6244 -12094
rect 6296 -12146 6540 -12094
rect 6000 -12414 6540 -12146
rect 6000 -12466 6244 -12414
rect 6296 -12466 6540 -12414
rect 6000 -12734 6540 -12466
rect 6000 -12786 6244 -12734
rect 6296 -12786 6540 -12734
rect 6000 -13054 6540 -12786
rect 6000 -13106 6244 -13054
rect 6296 -13106 6540 -13054
rect 6000 -13374 6540 -13106
rect 6000 -13426 6244 -13374
rect 6296 -13426 6540 -13374
rect 6000 -13694 6540 -13426
rect 6000 -13746 6244 -13694
rect 6296 -13746 6540 -13694
rect 6000 -14014 6540 -13746
rect 6000 -14066 6244 -14014
rect 6296 -14066 6540 -14014
rect 6000 -14334 6540 -14066
rect 6000 -14386 6244 -14334
rect 6296 -14386 6540 -14334
rect 6000 -14654 6540 -14386
rect 6000 -14706 6244 -14654
rect 6296 -14706 6540 -14654
rect 6000 -14974 6540 -14706
rect 6000 -15026 6244 -14974
rect 6296 -15026 6540 -14974
rect 6000 -15294 6540 -15026
rect 6000 -15346 6244 -15294
rect 6296 -15346 6540 -15294
rect 6000 -15614 6540 -15346
rect 6000 -15666 6244 -15614
rect 6296 -15666 6540 -15614
rect 6000 -15934 6540 -15666
rect 6000 -15986 6244 -15934
rect 6296 -15986 6540 -15934
rect 6000 -16254 6540 -15986
rect 6000 -16306 6244 -16254
rect 6296 -16306 6540 -16254
rect 6000 -16574 6540 -16306
rect 6000 -16626 6244 -16574
rect 6296 -16626 6540 -16574
rect 6000 -16894 6540 -16626
rect 6000 -16946 6244 -16894
rect 6296 -16946 6540 -16894
rect 6000 -17214 6540 -16946
rect 6000 -17266 6244 -17214
rect 6296 -17266 6540 -17214
rect 6000 -17534 6540 -17266
rect 6000 -17586 6244 -17534
rect 6296 -17586 6540 -17534
rect 6000 -17854 6540 -17586
rect 6000 -17906 6244 -17854
rect 6296 -17906 6540 -17854
rect 6000 -18174 6540 -17906
rect 6000 -18226 6244 -18174
rect 6296 -18226 6540 -18174
rect 6000 -18460 6540 -18226
rect 13460 -11774 14000 -11540
rect 13460 -11826 13710 -11774
rect 13762 -11826 14000 -11774
rect 13460 -12094 14000 -11826
rect 13460 -12146 13710 -12094
rect 13762 -12146 14000 -12094
rect 13460 -12414 14000 -12146
rect 13460 -12466 13710 -12414
rect 13762 -12466 14000 -12414
rect 13460 -12734 14000 -12466
rect 13460 -12786 13710 -12734
rect 13762 -12786 14000 -12734
rect 13460 -13054 14000 -12786
rect 13460 -13106 13710 -13054
rect 13762 -13106 14000 -13054
rect 13460 -13374 14000 -13106
rect 13460 -13426 13710 -13374
rect 13762 -13426 14000 -13374
rect 13460 -13694 14000 -13426
rect 13460 -13746 13710 -13694
rect 13762 -13746 14000 -13694
rect 13460 -14014 14000 -13746
rect 13460 -14066 13710 -14014
rect 13762 -14066 14000 -14014
rect 13460 -14334 14000 -14066
rect 13460 -14386 13710 -14334
rect 13762 -14386 14000 -14334
rect 13460 -14654 14000 -14386
rect 13460 -14706 13710 -14654
rect 13762 -14706 14000 -14654
rect 13460 -14974 14000 -14706
rect 13460 -15026 13710 -14974
rect 13762 -15026 14000 -14974
rect 13460 -15294 14000 -15026
rect 13460 -15346 13710 -15294
rect 13762 -15346 14000 -15294
rect 13460 -15614 14000 -15346
rect 13460 -15666 13710 -15614
rect 13762 -15666 14000 -15614
rect 13460 -15934 14000 -15666
rect 13460 -15986 13710 -15934
rect 13762 -15986 14000 -15934
rect 13460 -16254 14000 -15986
rect 13460 -16306 13710 -16254
rect 13762 -16306 14000 -16254
rect 13460 -16574 14000 -16306
rect 13460 -16626 13710 -16574
rect 13762 -16626 14000 -16574
rect 13460 -16894 14000 -16626
rect 13460 -16946 13710 -16894
rect 13762 -16946 14000 -16894
rect 13460 -17214 14000 -16946
rect 13460 -17266 13710 -17214
rect 13762 -17266 14000 -17214
rect 13460 -17534 14000 -17266
rect 13460 -17586 13710 -17534
rect 13762 -17586 14000 -17534
rect 13460 -17854 14000 -17586
rect 13460 -17906 13710 -17854
rect 13762 -17906 14000 -17854
rect 13460 -18174 14000 -17906
rect 13460 -18226 13710 -18174
rect 13762 -18226 14000 -18174
rect 13460 -18460 14000 -18226
rect 6000 -18494 14000 -18460
rect 6000 -18546 6244 -18494
rect 6296 -18546 13710 -18494
rect 13762 -18546 14000 -18494
rect 6000 -18704 14000 -18546
rect 6000 -18756 6614 -18704
rect 6666 -18756 6934 -18704
rect 6986 -18756 7254 -18704
rect 7306 -18756 7574 -18704
rect 7626 -18756 7894 -18704
rect 7946 -18756 8214 -18704
rect 8266 -18756 8534 -18704
rect 8586 -18756 8854 -18704
rect 8906 -18756 9174 -18704
rect 9226 -18756 9494 -18704
rect 9546 -18756 9814 -18704
rect 9866 -18756 10134 -18704
rect 10186 -18756 10454 -18704
rect 10506 -18756 10774 -18704
rect 10826 -18756 11094 -18704
rect 11146 -18756 11414 -18704
rect 11466 -18756 11734 -18704
rect 11786 -18756 12054 -18704
rect 12106 -18756 12374 -18704
rect 12426 -18756 12694 -18704
rect 12746 -18756 13014 -18704
rect 13066 -18756 13334 -18704
rect 13386 -18756 14000 -18704
rect 6000 -19000 14000 -18756
rect 18000 -11248 26000 -11000
rect 18000 -11300 18614 -11248
rect 18666 -11300 18934 -11248
rect 18986 -11300 19254 -11248
rect 19306 -11300 19574 -11248
rect 19626 -11300 19894 -11248
rect 19946 -11300 20214 -11248
rect 20266 -11300 20534 -11248
rect 20586 -11300 20854 -11248
rect 20906 -11300 21174 -11248
rect 21226 -11300 21494 -11248
rect 21546 -11300 21814 -11248
rect 21866 -11300 22134 -11248
rect 22186 -11300 22454 -11248
rect 22506 -11300 22774 -11248
rect 22826 -11300 23094 -11248
rect 23146 -11300 23414 -11248
rect 23466 -11300 23734 -11248
rect 23786 -11300 24054 -11248
rect 24106 -11300 24374 -11248
rect 24426 -11300 24694 -11248
rect 24746 -11300 25014 -11248
rect 25066 -11300 25334 -11248
rect 25386 -11300 26000 -11248
rect 18000 -11454 26000 -11300
rect 18000 -11506 18244 -11454
rect 18296 -11506 25710 -11454
rect 25762 -11506 26000 -11454
rect 18000 -11540 26000 -11506
rect 18000 -11774 18540 -11540
rect 18000 -11826 18244 -11774
rect 18296 -11826 18540 -11774
rect 18000 -12094 18540 -11826
rect 18000 -12146 18244 -12094
rect 18296 -12146 18540 -12094
rect 18000 -12414 18540 -12146
rect 18000 -12466 18244 -12414
rect 18296 -12466 18540 -12414
rect 18000 -12734 18540 -12466
rect 18000 -12786 18244 -12734
rect 18296 -12786 18540 -12734
rect 18000 -13054 18540 -12786
rect 18000 -13106 18244 -13054
rect 18296 -13106 18540 -13054
rect 18000 -13374 18540 -13106
rect 18000 -13426 18244 -13374
rect 18296 -13426 18540 -13374
rect 18000 -13694 18540 -13426
rect 18000 -13746 18244 -13694
rect 18296 -13746 18540 -13694
rect 18000 -14014 18540 -13746
rect 18000 -14066 18244 -14014
rect 18296 -14066 18540 -14014
rect 18000 -14334 18540 -14066
rect 18000 -14386 18244 -14334
rect 18296 -14386 18540 -14334
rect 18000 -14654 18540 -14386
rect 18000 -14706 18244 -14654
rect 18296 -14706 18540 -14654
rect 18000 -14974 18540 -14706
rect 18000 -15026 18244 -14974
rect 18296 -15026 18540 -14974
rect 18000 -15294 18540 -15026
rect 18000 -15346 18244 -15294
rect 18296 -15346 18540 -15294
rect 18000 -15614 18540 -15346
rect 18000 -15666 18244 -15614
rect 18296 -15666 18540 -15614
rect 18000 -15934 18540 -15666
rect 18000 -15986 18244 -15934
rect 18296 -15986 18540 -15934
rect 18000 -16254 18540 -15986
rect 18000 -16306 18244 -16254
rect 18296 -16306 18540 -16254
rect 18000 -16574 18540 -16306
rect 18000 -16626 18244 -16574
rect 18296 -16626 18540 -16574
rect 18000 -16894 18540 -16626
rect 18000 -16946 18244 -16894
rect 18296 -16946 18540 -16894
rect 18000 -17214 18540 -16946
rect 18000 -17266 18244 -17214
rect 18296 -17266 18540 -17214
rect 18000 -17534 18540 -17266
rect 18000 -17586 18244 -17534
rect 18296 -17586 18540 -17534
rect 18000 -17854 18540 -17586
rect 18000 -17906 18244 -17854
rect 18296 -17906 18540 -17854
rect 18000 -18174 18540 -17906
rect 18000 -18226 18244 -18174
rect 18296 -18226 18540 -18174
rect 18000 -18460 18540 -18226
rect 25460 -11774 26000 -11540
rect 25460 -11826 25710 -11774
rect 25762 -11826 26000 -11774
rect 25460 -12094 26000 -11826
rect 25460 -12146 25710 -12094
rect 25762 -12146 26000 -12094
rect 25460 -12414 26000 -12146
rect 25460 -12466 25710 -12414
rect 25762 -12466 26000 -12414
rect 25460 -12734 26000 -12466
rect 25460 -12786 25710 -12734
rect 25762 -12786 26000 -12734
rect 25460 -13054 26000 -12786
rect 25460 -13106 25710 -13054
rect 25762 -13106 26000 -13054
rect 25460 -13374 26000 -13106
rect 25460 -13426 25710 -13374
rect 25762 -13426 26000 -13374
rect 25460 -13694 26000 -13426
rect 25460 -13746 25710 -13694
rect 25762 -13746 26000 -13694
rect 25460 -14014 26000 -13746
rect 25460 -14066 25710 -14014
rect 25762 -14066 26000 -14014
rect 25460 -14334 26000 -14066
rect 25460 -14386 25710 -14334
rect 25762 -14386 26000 -14334
rect 25460 -14654 26000 -14386
rect 25460 -14706 25710 -14654
rect 25762 -14706 26000 -14654
rect 25460 -14974 26000 -14706
rect 25460 -15026 25710 -14974
rect 25762 -15026 26000 -14974
rect 25460 -15294 26000 -15026
rect 25460 -15346 25710 -15294
rect 25762 -15346 26000 -15294
rect 25460 -15614 26000 -15346
rect 25460 -15666 25710 -15614
rect 25762 -15666 26000 -15614
rect 25460 -15934 26000 -15666
rect 25460 -15986 25710 -15934
rect 25762 -15986 26000 -15934
rect 25460 -16254 26000 -15986
rect 25460 -16306 25710 -16254
rect 25762 -16306 26000 -16254
rect 25460 -16574 26000 -16306
rect 25460 -16626 25710 -16574
rect 25762 -16626 26000 -16574
rect 25460 -16894 26000 -16626
rect 25460 -16946 25710 -16894
rect 25762 -16946 26000 -16894
rect 25460 -17214 26000 -16946
rect 25460 -17266 25710 -17214
rect 25762 -17266 26000 -17214
rect 25460 -17534 26000 -17266
rect 25460 -17586 25710 -17534
rect 25762 -17586 26000 -17534
rect 25460 -17854 26000 -17586
rect 25460 -17906 25710 -17854
rect 25762 -17906 26000 -17854
rect 25460 -18174 26000 -17906
rect 25460 -18226 25710 -18174
rect 25762 -18226 26000 -18174
rect 25460 -18460 26000 -18226
rect 18000 -18494 26000 -18460
rect 18000 -18546 18244 -18494
rect 18296 -18546 25710 -18494
rect 25762 -18546 26000 -18494
rect 18000 -18704 26000 -18546
rect 18000 -18756 18614 -18704
rect 18666 -18756 18934 -18704
rect 18986 -18756 19254 -18704
rect 19306 -18756 19574 -18704
rect 19626 -18756 19894 -18704
rect 19946 -18756 20214 -18704
rect 20266 -18756 20534 -18704
rect 20586 -18756 20854 -18704
rect 20906 -18756 21174 -18704
rect 21226 -18756 21494 -18704
rect 21546 -18756 21814 -18704
rect 21866 -18756 22134 -18704
rect 22186 -18756 22454 -18704
rect 22506 -18756 22774 -18704
rect 22826 -18756 23094 -18704
rect 23146 -18756 23414 -18704
rect 23466 -18756 23734 -18704
rect 23786 -18756 24054 -18704
rect 24106 -18756 24374 -18704
rect 24426 -18756 24694 -18704
rect 24746 -18756 25014 -18704
rect 25066 -18756 25334 -18704
rect 25386 -18756 26000 -18704
rect 18000 -19000 26000 -18756
rect 30000 -11248 38000 -11000
rect 30000 -11300 30614 -11248
rect 30666 -11300 30934 -11248
rect 30986 -11300 31254 -11248
rect 31306 -11300 31574 -11248
rect 31626 -11300 31894 -11248
rect 31946 -11300 32214 -11248
rect 32266 -11300 32534 -11248
rect 32586 -11300 32854 -11248
rect 32906 -11300 33174 -11248
rect 33226 -11300 33494 -11248
rect 33546 -11300 33814 -11248
rect 33866 -11300 34134 -11248
rect 34186 -11300 34454 -11248
rect 34506 -11300 34774 -11248
rect 34826 -11300 35094 -11248
rect 35146 -11300 35414 -11248
rect 35466 -11300 35734 -11248
rect 35786 -11300 36054 -11248
rect 36106 -11300 36374 -11248
rect 36426 -11300 36694 -11248
rect 36746 -11300 37014 -11248
rect 37066 -11300 37334 -11248
rect 37386 -11300 38000 -11248
rect 30000 -11454 38000 -11300
rect 30000 -11506 30244 -11454
rect 30296 -11506 37710 -11454
rect 37762 -11506 38000 -11454
rect 30000 -11540 38000 -11506
rect 30000 -11774 30540 -11540
rect 30000 -11826 30244 -11774
rect 30296 -11826 30540 -11774
rect 30000 -12094 30540 -11826
rect 30000 -12146 30244 -12094
rect 30296 -12146 30540 -12094
rect 30000 -12414 30540 -12146
rect 30000 -12466 30244 -12414
rect 30296 -12466 30540 -12414
rect 30000 -12734 30540 -12466
rect 30000 -12786 30244 -12734
rect 30296 -12786 30540 -12734
rect 30000 -13054 30540 -12786
rect 30000 -13106 30244 -13054
rect 30296 -13106 30540 -13054
rect 30000 -13374 30540 -13106
rect 30000 -13426 30244 -13374
rect 30296 -13426 30540 -13374
rect 30000 -13694 30540 -13426
rect 30000 -13746 30244 -13694
rect 30296 -13746 30540 -13694
rect 30000 -14014 30540 -13746
rect 30000 -14066 30244 -14014
rect 30296 -14066 30540 -14014
rect 30000 -14334 30540 -14066
rect 30000 -14386 30244 -14334
rect 30296 -14386 30540 -14334
rect 30000 -14654 30540 -14386
rect 30000 -14706 30244 -14654
rect 30296 -14706 30540 -14654
rect 30000 -14974 30540 -14706
rect 30000 -15026 30244 -14974
rect 30296 -15026 30540 -14974
rect 30000 -15294 30540 -15026
rect 30000 -15346 30244 -15294
rect 30296 -15346 30540 -15294
rect 30000 -15614 30540 -15346
rect 30000 -15666 30244 -15614
rect 30296 -15666 30540 -15614
rect 30000 -15934 30540 -15666
rect 30000 -15986 30244 -15934
rect 30296 -15986 30540 -15934
rect 30000 -16254 30540 -15986
rect 30000 -16306 30244 -16254
rect 30296 -16306 30540 -16254
rect 30000 -16574 30540 -16306
rect 30000 -16626 30244 -16574
rect 30296 -16626 30540 -16574
rect 30000 -16894 30540 -16626
rect 30000 -16946 30244 -16894
rect 30296 -16946 30540 -16894
rect 30000 -17214 30540 -16946
rect 30000 -17266 30244 -17214
rect 30296 -17266 30540 -17214
rect 30000 -17534 30540 -17266
rect 30000 -17586 30244 -17534
rect 30296 -17586 30540 -17534
rect 30000 -17854 30540 -17586
rect 30000 -17906 30244 -17854
rect 30296 -17906 30540 -17854
rect 30000 -18174 30540 -17906
rect 30000 -18226 30244 -18174
rect 30296 -18226 30540 -18174
rect 30000 -18460 30540 -18226
rect 37460 -11774 38000 -11540
rect 37460 -11826 37710 -11774
rect 37762 -11826 38000 -11774
rect 37460 -12094 38000 -11826
rect 37460 -12146 37710 -12094
rect 37762 -12146 38000 -12094
rect 37460 -12414 38000 -12146
rect 37460 -12466 37710 -12414
rect 37762 -12466 38000 -12414
rect 37460 -12734 38000 -12466
rect 37460 -12786 37710 -12734
rect 37762 -12786 38000 -12734
rect 37460 -13054 38000 -12786
rect 37460 -13106 37710 -13054
rect 37762 -13106 38000 -13054
rect 37460 -13374 38000 -13106
rect 37460 -13426 37710 -13374
rect 37762 -13426 38000 -13374
rect 37460 -13694 38000 -13426
rect 37460 -13746 37710 -13694
rect 37762 -13746 38000 -13694
rect 37460 -14014 38000 -13746
rect 37460 -14066 37710 -14014
rect 37762 -14066 38000 -14014
rect 37460 -14334 38000 -14066
rect 37460 -14386 37710 -14334
rect 37762 -14386 38000 -14334
rect 37460 -14654 38000 -14386
rect 37460 -14706 37710 -14654
rect 37762 -14706 38000 -14654
rect 37460 -14974 38000 -14706
rect 37460 -15026 37710 -14974
rect 37762 -15026 38000 -14974
rect 37460 -15294 38000 -15026
rect 37460 -15346 37710 -15294
rect 37762 -15346 38000 -15294
rect 37460 -15614 38000 -15346
rect 37460 -15666 37710 -15614
rect 37762 -15666 38000 -15614
rect 37460 -15934 38000 -15666
rect 37460 -15986 37710 -15934
rect 37762 -15986 38000 -15934
rect 37460 -16254 38000 -15986
rect 37460 -16306 37710 -16254
rect 37762 -16306 38000 -16254
rect 37460 -16574 38000 -16306
rect 37460 -16626 37710 -16574
rect 37762 -16626 38000 -16574
rect 37460 -16894 38000 -16626
rect 37460 -16946 37710 -16894
rect 37762 -16946 38000 -16894
rect 37460 -17214 38000 -16946
rect 37460 -17266 37710 -17214
rect 37762 -17266 38000 -17214
rect 37460 -17534 38000 -17266
rect 37460 -17586 37710 -17534
rect 37762 -17586 38000 -17534
rect 37460 -17854 38000 -17586
rect 37460 -17906 37710 -17854
rect 37762 -17906 38000 -17854
rect 37460 -18174 38000 -17906
rect 37460 -18226 37710 -18174
rect 37762 -18226 38000 -18174
rect 37460 -18460 38000 -18226
rect 30000 -18494 38000 -18460
rect 30000 -18546 30244 -18494
rect 30296 -18546 37710 -18494
rect 37762 -18546 38000 -18494
rect 30000 -18704 38000 -18546
rect 30000 -18756 30614 -18704
rect 30666 -18756 30934 -18704
rect 30986 -18756 31254 -18704
rect 31306 -18756 31574 -18704
rect 31626 -18756 31894 -18704
rect 31946 -18756 32214 -18704
rect 32266 -18756 32534 -18704
rect 32586 -18756 32854 -18704
rect 32906 -18756 33174 -18704
rect 33226 -18756 33494 -18704
rect 33546 -18756 33814 -18704
rect 33866 -18756 34134 -18704
rect 34186 -18756 34454 -18704
rect 34506 -18756 34774 -18704
rect 34826 -18756 35094 -18704
rect 35146 -18756 35414 -18704
rect 35466 -18756 35734 -18704
rect 35786 -18756 36054 -18704
rect 36106 -18756 36374 -18704
rect 36426 -18756 36694 -18704
rect 36746 -18756 37014 -18704
rect 37066 -18756 37334 -18704
rect 37386 -18756 38000 -18704
rect 30000 -19000 38000 -18756
rect 42000 -11248 50000 -11000
rect 42000 -11300 42614 -11248
rect 42666 -11300 42934 -11248
rect 42986 -11300 43254 -11248
rect 43306 -11300 43574 -11248
rect 43626 -11300 43894 -11248
rect 43946 -11300 44214 -11248
rect 44266 -11300 44534 -11248
rect 44586 -11300 44854 -11248
rect 44906 -11300 45174 -11248
rect 45226 -11300 45494 -11248
rect 45546 -11300 45814 -11248
rect 45866 -11300 46134 -11248
rect 46186 -11300 46454 -11248
rect 46506 -11300 46774 -11248
rect 46826 -11300 47094 -11248
rect 47146 -11300 47414 -11248
rect 47466 -11300 47734 -11248
rect 47786 -11300 48054 -11248
rect 48106 -11300 48374 -11248
rect 48426 -11300 48694 -11248
rect 48746 -11300 49014 -11248
rect 49066 -11300 49334 -11248
rect 49386 -11300 50000 -11248
rect 42000 -11454 50000 -11300
rect 42000 -11506 42247 -11454
rect 42299 -11506 49701 -11454
rect 49753 -11506 50000 -11454
rect 42000 -11540 50000 -11506
rect 42000 -11774 42540 -11540
rect 42000 -11826 42247 -11774
rect 42299 -11826 42540 -11774
rect 42000 -12094 42540 -11826
rect 42000 -12146 42247 -12094
rect 42299 -12146 42540 -12094
rect 42000 -12414 42540 -12146
rect 42000 -12466 42247 -12414
rect 42299 -12466 42540 -12414
rect 42000 -12734 42540 -12466
rect 42000 -12786 42247 -12734
rect 42299 -12786 42540 -12734
rect 42000 -13054 42540 -12786
rect 42000 -13106 42247 -13054
rect 42299 -13106 42540 -13054
rect 42000 -13374 42540 -13106
rect 42000 -13426 42247 -13374
rect 42299 -13426 42540 -13374
rect 42000 -13694 42540 -13426
rect 42000 -13746 42247 -13694
rect 42299 -13746 42540 -13694
rect 42000 -14014 42540 -13746
rect 42000 -14066 42247 -14014
rect 42299 -14066 42540 -14014
rect 42000 -14334 42540 -14066
rect 42000 -14386 42247 -14334
rect 42299 -14386 42540 -14334
rect 42000 -14654 42540 -14386
rect 42000 -14706 42247 -14654
rect 42299 -14706 42540 -14654
rect 42000 -14974 42540 -14706
rect 42000 -15026 42247 -14974
rect 42299 -15026 42540 -14974
rect 42000 -15294 42540 -15026
rect 42000 -15346 42247 -15294
rect 42299 -15346 42540 -15294
rect 42000 -15614 42540 -15346
rect 42000 -15666 42247 -15614
rect 42299 -15666 42540 -15614
rect 42000 -15934 42540 -15666
rect 42000 -15986 42247 -15934
rect 42299 -15986 42540 -15934
rect 42000 -16254 42540 -15986
rect 42000 -16306 42247 -16254
rect 42299 -16306 42540 -16254
rect 42000 -16574 42540 -16306
rect 42000 -16626 42247 -16574
rect 42299 -16626 42540 -16574
rect 42000 -16894 42540 -16626
rect 42000 -16946 42247 -16894
rect 42299 -16946 42540 -16894
rect 42000 -17214 42540 -16946
rect 42000 -17266 42247 -17214
rect 42299 -17266 42540 -17214
rect 42000 -17534 42540 -17266
rect 42000 -17586 42247 -17534
rect 42299 -17586 42540 -17534
rect 42000 -17854 42540 -17586
rect 42000 -17906 42247 -17854
rect 42299 -17906 42540 -17854
rect 42000 -18174 42540 -17906
rect 42000 -18226 42247 -18174
rect 42299 -18226 42540 -18174
rect 42000 -18460 42540 -18226
rect 49460 -11774 50000 -11540
rect 49460 -11826 49701 -11774
rect 49753 -11826 50000 -11774
rect 49460 -12094 50000 -11826
rect 49460 -12146 49701 -12094
rect 49753 -12146 50000 -12094
rect 49460 -12414 50000 -12146
rect 49460 -12466 49701 -12414
rect 49753 -12466 50000 -12414
rect 49460 -12734 50000 -12466
rect 49460 -12786 49701 -12734
rect 49753 -12786 50000 -12734
rect 49460 -13054 50000 -12786
rect 49460 -13106 49701 -13054
rect 49753 -13106 50000 -13054
rect 49460 -13374 50000 -13106
rect 49460 -13426 49701 -13374
rect 49753 -13426 50000 -13374
rect 49460 -13694 50000 -13426
rect 49460 -13746 49701 -13694
rect 49753 -13746 50000 -13694
rect 49460 -14014 50000 -13746
rect 49460 -14066 49701 -14014
rect 49753 -14066 50000 -14014
rect 49460 -14334 50000 -14066
rect 49460 -14386 49701 -14334
rect 49753 -14386 50000 -14334
rect 49460 -14654 50000 -14386
rect 49460 -14706 49701 -14654
rect 49753 -14706 50000 -14654
rect 49460 -14974 50000 -14706
rect 49460 -15026 49701 -14974
rect 49753 -15026 50000 -14974
rect 49460 -15294 50000 -15026
rect 49460 -15346 49701 -15294
rect 49753 -15346 50000 -15294
rect 49460 -15614 50000 -15346
rect 49460 -15666 49701 -15614
rect 49753 -15666 50000 -15614
rect 49460 -15934 50000 -15666
rect 49460 -15986 49701 -15934
rect 49753 -15986 50000 -15934
rect 49460 -16254 50000 -15986
rect 49460 -16306 49701 -16254
rect 49753 -16306 50000 -16254
rect 49460 -16574 50000 -16306
rect 49460 -16626 49701 -16574
rect 49753 -16626 50000 -16574
rect 49460 -16894 50000 -16626
rect 49460 -16946 49701 -16894
rect 49753 -16946 50000 -16894
rect 49460 -17214 50000 -16946
rect 49460 -17266 49701 -17214
rect 49753 -17266 50000 -17214
rect 49460 -17534 50000 -17266
rect 49460 -17586 49701 -17534
rect 49753 -17586 50000 -17534
rect 49460 -17854 50000 -17586
rect 49460 -17906 49701 -17854
rect 49753 -17906 50000 -17854
rect 49460 -18174 50000 -17906
rect 49460 -18226 49701 -18174
rect 49753 -18226 50000 -18174
rect 49460 -18460 50000 -18226
rect 42000 -18494 50000 -18460
rect 42000 -18546 42247 -18494
rect 42299 -18546 49701 -18494
rect 49753 -18546 50000 -18494
rect 42000 -18704 50000 -18546
rect 42000 -18756 42614 -18704
rect 42666 -18756 42934 -18704
rect 42986 -18756 43254 -18704
rect 43306 -18756 43574 -18704
rect 43626 -18756 43894 -18704
rect 43946 -18756 44214 -18704
rect 44266 -18756 44534 -18704
rect 44586 -18756 44854 -18704
rect 44906 -18756 45174 -18704
rect 45226 -18756 45494 -18704
rect 45546 -18756 45814 -18704
rect 45866 -18756 46134 -18704
rect 46186 -18756 46454 -18704
rect 46506 -18756 46774 -18704
rect 46826 -18756 47094 -18704
rect 47146 -18756 47414 -18704
rect 47466 -18756 47734 -18704
rect 47786 -18756 48054 -18704
rect 48106 -18756 48374 -18704
rect 48426 -18756 48694 -18704
rect 48746 -18756 49014 -18704
rect 49066 -18756 49334 -18704
rect 49386 -18756 50000 -18704
rect 42000 -19000 50000 -18756
<< via1 >>
rect 20100 3227 20460 3260
rect 20100 3189 20460 3227
rect 20100 3160 20460 3189
rect 20940 3227 21340 3280
rect 20940 3189 21319 3227
rect 21319 3189 21340 3227
rect 20940 3140 21340 3189
rect 20020 1460 20260 1760
rect 14400 -1940 14460 -1880
rect 20380 -2200 20620 -1680
rect 21300 -3200 21540 -3060
rect 21200 -4500 21400 -4100
rect 21180 -5220 21260 -4860
rect 21360 -5220 21440 -4860
rect 6614 -11300 6666 -11248
rect 6934 -11300 6986 -11248
rect 7254 -11300 7306 -11248
rect 7574 -11300 7626 -11248
rect 7894 -11300 7946 -11248
rect 8214 -11300 8266 -11248
rect 8534 -11300 8586 -11248
rect 8854 -11300 8906 -11248
rect 9174 -11300 9226 -11248
rect 9494 -11300 9546 -11248
rect 9814 -11300 9866 -11248
rect 10134 -11300 10186 -11248
rect 10454 -11300 10506 -11248
rect 10774 -11300 10826 -11248
rect 11094 -11300 11146 -11248
rect 11414 -11300 11466 -11248
rect 11734 -11300 11786 -11248
rect 12054 -11300 12106 -11248
rect 12374 -11300 12426 -11248
rect 12694 -11300 12746 -11248
rect 13014 -11300 13066 -11248
rect 13334 -11300 13386 -11248
rect 6244 -11506 6296 -11454
rect 13710 -11506 13762 -11454
rect 6244 -11826 6296 -11774
rect 6244 -12146 6296 -12094
rect 6244 -12466 6296 -12414
rect 6244 -12786 6296 -12734
rect 6244 -13106 6296 -13054
rect 6244 -13426 6296 -13374
rect 6244 -13746 6296 -13694
rect 6244 -14066 6296 -14014
rect 6244 -14386 6296 -14334
rect 6244 -14706 6296 -14654
rect 6244 -15026 6296 -14974
rect 6244 -15346 6296 -15294
rect 6244 -15666 6296 -15614
rect 6244 -15986 6296 -15934
rect 6244 -16306 6296 -16254
rect 6244 -16626 6296 -16574
rect 6244 -16946 6296 -16894
rect 6244 -17266 6296 -17214
rect 6244 -17586 6296 -17534
rect 6244 -17906 6296 -17854
rect 6244 -18226 6296 -18174
rect 13710 -11826 13762 -11774
rect 13710 -12146 13762 -12094
rect 13710 -12466 13762 -12414
rect 13710 -12786 13762 -12734
rect 13710 -13106 13762 -13054
rect 13710 -13426 13762 -13374
rect 13710 -13746 13762 -13694
rect 13710 -14066 13762 -14014
rect 13710 -14386 13762 -14334
rect 13710 -14706 13762 -14654
rect 13710 -15026 13762 -14974
rect 13710 -15346 13762 -15294
rect 13710 -15666 13762 -15614
rect 13710 -15986 13762 -15934
rect 13710 -16306 13762 -16254
rect 13710 -16626 13762 -16574
rect 13710 -16946 13762 -16894
rect 13710 -17266 13762 -17214
rect 13710 -17586 13762 -17534
rect 13710 -17906 13762 -17854
rect 13710 -18226 13762 -18174
rect 6244 -18546 6296 -18494
rect 13710 -18546 13762 -18494
rect 6614 -18756 6666 -18704
rect 6934 -18756 6986 -18704
rect 7254 -18756 7306 -18704
rect 7574 -18756 7626 -18704
rect 7894 -18756 7946 -18704
rect 8214 -18756 8266 -18704
rect 8534 -18756 8586 -18704
rect 8854 -18756 8906 -18704
rect 9174 -18756 9226 -18704
rect 9494 -18756 9546 -18704
rect 9814 -18756 9866 -18704
rect 10134 -18756 10186 -18704
rect 10454 -18756 10506 -18704
rect 10774 -18756 10826 -18704
rect 11094 -18756 11146 -18704
rect 11414 -18756 11466 -18704
rect 11734 -18756 11786 -18704
rect 12054 -18756 12106 -18704
rect 12374 -18756 12426 -18704
rect 12694 -18756 12746 -18704
rect 13014 -18756 13066 -18704
rect 13334 -18756 13386 -18704
rect 18614 -11300 18666 -11248
rect 18934 -11300 18986 -11248
rect 19254 -11300 19306 -11248
rect 19574 -11300 19626 -11248
rect 19894 -11300 19946 -11248
rect 20214 -11300 20266 -11248
rect 20534 -11300 20586 -11248
rect 20854 -11300 20906 -11248
rect 21174 -11300 21226 -11248
rect 21494 -11300 21546 -11248
rect 21814 -11300 21866 -11248
rect 22134 -11300 22186 -11248
rect 22454 -11300 22506 -11248
rect 22774 -11300 22826 -11248
rect 23094 -11300 23146 -11248
rect 23414 -11300 23466 -11248
rect 23734 -11300 23786 -11248
rect 24054 -11300 24106 -11248
rect 24374 -11300 24426 -11248
rect 24694 -11300 24746 -11248
rect 25014 -11300 25066 -11248
rect 25334 -11300 25386 -11248
rect 18244 -11506 18296 -11454
rect 25710 -11506 25762 -11454
rect 18244 -11826 18296 -11774
rect 18244 -12146 18296 -12094
rect 18244 -12466 18296 -12414
rect 18244 -12786 18296 -12734
rect 18244 -13106 18296 -13054
rect 18244 -13426 18296 -13374
rect 18244 -13746 18296 -13694
rect 18244 -14066 18296 -14014
rect 18244 -14386 18296 -14334
rect 18244 -14706 18296 -14654
rect 18244 -15026 18296 -14974
rect 18244 -15346 18296 -15294
rect 18244 -15666 18296 -15614
rect 18244 -15986 18296 -15934
rect 18244 -16306 18296 -16254
rect 18244 -16626 18296 -16574
rect 18244 -16946 18296 -16894
rect 18244 -17266 18296 -17214
rect 18244 -17586 18296 -17534
rect 18244 -17906 18296 -17854
rect 18244 -18226 18296 -18174
rect 25710 -11826 25762 -11774
rect 25710 -12146 25762 -12094
rect 25710 -12466 25762 -12414
rect 25710 -12786 25762 -12734
rect 25710 -13106 25762 -13054
rect 25710 -13426 25762 -13374
rect 25710 -13746 25762 -13694
rect 25710 -14066 25762 -14014
rect 25710 -14386 25762 -14334
rect 25710 -14706 25762 -14654
rect 25710 -15026 25762 -14974
rect 25710 -15346 25762 -15294
rect 25710 -15666 25762 -15614
rect 25710 -15986 25762 -15934
rect 25710 -16306 25762 -16254
rect 25710 -16626 25762 -16574
rect 25710 -16946 25762 -16894
rect 25710 -17266 25762 -17214
rect 25710 -17586 25762 -17534
rect 25710 -17906 25762 -17854
rect 25710 -18226 25762 -18174
rect 18244 -18546 18296 -18494
rect 25710 -18546 25762 -18494
rect 18614 -18756 18666 -18704
rect 18934 -18756 18986 -18704
rect 19254 -18756 19306 -18704
rect 19574 -18756 19626 -18704
rect 19894 -18756 19946 -18704
rect 20214 -18756 20266 -18704
rect 20534 -18756 20586 -18704
rect 20854 -18756 20906 -18704
rect 21174 -18756 21226 -18704
rect 21494 -18756 21546 -18704
rect 21814 -18756 21866 -18704
rect 22134 -18756 22186 -18704
rect 22454 -18756 22506 -18704
rect 22774 -18756 22826 -18704
rect 23094 -18756 23146 -18704
rect 23414 -18756 23466 -18704
rect 23734 -18756 23786 -18704
rect 24054 -18756 24106 -18704
rect 24374 -18756 24426 -18704
rect 24694 -18756 24746 -18704
rect 25014 -18756 25066 -18704
rect 25334 -18756 25386 -18704
rect 30614 -11300 30666 -11248
rect 30934 -11300 30986 -11248
rect 31254 -11300 31306 -11248
rect 31574 -11300 31626 -11248
rect 31894 -11300 31946 -11248
rect 32214 -11300 32266 -11248
rect 32534 -11300 32586 -11248
rect 32854 -11300 32906 -11248
rect 33174 -11300 33226 -11248
rect 33494 -11300 33546 -11248
rect 33814 -11300 33866 -11248
rect 34134 -11300 34186 -11248
rect 34454 -11300 34506 -11248
rect 34774 -11300 34826 -11248
rect 35094 -11300 35146 -11248
rect 35414 -11300 35466 -11248
rect 35734 -11300 35786 -11248
rect 36054 -11300 36106 -11248
rect 36374 -11300 36426 -11248
rect 36694 -11300 36746 -11248
rect 37014 -11300 37066 -11248
rect 37334 -11300 37386 -11248
rect 30244 -11506 30296 -11454
rect 37710 -11506 37762 -11454
rect 30244 -11826 30296 -11774
rect 30244 -12146 30296 -12094
rect 30244 -12466 30296 -12414
rect 30244 -12786 30296 -12734
rect 30244 -13106 30296 -13054
rect 30244 -13426 30296 -13374
rect 30244 -13746 30296 -13694
rect 30244 -14066 30296 -14014
rect 30244 -14386 30296 -14334
rect 30244 -14706 30296 -14654
rect 30244 -15026 30296 -14974
rect 30244 -15346 30296 -15294
rect 30244 -15666 30296 -15614
rect 30244 -15986 30296 -15934
rect 30244 -16306 30296 -16254
rect 30244 -16626 30296 -16574
rect 30244 -16946 30296 -16894
rect 30244 -17266 30296 -17214
rect 30244 -17586 30296 -17534
rect 30244 -17906 30296 -17854
rect 30244 -18226 30296 -18174
rect 37710 -11826 37762 -11774
rect 37710 -12146 37762 -12094
rect 37710 -12466 37762 -12414
rect 37710 -12786 37762 -12734
rect 37710 -13106 37762 -13054
rect 37710 -13426 37762 -13374
rect 37710 -13746 37762 -13694
rect 37710 -14066 37762 -14014
rect 37710 -14386 37762 -14334
rect 37710 -14706 37762 -14654
rect 37710 -15026 37762 -14974
rect 37710 -15346 37762 -15294
rect 37710 -15666 37762 -15614
rect 37710 -15986 37762 -15934
rect 37710 -16306 37762 -16254
rect 37710 -16626 37762 -16574
rect 37710 -16946 37762 -16894
rect 37710 -17266 37762 -17214
rect 37710 -17586 37762 -17534
rect 37710 -17906 37762 -17854
rect 37710 -18226 37762 -18174
rect 30244 -18546 30296 -18494
rect 37710 -18546 37762 -18494
rect 30614 -18756 30666 -18704
rect 30934 -18756 30986 -18704
rect 31254 -18756 31306 -18704
rect 31574 -18756 31626 -18704
rect 31894 -18756 31946 -18704
rect 32214 -18756 32266 -18704
rect 32534 -18756 32586 -18704
rect 32854 -18756 32906 -18704
rect 33174 -18756 33226 -18704
rect 33494 -18756 33546 -18704
rect 33814 -18756 33866 -18704
rect 34134 -18756 34186 -18704
rect 34454 -18756 34506 -18704
rect 34774 -18756 34826 -18704
rect 35094 -18756 35146 -18704
rect 35414 -18756 35466 -18704
rect 35734 -18756 35786 -18704
rect 36054 -18756 36106 -18704
rect 36374 -18756 36426 -18704
rect 36694 -18756 36746 -18704
rect 37014 -18756 37066 -18704
rect 37334 -18756 37386 -18704
rect 42614 -11300 42666 -11248
rect 42934 -11300 42986 -11248
rect 43254 -11300 43306 -11248
rect 43574 -11300 43626 -11248
rect 43894 -11300 43946 -11248
rect 44214 -11300 44266 -11248
rect 44534 -11300 44586 -11248
rect 44854 -11300 44906 -11248
rect 45174 -11300 45226 -11248
rect 45494 -11300 45546 -11248
rect 45814 -11300 45866 -11248
rect 46134 -11300 46186 -11248
rect 46454 -11300 46506 -11248
rect 46774 -11300 46826 -11248
rect 47094 -11300 47146 -11248
rect 47414 -11300 47466 -11248
rect 47734 -11300 47786 -11248
rect 48054 -11300 48106 -11248
rect 48374 -11300 48426 -11248
rect 48694 -11300 48746 -11248
rect 49014 -11300 49066 -11248
rect 49334 -11300 49386 -11248
rect 42247 -11506 42299 -11454
rect 49701 -11506 49753 -11454
rect 42247 -11826 42299 -11774
rect 42247 -12146 42299 -12094
rect 42247 -12466 42299 -12414
rect 42247 -12786 42299 -12734
rect 42247 -13106 42299 -13054
rect 42247 -13426 42299 -13374
rect 42247 -13746 42299 -13694
rect 42247 -14066 42299 -14014
rect 42247 -14386 42299 -14334
rect 42247 -14706 42299 -14654
rect 42247 -15026 42299 -14974
rect 42247 -15346 42299 -15294
rect 42247 -15666 42299 -15614
rect 42247 -15986 42299 -15934
rect 42247 -16306 42299 -16254
rect 42247 -16626 42299 -16574
rect 42247 -16946 42299 -16894
rect 42247 -17266 42299 -17214
rect 42247 -17586 42299 -17534
rect 42247 -17906 42299 -17854
rect 42247 -18226 42299 -18174
rect 49701 -11826 49753 -11774
rect 49701 -12146 49753 -12094
rect 49701 -12466 49753 -12414
rect 49701 -12786 49753 -12734
rect 49701 -13106 49753 -13054
rect 49701 -13426 49753 -13374
rect 49701 -13746 49753 -13694
rect 49701 -14066 49753 -14014
rect 49701 -14386 49753 -14334
rect 49701 -14706 49753 -14654
rect 49701 -15026 49753 -14974
rect 49701 -15346 49753 -15294
rect 49701 -15666 49753 -15614
rect 49701 -15986 49753 -15934
rect 49701 -16306 49753 -16254
rect 49701 -16626 49753 -16574
rect 49701 -16946 49753 -16894
rect 49701 -17266 49753 -17214
rect 49701 -17586 49753 -17534
rect 49701 -17906 49753 -17854
rect 49701 -18226 49753 -18174
rect 42247 -18546 42299 -18494
rect 49701 -18546 49753 -18494
rect 42614 -18756 42666 -18704
rect 42934 -18756 42986 -18704
rect 43254 -18756 43306 -18704
rect 43574 -18756 43626 -18704
rect 43894 -18756 43946 -18704
rect 44214 -18756 44266 -18704
rect 44534 -18756 44586 -18704
rect 44854 -18756 44906 -18704
rect 45174 -18756 45226 -18704
rect 45494 -18756 45546 -18704
rect 45814 -18756 45866 -18704
rect 46134 -18756 46186 -18704
rect 46454 -18756 46506 -18704
rect 46774 -18756 46826 -18704
rect 47094 -18756 47146 -18704
rect 47414 -18756 47466 -18704
rect 47734 -18756 47786 -18704
rect 48054 -18756 48106 -18704
rect 48374 -18756 48426 -18704
rect 48694 -18756 48746 -18704
rect 49014 -18756 49066 -18704
rect 49334 -18756 49386 -18704
<< metal2 >>
rect 20060 3280 20500 3300
rect 20060 3140 20080 3280
rect 20480 3140 20500 3280
rect 20060 3120 20500 3140
rect 20920 3280 21360 3300
rect 20920 3140 20940 3280
rect 21340 3140 21360 3280
rect 20920 3120 21360 3140
rect 15160 2940 15380 2960
rect 15160 2680 15180 2940
rect 15360 2680 15380 2940
rect 15160 2660 15380 2680
rect 13920 320 14120 340
rect 13920 -80 13940 320
rect 14100 -80 14120 320
rect 13920 -100 14120 -80
rect 14180 320 14520 340
rect 14180 -80 14200 320
rect 14500 -45 14520 320
rect 14500 -75 14690 -45
rect 14500 -80 14520 -75
rect 14180 -100 14520 -80
rect 14055 -195 14085 -100
rect 14055 -225 14479 -195
rect 14449 -445 14479 -225
rect 14390 -1100 14550 -1060
rect 14390 -1860 14430 -1100
rect 14520 -1620 14560 -1580
rect 14660 -1755 14690 -75
rect 14515 -1785 14690 -1755
rect 14390 -1880 14460 -1860
rect 14390 -1940 14400 -1880
rect 14390 -1960 14460 -1940
rect 14515 -2095 14545 -1785
rect 15300 -1840 15380 2660
rect 19980 1760 20800 1800
rect 19980 1460 20020 1760
rect 20260 1460 20800 1760
rect 19980 1420 20800 1460
rect 20780 -1220 23000 -1200
rect 20780 -1580 22820 -1220
rect 22980 -1580 23000 -1220
rect 20780 -1600 23000 -1580
rect 14600 -1920 15380 -1840
rect 20340 -1680 20660 -1640
rect 14600 -2000 14680 -1920
rect 14205 -2100 14545 -2095
rect 14200 -2125 14545 -2100
rect 14200 -2900 14400 -2125
rect 20340 -2200 20380 -1680
rect 20620 -2200 20660 -1680
rect 20340 -2240 20660 -2200
rect 20780 -2240 21000 -1600
rect 14200 -11000 14500 -2900
rect 20880 -3890 21000 -2240
rect 21280 -3060 21560 -3040
rect 21280 -3200 21300 -3060
rect 21540 -3200 21560 -3060
rect 21280 -3220 21560 -3200
rect 20880 -3960 21569 -3890
rect 21180 -4100 21420 -4080
rect 21180 -4500 21200 -4100
rect 21400 -4500 21420 -4100
rect 21180 -4520 21420 -4500
rect 20340 -4660 21240 -4620
rect 20340 -4840 20380 -4660
rect 21200 -4820 21240 -4660
rect 20280 -4860 20380 -4840
rect 20280 -4980 20300 -4860
rect 20360 -4980 20380 -4860
rect 20280 -5000 20380 -4980
rect 21180 -4860 21260 -4820
rect 21180 -5260 21260 -5220
rect 21360 -4860 21440 -4820
rect 21510 -4890 21569 -3960
rect 21440 -4920 21569 -4890
rect 21540 -4949 21569 -4920
rect 21360 -5480 21380 -5220
rect 21540 -5480 21560 -4949
rect 21360 -5500 21560 -5480
rect 6000 -11246 14000 -11000
rect 6000 -11302 6612 -11246
rect 6668 -11302 6932 -11246
rect 6988 -11302 7252 -11246
rect 7308 -11302 7572 -11246
rect 7628 -11302 7892 -11246
rect 7948 -11302 8212 -11246
rect 8268 -11302 8532 -11246
rect 8588 -11302 8852 -11246
rect 8908 -11302 9172 -11246
rect 9228 -11302 9492 -11246
rect 9548 -11302 9812 -11246
rect 9868 -11302 10132 -11246
rect 10188 -11302 10452 -11246
rect 10508 -11302 10772 -11246
rect 10828 -11302 11092 -11246
rect 11148 -11302 11412 -11246
rect 11468 -11302 11732 -11246
rect 11788 -11302 12052 -11246
rect 12108 -11302 12372 -11246
rect 12428 -11302 12692 -11246
rect 12748 -11302 13012 -11246
rect 13068 -11302 13332 -11246
rect 13388 -11302 14000 -11246
rect 6000 -11452 14000 -11302
rect 6000 -11508 6242 -11452
rect 6298 -11508 13708 -11452
rect 13764 -11508 14000 -11452
rect 6000 -11540 14000 -11508
rect 14180 -11100 14520 -11000
rect 14180 -11500 14200 -11100
rect 14500 -11500 14520 -11100
rect 14180 -11520 14520 -11500
rect 18000 -11246 26000 -11000
rect 18000 -11302 18612 -11246
rect 18668 -11302 18932 -11246
rect 18988 -11302 19252 -11246
rect 19308 -11302 19572 -11246
rect 19628 -11302 19892 -11246
rect 19948 -11302 20212 -11246
rect 20268 -11302 20532 -11246
rect 20588 -11302 20852 -11246
rect 20908 -11302 21172 -11246
rect 21228 -11302 21492 -11246
rect 21548 -11302 21812 -11246
rect 21868 -11302 22132 -11246
rect 22188 -11302 22452 -11246
rect 22508 -11302 22772 -11246
rect 22828 -11302 23092 -11246
rect 23148 -11302 23412 -11246
rect 23468 -11302 23732 -11246
rect 23788 -11302 24052 -11246
rect 24108 -11302 24372 -11246
rect 24428 -11302 24692 -11246
rect 24748 -11302 25012 -11246
rect 25068 -11302 25332 -11246
rect 25388 -11302 26000 -11246
rect 18000 -11452 26000 -11302
rect 18000 -11508 18242 -11452
rect 18298 -11508 25708 -11452
rect 25764 -11508 26000 -11452
rect 6000 -11772 6540 -11540
rect 6000 -11828 6242 -11772
rect 6298 -11828 6540 -11772
rect 6000 -12092 6540 -11828
rect 6000 -12148 6242 -12092
rect 6298 -12148 6540 -12092
rect 6000 -12412 6540 -12148
rect 6000 -12468 6242 -12412
rect 6298 -12468 6540 -12412
rect 6000 -12732 6540 -12468
rect 6000 -12788 6242 -12732
rect 6298 -12788 6540 -12732
rect 6000 -13052 6540 -12788
rect 6000 -13108 6242 -13052
rect 6298 -13108 6540 -13052
rect 6000 -13372 6540 -13108
rect 6000 -13428 6242 -13372
rect 6298 -13428 6540 -13372
rect 6000 -13692 6540 -13428
rect 6000 -13748 6242 -13692
rect 6298 -13748 6540 -13692
rect 6000 -14012 6540 -13748
rect 6000 -14068 6242 -14012
rect 6298 -14068 6540 -14012
rect 6000 -14332 6540 -14068
rect 6000 -14388 6242 -14332
rect 6298 -14388 6540 -14332
rect 6000 -14652 6540 -14388
rect 6000 -14708 6242 -14652
rect 6298 -14708 6540 -14652
rect 6000 -14972 6540 -14708
rect 6000 -15028 6242 -14972
rect 6298 -15028 6540 -14972
rect 6000 -15292 6540 -15028
rect 6000 -15348 6242 -15292
rect 6298 -15348 6540 -15292
rect 6000 -15612 6540 -15348
rect 6000 -15668 6242 -15612
rect 6298 -15668 6540 -15612
rect 6000 -15932 6540 -15668
rect 6000 -15988 6242 -15932
rect 6298 -15988 6540 -15932
rect 6000 -16252 6540 -15988
rect 6000 -16308 6242 -16252
rect 6298 -16308 6540 -16252
rect 6000 -16572 6540 -16308
rect 6000 -16628 6242 -16572
rect 6298 -16628 6540 -16572
rect 6000 -16892 6540 -16628
rect 6000 -16948 6242 -16892
rect 6298 -16948 6540 -16892
rect 6000 -17212 6540 -16948
rect 6000 -17268 6242 -17212
rect 6298 -17268 6540 -17212
rect 6000 -17532 6540 -17268
rect 6000 -17588 6242 -17532
rect 6298 -17588 6540 -17532
rect 6000 -17852 6540 -17588
rect 6000 -17908 6242 -17852
rect 6298 -17908 6540 -17852
rect 6000 -18172 6540 -17908
rect 6000 -18228 6242 -18172
rect 6298 -18228 6540 -18172
rect 6000 -18460 6540 -18228
rect 13460 -11772 14000 -11540
rect 13460 -11828 13708 -11772
rect 13764 -11828 14000 -11772
rect 13460 -12092 14000 -11828
rect 13460 -12148 13708 -12092
rect 13764 -12148 14000 -12092
rect 13460 -12412 14000 -12148
rect 13460 -12468 13708 -12412
rect 13764 -12468 14000 -12412
rect 13460 -12732 14000 -12468
rect 13460 -12788 13708 -12732
rect 13764 -12788 14000 -12732
rect 13460 -13052 14000 -12788
rect 13460 -13108 13708 -13052
rect 13764 -13108 14000 -13052
rect 13460 -13372 14000 -13108
rect 13460 -13428 13708 -13372
rect 13764 -13428 14000 -13372
rect 13460 -13692 14000 -13428
rect 13460 -13748 13708 -13692
rect 13764 -13748 14000 -13692
rect 13460 -14012 14000 -13748
rect 13460 -14068 13708 -14012
rect 13764 -14068 14000 -14012
rect 13460 -14332 14000 -14068
rect 13460 -14388 13708 -14332
rect 13764 -14388 14000 -14332
rect 13460 -14652 14000 -14388
rect 13460 -14708 13708 -14652
rect 13764 -14708 14000 -14652
rect 13460 -14972 14000 -14708
rect 13460 -15028 13708 -14972
rect 13764 -15028 14000 -14972
rect 13460 -15292 14000 -15028
rect 13460 -15348 13708 -15292
rect 13764 -15348 14000 -15292
rect 13460 -15612 14000 -15348
rect 13460 -15668 13708 -15612
rect 13764 -15668 14000 -15612
rect 13460 -15932 14000 -15668
rect 13460 -15988 13708 -15932
rect 13764 -15988 14000 -15932
rect 13460 -16252 14000 -15988
rect 13460 -16308 13708 -16252
rect 13764 -16308 14000 -16252
rect 13460 -16572 14000 -16308
rect 13460 -16628 13708 -16572
rect 13764 -16628 14000 -16572
rect 13460 -16892 14000 -16628
rect 13460 -16948 13708 -16892
rect 13764 -16948 14000 -16892
rect 13460 -17212 14000 -16948
rect 13460 -17268 13708 -17212
rect 13764 -17268 14000 -17212
rect 13460 -17532 14000 -17268
rect 13460 -17588 13708 -17532
rect 13764 -17588 14000 -17532
rect 13460 -17852 14000 -17588
rect 13460 -17908 13708 -17852
rect 13764 -17908 14000 -17852
rect 13460 -18172 14000 -17908
rect 13460 -18228 13708 -18172
rect 13764 -18228 14000 -18172
rect 13460 -18460 14000 -18228
rect 6000 -18492 14000 -18460
rect 6000 -18548 6242 -18492
rect 6298 -18548 13708 -18492
rect 13764 -18548 14000 -18492
rect 6000 -18702 14000 -18548
rect 6000 -18758 6612 -18702
rect 6668 -18758 6932 -18702
rect 6988 -18758 7252 -18702
rect 7308 -18758 7572 -18702
rect 7628 -18758 7892 -18702
rect 7948 -18758 8212 -18702
rect 8268 -18758 8532 -18702
rect 8588 -18758 8852 -18702
rect 8908 -18758 9172 -18702
rect 9228 -18758 9492 -18702
rect 9548 -18758 9812 -18702
rect 9868 -18758 10132 -18702
rect 10188 -18758 10452 -18702
rect 10508 -18758 10772 -18702
rect 10828 -18758 11092 -18702
rect 11148 -18758 11412 -18702
rect 11468 -18758 11732 -18702
rect 11788 -18758 12052 -18702
rect 12108 -18758 12372 -18702
rect 12428 -18758 12692 -18702
rect 12748 -18758 13012 -18702
rect 13068 -18758 13332 -18702
rect 13388 -18758 14000 -18702
rect 6000 -19000 14000 -18758
rect 18000 -11540 26000 -11508
rect 18000 -11772 18540 -11540
rect 18000 -11828 18242 -11772
rect 18298 -11828 18540 -11772
rect 18000 -12092 18540 -11828
rect 18000 -12148 18242 -12092
rect 18298 -12148 18540 -12092
rect 18000 -12412 18540 -12148
rect 18000 -12468 18242 -12412
rect 18298 -12468 18540 -12412
rect 18000 -12732 18540 -12468
rect 18000 -12788 18242 -12732
rect 18298 -12788 18540 -12732
rect 18000 -13052 18540 -12788
rect 18000 -13108 18242 -13052
rect 18298 -13108 18540 -13052
rect 18000 -13372 18540 -13108
rect 18000 -13428 18242 -13372
rect 18298 -13428 18540 -13372
rect 18000 -13692 18540 -13428
rect 18000 -13748 18242 -13692
rect 18298 -13748 18540 -13692
rect 18000 -14012 18540 -13748
rect 18000 -14068 18242 -14012
rect 18298 -14068 18540 -14012
rect 18000 -14332 18540 -14068
rect 18000 -14388 18242 -14332
rect 18298 -14388 18540 -14332
rect 18000 -14652 18540 -14388
rect 18000 -14708 18242 -14652
rect 18298 -14708 18540 -14652
rect 18000 -14972 18540 -14708
rect 18000 -15028 18242 -14972
rect 18298 -15028 18540 -14972
rect 18000 -15292 18540 -15028
rect 18000 -15348 18242 -15292
rect 18298 -15348 18540 -15292
rect 18000 -15612 18540 -15348
rect 18000 -15668 18242 -15612
rect 18298 -15668 18540 -15612
rect 18000 -15932 18540 -15668
rect 18000 -15988 18242 -15932
rect 18298 -15988 18540 -15932
rect 18000 -16252 18540 -15988
rect 18000 -16308 18242 -16252
rect 18298 -16308 18540 -16252
rect 18000 -16572 18540 -16308
rect 18000 -16628 18242 -16572
rect 18298 -16628 18540 -16572
rect 18000 -16892 18540 -16628
rect 18000 -16948 18242 -16892
rect 18298 -16948 18540 -16892
rect 18000 -17212 18540 -16948
rect 18000 -17268 18242 -17212
rect 18298 -17268 18540 -17212
rect 18000 -17532 18540 -17268
rect 18000 -17588 18242 -17532
rect 18298 -17588 18540 -17532
rect 18000 -17852 18540 -17588
rect 18000 -17908 18242 -17852
rect 18298 -17908 18540 -17852
rect 18000 -18172 18540 -17908
rect 18000 -18228 18242 -18172
rect 18298 -18228 18540 -18172
rect 18000 -18460 18540 -18228
rect 25460 -11772 26000 -11540
rect 25460 -11828 25708 -11772
rect 25764 -11828 26000 -11772
rect 25460 -12092 26000 -11828
rect 25460 -12148 25708 -12092
rect 25764 -12148 26000 -12092
rect 25460 -12412 26000 -12148
rect 25460 -12468 25708 -12412
rect 25764 -12468 26000 -12412
rect 25460 -12732 26000 -12468
rect 25460 -12788 25708 -12732
rect 25764 -12788 26000 -12732
rect 25460 -13052 26000 -12788
rect 25460 -13108 25708 -13052
rect 25764 -13108 26000 -13052
rect 25460 -13372 26000 -13108
rect 25460 -13428 25708 -13372
rect 25764 -13428 26000 -13372
rect 25460 -13692 26000 -13428
rect 25460 -13748 25708 -13692
rect 25764 -13748 26000 -13692
rect 25460 -14012 26000 -13748
rect 25460 -14068 25708 -14012
rect 25764 -14068 26000 -14012
rect 25460 -14332 26000 -14068
rect 25460 -14388 25708 -14332
rect 25764 -14388 26000 -14332
rect 25460 -14652 26000 -14388
rect 25460 -14708 25708 -14652
rect 25764 -14708 26000 -14652
rect 25460 -14972 26000 -14708
rect 25460 -15028 25708 -14972
rect 25764 -15028 26000 -14972
rect 25460 -15292 26000 -15028
rect 25460 -15348 25708 -15292
rect 25764 -15348 26000 -15292
rect 25460 -15612 26000 -15348
rect 25460 -15668 25708 -15612
rect 25764 -15668 26000 -15612
rect 25460 -15932 26000 -15668
rect 25460 -15988 25708 -15932
rect 25764 -15988 26000 -15932
rect 25460 -16252 26000 -15988
rect 25460 -16308 25708 -16252
rect 25764 -16308 26000 -16252
rect 25460 -16572 26000 -16308
rect 25460 -16628 25708 -16572
rect 25764 -16628 26000 -16572
rect 25460 -16892 26000 -16628
rect 25460 -16948 25708 -16892
rect 25764 -16948 26000 -16892
rect 25460 -17212 26000 -16948
rect 25460 -17268 25708 -17212
rect 25764 -17268 26000 -17212
rect 25460 -17532 26000 -17268
rect 25460 -17588 25708 -17532
rect 25764 -17588 26000 -17532
rect 25460 -17852 26000 -17588
rect 25460 -17908 25708 -17852
rect 25764 -17908 26000 -17852
rect 25460 -18172 26000 -17908
rect 25460 -18228 25708 -18172
rect 25764 -18228 26000 -18172
rect 25460 -18460 26000 -18228
rect 18000 -18492 26000 -18460
rect 18000 -18548 18242 -18492
rect 18298 -18548 25708 -18492
rect 25764 -18548 26000 -18492
rect 18000 -18702 26000 -18548
rect 18000 -18758 18612 -18702
rect 18668 -18758 18932 -18702
rect 18988 -18758 19252 -18702
rect 19308 -18758 19572 -18702
rect 19628 -18758 19892 -18702
rect 19948 -18758 20212 -18702
rect 20268 -18758 20532 -18702
rect 20588 -18758 20852 -18702
rect 20908 -18758 21172 -18702
rect 21228 -18758 21492 -18702
rect 21548 -18758 21812 -18702
rect 21868 -18758 22132 -18702
rect 22188 -18758 22452 -18702
rect 22508 -18758 22772 -18702
rect 22828 -18758 23092 -18702
rect 23148 -18758 23412 -18702
rect 23468 -18758 23732 -18702
rect 23788 -18758 24052 -18702
rect 24108 -18758 24372 -18702
rect 24428 -18758 24692 -18702
rect 24748 -18758 25012 -18702
rect 25068 -18758 25332 -18702
rect 25388 -18758 26000 -18702
rect 18000 -19000 26000 -18758
rect 30000 -11246 38000 -11000
rect 30000 -11302 30612 -11246
rect 30668 -11302 30932 -11246
rect 30988 -11302 31252 -11246
rect 31308 -11302 31572 -11246
rect 31628 -11302 31892 -11246
rect 31948 -11302 32212 -11246
rect 32268 -11302 32532 -11246
rect 32588 -11302 32852 -11246
rect 32908 -11302 33172 -11246
rect 33228 -11302 33492 -11246
rect 33548 -11302 33812 -11246
rect 33868 -11302 34132 -11246
rect 34188 -11302 34452 -11246
rect 34508 -11302 34772 -11246
rect 34828 -11302 35092 -11246
rect 35148 -11302 35412 -11246
rect 35468 -11302 35732 -11246
rect 35788 -11302 36052 -11246
rect 36108 -11302 36372 -11246
rect 36428 -11302 36692 -11246
rect 36748 -11302 37012 -11246
rect 37068 -11302 37332 -11246
rect 37388 -11302 38000 -11246
rect 30000 -11452 38000 -11302
rect 30000 -11508 30242 -11452
rect 30298 -11508 37708 -11452
rect 37764 -11508 38000 -11452
rect 30000 -11540 38000 -11508
rect 30000 -11772 30540 -11540
rect 30000 -11828 30242 -11772
rect 30298 -11828 30540 -11772
rect 30000 -12092 30540 -11828
rect 30000 -12148 30242 -12092
rect 30298 -12148 30540 -12092
rect 30000 -12412 30540 -12148
rect 30000 -12468 30242 -12412
rect 30298 -12468 30540 -12412
rect 30000 -12732 30540 -12468
rect 30000 -12788 30242 -12732
rect 30298 -12788 30540 -12732
rect 30000 -13052 30540 -12788
rect 30000 -13108 30242 -13052
rect 30298 -13108 30540 -13052
rect 30000 -13372 30540 -13108
rect 30000 -13428 30242 -13372
rect 30298 -13428 30540 -13372
rect 30000 -13692 30540 -13428
rect 30000 -13748 30242 -13692
rect 30298 -13748 30540 -13692
rect 30000 -14012 30540 -13748
rect 30000 -14068 30242 -14012
rect 30298 -14068 30540 -14012
rect 30000 -14332 30540 -14068
rect 30000 -14388 30242 -14332
rect 30298 -14388 30540 -14332
rect 30000 -14652 30540 -14388
rect 30000 -14708 30242 -14652
rect 30298 -14708 30540 -14652
rect 30000 -14972 30540 -14708
rect 30000 -15028 30242 -14972
rect 30298 -15028 30540 -14972
rect 30000 -15292 30540 -15028
rect 30000 -15348 30242 -15292
rect 30298 -15348 30540 -15292
rect 30000 -15612 30540 -15348
rect 30000 -15668 30242 -15612
rect 30298 -15668 30540 -15612
rect 30000 -15932 30540 -15668
rect 30000 -15988 30242 -15932
rect 30298 -15988 30540 -15932
rect 30000 -16252 30540 -15988
rect 30000 -16308 30242 -16252
rect 30298 -16308 30540 -16252
rect 30000 -16572 30540 -16308
rect 30000 -16628 30242 -16572
rect 30298 -16628 30540 -16572
rect 30000 -16892 30540 -16628
rect 30000 -16948 30242 -16892
rect 30298 -16948 30540 -16892
rect 30000 -17212 30540 -16948
rect 30000 -17268 30242 -17212
rect 30298 -17268 30540 -17212
rect 30000 -17532 30540 -17268
rect 30000 -17588 30242 -17532
rect 30298 -17588 30540 -17532
rect 30000 -17852 30540 -17588
rect 30000 -17908 30242 -17852
rect 30298 -17908 30540 -17852
rect 30000 -18172 30540 -17908
rect 30000 -18228 30242 -18172
rect 30298 -18228 30540 -18172
rect 30000 -18460 30540 -18228
rect 37460 -11772 38000 -11540
rect 37460 -11828 37708 -11772
rect 37764 -11828 38000 -11772
rect 37460 -12092 38000 -11828
rect 37460 -12148 37708 -12092
rect 37764 -12148 38000 -12092
rect 37460 -12412 38000 -12148
rect 37460 -12468 37708 -12412
rect 37764 -12468 38000 -12412
rect 37460 -12732 38000 -12468
rect 37460 -12788 37708 -12732
rect 37764 -12788 38000 -12732
rect 37460 -13052 38000 -12788
rect 37460 -13108 37708 -13052
rect 37764 -13108 38000 -13052
rect 37460 -13372 38000 -13108
rect 37460 -13428 37708 -13372
rect 37764 -13428 38000 -13372
rect 37460 -13692 38000 -13428
rect 37460 -13748 37708 -13692
rect 37764 -13748 38000 -13692
rect 37460 -14012 38000 -13748
rect 37460 -14068 37708 -14012
rect 37764 -14068 38000 -14012
rect 37460 -14332 38000 -14068
rect 37460 -14388 37708 -14332
rect 37764 -14388 38000 -14332
rect 37460 -14652 38000 -14388
rect 37460 -14708 37708 -14652
rect 37764 -14708 38000 -14652
rect 37460 -14972 38000 -14708
rect 37460 -15028 37708 -14972
rect 37764 -15028 38000 -14972
rect 37460 -15292 38000 -15028
rect 37460 -15348 37708 -15292
rect 37764 -15348 38000 -15292
rect 37460 -15612 38000 -15348
rect 37460 -15668 37708 -15612
rect 37764 -15668 38000 -15612
rect 37460 -15932 38000 -15668
rect 37460 -15988 37708 -15932
rect 37764 -15988 38000 -15932
rect 37460 -16252 38000 -15988
rect 37460 -16308 37708 -16252
rect 37764 -16308 38000 -16252
rect 37460 -16572 38000 -16308
rect 37460 -16628 37708 -16572
rect 37764 -16628 38000 -16572
rect 37460 -16892 38000 -16628
rect 37460 -16948 37708 -16892
rect 37764 -16948 38000 -16892
rect 37460 -17212 38000 -16948
rect 37460 -17268 37708 -17212
rect 37764 -17268 38000 -17212
rect 37460 -17532 38000 -17268
rect 37460 -17588 37708 -17532
rect 37764 -17588 38000 -17532
rect 37460 -17852 38000 -17588
rect 37460 -17908 37708 -17852
rect 37764 -17908 38000 -17852
rect 37460 -18172 38000 -17908
rect 37460 -18228 37708 -18172
rect 37764 -18228 38000 -18172
rect 37460 -18460 38000 -18228
rect 30000 -18492 38000 -18460
rect 30000 -18548 30242 -18492
rect 30298 -18548 37708 -18492
rect 37764 -18548 38000 -18492
rect 30000 -18702 38000 -18548
rect 30000 -18758 30612 -18702
rect 30668 -18758 30932 -18702
rect 30988 -18758 31252 -18702
rect 31308 -18758 31572 -18702
rect 31628 -18758 31892 -18702
rect 31948 -18758 32212 -18702
rect 32268 -18758 32532 -18702
rect 32588 -18758 32852 -18702
rect 32908 -18758 33172 -18702
rect 33228 -18758 33492 -18702
rect 33548 -18758 33812 -18702
rect 33868 -18758 34132 -18702
rect 34188 -18758 34452 -18702
rect 34508 -18758 34772 -18702
rect 34828 -18758 35092 -18702
rect 35148 -18758 35412 -18702
rect 35468 -18758 35732 -18702
rect 35788 -18758 36052 -18702
rect 36108 -18758 36372 -18702
rect 36428 -18758 36692 -18702
rect 36748 -18758 37012 -18702
rect 37068 -18758 37332 -18702
rect 37388 -18758 38000 -18702
rect 30000 -19000 38000 -18758
rect 42000 -11246 50000 -11000
rect 42000 -11302 42612 -11246
rect 42668 -11302 42932 -11246
rect 42988 -11302 43252 -11246
rect 43308 -11302 43572 -11246
rect 43628 -11302 43892 -11246
rect 43948 -11302 44212 -11246
rect 44268 -11302 44532 -11246
rect 44588 -11302 44852 -11246
rect 44908 -11302 45172 -11246
rect 45228 -11302 45492 -11246
rect 45548 -11302 45812 -11246
rect 45868 -11302 46132 -11246
rect 46188 -11302 46452 -11246
rect 46508 -11302 46772 -11246
rect 46828 -11302 47092 -11246
rect 47148 -11302 47412 -11246
rect 47468 -11302 47732 -11246
rect 47788 -11302 48052 -11246
rect 48108 -11302 48372 -11246
rect 48428 -11302 48692 -11246
rect 48748 -11302 49012 -11246
rect 49068 -11302 49332 -11246
rect 49388 -11302 50000 -11246
rect 42000 -11452 50000 -11302
rect 42000 -11508 42245 -11452
rect 42301 -11508 49699 -11452
rect 49755 -11508 50000 -11452
rect 42000 -11540 50000 -11508
rect 42000 -11772 42540 -11540
rect 42000 -11828 42245 -11772
rect 42301 -11828 42540 -11772
rect 42000 -12092 42540 -11828
rect 42000 -12148 42245 -12092
rect 42301 -12148 42540 -12092
rect 42000 -12412 42540 -12148
rect 42000 -12468 42245 -12412
rect 42301 -12468 42540 -12412
rect 42000 -12732 42540 -12468
rect 42000 -12788 42245 -12732
rect 42301 -12788 42540 -12732
rect 42000 -13052 42540 -12788
rect 42000 -13108 42245 -13052
rect 42301 -13108 42540 -13052
rect 42000 -13372 42540 -13108
rect 42000 -13428 42245 -13372
rect 42301 -13428 42540 -13372
rect 42000 -13692 42540 -13428
rect 42000 -13748 42245 -13692
rect 42301 -13748 42540 -13692
rect 42000 -14012 42540 -13748
rect 42000 -14068 42245 -14012
rect 42301 -14068 42540 -14012
rect 42000 -14332 42540 -14068
rect 42000 -14388 42245 -14332
rect 42301 -14388 42540 -14332
rect 42000 -14652 42540 -14388
rect 42000 -14708 42245 -14652
rect 42301 -14708 42540 -14652
rect 42000 -14972 42540 -14708
rect 42000 -15028 42245 -14972
rect 42301 -15028 42540 -14972
rect 42000 -15292 42540 -15028
rect 42000 -15348 42245 -15292
rect 42301 -15348 42540 -15292
rect 42000 -15612 42540 -15348
rect 42000 -15668 42245 -15612
rect 42301 -15668 42540 -15612
rect 42000 -15932 42540 -15668
rect 42000 -15988 42245 -15932
rect 42301 -15988 42540 -15932
rect 42000 -16252 42540 -15988
rect 42000 -16308 42245 -16252
rect 42301 -16308 42540 -16252
rect 42000 -16572 42540 -16308
rect 42000 -16628 42245 -16572
rect 42301 -16628 42540 -16572
rect 42000 -16892 42540 -16628
rect 42000 -16948 42245 -16892
rect 42301 -16948 42540 -16892
rect 42000 -17212 42540 -16948
rect 42000 -17268 42245 -17212
rect 42301 -17268 42540 -17212
rect 42000 -17532 42540 -17268
rect 42000 -17588 42245 -17532
rect 42301 -17588 42540 -17532
rect 42000 -17852 42540 -17588
rect 42000 -17908 42245 -17852
rect 42301 -17908 42540 -17852
rect 42000 -18172 42540 -17908
rect 42000 -18228 42245 -18172
rect 42301 -18228 42540 -18172
rect 42000 -18460 42540 -18228
rect 49460 -11772 50000 -11540
rect 49460 -11828 49699 -11772
rect 49755 -11828 50000 -11772
rect 49460 -12092 50000 -11828
rect 49460 -12148 49699 -12092
rect 49755 -12148 50000 -12092
rect 49460 -12412 50000 -12148
rect 49460 -12468 49699 -12412
rect 49755 -12468 50000 -12412
rect 49460 -12732 50000 -12468
rect 49460 -12788 49699 -12732
rect 49755 -12788 50000 -12732
rect 49460 -13052 50000 -12788
rect 49460 -13108 49699 -13052
rect 49755 -13108 50000 -13052
rect 49460 -13372 50000 -13108
rect 49460 -13428 49699 -13372
rect 49755 -13428 50000 -13372
rect 49460 -13692 50000 -13428
rect 49460 -13748 49699 -13692
rect 49755 -13748 50000 -13692
rect 49460 -14012 50000 -13748
rect 49460 -14068 49699 -14012
rect 49755 -14068 50000 -14012
rect 49460 -14332 50000 -14068
rect 49460 -14388 49699 -14332
rect 49755 -14388 50000 -14332
rect 49460 -14652 50000 -14388
rect 49460 -14708 49699 -14652
rect 49755 -14708 50000 -14652
rect 49460 -14972 50000 -14708
rect 49460 -15028 49699 -14972
rect 49755 -15028 50000 -14972
rect 49460 -15292 50000 -15028
rect 49460 -15348 49699 -15292
rect 49755 -15348 50000 -15292
rect 49460 -15612 50000 -15348
rect 49460 -15668 49699 -15612
rect 49755 -15668 50000 -15612
rect 49460 -15932 50000 -15668
rect 49460 -15988 49699 -15932
rect 49755 -15988 50000 -15932
rect 49460 -16252 50000 -15988
rect 49460 -16308 49699 -16252
rect 49755 -16308 50000 -16252
rect 49460 -16572 50000 -16308
rect 49460 -16628 49699 -16572
rect 49755 -16628 50000 -16572
rect 49460 -16892 50000 -16628
rect 49460 -16948 49699 -16892
rect 49755 -16948 50000 -16892
rect 49460 -17212 50000 -16948
rect 49460 -17268 49699 -17212
rect 49755 -17268 50000 -17212
rect 49460 -17532 50000 -17268
rect 49460 -17588 49699 -17532
rect 49755 -17588 50000 -17532
rect 49460 -17852 50000 -17588
rect 49460 -17908 49699 -17852
rect 49755 -17908 50000 -17852
rect 49460 -18172 50000 -17908
rect 49460 -18228 49699 -18172
rect 49755 -18228 50000 -18172
rect 49460 -18460 50000 -18228
rect 42000 -18492 50000 -18460
rect 42000 -18548 42245 -18492
rect 42301 -18548 49699 -18492
rect 49755 -18548 50000 -18492
rect 42000 -18702 50000 -18548
rect 42000 -18758 42612 -18702
rect 42668 -18758 42932 -18702
rect 42988 -18758 43252 -18702
rect 43308 -18758 43572 -18702
rect 43628 -18758 43892 -18702
rect 43948 -18758 44212 -18702
rect 44268 -18758 44532 -18702
rect 44588 -18758 44852 -18702
rect 44908 -18758 45172 -18702
rect 45228 -18758 45492 -18702
rect 45548 -18758 45812 -18702
rect 45868 -18758 46132 -18702
rect 46188 -18758 46452 -18702
rect 46508 -18758 46772 -18702
rect 46828 -18758 47092 -18702
rect 47148 -18758 47412 -18702
rect 47468 -18758 47732 -18702
rect 47788 -18758 48052 -18702
rect 48108 -18758 48372 -18702
rect 48428 -18758 48692 -18702
rect 48748 -18758 49012 -18702
rect 49068 -18758 49332 -18702
rect 49388 -18758 50000 -18702
rect 42000 -19000 50000 -18758
rect 14200 -19400 15000 -19300
rect 14200 -19700 14300 -19400
rect 14900 -19700 15000 -19400
rect 14200 -19800 15000 -19700
<< via2 >>
rect 20080 3260 20480 3280
rect 20080 3160 20100 3260
rect 20100 3160 20460 3260
rect 20460 3160 20480 3260
rect 20080 3140 20480 3160
rect 20940 3140 21340 3280
rect 15180 2680 15360 2940
rect 13940 -80 14100 320
rect 14200 -80 14500 320
rect 20020 1460 20260 1760
rect 22820 -1580 22980 -1220
rect 20380 -2200 20620 -1680
rect 21300 -3200 21540 -3060
rect 21200 -4500 21400 -4100
rect 20300 -4980 20360 -4860
rect 21380 -5220 21440 -4920
rect 21440 -5220 21540 -4920
rect 21380 -5480 21540 -5220
rect 6612 -11248 6668 -11246
rect 6612 -11300 6614 -11248
rect 6614 -11300 6666 -11248
rect 6666 -11300 6668 -11248
rect 6612 -11302 6668 -11300
rect 6932 -11248 6988 -11246
rect 6932 -11300 6934 -11248
rect 6934 -11300 6986 -11248
rect 6986 -11300 6988 -11248
rect 6932 -11302 6988 -11300
rect 7252 -11248 7308 -11246
rect 7252 -11300 7254 -11248
rect 7254 -11300 7306 -11248
rect 7306 -11300 7308 -11248
rect 7252 -11302 7308 -11300
rect 7572 -11248 7628 -11246
rect 7572 -11300 7574 -11248
rect 7574 -11300 7626 -11248
rect 7626 -11300 7628 -11248
rect 7572 -11302 7628 -11300
rect 7892 -11248 7948 -11246
rect 7892 -11300 7894 -11248
rect 7894 -11300 7946 -11248
rect 7946 -11300 7948 -11248
rect 7892 -11302 7948 -11300
rect 8212 -11248 8268 -11246
rect 8212 -11300 8214 -11248
rect 8214 -11300 8266 -11248
rect 8266 -11300 8268 -11248
rect 8212 -11302 8268 -11300
rect 8532 -11248 8588 -11246
rect 8532 -11300 8534 -11248
rect 8534 -11300 8586 -11248
rect 8586 -11300 8588 -11248
rect 8532 -11302 8588 -11300
rect 8852 -11248 8908 -11246
rect 8852 -11300 8854 -11248
rect 8854 -11300 8906 -11248
rect 8906 -11300 8908 -11248
rect 8852 -11302 8908 -11300
rect 9172 -11248 9228 -11246
rect 9172 -11300 9174 -11248
rect 9174 -11300 9226 -11248
rect 9226 -11300 9228 -11248
rect 9172 -11302 9228 -11300
rect 9492 -11248 9548 -11246
rect 9492 -11300 9494 -11248
rect 9494 -11300 9546 -11248
rect 9546 -11300 9548 -11248
rect 9492 -11302 9548 -11300
rect 9812 -11248 9868 -11246
rect 9812 -11300 9814 -11248
rect 9814 -11300 9866 -11248
rect 9866 -11300 9868 -11248
rect 9812 -11302 9868 -11300
rect 10132 -11248 10188 -11246
rect 10132 -11300 10134 -11248
rect 10134 -11300 10186 -11248
rect 10186 -11300 10188 -11248
rect 10132 -11302 10188 -11300
rect 10452 -11248 10508 -11246
rect 10452 -11300 10454 -11248
rect 10454 -11300 10506 -11248
rect 10506 -11300 10508 -11248
rect 10452 -11302 10508 -11300
rect 10772 -11248 10828 -11246
rect 10772 -11300 10774 -11248
rect 10774 -11300 10826 -11248
rect 10826 -11300 10828 -11248
rect 10772 -11302 10828 -11300
rect 11092 -11248 11148 -11246
rect 11092 -11300 11094 -11248
rect 11094 -11300 11146 -11248
rect 11146 -11300 11148 -11248
rect 11092 -11302 11148 -11300
rect 11412 -11248 11468 -11246
rect 11412 -11300 11414 -11248
rect 11414 -11300 11466 -11248
rect 11466 -11300 11468 -11248
rect 11412 -11302 11468 -11300
rect 11732 -11248 11788 -11246
rect 11732 -11300 11734 -11248
rect 11734 -11300 11786 -11248
rect 11786 -11300 11788 -11248
rect 11732 -11302 11788 -11300
rect 12052 -11248 12108 -11246
rect 12052 -11300 12054 -11248
rect 12054 -11300 12106 -11248
rect 12106 -11300 12108 -11248
rect 12052 -11302 12108 -11300
rect 12372 -11248 12428 -11246
rect 12372 -11300 12374 -11248
rect 12374 -11300 12426 -11248
rect 12426 -11300 12428 -11248
rect 12372 -11302 12428 -11300
rect 12692 -11248 12748 -11246
rect 12692 -11300 12694 -11248
rect 12694 -11300 12746 -11248
rect 12746 -11300 12748 -11248
rect 12692 -11302 12748 -11300
rect 13012 -11248 13068 -11246
rect 13012 -11300 13014 -11248
rect 13014 -11300 13066 -11248
rect 13066 -11300 13068 -11248
rect 13012 -11302 13068 -11300
rect 13332 -11248 13388 -11246
rect 13332 -11300 13334 -11248
rect 13334 -11300 13386 -11248
rect 13386 -11300 13388 -11248
rect 13332 -11302 13388 -11300
rect 6242 -11454 6298 -11452
rect 6242 -11506 6244 -11454
rect 6244 -11506 6296 -11454
rect 6296 -11506 6298 -11454
rect 6242 -11508 6298 -11506
rect 13708 -11454 13764 -11452
rect 13708 -11506 13710 -11454
rect 13710 -11506 13762 -11454
rect 13762 -11506 13764 -11454
rect 13708 -11508 13764 -11506
rect 14200 -11500 14500 -11100
rect 18612 -11248 18668 -11246
rect 18612 -11300 18614 -11248
rect 18614 -11300 18666 -11248
rect 18666 -11300 18668 -11248
rect 18612 -11302 18668 -11300
rect 18932 -11248 18988 -11246
rect 18932 -11300 18934 -11248
rect 18934 -11300 18986 -11248
rect 18986 -11300 18988 -11248
rect 18932 -11302 18988 -11300
rect 19252 -11248 19308 -11246
rect 19252 -11300 19254 -11248
rect 19254 -11300 19306 -11248
rect 19306 -11300 19308 -11248
rect 19252 -11302 19308 -11300
rect 19572 -11248 19628 -11246
rect 19572 -11300 19574 -11248
rect 19574 -11300 19626 -11248
rect 19626 -11300 19628 -11248
rect 19572 -11302 19628 -11300
rect 19892 -11248 19948 -11246
rect 19892 -11300 19894 -11248
rect 19894 -11300 19946 -11248
rect 19946 -11300 19948 -11248
rect 19892 -11302 19948 -11300
rect 20212 -11248 20268 -11246
rect 20212 -11300 20214 -11248
rect 20214 -11300 20266 -11248
rect 20266 -11300 20268 -11248
rect 20212 -11302 20268 -11300
rect 20532 -11248 20588 -11246
rect 20532 -11300 20534 -11248
rect 20534 -11300 20586 -11248
rect 20586 -11300 20588 -11248
rect 20532 -11302 20588 -11300
rect 20852 -11248 20908 -11246
rect 20852 -11300 20854 -11248
rect 20854 -11300 20906 -11248
rect 20906 -11300 20908 -11248
rect 20852 -11302 20908 -11300
rect 21172 -11248 21228 -11246
rect 21172 -11300 21174 -11248
rect 21174 -11300 21226 -11248
rect 21226 -11300 21228 -11248
rect 21172 -11302 21228 -11300
rect 21492 -11248 21548 -11246
rect 21492 -11300 21494 -11248
rect 21494 -11300 21546 -11248
rect 21546 -11300 21548 -11248
rect 21492 -11302 21548 -11300
rect 21812 -11248 21868 -11246
rect 21812 -11300 21814 -11248
rect 21814 -11300 21866 -11248
rect 21866 -11300 21868 -11248
rect 21812 -11302 21868 -11300
rect 22132 -11248 22188 -11246
rect 22132 -11300 22134 -11248
rect 22134 -11300 22186 -11248
rect 22186 -11300 22188 -11248
rect 22132 -11302 22188 -11300
rect 22452 -11248 22508 -11246
rect 22452 -11300 22454 -11248
rect 22454 -11300 22506 -11248
rect 22506 -11300 22508 -11248
rect 22452 -11302 22508 -11300
rect 22772 -11248 22828 -11246
rect 22772 -11300 22774 -11248
rect 22774 -11300 22826 -11248
rect 22826 -11300 22828 -11248
rect 22772 -11302 22828 -11300
rect 23092 -11248 23148 -11246
rect 23092 -11300 23094 -11248
rect 23094 -11300 23146 -11248
rect 23146 -11300 23148 -11248
rect 23092 -11302 23148 -11300
rect 23412 -11248 23468 -11246
rect 23412 -11300 23414 -11248
rect 23414 -11300 23466 -11248
rect 23466 -11300 23468 -11248
rect 23412 -11302 23468 -11300
rect 23732 -11248 23788 -11246
rect 23732 -11300 23734 -11248
rect 23734 -11300 23786 -11248
rect 23786 -11300 23788 -11248
rect 23732 -11302 23788 -11300
rect 24052 -11248 24108 -11246
rect 24052 -11300 24054 -11248
rect 24054 -11300 24106 -11248
rect 24106 -11300 24108 -11248
rect 24052 -11302 24108 -11300
rect 24372 -11248 24428 -11246
rect 24372 -11300 24374 -11248
rect 24374 -11300 24426 -11248
rect 24426 -11300 24428 -11248
rect 24372 -11302 24428 -11300
rect 24692 -11248 24748 -11246
rect 24692 -11300 24694 -11248
rect 24694 -11300 24746 -11248
rect 24746 -11300 24748 -11248
rect 24692 -11302 24748 -11300
rect 25012 -11248 25068 -11246
rect 25012 -11300 25014 -11248
rect 25014 -11300 25066 -11248
rect 25066 -11300 25068 -11248
rect 25012 -11302 25068 -11300
rect 25332 -11248 25388 -11246
rect 25332 -11300 25334 -11248
rect 25334 -11300 25386 -11248
rect 25386 -11300 25388 -11248
rect 25332 -11302 25388 -11300
rect 18242 -11454 18298 -11452
rect 18242 -11506 18244 -11454
rect 18244 -11506 18296 -11454
rect 18296 -11506 18298 -11454
rect 18242 -11508 18298 -11506
rect 25708 -11454 25764 -11452
rect 25708 -11506 25710 -11454
rect 25710 -11506 25762 -11454
rect 25762 -11506 25764 -11454
rect 25708 -11508 25764 -11506
rect 6242 -11774 6298 -11772
rect 6242 -11826 6244 -11774
rect 6244 -11826 6296 -11774
rect 6296 -11826 6298 -11774
rect 6242 -11828 6298 -11826
rect 6242 -12094 6298 -12092
rect 6242 -12146 6244 -12094
rect 6244 -12146 6296 -12094
rect 6296 -12146 6298 -12094
rect 6242 -12148 6298 -12146
rect 6242 -12414 6298 -12412
rect 6242 -12466 6244 -12414
rect 6244 -12466 6296 -12414
rect 6296 -12466 6298 -12414
rect 6242 -12468 6298 -12466
rect 6242 -12734 6298 -12732
rect 6242 -12786 6244 -12734
rect 6244 -12786 6296 -12734
rect 6296 -12786 6298 -12734
rect 6242 -12788 6298 -12786
rect 6242 -13054 6298 -13052
rect 6242 -13106 6244 -13054
rect 6244 -13106 6296 -13054
rect 6296 -13106 6298 -13054
rect 6242 -13108 6298 -13106
rect 6242 -13374 6298 -13372
rect 6242 -13426 6244 -13374
rect 6244 -13426 6296 -13374
rect 6296 -13426 6298 -13374
rect 6242 -13428 6298 -13426
rect 6242 -13694 6298 -13692
rect 6242 -13746 6244 -13694
rect 6244 -13746 6296 -13694
rect 6296 -13746 6298 -13694
rect 6242 -13748 6298 -13746
rect 6242 -14014 6298 -14012
rect 6242 -14066 6244 -14014
rect 6244 -14066 6296 -14014
rect 6296 -14066 6298 -14014
rect 6242 -14068 6298 -14066
rect 6242 -14334 6298 -14332
rect 6242 -14386 6244 -14334
rect 6244 -14386 6296 -14334
rect 6296 -14386 6298 -14334
rect 6242 -14388 6298 -14386
rect 6242 -14654 6298 -14652
rect 6242 -14706 6244 -14654
rect 6244 -14706 6296 -14654
rect 6296 -14706 6298 -14654
rect 6242 -14708 6298 -14706
rect 6242 -14974 6298 -14972
rect 6242 -15026 6244 -14974
rect 6244 -15026 6296 -14974
rect 6296 -15026 6298 -14974
rect 6242 -15028 6298 -15026
rect 6242 -15294 6298 -15292
rect 6242 -15346 6244 -15294
rect 6244 -15346 6296 -15294
rect 6296 -15346 6298 -15294
rect 6242 -15348 6298 -15346
rect 6242 -15614 6298 -15612
rect 6242 -15666 6244 -15614
rect 6244 -15666 6296 -15614
rect 6296 -15666 6298 -15614
rect 6242 -15668 6298 -15666
rect 6242 -15934 6298 -15932
rect 6242 -15986 6244 -15934
rect 6244 -15986 6296 -15934
rect 6296 -15986 6298 -15934
rect 6242 -15988 6298 -15986
rect 6242 -16254 6298 -16252
rect 6242 -16306 6244 -16254
rect 6244 -16306 6296 -16254
rect 6296 -16306 6298 -16254
rect 6242 -16308 6298 -16306
rect 6242 -16574 6298 -16572
rect 6242 -16626 6244 -16574
rect 6244 -16626 6296 -16574
rect 6296 -16626 6298 -16574
rect 6242 -16628 6298 -16626
rect 6242 -16894 6298 -16892
rect 6242 -16946 6244 -16894
rect 6244 -16946 6296 -16894
rect 6296 -16946 6298 -16894
rect 6242 -16948 6298 -16946
rect 6242 -17214 6298 -17212
rect 6242 -17266 6244 -17214
rect 6244 -17266 6296 -17214
rect 6296 -17266 6298 -17214
rect 6242 -17268 6298 -17266
rect 6242 -17534 6298 -17532
rect 6242 -17586 6244 -17534
rect 6244 -17586 6296 -17534
rect 6296 -17586 6298 -17534
rect 6242 -17588 6298 -17586
rect 6242 -17854 6298 -17852
rect 6242 -17906 6244 -17854
rect 6244 -17906 6296 -17854
rect 6296 -17906 6298 -17854
rect 6242 -17908 6298 -17906
rect 6242 -18174 6298 -18172
rect 6242 -18226 6244 -18174
rect 6244 -18226 6296 -18174
rect 6296 -18226 6298 -18174
rect 6242 -18228 6298 -18226
rect 13708 -11774 13764 -11772
rect 13708 -11826 13710 -11774
rect 13710 -11826 13762 -11774
rect 13762 -11826 13764 -11774
rect 13708 -11828 13764 -11826
rect 13708 -12094 13764 -12092
rect 13708 -12146 13710 -12094
rect 13710 -12146 13762 -12094
rect 13762 -12146 13764 -12094
rect 13708 -12148 13764 -12146
rect 13708 -12414 13764 -12412
rect 13708 -12466 13710 -12414
rect 13710 -12466 13762 -12414
rect 13762 -12466 13764 -12414
rect 13708 -12468 13764 -12466
rect 13708 -12734 13764 -12732
rect 13708 -12786 13710 -12734
rect 13710 -12786 13762 -12734
rect 13762 -12786 13764 -12734
rect 13708 -12788 13764 -12786
rect 13708 -13054 13764 -13052
rect 13708 -13106 13710 -13054
rect 13710 -13106 13762 -13054
rect 13762 -13106 13764 -13054
rect 13708 -13108 13764 -13106
rect 13708 -13374 13764 -13372
rect 13708 -13426 13710 -13374
rect 13710 -13426 13762 -13374
rect 13762 -13426 13764 -13374
rect 13708 -13428 13764 -13426
rect 13708 -13694 13764 -13692
rect 13708 -13746 13710 -13694
rect 13710 -13746 13762 -13694
rect 13762 -13746 13764 -13694
rect 13708 -13748 13764 -13746
rect 13708 -14014 13764 -14012
rect 13708 -14066 13710 -14014
rect 13710 -14066 13762 -14014
rect 13762 -14066 13764 -14014
rect 13708 -14068 13764 -14066
rect 13708 -14334 13764 -14332
rect 13708 -14386 13710 -14334
rect 13710 -14386 13762 -14334
rect 13762 -14386 13764 -14334
rect 13708 -14388 13764 -14386
rect 13708 -14654 13764 -14652
rect 13708 -14706 13710 -14654
rect 13710 -14706 13762 -14654
rect 13762 -14706 13764 -14654
rect 13708 -14708 13764 -14706
rect 13708 -14974 13764 -14972
rect 13708 -15026 13710 -14974
rect 13710 -15026 13762 -14974
rect 13762 -15026 13764 -14974
rect 13708 -15028 13764 -15026
rect 13708 -15294 13764 -15292
rect 13708 -15346 13710 -15294
rect 13710 -15346 13762 -15294
rect 13762 -15346 13764 -15294
rect 13708 -15348 13764 -15346
rect 13708 -15614 13764 -15612
rect 13708 -15666 13710 -15614
rect 13710 -15666 13762 -15614
rect 13762 -15666 13764 -15614
rect 13708 -15668 13764 -15666
rect 13708 -15934 13764 -15932
rect 13708 -15986 13710 -15934
rect 13710 -15986 13762 -15934
rect 13762 -15986 13764 -15934
rect 13708 -15988 13764 -15986
rect 13708 -16254 13764 -16252
rect 13708 -16306 13710 -16254
rect 13710 -16306 13762 -16254
rect 13762 -16306 13764 -16254
rect 13708 -16308 13764 -16306
rect 13708 -16574 13764 -16572
rect 13708 -16626 13710 -16574
rect 13710 -16626 13762 -16574
rect 13762 -16626 13764 -16574
rect 13708 -16628 13764 -16626
rect 13708 -16894 13764 -16892
rect 13708 -16946 13710 -16894
rect 13710 -16946 13762 -16894
rect 13762 -16946 13764 -16894
rect 13708 -16948 13764 -16946
rect 13708 -17214 13764 -17212
rect 13708 -17266 13710 -17214
rect 13710 -17266 13762 -17214
rect 13762 -17266 13764 -17214
rect 13708 -17268 13764 -17266
rect 13708 -17534 13764 -17532
rect 13708 -17586 13710 -17534
rect 13710 -17586 13762 -17534
rect 13762 -17586 13764 -17534
rect 13708 -17588 13764 -17586
rect 13708 -17854 13764 -17852
rect 13708 -17906 13710 -17854
rect 13710 -17906 13762 -17854
rect 13762 -17906 13764 -17854
rect 13708 -17908 13764 -17906
rect 13708 -18174 13764 -18172
rect 13708 -18226 13710 -18174
rect 13710 -18226 13762 -18174
rect 13762 -18226 13764 -18174
rect 13708 -18228 13764 -18226
rect 6242 -18494 6298 -18492
rect 6242 -18546 6244 -18494
rect 6244 -18546 6296 -18494
rect 6296 -18546 6298 -18494
rect 6242 -18548 6298 -18546
rect 13708 -18494 13764 -18492
rect 13708 -18546 13710 -18494
rect 13710 -18546 13762 -18494
rect 13762 -18546 13764 -18494
rect 13708 -18548 13764 -18546
rect 6612 -18704 6668 -18702
rect 6612 -18756 6614 -18704
rect 6614 -18756 6666 -18704
rect 6666 -18756 6668 -18704
rect 6612 -18758 6668 -18756
rect 6932 -18704 6988 -18702
rect 6932 -18756 6934 -18704
rect 6934 -18756 6986 -18704
rect 6986 -18756 6988 -18704
rect 6932 -18758 6988 -18756
rect 7252 -18704 7308 -18702
rect 7252 -18756 7254 -18704
rect 7254 -18756 7306 -18704
rect 7306 -18756 7308 -18704
rect 7252 -18758 7308 -18756
rect 7572 -18704 7628 -18702
rect 7572 -18756 7574 -18704
rect 7574 -18756 7626 -18704
rect 7626 -18756 7628 -18704
rect 7572 -18758 7628 -18756
rect 7892 -18704 7948 -18702
rect 7892 -18756 7894 -18704
rect 7894 -18756 7946 -18704
rect 7946 -18756 7948 -18704
rect 7892 -18758 7948 -18756
rect 8212 -18704 8268 -18702
rect 8212 -18756 8214 -18704
rect 8214 -18756 8266 -18704
rect 8266 -18756 8268 -18704
rect 8212 -18758 8268 -18756
rect 8532 -18704 8588 -18702
rect 8532 -18756 8534 -18704
rect 8534 -18756 8586 -18704
rect 8586 -18756 8588 -18704
rect 8532 -18758 8588 -18756
rect 8852 -18704 8908 -18702
rect 8852 -18756 8854 -18704
rect 8854 -18756 8906 -18704
rect 8906 -18756 8908 -18704
rect 8852 -18758 8908 -18756
rect 9172 -18704 9228 -18702
rect 9172 -18756 9174 -18704
rect 9174 -18756 9226 -18704
rect 9226 -18756 9228 -18704
rect 9172 -18758 9228 -18756
rect 9492 -18704 9548 -18702
rect 9492 -18756 9494 -18704
rect 9494 -18756 9546 -18704
rect 9546 -18756 9548 -18704
rect 9492 -18758 9548 -18756
rect 9812 -18704 9868 -18702
rect 9812 -18756 9814 -18704
rect 9814 -18756 9866 -18704
rect 9866 -18756 9868 -18704
rect 9812 -18758 9868 -18756
rect 10132 -18704 10188 -18702
rect 10132 -18756 10134 -18704
rect 10134 -18756 10186 -18704
rect 10186 -18756 10188 -18704
rect 10132 -18758 10188 -18756
rect 10452 -18704 10508 -18702
rect 10452 -18756 10454 -18704
rect 10454 -18756 10506 -18704
rect 10506 -18756 10508 -18704
rect 10452 -18758 10508 -18756
rect 10772 -18704 10828 -18702
rect 10772 -18756 10774 -18704
rect 10774 -18756 10826 -18704
rect 10826 -18756 10828 -18704
rect 10772 -18758 10828 -18756
rect 11092 -18704 11148 -18702
rect 11092 -18756 11094 -18704
rect 11094 -18756 11146 -18704
rect 11146 -18756 11148 -18704
rect 11092 -18758 11148 -18756
rect 11412 -18704 11468 -18702
rect 11412 -18756 11414 -18704
rect 11414 -18756 11466 -18704
rect 11466 -18756 11468 -18704
rect 11412 -18758 11468 -18756
rect 11732 -18704 11788 -18702
rect 11732 -18756 11734 -18704
rect 11734 -18756 11786 -18704
rect 11786 -18756 11788 -18704
rect 11732 -18758 11788 -18756
rect 12052 -18704 12108 -18702
rect 12052 -18756 12054 -18704
rect 12054 -18756 12106 -18704
rect 12106 -18756 12108 -18704
rect 12052 -18758 12108 -18756
rect 12372 -18704 12428 -18702
rect 12372 -18756 12374 -18704
rect 12374 -18756 12426 -18704
rect 12426 -18756 12428 -18704
rect 12372 -18758 12428 -18756
rect 12692 -18704 12748 -18702
rect 12692 -18756 12694 -18704
rect 12694 -18756 12746 -18704
rect 12746 -18756 12748 -18704
rect 12692 -18758 12748 -18756
rect 13012 -18704 13068 -18702
rect 13012 -18756 13014 -18704
rect 13014 -18756 13066 -18704
rect 13066 -18756 13068 -18704
rect 13012 -18758 13068 -18756
rect 13332 -18704 13388 -18702
rect 13332 -18756 13334 -18704
rect 13334 -18756 13386 -18704
rect 13386 -18756 13388 -18704
rect 13332 -18758 13388 -18756
rect 18242 -11774 18298 -11772
rect 18242 -11826 18244 -11774
rect 18244 -11826 18296 -11774
rect 18296 -11826 18298 -11774
rect 18242 -11828 18298 -11826
rect 18242 -12094 18298 -12092
rect 18242 -12146 18244 -12094
rect 18244 -12146 18296 -12094
rect 18296 -12146 18298 -12094
rect 18242 -12148 18298 -12146
rect 18242 -12414 18298 -12412
rect 18242 -12466 18244 -12414
rect 18244 -12466 18296 -12414
rect 18296 -12466 18298 -12414
rect 18242 -12468 18298 -12466
rect 18242 -12734 18298 -12732
rect 18242 -12786 18244 -12734
rect 18244 -12786 18296 -12734
rect 18296 -12786 18298 -12734
rect 18242 -12788 18298 -12786
rect 18242 -13054 18298 -13052
rect 18242 -13106 18244 -13054
rect 18244 -13106 18296 -13054
rect 18296 -13106 18298 -13054
rect 18242 -13108 18298 -13106
rect 18242 -13374 18298 -13372
rect 18242 -13426 18244 -13374
rect 18244 -13426 18296 -13374
rect 18296 -13426 18298 -13374
rect 18242 -13428 18298 -13426
rect 18242 -13694 18298 -13692
rect 18242 -13746 18244 -13694
rect 18244 -13746 18296 -13694
rect 18296 -13746 18298 -13694
rect 18242 -13748 18298 -13746
rect 18242 -14014 18298 -14012
rect 18242 -14066 18244 -14014
rect 18244 -14066 18296 -14014
rect 18296 -14066 18298 -14014
rect 18242 -14068 18298 -14066
rect 18242 -14334 18298 -14332
rect 18242 -14386 18244 -14334
rect 18244 -14386 18296 -14334
rect 18296 -14386 18298 -14334
rect 18242 -14388 18298 -14386
rect 18242 -14654 18298 -14652
rect 18242 -14706 18244 -14654
rect 18244 -14706 18296 -14654
rect 18296 -14706 18298 -14654
rect 18242 -14708 18298 -14706
rect 18242 -14974 18298 -14972
rect 18242 -15026 18244 -14974
rect 18244 -15026 18296 -14974
rect 18296 -15026 18298 -14974
rect 18242 -15028 18298 -15026
rect 18242 -15294 18298 -15292
rect 18242 -15346 18244 -15294
rect 18244 -15346 18296 -15294
rect 18296 -15346 18298 -15294
rect 18242 -15348 18298 -15346
rect 18242 -15614 18298 -15612
rect 18242 -15666 18244 -15614
rect 18244 -15666 18296 -15614
rect 18296 -15666 18298 -15614
rect 18242 -15668 18298 -15666
rect 18242 -15934 18298 -15932
rect 18242 -15986 18244 -15934
rect 18244 -15986 18296 -15934
rect 18296 -15986 18298 -15934
rect 18242 -15988 18298 -15986
rect 18242 -16254 18298 -16252
rect 18242 -16306 18244 -16254
rect 18244 -16306 18296 -16254
rect 18296 -16306 18298 -16254
rect 18242 -16308 18298 -16306
rect 18242 -16574 18298 -16572
rect 18242 -16626 18244 -16574
rect 18244 -16626 18296 -16574
rect 18296 -16626 18298 -16574
rect 18242 -16628 18298 -16626
rect 18242 -16894 18298 -16892
rect 18242 -16946 18244 -16894
rect 18244 -16946 18296 -16894
rect 18296 -16946 18298 -16894
rect 18242 -16948 18298 -16946
rect 18242 -17214 18298 -17212
rect 18242 -17266 18244 -17214
rect 18244 -17266 18296 -17214
rect 18296 -17266 18298 -17214
rect 18242 -17268 18298 -17266
rect 18242 -17534 18298 -17532
rect 18242 -17586 18244 -17534
rect 18244 -17586 18296 -17534
rect 18296 -17586 18298 -17534
rect 18242 -17588 18298 -17586
rect 18242 -17854 18298 -17852
rect 18242 -17906 18244 -17854
rect 18244 -17906 18296 -17854
rect 18296 -17906 18298 -17854
rect 18242 -17908 18298 -17906
rect 18242 -18174 18298 -18172
rect 18242 -18226 18244 -18174
rect 18244 -18226 18296 -18174
rect 18296 -18226 18298 -18174
rect 18242 -18228 18298 -18226
rect 25708 -11774 25764 -11772
rect 25708 -11826 25710 -11774
rect 25710 -11826 25762 -11774
rect 25762 -11826 25764 -11774
rect 25708 -11828 25764 -11826
rect 25708 -12094 25764 -12092
rect 25708 -12146 25710 -12094
rect 25710 -12146 25762 -12094
rect 25762 -12146 25764 -12094
rect 25708 -12148 25764 -12146
rect 25708 -12414 25764 -12412
rect 25708 -12466 25710 -12414
rect 25710 -12466 25762 -12414
rect 25762 -12466 25764 -12414
rect 25708 -12468 25764 -12466
rect 25708 -12734 25764 -12732
rect 25708 -12786 25710 -12734
rect 25710 -12786 25762 -12734
rect 25762 -12786 25764 -12734
rect 25708 -12788 25764 -12786
rect 25708 -13054 25764 -13052
rect 25708 -13106 25710 -13054
rect 25710 -13106 25762 -13054
rect 25762 -13106 25764 -13054
rect 25708 -13108 25764 -13106
rect 25708 -13374 25764 -13372
rect 25708 -13426 25710 -13374
rect 25710 -13426 25762 -13374
rect 25762 -13426 25764 -13374
rect 25708 -13428 25764 -13426
rect 25708 -13694 25764 -13692
rect 25708 -13746 25710 -13694
rect 25710 -13746 25762 -13694
rect 25762 -13746 25764 -13694
rect 25708 -13748 25764 -13746
rect 25708 -14014 25764 -14012
rect 25708 -14066 25710 -14014
rect 25710 -14066 25762 -14014
rect 25762 -14066 25764 -14014
rect 25708 -14068 25764 -14066
rect 25708 -14334 25764 -14332
rect 25708 -14386 25710 -14334
rect 25710 -14386 25762 -14334
rect 25762 -14386 25764 -14334
rect 25708 -14388 25764 -14386
rect 25708 -14654 25764 -14652
rect 25708 -14706 25710 -14654
rect 25710 -14706 25762 -14654
rect 25762 -14706 25764 -14654
rect 25708 -14708 25764 -14706
rect 25708 -14974 25764 -14972
rect 25708 -15026 25710 -14974
rect 25710 -15026 25762 -14974
rect 25762 -15026 25764 -14974
rect 25708 -15028 25764 -15026
rect 25708 -15294 25764 -15292
rect 25708 -15346 25710 -15294
rect 25710 -15346 25762 -15294
rect 25762 -15346 25764 -15294
rect 25708 -15348 25764 -15346
rect 25708 -15614 25764 -15612
rect 25708 -15666 25710 -15614
rect 25710 -15666 25762 -15614
rect 25762 -15666 25764 -15614
rect 25708 -15668 25764 -15666
rect 25708 -15934 25764 -15932
rect 25708 -15986 25710 -15934
rect 25710 -15986 25762 -15934
rect 25762 -15986 25764 -15934
rect 25708 -15988 25764 -15986
rect 25708 -16254 25764 -16252
rect 25708 -16306 25710 -16254
rect 25710 -16306 25762 -16254
rect 25762 -16306 25764 -16254
rect 25708 -16308 25764 -16306
rect 25708 -16574 25764 -16572
rect 25708 -16626 25710 -16574
rect 25710 -16626 25762 -16574
rect 25762 -16626 25764 -16574
rect 25708 -16628 25764 -16626
rect 25708 -16894 25764 -16892
rect 25708 -16946 25710 -16894
rect 25710 -16946 25762 -16894
rect 25762 -16946 25764 -16894
rect 25708 -16948 25764 -16946
rect 25708 -17214 25764 -17212
rect 25708 -17266 25710 -17214
rect 25710 -17266 25762 -17214
rect 25762 -17266 25764 -17214
rect 25708 -17268 25764 -17266
rect 25708 -17534 25764 -17532
rect 25708 -17586 25710 -17534
rect 25710 -17586 25762 -17534
rect 25762 -17586 25764 -17534
rect 25708 -17588 25764 -17586
rect 25708 -17854 25764 -17852
rect 25708 -17906 25710 -17854
rect 25710 -17906 25762 -17854
rect 25762 -17906 25764 -17854
rect 25708 -17908 25764 -17906
rect 25708 -18174 25764 -18172
rect 25708 -18226 25710 -18174
rect 25710 -18226 25762 -18174
rect 25762 -18226 25764 -18174
rect 25708 -18228 25764 -18226
rect 18242 -18494 18298 -18492
rect 18242 -18546 18244 -18494
rect 18244 -18546 18296 -18494
rect 18296 -18546 18298 -18494
rect 18242 -18548 18298 -18546
rect 25708 -18494 25764 -18492
rect 25708 -18546 25710 -18494
rect 25710 -18546 25762 -18494
rect 25762 -18546 25764 -18494
rect 25708 -18548 25764 -18546
rect 18612 -18704 18668 -18702
rect 18612 -18756 18614 -18704
rect 18614 -18756 18666 -18704
rect 18666 -18756 18668 -18704
rect 18612 -18758 18668 -18756
rect 18932 -18704 18988 -18702
rect 18932 -18756 18934 -18704
rect 18934 -18756 18986 -18704
rect 18986 -18756 18988 -18704
rect 18932 -18758 18988 -18756
rect 19252 -18704 19308 -18702
rect 19252 -18756 19254 -18704
rect 19254 -18756 19306 -18704
rect 19306 -18756 19308 -18704
rect 19252 -18758 19308 -18756
rect 19572 -18704 19628 -18702
rect 19572 -18756 19574 -18704
rect 19574 -18756 19626 -18704
rect 19626 -18756 19628 -18704
rect 19572 -18758 19628 -18756
rect 19892 -18704 19948 -18702
rect 19892 -18756 19894 -18704
rect 19894 -18756 19946 -18704
rect 19946 -18756 19948 -18704
rect 19892 -18758 19948 -18756
rect 20212 -18704 20268 -18702
rect 20212 -18756 20214 -18704
rect 20214 -18756 20266 -18704
rect 20266 -18756 20268 -18704
rect 20212 -18758 20268 -18756
rect 20532 -18704 20588 -18702
rect 20532 -18756 20534 -18704
rect 20534 -18756 20586 -18704
rect 20586 -18756 20588 -18704
rect 20532 -18758 20588 -18756
rect 20852 -18704 20908 -18702
rect 20852 -18756 20854 -18704
rect 20854 -18756 20906 -18704
rect 20906 -18756 20908 -18704
rect 20852 -18758 20908 -18756
rect 21172 -18704 21228 -18702
rect 21172 -18756 21174 -18704
rect 21174 -18756 21226 -18704
rect 21226 -18756 21228 -18704
rect 21172 -18758 21228 -18756
rect 21492 -18704 21548 -18702
rect 21492 -18756 21494 -18704
rect 21494 -18756 21546 -18704
rect 21546 -18756 21548 -18704
rect 21492 -18758 21548 -18756
rect 21812 -18704 21868 -18702
rect 21812 -18756 21814 -18704
rect 21814 -18756 21866 -18704
rect 21866 -18756 21868 -18704
rect 21812 -18758 21868 -18756
rect 22132 -18704 22188 -18702
rect 22132 -18756 22134 -18704
rect 22134 -18756 22186 -18704
rect 22186 -18756 22188 -18704
rect 22132 -18758 22188 -18756
rect 22452 -18704 22508 -18702
rect 22452 -18756 22454 -18704
rect 22454 -18756 22506 -18704
rect 22506 -18756 22508 -18704
rect 22452 -18758 22508 -18756
rect 22772 -18704 22828 -18702
rect 22772 -18756 22774 -18704
rect 22774 -18756 22826 -18704
rect 22826 -18756 22828 -18704
rect 22772 -18758 22828 -18756
rect 23092 -18704 23148 -18702
rect 23092 -18756 23094 -18704
rect 23094 -18756 23146 -18704
rect 23146 -18756 23148 -18704
rect 23092 -18758 23148 -18756
rect 23412 -18704 23468 -18702
rect 23412 -18756 23414 -18704
rect 23414 -18756 23466 -18704
rect 23466 -18756 23468 -18704
rect 23412 -18758 23468 -18756
rect 23732 -18704 23788 -18702
rect 23732 -18756 23734 -18704
rect 23734 -18756 23786 -18704
rect 23786 -18756 23788 -18704
rect 23732 -18758 23788 -18756
rect 24052 -18704 24108 -18702
rect 24052 -18756 24054 -18704
rect 24054 -18756 24106 -18704
rect 24106 -18756 24108 -18704
rect 24052 -18758 24108 -18756
rect 24372 -18704 24428 -18702
rect 24372 -18756 24374 -18704
rect 24374 -18756 24426 -18704
rect 24426 -18756 24428 -18704
rect 24372 -18758 24428 -18756
rect 24692 -18704 24748 -18702
rect 24692 -18756 24694 -18704
rect 24694 -18756 24746 -18704
rect 24746 -18756 24748 -18704
rect 24692 -18758 24748 -18756
rect 25012 -18704 25068 -18702
rect 25012 -18756 25014 -18704
rect 25014 -18756 25066 -18704
rect 25066 -18756 25068 -18704
rect 25012 -18758 25068 -18756
rect 25332 -18704 25388 -18702
rect 25332 -18756 25334 -18704
rect 25334 -18756 25386 -18704
rect 25386 -18756 25388 -18704
rect 25332 -18758 25388 -18756
rect 30612 -11248 30668 -11246
rect 30612 -11300 30614 -11248
rect 30614 -11300 30666 -11248
rect 30666 -11300 30668 -11248
rect 30612 -11302 30668 -11300
rect 30932 -11248 30988 -11246
rect 30932 -11300 30934 -11248
rect 30934 -11300 30986 -11248
rect 30986 -11300 30988 -11248
rect 30932 -11302 30988 -11300
rect 31252 -11248 31308 -11246
rect 31252 -11300 31254 -11248
rect 31254 -11300 31306 -11248
rect 31306 -11300 31308 -11248
rect 31252 -11302 31308 -11300
rect 31572 -11248 31628 -11246
rect 31572 -11300 31574 -11248
rect 31574 -11300 31626 -11248
rect 31626 -11300 31628 -11248
rect 31572 -11302 31628 -11300
rect 31892 -11248 31948 -11246
rect 31892 -11300 31894 -11248
rect 31894 -11300 31946 -11248
rect 31946 -11300 31948 -11248
rect 31892 -11302 31948 -11300
rect 32212 -11248 32268 -11246
rect 32212 -11300 32214 -11248
rect 32214 -11300 32266 -11248
rect 32266 -11300 32268 -11248
rect 32212 -11302 32268 -11300
rect 32532 -11248 32588 -11246
rect 32532 -11300 32534 -11248
rect 32534 -11300 32586 -11248
rect 32586 -11300 32588 -11248
rect 32532 -11302 32588 -11300
rect 32852 -11248 32908 -11246
rect 32852 -11300 32854 -11248
rect 32854 -11300 32906 -11248
rect 32906 -11300 32908 -11248
rect 32852 -11302 32908 -11300
rect 33172 -11248 33228 -11246
rect 33172 -11300 33174 -11248
rect 33174 -11300 33226 -11248
rect 33226 -11300 33228 -11248
rect 33172 -11302 33228 -11300
rect 33492 -11248 33548 -11246
rect 33492 -11300 33494 -11248
rect 33494 -11300 33546 -11248
rect 33546 -11300 33548 -11248
rect 33492 -11302 33548 -11300
rect 33812 -11248 33868 -11246
rect 33812 -11300 33814 -11248
rect 33814 -11300 33866 -11248
rect 33866 -11300 33868 -11248
rect 33812 -11302 33868 -11300
rect 34132 -11248 34188 -11246
rect 34132 -11300 34134 -11248
rect 34134 -11300 34186 -11248
rect 34186 -11300 34188 -11248
rect 34132 -11302 34188 -11300
rect 34452 -11248 34508 -11246
rect 34452 -11300 34454 -11248
rect 34454 -11300 34506 -11248
rect 34506 -11300 34508 -11248
rect 34452 -11302 34508 -11300
rect 34772 -11248 34828 -11246
rect 34772 -11300 34774 -11248
rect 34774 -11300 34826 -11248
rect 34826 -11300 34828 -11248
rect 34772 -11302 34828 -11300
rect 35092 -11248 35148 -11246
rect 35092 -11300 35094 -11248
rect 35094 -11300 35146 -11248
rect 35146 -11300 35148 -11248
rect 35092 -11302 35148 -11300
rect 35412 -11248 35468 -11246
rect 35412 -11300 35414 -11248
rect 35414 -11300 35466 -11248
rect 35466 -11300 35468 -11248
rect 35412 -11302 35468 -11300
rect 35732 -11248 35788 -11246
rect 35732 -11300 35734 -11248
rect 35734 -11300 35786 -11248
rect 35786 -11300 35788 -11248
rect 35732 -11302 35788 -11300
rect 36052 -11248 36108 -11246
rect 36052 -11300 36054 -11248
rect 36054 -11300 36106 -11248
rect 36106 -11300 36108 -11248
rect 36052 -11302 36108 -11300
rect 36372 -11248 36428 -11246
rect 36372 -11300 36374 -11248
rect 36374 -11300 36426 -11248
rect 36426 -11300 36428 -11248
rect 36372 -11302 36428 -11300
rect 36692 -11248 36748 -11246
rect 36692 -11300 36694 -11248
rect 36694 -11300 36746 -11248
rect 36746 -11300 36748 -11248
rect 36692 -11302 36748 -11300
rect 37012 -11248 37068 -11246
rect 37012 -11300 37014 -11248
rect 37014 -11300 37066 -11248
rect 37066 -11300 37068 -11248
rect 37012 -11302 37068 -11300
rect 37332 -11248 37388 -11246
rect 37332 -11300 37334 -11248
rect 37334 -11300 37386 -11248
rect 37386 -11300 37388 -11248
rect 37332 -11302 37388 -11300
rect 30242 -11454 30298 -11452
rect 30242 -11506 30244 -11454
rect 30244 -11506 30296 -11454
rect 30296 -11506 30298 -11454
rect 30242 -11508 30298 -11506
rect 37708 -11454 37764 -11452
rect 37708 -11506 37710 -11454
rect 37710 -11506 37762 -11454
rect 37762 -11506 37764 -11454
rect 37708 -11508 37764 -11506
rect 30242 -11774 30298 -11772
rect 30242 -11826 30244 -11774
rect 30244 -11826 30296 -11774
rect 30296 -11826 30298 -11774
rect 30242 -11828 30298 -11826
rect 30242 -12094 30298 -12092
rect 30242 -12146 30244 -12094
rect 30244 -12146 30296 -12094
rect 30296 -12146 30298 -12094
rect 30242 -12148 30298 -12146
rect 30242 -12414 30298 -12412
rect 30242 -12466 30244 -12414
rect 30244 -12466 30296 -12414
rect 30296 -12466 30298 -12414
rect 30242 -12468 30298 -12466
rect 30242 -12734 30298 -12732
rect 30242 -12786 30244 -12734
rect 30244 -12786 30296 -12734
rect 30296 -12786 30298 -12734
rect 30242 -12788 30298 -12786
rect 30242 -13054 30298 -13052
rect 30242 -13106 30244 -13054
rect 30244 -13106 30296 -13054
rect 30296 -13106 30298 -13054
rect 30242 -13108 30298 -13106
rect 30242 -13374 30298 -13372
rect 30242 -13426 30244 -13374
rect 30244 -13426 30296 -13374
rect 30296 -13426 30298 -13374
rect 30242 -13428 30298 -13426
rect 30242 -13694 30298 -13692
rect 30242 -13746 30244 -13694
rect 30244 -13746 30296 -13694
rect 30296 -13746 30298 -13694
rect 30242 -13748 30298 -13746
rect 30242 -14014 30298 -14012
rect 30242 -14066 30244 -14014
rect 30244 -14066 30296 -14014
rect 30296 -14066 30298 -14014
rect 30242 -14068 30298 -14066
rect 30242 -14334 30298 -14332
rect 30242 -14386 30244 -14334
rect 30244 -14386 30296 -14334
rect 30296 -14386 30298 -14334
rect 30242 -14388 30298 -14386
rect 30242 -14654 30298 -14652
rect 30242 -14706 30244 -14654
rect 30244 -14706 30296 -14654
rect 30296 -14706 30298 -14654
rect 30242 -14708 30298 -14706
rect 30242 -14974 30298 -14972
rect 30242 -15026 30244 -14974
rect 30244 -15026 30296 -14974
rect 30296 -15026 30298 -14974
rect 30242 -15028 30298 -15026
rect 30242 -15294 30298 -15292
rect 30242 -15346 30244 -15294
rect 30244 -15346 30296 -15294
rect 30296 -15346 30298 -15294
rect 30242 -15348 30298 -15346
rect 30242 -15614 30298 -15612
rect 30242 -15666 30244 -15614
rect 30244 -15666 30296 -15614
rect 30296 -15666 30298 -15614
rect 30242 -15668 30298 -15666
rect 30242 -15934 30298 -15932
rect 30242 -15986 30244 -15934
rect 30244 -15986 30296 -15934
rect 30296 -15986 30298 -15934
rect 30242 -15988 30298 -15986
rect 30242 -16254 30298 -16252
rect 30242 -16306 30244 -16254
rect 30244 -16306 30296 -16254
rect 30296 -16306 30298 -16254
rect 30242 -16308 30298 -16306
rect 30242 -16574 30298 -16572
rect 30242 -16626 30244 -16574
rect 30244 -16626 30296 -16574
rect 30296 -16626 30298 -16574
rect 30242 -16628 30298 -16626
rect 30242 -16894 30298 -16892
rect 30242 -16946 30244 -16894
rect 30244 -16946 30296 -16894
rect 30296 -16946 30298 -16894
rect 30242 -16948 30298 -16946
rect 30242 -17214 30298 -17212
rect 30242 -17266 30244 -17214
rect 30244 -17266 30296 -17214
rect 30296 -17266 30298 -17214
rect 30242 -17268 30298 -17266
rect 30242 -17534 30298 -17532
rect 30242 -17586 30244 -17534
rect 30244 -17586 30296 -17534
rect 30296 -17586 30298 -17534
rect 30242 -17588 30298 -17586
rect 30242 -17854 30298 -17852
rect 30242 -17906 30244 -17854
rect 30244 -17906 30296 -17854
rect 30296 -17906 30298 -17854
rect 30242 -17908 30298 -17906
rect 30242 -18174 30298 -18172
rect 30242 -18226 30244 -18174
rect 30244 -18226 30296 -18174
rect 30296 -18226 30298 -18174
rect 30242 -18228 30298 -18226
rect 37708 -11774 37764 -11772
rect 37708 -11826 37710 -11774
rect 37710 -11826 37762 -11774
rect 37762 -11826 37764 -11774
rect 37708 -11828 37764 -11826
rect 37708 -12094 37764 -12092
rect 37708 -12146 37710 -12094
rect 37710 -12146 37762 -12094
rect 37762 -12146 37764 -12094
rect 37708 -12148 37764 -12146
rect 37708 -12414 37764 -12412
rect 37708 -12466 37710 -12414
rect 37710 -12466 37762 -12414
rect 37762 -12466 37764 -12414
rect 37708 -12468 37764 -12466
rect 37708 -12734 37764 -12732
rect 37708 -12786 37710 -12734
rect 37710 -12786 37762 -12734
rect 37762 -12786 37764 -12734
rect 37708 -12788 37764 -12786
rect 37708 -13054 37764 -13052
rect 37708 -13106 37710 -13054
rect 37710 -13106 37762 -13054
rect 37762 -13106 37764 -13054
rect 37708 -13108 37764 -13106
rect 37708 -13374 37764 -13372
rect 37708 -13426 37710 -13374
rect 37710 -13426 37762 -13374
rect 37762 -13426 37764 -13374
rect 37708 -13428 37764 -13426
rect 37708 -13694 37764 -13692
rect 37708 -13746 37710 -13694
rect 37710 -13746 37762 -13694
rect 37762 -13746 37764 -13694
rect 37708 -13748 37764 -13746
rect 37708 -14014 37764 -14012
rect 37708 -14066 37710 -14014
rect 37710 -14066 37762 -14014
rect 37762 -14066 37764 -14014
rect 37708 -14068 37764 -14066
rect 37708 -14334 37764 -14332
rect 37708 -14386 37710 -14334
rect 37710 -14386 37762 -14334
rect 37762 -14386 37764 -14334
rect 37708 -14388 37764 -14386
rect 37708 -14654 37764 -14652
rect 37708 -14706 37710 -14654
rect 37710 -14706 37762 -14654
rect 37762 -14706 37764 -14654
rect 37708 -14708 37764 -14706
rect 37708 -14974 37764 -14972
rect 37708 -15026 37710 -14974
rect 37710 -15026 37762 -14974
rect 37762 -15026 37764 -14974
rect 37708 -15028 37764 -15026
rect 37708 -15294 37764 -15292
rect 37708 -15346 37710 -15294
rect 37710 -15346 37762 -15294
rect 37762 -15346 37764 -15294
rect 37708 -15348 37764 -15346
rect 37708 -15614 37764 -15612
rect 37708 -15666 37710 -15614
rect 37710 -15666 37762 -15614
rect 37762 -15666 37764 -15614
rect 37708 -15668 37764 -15666
rect 37708 -15934 37764 -15932
rect 37708 -15986 37710 -15934
rect 37710 -15986 37762 -15934
rect 37762 -15986 37764 -15934
rect 37708 -15988 37764 -15986
rect 37708 -16254 37764 -16252
rect 37708 -16306 37710 -16254
rect 37710 -16306 37762 -16254
rect 37762 -16306 37764 -16254
rect 37708 -16308 37764 -16306
rect 37708 -16574 37764 -16572
rect 37708 -16626 37710 -16574
rect 37710 -16626 37762 -16574
rect 37762 -16626 37764 -16574
rect 37708 -16628 37764 -16626
rect 37708 -16894 37764 -16892
rect 37708 -16946 37710 -16894
rect 37710 -16946 37762 -16894
rect 37762 -16946 37764 -16894
rect 37708 -16948 37764 -16946
rect 37708 -17214 37764 -17212
rect 37708 -17266 37710 -17214
rect 37710 -17266 37762 -17214
rect 37762 -17266 37764 -17214
rect 37708 -17268 37764 -17266
rect 37708 -17534 37764 -17532
rect 37708 -17586 37710 -17534
rect 37710 -17586 37762 -17534
rect 37762 -17586 37764 -17534
rect 37708 -17588 37764 -17586
rect 37708 -17854 37764 -17852
rect 37708 -17906 37710 -17854
rect 37710 -17906 37762 -17854
rect 37762 -17906 37764 -17854
rect 37708 -17908 37764 -17906
rect 37708 -18174 37764 -18172
rect 37708 -18226 37710 -18174
rect 37710 -18226 37762 -18174
rect 37762 -18226 37764 -18174
rect 37708 -18228 37764 -18226
rect 30242 -18494 30298 -18492
rect 30242 -18546 30244 -18494
rect 30244 -18546 30296 -18494
rect 30296 -18546 30298 -18494
rect 30242 -18548 30298 -18546
rect 37708 -18494 37764 -18492
rect 37708 -18546 37710 -18494
rect 37710 -18546 37762 -18494
rect 37762 -18546 37764 -18494
rect 37708 -18548 37764 -18546
rect 30612 -18704 30668 -18702
rect 30612 -18756 30614 -18704
rect 30614 -18756 30666 -18704
rect 30666 -18756 30668 -18704
rect 30612 -18758 30668 -18756
rect 30932 -18704 30988 -18702
rect 30932 -18756 30934 -18704
rect 30934 -18756 30986 -18704
rect 30986 -18756 30988 -18704
rect 30932 -18758 30988 -18756
rect 31252 -18704 31308 -18702
rect 31252 -18756 31254 -18704
rect 31254 -18756 31306 -18704
rect 31306 -18756 31308 -18704
rect 31252 -18758 31308 -18756
rect 31572 -18704 31628 -18702
rect 31572 -18756 31574 -18704
rect 31574 -18756 31626 -18704
rect 31626 -18756 31628 -18704
rect 31572 -18758 31628 -18756
rect 31892 -18704 31948 -18702
rect 31892 -18756 31894 -18704
rect 31894 -18756 31946 -18704
rect 31946 -18756 31948 -18704
rect 31892 -18758 31948 -18756
rect 32212 -18704 32268 -18702
rect 32212 -18756 32214 -18704
rect 32214 -18756 32266 -18704
rect 32266 -18756 32268 -18704
rect 32212 -18758 32268 -18756
rect 32532 -18704 32588 -18702
rect 32532 -18756 32534 -18704
rect 32534 -18756 32586 -18704
rect 32586 -18756 32588 -18704
rect 32532 -18758 32588 -18756
rect 32852 -18704 32908 -18702
rect 32852 -18756 32854 -18704
rect 32854 -18756 32906 -18704
rect 32906 -18756 32908 -18704
rect 32852 -18758 32908 -18756
rect 33172 -18704 33228 -18702
rect 33172 -18756 33174 -18704
rect 33174 -18756 33226 -18704
rect 33226 -18756 33228 -18704
rect 33172 -18758 33228 -18756
rect 33492 -18704 33548 -18702
rect 33492 -18756 33494 -18704
rect 33494 -18756 33546 -18704
rect 33546 -18756 33548 -18704
rect 33492 -18758 33548 -18756
rect 33812 -18704 33868 -18702
rect 33812 -18756 33814 -18704
rect 33814 -18756 33866 -18704
rect 33866 -18756 33868 -18704
rect 33812 -18758 33868 -18756
rect 34132 -18704 34188 -18702
rect 34132 -18756 34134 -18704
rect 34134 -18756 34186 -18704
rect 34186 -18756 34188 -18704
rect 34132 -18758 34188 -18756
rect 34452 -18704 34508 -18702
rect 34452 -18756 34454 -18704
rect 34454 -18756 34506 -18704
rect 34506 -18756 34508 -18704
rect 34452 -18758 34508 -18756
rect 34772 -18704 34828 -18702
rect 34772 -18756 34774 -18704
rect 34774 -18756 34826 -18704
rect 34826 -18756 34828 -18704
rect 34772 -18758 34828 -18756
rect 35092 -18704 35148 -18702
rect 35092 -18756 35094 -18704
rect 35094 -18756 35146 -18704
rect 35146 -18756 35148 -18704
rect 35092 -18758 35148 -18756
rect 35412 -18704 35468 -18702
rect 35412 -18756 35414 -18704
rect 35414 -18756 35466 -18704
rect 35466 -18756 35468 -18704
rect 35412 -18758 35468 -18756
rect 35732 -18704 35788 -18702
rect 35732 -18756 35734 -18704
rect 35734 -18756 35786 -18704
rect 35786 -18756 35788 -18704
rect 35732 -18758 35788 -18756
rect 36052 -18704 36108 -18702
rect 36052 -18756 36054 -18704
rect 36054 -18756 36106 -18704
rect 36106 -18756 36108 -18704
rect 36052 -18758 36108 -18756
rect 36372 -18704 36428 -18702
rect 36372 -18756 36374 -18704
rect 36374 -18756 36426 -18704
rect 36426 -18756 36428 -18704
rect 36372 -18758 36428 -18756
rect 36692 -18704 36748 -18702
rect 36692 -18756 36694 -18704
rect 36694 -18756 36746 -18704
rect 36746 -18756 36748 -18704
rect 36692 -18758 36748 -18756
rect 37012 -18704 37068 -18702
rect 37012 -18756 37014 -18704
rect 37014 -18756 37066 -18704
rect 37066 -18756 37068 -18704
rect 37012 -18758 37068 -18756
rect 37332 -18704 37388 -18702
rect 37332 -18756 37334 -18704
rect 37334 -18756 37386 -18704
rect 37386 -18756 37388 -18704
rect 37332 -18758 37388 -18756
rect 42612 -11248 42668 -11246
rect 42612 -11300 42614 -11248
rect 42614 -11300 42666 -11248
rect 42666 -11300 42668 -11248
rect 42612 -11302 42668 -11300
rect 42932 -11248 42988 -11246
rect 42932 -11300 42934 -11248
rect 42934 -11300 42986 -11248
rect 42986 -11300 42988 -11248
rect 42932 -11302 42988 -11300
rect 43252 -11248 43308 -11246
rect 43252 -11300 43254 -11248
rect 43254 -11300 43306 -11248
rect 43306 -11300 43308 -11248
rect 43252 -11302 43308 -11300
rect 43572 -11248 43628 -11246
rect 43572 -11300 43574 -11248
rect 43574 -11300 43626 -11248
rect 43626 -11300 43628 -11248
rect 43572 -11302 43628 -11300
rect 43892 -11248 43948 -11246
rect 43892 -11300 43894 -11248
rect 43894 -11300 43946 -11248
rect 43946 -11300 43948 -11248
rect 43892 -11302 43948 -11300
rect 44212 -11248 44268 -11246
rect 44212 -11300 44214 -11248
rect 44214 -11300 44266 -11248
rect 44266 -11300 44268 -11248
rect 44212 -11302 44268 -11300
rect 44532 -11248 44588 -11246
rect 44532 -11300 44534 -11248
rect 44534 -11300 44586 -11248
rect 44586 -11300 44588 -11248
rect 44532 -11302 44588 -11300
rect 44852 -11248 44908 -11246
rect 44852 -11300 44854 -11248
rect 44854 -11300 44906 -11248
rect 44906 -11300 44908 -11248
rect 44852 -11302 44908 -11300
rect 45172 -11248 45228 -11246
rect 45172 -11300 45174 -11248
rect 45174 -11300 45226 -11248
rect 45226 -11300 45228 -11248
rect 45172 -11302 45228 -11300
rect 45492 -11248 45548 -11246
rect 45492 -11300 45494 -11248
rect 45494 -11300 45546 -11248
rect 45546 -11300 45548 -11248
rect 45492 -11302 45548 -11300
rect 45812 -11248 45868 -11246
rect 45812 -11300 45814 -11248
rect 45814 -11300 45866 -11248
rect 45866 -11300 45868 -11248
rect 45812 -11302 45868 -11300
rect 46132 -11248 46188 -11246
rect 46132 -11300 46134 -11248
rect 46134 -11300 46186 -11248
rect 46186 -11300 46188 -11248
rect 46132 -11302 46188 -11300
rect 46452 -11248 46508 -11246
rect 46452 -11300 46454 -11248
rect 46454 -11300 46506 -11248
rect 46506 -11300 46508 -11248
rect 46452 -11302 46508 -11300
rect 46772 -11248 46828 -11246
rect 46772 -11300 46774 -11248
rect 46774 -11300 46826 -11248
rect 46826 -11300 46828 -11248
rect 46772 -11302 46828 -11300
rect 47092 -11248 47148 -11246
rect 47092 -11300 47094 -11248
rect 47094 -11300 47146 -11248
rect 47146 -11300 47148 -11248
rect 47092 -11302 47148 -11300
rect 47412 -11248 47468 -11246
rect 47412 -11300 47414 -11248
rect 47414 -11300 47466 -11248
rect 47466 -11300 47468 -11248
rect 47412 -11302 47468 -11300
rect 47732 -11248 47788 -11246
rect 47732 -11300 47734 -11248
rect 47734 -11300 47786 -11248
rect 47786 -11300 47788 -11248
rect 47732 -11302 47788 -11300
rect 48052 -11248 48108 -11246
rect 48052 -11300 48054 -11248
rect 48054 -11300 48106 -11248
rect 48106 -11300 48108 -11248
rect 48052 -11302 48108 -11300
rect 48372 -11248 48428 -11246
rect 48372 -11300 48374 -11248
rect 48374 -11300 48426 -11248
rect 48426 -11300 48428 -11248
rect 48372 -11302 48428 -11300
rect 48692 -11248 48748 -11246
rect 48692 -11300 48694 -11248
rect 48694 -11300 48746 -11248
rect 48746 -11300 48748 -11248
rect 48692 -11302 48748 -11300
rect 49012 -11248 49068 -11246
rect 49012 -11300 49014 -11248
rect 49014 -11300 49066 -11248
rect 49066 -11300 49068 -11248
rect 49012 -11302 49068 -11300
rect 49332 -11248 49388 -11246
rect 49332 -11300 49334 -11248
rect 49334 -11300 49386 -11248
rect 49386 -11300 49388 -11248
rect 49332 -11302 49388 -11300
rect 42245 -11454 42301 -11452
rect 42245 -11506 42247 -11454
rect 42247 -11506 42299 -11454
rect 42299 -11506 42301 -11454
rect 42245 -11508 42301 -11506
rect 49699 -11454 49755 -11452
rect 49699 -11506 49701 -11454
rect 49701 -11506 49753 -11454
rect 49753 -11506 49755 -11454
rect 49699 -11508 49755 -11506
rect 42245 -11774 42301 -11772
rect 42245 -11826 42247 -11774
rect 42247 -11826 42299 -11774
rect 42299 -11826 42301 -11774
rect 42245 -11828 42301 -11826
rect 42245 -12094 42301 -12092
rect 42245 -12146 42247 -12094
rect 42247 -12146 42299 -12094
rect 42299 -12146 42301 -12094
rect 42245 -12148 42301 -12146
rect 42245 -12414 42301 -12412
rect 42245 -12466 42247 -12414
rect 42247 -12466 42299 -12414
rect 42299 -12466 42301 -12414
rect 42245 -12468 42301 -12466
rect 42245 -12734 42301 -12732
rect 42245 -12786 42247 -12734
rect 42247 -12786 42299 -12734
rect 42299 -12786 42301 -12734
rect 42245 -12788 42301 -12786
rect 42245 -13054 42301 -13052
rect 42245 -13106 42247 -13054
rect 42247 -13106 42299 -13054
rect 42299 -13106 42301 -13054
rect 42245 -13108 42301 -13106
rect 42245 -13374 42301 -13372
rect 42245 -13426 42247 -13374
rect 42247 -13426 42299 -13374
rect 42299 -13426 42301 -13374
rect 42245 -13428 42301 -13426
rect 42245 -13694 42301 -13692
rect 42245 -13746 42247 -13694
rect 42247 -13746 42299 -13694
rect 42299 -13746 42301 -13694
rect 42245 -13748 42301 -13746
rect 42245 -14014 42301 -14012
rect 42245 -14066 42247 -14014
rect 42247 -14066 42299 -14014
rect 42299 -14066 42301 -14014
rect 42245 -14068 42301 -14066
rect 42245 -14334 42301 -14332
rect 42245 -14386 42247 -14334
rect 42247 -14386 42299 -14334
rect 42299 -14386 42301 -14334
rect 42245 -14388 42301 -14386
rect 42245 -14654 42301 -14652
rect 42245 -14706 42247 -14654
rect 42247 -14706 42299 -14654
rect 42299 -14706 42301 -14654
rect 42245 -14708 42301 -14706
rect 42245 -14974 42301 -14972
rect 42245 -15026 42247 -14974
rect 42247 -15026 42299 -14974
rect 42299 -15026 42301 -14974
rect 42245 -15028 42301 -15026
rect 42245 -15294 42301 -15292
rect 42245 -15346 42247 -15294
rect 42247 -15346 42299 -15294
rect 42299 -15346 42301 -15294
rect 42245 -15348 42301 -15346
rect 42245 -15614 42301 -15612
rect 42245 -15666 42247 -15614
rect 42247 -15666 42299 -15614
rect 42299 -15666 42301 -15614
rect 42245 -15668 42301 -15666
rect 42245 -15934 42301 -15932
rect 42245 -15986 42247 -15934
rect 42247 -15986 42299 -15934
rect 42299 -15986 42301 -15934
rect 42245 -15988 42301 -15986
rect 42245 -16254 42301 -16252
rect 42245 -16306 42247 -16254
rect 42247 -16306 42299 -16254
rect 42299 -16306 42301 -16254
rect 42245 -16308 42301 -16306
rect 42245 -16574 42301 -16572
rect 42245 -16626 42247 -16574
rect 42247 -16626 42299 -16574
rect 42299 -16626 42301 -16574
rect 42245 -16628 42301 -16626
rect 42245 -16894 42301 -16892
rect 42245 -16946 42247 -16894
rect 42247 -16946 42299 -16894
rect 42299 -16946 42301 -16894
rect 42245 -16948 42301 -16946
rect 42245 -17214 42301 -17212
rect 42245 -17266 42247 -17214
rect 42247 -17266 42299 -17214
rect 42299 -17266 42301 -17214
rect 42245 -17268 42301 -17266
rect 42245 -17534 42301 -17532
rect 42245 -17586 42247 -17534
rect 42247 -17586 42299 -17534
rect 42299 -17586 42301 -17534
rect 42245 -17588 42301 -17586
rect 42245 -17854 42301 -17852
rect 42245 -17906 42247 -17854
rect 42247 -17906 42299 -17854
rect 42299 -17906 42301 -17854
rect 42245 -17908 42301 -17906
rect 42245 -18174 42301 -18172
rect 42245 -18226 42247 -18174
rect 42247 -18226 42299 -18174
rect 42299 -18226 42301 -18174
rect 42245 -18228 42301 -18226
rect 49699 -11774 49755 -11772
rect 49699 -11826 49701 -11774
rect 49701 -11826 49753 -11774
rect 49753 -11826 49755 -11774
rect 49699 -11828 49755 -11826
rect 49699 -12094 49755 -12092
rect 49699 -12146 49701 -12094
rect 49701 -12146 49753 -12094
rect 49753 -12146 49755 -12094
rect 49699 -12148 49755 -12146
rect 49699 -12414 49755 -12412
rect 49699 -12466 49701 -12414
rect 49701 -12466 49753 -12414
rect 49753 -12466 49755 -12414
rect 49699 -12468 49755 -12466
rect 49699 -12734 49755 -12732
rect 49699 -12786 49701 -12734
rect 49701 -12786 49753 -12734
rect 49753 -12786 49755 -12734
rect 49699 -12788 49755 -12786
rect 49699 -13054 49755 -13052
rect 49699 -13106 49701 -13054
rect 49701 -13106 49753 -13054
rect 49753 -13106 49755 -13054
rect 49699 -13108 49755 -13106
rect 49699 -13374 49755 -13372
rect 49699 -13426 49701 -13374
rect 49701 -13426 49753 -13374
rect 49753 -13426 49755 -13374
rect 49699 -13428 49755 -13426
rect 49699 -13694 49755 -13692
rect 49699 -13746 49701 -13694
rect 49701 -13746 49753 -13694
rect 49753 -13746 49755 -13694
rect 49699 -13748 49755 -13746
rect 49699 -14014 49755 -14012
rect 49699 -14066 49701 -14014
rect 49701 -14066 49753 -14014
rect 49753 -14066 49755 -14014
rect 49699 -14068 49755 -14066
rect 49699 -14334 49755 -14332
rect 49699 -14386 49701 -14334
rect 49701 -14386 49753 -14334
rect 49753 -14386 49755 -14334
rect 49699 -14388 49755 -14386
rect 49699 -14654 49755 -14652
rect 49699 -14706 49701 -14654
rect 49701 -14706 49753 -14654
rect 49753 -14706 49755 -14654
rect 49699 -14708 49755 -14706
rect 49699 -14974 49755 -14972
rect 49699 -15026 49701 -14974
rect 49701 -15026 49753 -14974
rect 49753 -15026 49755 -14974
rect 49699 -15028 49755 -15026
rect 49699 -15294 49755 -15292
rect 49699 -15346 49701 -15294
rect 49701 -15346 49753 -15294
rect 49753 -15346 49755 -15294
rect 49699 -15348 49755 -15346
rect 49699 -15614 49755 -15612
rect 49699 -15666 49701 -15614
rect 49701 -15666 49753 -15614
rect 49753 -15666 49755 -15614
rect 49699 -15668 49755 -15666
rect 49699 -15934 49755 -15932
rect 49699 -15986 49701 -15934
rect 49701 -15986 49753 -15934
rect 49753 -15986 49755 -15934
rect 49699 -15988 49755 -15986
rect 49699 -16254 49755 -16252
rect 49699 -16306 49701 -16254
rect 49701 -16306 49753 -16254
rect 49753 -16306 49755 -16254
rect 49699 -16308 49755 -16306
rect 49699 -16574 49755 -16572
rect 49699 -16626 49701 -16574
rect 49701 -16626 49753 -16574
rect 49753 -16626 49755 -16574
rect 49699 -16628 49755 -16626
rect 49699 -16894 49755 -16892
rect 49699 -16946 49701 -16894
rect 49701 -16946 49753 -16894
rect 49753 -16946 49755 -16894
rect 49699 -16948 49755 -16946
rect 49699 -17214 49755 -17212
rect 49699 -17266 49701 -17214
rect 49701 -17266 49753 -17214
rect 49753 -17266 49755 -17214
rect 49699 -17268 49755 -17266
rect 49699 -17534 49755 -17532
rect 49699 -17586 49701 -17534
rect 49701 -17586 49753 -17534
rect 49753 -17586 49755 -17534
rect 49699 -17588 49755 -17586
rect 49699 -17854 49755 -17852
rect 49699 -17906 49701 -17854
rect 49701 -17906 49753 -17854
rect 49753 -17906 49755 -17854
rect 49699 -17908 49755 -17906
rect 49699 -18174 49755 -18172
rect 49699 -18226 49701 -18174
rect 49701 -18226 49753 -18174
rect 49753 -18226 49755 -18174
rect 49699 -18228 49755 -18226
rect 42245 -18494 42301 -18492
rect 42245 -18546 42247 -18494
rect 42247 -18546 42299 -18494
rect 42299 -18546 42301 -18494
rect 42245 -18548 42301 -18546
rect 49699 -18494 49755 -18492
rect 49699 -18546 49701 -18494
rect 49701 -18546 49753 -18494
rect 49753 -18546 49755 -18494
rect 49699 -18548 49755 -18546
rect 42612 -18704 42668 -18702
rect 42612 -18756 42614 -18704
rect 42614 -18756 42666 -18704
rect 42666 -18756 42668 -18704
rect 42612 -18758 42668 -18756
rect 42932 -18704 42988 -18702
rect 42932 -18756 42934 -18704
rect 42934 -18756 42986 -18704
rect 42986 -18756 42988 -18704
rect 42932 -18758 42988 -18756
rect 43252 -18704 43308 -18702
rect 43252 -18756 43254 -18704
rect 43254 -18756 43306 -18704
rect 43306 -18756 43308 -18704
rect 43252 -18758 43308 -18756
rect 43572 -18704 43628 -18702
rect 43572 -18756 43574 -18704
rect 43574 -18756 43626 -18704
rect 43626 -18756 43628 -18704
rect 43572 -18758 43628 -18756
rect 43892 -18704 43948 -18702
rect 43892 -18756 43894 -18704
rect 43894 -18756 43946 -18704
rect 43946 -18756 43948 -18704
rect 43892 -18758 43948 -18756
rect 44212 -18704 44268 -18702
rect 44212 -18756 44214 -18704
rect 44214 -18756 44266 -18704
rect 44266 -18756 44268 -18704
rect 44212 -18758 44268 -18756
rect 44532 -18704 44588 -18702
rect 44532 -18756 44534 -18704
rect 44534 -18756 44586 -18704
rect 44586 -18756 44588 -18704
rect 44532 -18758 44588 -18756
rect 44852 -18704 44908 -18702
rect 44852 -18756 44854 -18704
rect 44854 -18756 44906 -18704
rect 44906 -18756 44908 -18704
rect 44852 -18758 44908 -18756
rect 45172 -18704 45228 -18702
rect 45172 -18756 45174 -18704
rect 45174 -18756 45226 -18704
rect 45226 -18756 45228 -18704
rect 45172 -18758 45228 -18756
rect 45492 -18704 45548 -18702
rect 45492 -18756 45494 -18704
rect 45494 -18756 45546 -18704
rect 45546 -18756 45548 -18704
rect 45492 -18758 45548 -18756
rect 45812 -18704 45868 -18702
rect 45812 -18756 45814 -18704
rect 45814 -18756 45866 -18704
rect 45866 -18756 45868 -18704
rect 45812 -18758 45868 -18756
rect 46132 -18704 46188 -18702
rect 46132 -18756 46134 -18704
rect 46134 -18756 46186 -18704
rect 46186 -18756 46188 -18704
rect 46132 -18758 46188 -18756
rect 46452 -18704 46508 -18702
rect 46452 -18756 46454 -18704
rect 46454 -18756 46506 -18704
rect 46506 -18756 46508 -18704
rect 46452 -18758 46508 -18756
rect 46772 -18704 46828 -18702
rect 46772 -18756 46774 -18704
rect 46774 -18756 46826 -18704
rect 46826 -18756 46828 -18704
rect 46772 -18758 46828 -18756
rect 47092 -18704 47148 -18702
rect 47092 -18756 47094 -18704
rect 47094 -18756 47146 -18704
rect 47146 -18756 47148 -18704
rect 47092 -18758 47148 -18756
rect 47412 -18704 47468 -18702
rect 47412 -18756 47414 -18704
rect 47414 -18756 47466 -18704
rect 47466 -18756 47468 -18704
rect 47412 -18758 47468 -18756
rect 47732 -18704 47788 -18702
rect 47732 -18756 47734 -18704
rect 47734 -18756 47786 -18704
rect 47786 -18756 47788 -18704
rect 47732 -18758 47788 -18756
rect 48052 -18704 48108 -18702
rect 48052 -18756 48054 -18704
rect 48054 -18756 48106 -18704
rect 48106 -18756 48108 -18704
rect 48052 -18758 48108 -18756
rect 48372 -18704 48428 -18702
rect 48372 -18756 48374 -18704
rect 48374 -18756 48426 -18704
rect 48426 -18756 48428 -18704
rect 48372 -18758 48428 -18756
rect 48692 -18704 48748 -18702
rect 48692 -18756 48694 -18704
rect 48694 -18756 48746 -18704
rect 48746 -18756 48748 -18704
rect 48692 -18758 48748 -18756
rect 49012 -18704 49068 -18702
rect 49012 -18756 49014 -18704
rect 49014 -18756 49066 -18704
rect 49066 -18756 49068 -18704
rect 49012 -18758 49068 -18756
rect 49332 -18704 49388 -18702
rect 49332 -18756 49334 -18704
rect 49334 -18756 49386 -18704
rect 49386 -18756 49388 -18704
rect 49332 -18758 49388 -18756
rect 14300 -19700 14900 -19400
<< metal3 >>
rect 14200 4000 15000 7000
rect 13940 3720 14080 3740
rect 13940 3480 13960 3720
rect 14060 3480 14080 3720
rect 13940 2600 14080 3480
rect 13940 340 14100 2600
rect 14200 340 14500 4000
rect 20060 3280 20500 3300
rect 20060 3140 20080 3280
rect 20480 3140 20500 3280
rect 20060 3120 20500 3140
rect 20920 3280 23040 3300
rect 20920 3140 20940 3280
rect 21340 3140 23040 3280
rect 20920 3120 23040 3140
rect 15160 2940 15380 2960
rect 15160 2680 15180 2940
rect 15360 2680 15380 2940
rect 15160 2660 15380 2680
rect 22840 1800 23040 3120
rect 19980 1760 20300 1800
rect 19980 1460 20020 1760
rect 20260 1460 20300 1760
rect 19980 1420 20300 1460
rect 13920 320 14120 340
rect 13920 -80 13940 320
rect 14100 -80 14120 320
rect 13920 -100 14120 -80
rect 14180 320 14520 340
rect 14180 -80 14200 320
rect 14500 -80 14520 320
rect 14180 -100 14520 -80
rect 14920 -200 15160 -180
rect 14920 -580 14940 -200
rect 15140 -580 15160 -200
rect 14920 -600 15160 -580
rect 22800 -600 24440 1800
rect 14100 -1100 14280 -1080
rect 14100 -1620 14120 -1100
rect 14260 -1620 14280 -1100
rect 22800 -1220 23100 -600
rect 22800 -1580 22820 -1220
rect 22980 -1580 23100 -1220
rect 22800 -1600 23100 -1580
rect 14100 -1640 14280 -1620
rect 20340 -1680 20660 -1640
rect 20340 -2200 20380 -1680
rect 20620 -2200 20660 -1680
rect 20340 -2240 20660 -2200
rect 20740 -2570 21680 -2510
rect 20740 -4120 20800 -2570
rect 21720 -2780 23000 -2720
rect 21280 -3060 21560 -3040
rect 21650 -3050 21720 -2920
rect 21280 -3200 21300 -3060
rect 21540 -3200 21560 -3060
rect 21280 -3220 21560 -3200
rect 21440 -3680 21560 -3220
rect 21630 -3355 21740 -3050
rect 21630 -3500 22560 -3355
rect 21440 -3800 22080 -3680
rect 21180 -4100 21420 -4080
rect 21180 -4120 21200 -4100
rect 20740 -4200 21200 -4120
rect 17820 -4940 17900 -4800
rect 20280 -4860 20380 -4840
rect 20280 -4940 20300 -4860
rect 17820 -4980 20300 -4940
rect 20360 -4980 20380 -4860
rect 17820 -5000 20380 -4980
rect 20740 -4980 20800 -4200
rect 21180 -4500 21200 -4200
rect 21400 -4500 21420 -4100
rect 21180 -4520 21420 -4500
rect 21360 -4920 21560 -4900
rect 20740 -4990 20780 -4980
rect 21360 -5480 21380 -4920
rect 21540 -5480 21560 -4920
rect 21360 -5500 21560 -5480
rect 21260 -8780 21700 -5500
rect 21260 -8840 21860 -8780
rect 21340 -9260 21860 -8840
rect 21340 -9380 21360 -9260
rect 21840 -9380 21860 -9260
rect 21340 -9400 21860 -9380
rect 21960 -10740 22080 -3800
rect 13680 -10860 22080 -10740
rect 13680 -11000 13800 -10860
rect 22440 -11000 22560 -3500
rect 22880 -10440 23000 -2780
rect 22880 -10560 30440 -10440
rect 30320 -11000 30440 -10560
rect 6000 -11242 14000 -11000
rect 6000 -11306 6608 -11242
rect 6672 -11306 6928 -11242
rect 6992 -11306 7248 -11242
rect 7312 -11306 7568 -11242
rect 7632 -11306 7888 -11242
rect 7952 -11306 8208 -11242
rect 8272 -11306 8528 -11242
rect 8592 -11306 8848 -11242
rect 8912 -11306 9168 -11242
rect 9232 -11306 9488 -11242
rect 9552 -11306 9808 -11242
rect 9872 -11306 10128 -11242
rect 10192 -11306 10448 -11242
rect 10512 -11306 10768 -11242
rect 10832 -11306 11088 -11242
rect 11152 -11306 11408 -11242
rect 11472 -11306 11728 -11242
rect 11792 -11306 12048 -11242
rect 12112 -11306 12368 -11242
rect 12432 -11306 12688 -11242
rect 12752 -11306 13008 -11242
rect 13072 -11306 13328 -11242
rect 13392 -11306 14000 -11242
rect 6000 -11448 14000 -11306
rect 6000 -11512 6238 -11448
rect 6302 -11512 13704 -11448
rect 13768 -11512 14000 -11448
rect 6000 -11540 14000 -11512
rect 14180 -11100 14520 -11000
rect 14180 -11500 14200 -11100
rect 14500 -11500 14520 -11100
rect 14180 -11520 14520 -11500
rect 18000 -11242 26000 -11000
rect 18000 -11306 18608 -11242
rect 18672 -11306 18928 -11242
rect 18992 -11306 19248 -11242
rect 19312 -11306 19568 -11242
rect 19632 -11306 19888 -11242
rect 19952 -11306 20208 -11242
rect 20272 -11306 20528 -11242
rect 20592 -11306 20848 -11242
rect 20912 -11306 21168 -11242
rect 21232 -11306 21488 -11242
rect 21552 -11306 21808 -11242
rect 21872 -11306 22128 -11242
rect 22192 -11306 22448 -11242
rect 22512 -11306 22768 -11242
rect 22832 -11306 23088 -11242
rect 23152 -11306 23408 -11242
rect 23472 -11306 23728 -11242
rect 23792 -11306 24048 -11242
rect 24112 -11306 24368 -11242
rect 24432 -11306 24688 -11242
rect 24752 -11306 25008 -11242
rect 25072 -11306 25328 -11242
rect 25392 -11306 26000 -11242
rect 18000 -11448 26000 -11306
rect 18000 -11512 18238 -11448
rect 18302 -11512 25704 -11448
rect 25768 -11512 26000 -11448
rect 6000 -11768 6540 -11540
rect 6000 -11832 6238 -11768
rect 6302 -11832 6540 -11768
rect 6000 -12088 6540 -11832
rect 6000 -12152 6238 -12088
rect 6302 -12152 6540 -12088
rect 6000 -12408 6540 -12152
rect 6000 -12472 6238 -12408
rect 6302 -12472 6540 -12408
rect 6000 -12728 6540 -12472
rect 6000 -12792 6238 -12728
rect 6302 -12792 6540 -12728
rect 6000 -13048 6540 -12792
rect 6000 -13112 6238 -13048
rect 6302 -13112 6540 -13048
rect 6000 -13368 6540 -13112
rect 6000 -13432 6238 -13368
rect 6302 -13432 6540 -13368
rect 6000 -13688 6540 -13432
rect 6000 -13752 6238 -13688
rect 6302 -13752 6540 -13688
rect 6000 -14008 6540 -13752
rect 6000 -14072 6238 -14008
rect 6302 -14072 6540 -14008
rect 6000 -14328 6540 -14072
rect 6000 -14392 6238 -14328
rect 6302 -14392 6540 -14328
rect 6000 -14648 6540 -14392
rect 6000 -14712 6238 -14648
rect 6302 -14712 6540 -14648
rect 6000 -14968 6540 -14712
rect 6000 -15032 6238 -14968
rect 6302 -15032 6540 -14968
rect 6000 -15288 6540 -15032
rect 6000 -15352 6238 -15288
rect 6302 -15352 6540 -15288
rect 6000 -15608 6540 -15352
rect 6000 -15672 6238 -15608
rect 6302 -15672 6540 -15608
rect 6000 -15928 6540 -15672
rect 6000 -15992 6238 -15928
rect 6302 -15992 6540 -15928
rect 6000 -16248 6540 -15992
rect 6000 -16312 6238 -16248
rect 6302 -16312 6540 -16248
rect 6000 -16568 6540 -16312
rect 6000 -16632 6238 -16568
rect 6302 -16632 6540 -16568
rect 6000 -16888 6540 -16632
rect 6000 -16952 6238 -16888
rect 6302 -16952 6540 -16888
rect 6000 -17208 6540 -16952
rect 6000 -17272 6238 -17208
rect 6302 -17272 6540 -17208
rect 6000 -17528 6540 -17272
rect 6000 -17592 6238 -17528
rect 6302 -17592 6540 -17528
rect 6000 -17848 6540 -17592
rect 6000 -17912 6238 -17848
rect 6302 -17912 6540 -17848
rect 6000 -18168 6540 -17912
rect 6000 -18232 6238 -18168
rect 6302 -18232 6540 -18168
rect 6000 -18460 6540 -18232
rect 13460 -11768 14000 -11540
rect 13460 -11832 13704 -11768
rect 13768 -11832 14000 -11768
rect 13460 -12088 14000 -11832
rect 13460 -12152 13704 -12088
rect 13768 -12152 14000 -12088
rect 13460 -12408 14000 -12152
rect 13460 -12472 13704 -12408
rect 13768 -12472 14000 -12408
rect 13460 -12728 14000 -12472
rect 13460 -12792 13704 -12728
rect 13768 -12792 14000 -12728
rect 13460 -13048 14000 -12792
rect 13460 -13112 13704 -13048
rect 13768 -13112 14000 -13048
rect 13460 -13368 14000 -13112
rect 13460 -13432 13704 -13368
rect 13768 -13432 14000 -13368
rect 13460 -13688 14000 -13432
rect 13460 -13752 13704 -13688
rect 13768 -13752 14000 -13688
rect 13460 -14008 14000 -13752
rect 13460 -14072 13704 -14008
rect 13768 -14072 14000 -14008
rect 13460 -14328 14000 -14072
rect 13460 -14392 13704 -14328
rect 13768 -14392 14000 -14328
rect 13460 -14648 14000 -14392
rect 13460 -14712 13704 -14648
rect 13768 -14712 14000 -14648
rect 13460 -14968 14000 -14712
rect 13460 -15032 13704 -14968
rect 13768 -15032 14000 -14968
rect 13460 -15288 14000 -15032
rect 13460 -15352 13704 -15288
rect 13768 -15352 14000 -15288
rect 13460 -15608 14000 -15352
rect 13460 -15672 13704 -15608
rect 13768 -15672 14000 -15608
rect 13460 -15928 14000 -15672
rect 13460 -15992 13704 -15928
rect 13768 -15992 14000 -15928
rect 13460 -16248 14000 -15992
rect 13460 -16312 13704 -16248
rect 13768 -16312 14000 -16248
rect 13460 -16568 14000 -16312
rect 13460 -16632 13704 -16568
rect 13768 -16632 14000 -16568
rect 13460 -16888 14000 -16632
rect 13460 -16952 13704 -16888
rect 13768 -16952 14000 -16888
rect 13460 -17208 14000 -16952
rect 13460 -17272 13704 -17208
rect 13768 -17272 14000 -17208
rect 13460 -17528 14000 -17272
rect 13460 -17592 13704 -17528
rect 13768 -17592 14000 -17528
rect 13460 -17848 14000 -17592
rect 13460 -17912 13704 -17848
rect 13768 -17912 14000 -17848
rect 13460 -18168 14000 -17912
rect 13460 -18232 13704 -18168
rect 13768 -18232 14000 -18168
rect 13460 -18460 14000 -18232
rect 6000 -18488 14000 -18460
rect 6000 -18552 6238 -18488
rect 6302 -18552 13704 -18488
rect 13768 -18552 14000 -18488
rect 6000 -18698 14000 -18552
rect 6000 -18762 6608 -18698
rect 6672 -18762 6928 -18698
rect 6992 -18762 7248 -18698
rect 7312 -18762 7568 -18698
rect 7632 -18762 7888 -18698
rect 7952 -18762 8208 -18698
rect 8272 -18762 8528 -18698
rect 8592 -18762 8848 -18698
rect 8912 -18762 9168 -18698
rect 9232 -18762 9488 -18698
rect 9552 -18762 9808 -18698
rect 9872 -18762 10128 -18698
rect 10192 -18762 10448 -18698
rect 10512 -18762 10768 -18698
rect 10832 -18762 11088 -18698
rect 11152 -18762 11408 -18698
rect 11472 -18762 11728 -18698
rect 11792 -18762 12048 -18698
rect 12112 -18762 12368 -18698
rect 12432 -18762 12688 -18698
rect 12752 -18762 13008 -18698
rect 13072 -18762 13328 -18698
rect 13392 -18762 14000 -18698
rect 6000 -19000 14000 -18762
rect 14200 -12200 14500 -11520
rect 18000 -11540 26000 -11512
rect 18000 -11768 18540 -11540
rect 18000 -11832 18238 -11768
rect 18302 -11832 18540 -11768
rect 18000 -12088 18540 -11832
rect 18000 -12152 18238 -12088
rect 18302 -12152 18540 -12088
rect 14200 -19400 15000 -12200
rect 18000 -12408 18540 -12152
rect 18000 -12472 18238 -12408
rect 18302 -12472 18540 -12408
rect 18000 -12728 18540 -12472
rect 18000 -12792 18238 -12728
rect 18302 -12792 18540 -12728
rect 18000 -13048 18540 -12792
rect 18000 -13112 18238 -13048
rect 18302 -13112 18540 -13048
rect 18000 -13368 18540 -13112
rect 18000 -13432 18238 -13368
rect 18302 -13432 18540 -13368
rect 18000 -13688 18540 -13432
rect 18000 -13752 18238 -13688
rect 18302 -13752 18540 -13688
rect 18000 -14008 18540 -13752
rect 18000 -14072 18238 -14008
rect 18302 -14072 18540 -14008
rect 18000 -14328 18540 -14072
rect 18000 -14392 18238 -14328
rect 18302 -14392 18540 -14328
rect 18000 -14648 18540 -14392
rect 18000 -14712 18238 -14648
rect 18302 -14712 18540 -14648
rect 18000 -14968 18540 -14712
rect 18000 -15032 18238 -14968
rect 18302 -15032 18540 -14968
rect 18000 -15288 18540 -15032
rect 18000 -15352 18238 -15288
rect 18302 -15352 18540 -15288
rect 18000 -15608 18540 -15352
rect 18000 -15672 18238 -15608
rect 18302 -15672 18540 -15608
rect 18000 -15928 18540 -15672
rect 18000 -15992 18238 -15928
rect 18302 -15992 18540 -15928
rect 18000 -16248 18540 -15992
rect 18000 -16312 18238 -16248
rect 18302 -16312 18540 -16248
rect 18000 -16568 18540 -16312
rect 18000 -16632 18238 -16568
rect 18302 -16632 18540 -16568
rect 18000 -16888 18540 -16632
rect 18000 -16952 18238 -16888
rect 18302 -16952 18540 -16888
rect 18000 -17208 18540 -16952
rect 18000 -17272 18238 -17208
rect 18302 -17272 18540 -17208
rect 18000 -17528 18540 -17272
rect 18000 -17592 18238 -17528
rect 18302 -17592 18540 -17528
rect 18000 -17848 18540 -17592
rect 18000 -17912 18238 -17848
rect 18302 -17912 18540 -17848
rect 18000 -18168 18540 -17912
rect 18000 -18232 18238 -18168
rect 18302 -18232 18540 -18168
rect 18000 -18460 18540 -18232
rect 25460 -11768 26000 -11540
rect 25460 -11832 25704 -11768
rect 25768 -11832 26000 -11768
rect 25460 -12088 26000 -11832
rect 25460 -12152 25704 -12088
rect 25768 -12152 26000 -12088
rect 25460 -12408 26000 -12152
rect 25460 -12472 25704 -12408
rect 25768 -12472 26000 -12408
rect 25460 -12728 26000 -12472
rect 25460 -12792 25704 -12728
rect 25768 -12792 26000 -12728
rect 25460 -13048 26000 -12792
rect 25460 -13112 25704 -13048
rect 25768 -13112 26000 -13048
rect 25460 -13368 26000 -13112
rect 25460 -13432 25704 -13368
rect 25768 -13432 26000 -13368
rect 25460 -13688 26000 -13432
rect 25460 -13752 25704 -13688
rect 25768 -13752 26000 -13688
rect 25460 -14008 26000 -13752
rect 25460 -14072 25704 -14008
rect 25768 -14072 26000 -14008
rect 25460 -14328 26000 -14072
rect 25460 -14392 25704 -14328
rect 25768 -14392 26000 -14328
rect 25460 -14648 26000 -14392
rect 25460 -14712 25704 -14648
rect 25768 -14712 26000 -14648
rect 25460 -14968 26000 -14712
rect 25460 -15032 25704 -14968
rect 25768 -15032 26000 -14968
rect 25460 -15288 26000 -15032
rect 25460 -15352 25704 -15288
rect 25768 -15352 26000 -15288
rect 25460 -15608 26000 -15352
rect 25460 -15672 25704 -15608
rect 25768 -15672 26000 -15608
rect 25460 -15928 26000 -15672
rect 25460 -15992 25704 -15928
rect 25768 -15992 26000 -15928
rect 25460 -16248 26000 -15992
rect 25460 -16312 25704 -16248
rect 25768 -16312 26000 -16248
rect 25460 -16568 26000 -16312
rect 25460 -16632 25704 -16568
rect 25768 -16632 26000 -16568
rect 25460 -16888 26000 -16632
rect 25460 -16952 25704 -16888
rect 25768 -16952 26000 -16888
rect 25460 -17208 26000 -16952
rect 25460 -17272 25704 -17208
rect 25768 -17272 26000 -17208
rect 25460 -17528 26000 -17272
rect 25460 -17592 25704 -17528
rect 25768 -17592 26000 -17528
rect 25460 -17848 26000 -17592
rect 25460 -17912 25704 -17848
rect 25768 -17912 26000 -17848
rect 25460 -18168 26000 -17912
rect 25460 -18232 25704 -18168
rect 25768 -18232 26000 -18168
rect 25460 -18460 26000 -18232
rect 18000 -18488 26000 -18460
rect 18000 -18552 18238 -18488
rect 18302 -18552 25704 -18488
rect 25768 -18552 26000 -18488
rect 18000 -18698 26000 -18552
rect 18000 -18762 18608 -18698
rect 18672 -18762 18928 -18698
rect 18992 -18762 19248 -18698
rect 19312 -18762 19568 -18698
rect 19632 -18762 19888 -18698
rect 19952 -18762 20208 -18698
rect 20272 -18762 20528 -18698
rect 20592 -18762 20848 -18698
rect 20912 -18762 21168 -18698
rect 21232 -18762 21488 -18698
rect 21552 -18762 21808 -18698
rect 21872 -18762 22128 -18698
rect 22192 -18762 22448 -18698
rect 22512 -18762 22768 -18698
rect 22832 -18762 23088 -18698
rect 23152 -18762 23408 -18698
rect 23472 -18762 23728 -18698
rect 23792 -18762 24048 -18698
rect 24112 -18762 24368 -18698
rect 24432 -18762 24688 -18698
rect 24752 -18762 25008 -18698
rect 25072 -18762 25328 -18698
rect 25392 -18762 26000 -18698
rect 18000 -19000 26000 -18762
rect 30000 -11242 38000 -11000
rect 30000 -11306 30608 -11242
rect 30672 -11306 30928 -11242
rect 30992 -11306 31248 -11242
rect 31312 -11306 31568 -11242
rect 31632 -11306 31888 -11242
rect 31952 -11306 32208 -11242
rect 32272 -11306 32528 -11242
rect 32592 -11306 32848 -11242
rect 32912 -11306 33168 -11242
rect 33232 -11306 33488 -11242
rect 33552 -11306 33808 -11242
rect 33872 -11306 34128 -11242
rect 34192 -11306 34448 -11242
rect 34512 -11306 34768 -11242
rect 34832 -11306 35088 -11242
rect 35152 -11306 35408 -11242
rect 35472 -11306 35728 -11242
rect 35792 -11306 36048 -11242
rect 36112 -11306 36368 -11242
rect 36432 -11306 36688 -11242
rect 36752 -11306 37008 -11242
rect 37072 -11306 37328 -11242
rect 37392 -11306 38000 -11242
rect 30000 -11448 38000 -11306
rect 30000 -11512 30238 -11448
rect 30302 -11512 37704 -11448
rect 37768 -11512 38000 -11448
rect 30000 -11540 38000 -11512
rect 30000 -11768 30540 -11540
rect 30000 -11832 30238 -11768
rect 30302 -11832 30540 -11768
rect 30000 -12088 30540 -11832
rect 30000 -12152 30238 -12088
rect 30302 -12152 30540 -12088
rect 30000 -12408 30540 -12152
rect 30000 -12472 30238 -12408
rect 30302 -12472 30540 -12408
rect 30000 -12728 30540 -12472
rect 30000 -12792 30238 -12728
rect 30302 -12792 30540 -12728
rect 30000 -13048 30540 -12792
rect 30000 -13112 30238 -13048
rect 30302 -13112 30540 -13048
rect 30000 -13368 30540 -13112
rect 30000 -13432 30238 -13368
rect 30302 -13432 30540 -13368
rect 30000 -13688 30540 -13432
rect 30000 -13752 30238 -13688
rect 30302 -13752 30540 -13688
rect 30000 -14008 30540 -13752
rect 30000 -14072 30238 -14008
rect 30302 -14072 30540 -14008
rect 30000 -14328 30540 -14072
rect 30000 -14392 30238 -14328
rect 30302 -14392 30540 -14328
rect 30000 -14648 30540 -14392
rect 30000 -14712 30238 -14648
rect 30302 -14712 30540 -14648
rect 30000 -14968 30540 -14712
rect 30000 -15032 30238 -14968
rect 30302 -15032 30540 -14968
rect 30000 -15288 30540 -15032
rect 30000 -15352 30238 -15288
rect 30302 -15352 30540 -15288
rect 30000 -15608 30540 -15352
rect 30000 -15672 30238 -15608
rect 30302 -15672 30540 -15608
rect 30000 -15928 30540 -15672
rect 30000 -15992 30238 -15928
rect 30302 -15992 30540 -15928
rect 30000 -16248 30540 -15992
rect 30000 -16312 30238 -16248
rect 30302 -16312 30540 -16248
rect 30000 -16568 30540 -16312
rect 30000 -16632 30238 -16568
rect 30302 -16632 30540 -16568
rect 30000 -16888 30540 -16632
rect 30000 -16952 30238 -16888
rect 30302 -16952 30540 -16888
rect 30000 -17208 30540 -16952
rect 30000 -17272 30238 -17208
rect 30302 -17272 30540 -17208
rect 30000 -17528 30540 -17272
rect 30000 -17592 30238 -17528
rect 30302 -17592 30540 -17528
rect 30000 -17848 30540 -17592
rect 30000 -17912 30238 -17848
rect 30302 -17912 30540 -17848
rect 30000 -18168 30540 -17912
rect 30000 -18232 30238 -18168
rect 30302 -18232 30540 -18168
rect 30000 -18460 30540 -18232
rect 37460 -11768 38000 -11540
rect 37460 -11832 37704 -11768
rect 37768 -11832 38000 -11768
rect 37460 -12088 38000 -11832
rect 37460 -12152 37704 -12088
rect 37768 -12152 38000 -12088
rect 37460 -12408 38000 -12152
rect 37460 -12472 37704 -12408
rect 37768 -12472 38000 -12408
rect 37460 -12728 38000 -12472
rect 37460 -12792 37704 -12728
rect 37768 -12792 38000 -12728
rect 37460 -13048 38000 -12792
rect 37460 -13112 37704 -13048
rect 37768 -13112 38000 -13048
rect 37460 -13368 38000 -13112
rect 37460 -13432 37704 -13368
rect 37768 -13432 38000 -13368
rect 37460 -13688 38000 -13432
rect 37460 -13752 37704 -13688
rect 37768 -13752 38000 -13688
rect 37460 -14008 38000 -13752
rect 37460 -14072 37704 -14008
rect 37768 -14072 38000 -14008
rect 37460 -14328 38000 -14072
rect 37460 -14392 37704 -14328
rect 37768 -14392 38000 -14328
rect 37460 -14648 38000 -14392
rect 37460 -14712 37704 -14648
rect 37768 -14712 38000 -14648
rect 37460 -14968 38000 -14712
rect 37460 -15032 37704 -14968
rect 37768 -15032 38000 -14968
rect 37460 -15288 38000 -15032
rect 37460 -15352 37704 -15288
rect 37768 -15352 38000 -15288
rect 37460 -15608 38000 -15352
rect 37460 -15672 37704 -15608
rect 37768 -15672 38000 -15608
rect 37460 -15928 38000 -15672
rect 37460 -15992 37704 -15928
rect 37768 -15992 38000 -15928
rect 37460 -16248 38000 -15992
rect 37460 -16312 37704 -16248
rect 37768 -16312 38000 -16248
rect 37460 -16568 38000 -16312
rect 37460 -16632 37704 -16568
rect 37768 -16632 38000 -16568
rect 37460 -16888 38000 -16632
rect 37460 -16952 37704 -16888
rect 37768 -16952 38000 -16888
rect 37460 -17208 38000 -16952
rect 37460 -17272 37704 -17208
rect 37768 -17272 38000 -17208
rect 37460 -17528 38000 -17272
rect 37460 -17592 37704 -17528
rect 37768 -17592 38000 -17528
rect 37460 -17848 38000 -17592
rect 37460 -17912 37704 -17848
rect 37768 -17912 38000 -17848
rect 37460 -18168 38000 -17912
rect 37460 -18232 37704 -18168
rect 37768 -18232 38000 -18168
rect 37460 -18460 38000 -18232
rect 30000 -18488 38000 -18460
rect 30000 -18552 30238 -18488
rect 30302 -18552 37704 -18488
rect 37768 -18552 38000 -18488
rect 30000 -18698 38000 -18552
rect 30000 -18762 30608 -18698
rect 30672 -18762 30928 -18698
rect 30992 -18762 31248 -18698
rect 31312 -18762 31568 -18698
rect 31632 -18762 31888 -18698
rect 31952 -18762 32208 -18698
rect 32272 -18762 32528 -18698
rect 32592 -18762 32848 -18698
rect 32912 -18762 33168 -18698
rect 33232 -18762 33488 -18698
rect 33552 -18762 33808 -18698
rect 33872 -18762 34128 -18698
rect 34192 -18762 34448 -18698
rect 34512 -18762 34768 -18698
rect 34832 -18762 35088 -18698
rect 35152 -18762 35408 -18698
rect 35472 -18762 35728 -18698
rect 35792 -18762 36048 -18698
rect 36112 -18762 36368 -18698
rect 36432 -18762 36688 -18698
rect 36752 -18762 37008 -18698
rect 37072 -18762 37328 -18698
rect 37392 -18762 38000 -18698
rect 30000 -19000 38000 -18762
rect 42000 -11242 50000 -11000
rect 42000 -11306 42608 -11242
rect 42672 -11306 42928 -11242
rect 42992 -11306 43248 -11242
rect 43312 -11306 43568 -11242
rect 43632 -11306 43888 -11242
rect 43952 -11306 44208 -11242
rect 44272 -11306 44528 -11242
rect 44592 -11306 44848 -11242
rect 44912 -11306 45168 -11242
rect 45232 -11306 45488 -11242
rect 45552 -11306 45808 -11242
rect 45872 -11306 46128 -11242
rect 46192 -11306 46448 -11242
rect 46512 -11306 46768 -11242
rect 46832 -11306 47088 -11242
rect 47152 -11306 47408 -11242
rect 47472 -11306 47728 -11242
rect 47792 -11306 48048 -11242
rect 48112 -11306 48368 -11242
rect 48432 -11306 48688 -11242
rect 48752 -11306 49008 -11242
rect 49072 -11306 49328 -11242
rect 49392 -11306 50000 -11242
rect 42000 -11448 50000 -11306
rect 42000 -11512 42241 -11448
rect 42305 -11512 49695 -11448
rect 49759 -11512 50000 -11448
rect 42000 -11540 50000 -11512
rect 42000 -11768 42540 -11540
rect 42000 -11832 42241 -11768
rect 42305 -11832 42540 -11768
rect 42000 -12088 42540 -11832
rect 42000 -12152 42241 -12088
rect 42305 -12152 42540 -12088
rect 42000 -12408 42540 -12152
rect 42000 -12472 42241 -12408
rect 42305 -12472 42540 -12408
rect 42000 -12728 42540 -12472
rect 42000 -12792 42241 -12728
rect 42305 -12792 42540 -12728
rect 42000 -13048 42540 -12792
rect 42000 -13112 42241 -13048
rect 42305 -13112 42540 -13048
rect 42000 -13368 42540 -13112
rect 42000 -13432 42241 -13368
rect 42305 -13432 42540 -13368
rect 42000 -13688 42540 -13432
rect 42000 -13752 42241 -13688
rect 42305 -13752 42540 -13688
rect 42000 -14008 42540 -13752
rect 42000 -14072 42241 -14008
rect 42305 -14072 42540 -14008
rect 42000 -14328 42540 -14072
rect 42000 -14392 42241 -14328
rect 42305 -14392 42540 -14328
rect 42000 -14648 42540 -14392
rect 42000 -14712 42241 -14648
rect 42305 -14712 42540 -14648
rect 42000 -14968 42540 -14712
rect 42000 -15032 42241 -14968
rect 42305 -15032 42540 -14968
rect 42000 -15288 42540 -15032
rect 42000 -15352 42241 -15288
rect 42305 -15352 42540 -15288
rect 42000 -15608 42540 -15352
rect 42000 -15672 42241 -15608
rect 42305 -15672 42540 -15608
rect 42000 -15928 42540 -15672
rect 42000 -15992 42241 -15928
rect 42305 -15992 42540 -15928
rect 42000 -16248 42540 -15992
rect 42000 -16312 42241 -16248
rect 42305 -16312 42540 -16248
rect 42000 -16568 42540 -16312
rect 42000 -16632 42241 -16568
rect 42305 -16632 42540 -16568
rect 42000 -16888 42540 -16632
rect 42000 -16952 42241 -16888
rect 42305 -16952 42540 -16888
rect 42000 -17208 42540 -16952
rect 42000 -17272 42241 -17208
rect 42305 -17272 42540 -17208
rect 42000 -17528 42540 -17272
rect 42000 -17592 42241 -17528
rect 42305 -17592 42540 -17528
rect 42000 -17848 42540 -17592
rect 42000 -17912 42241 -17848
rect 42305 -17912 42540 -17848
rect 42000 -18168 42540 -17912
rect 42000 -18232 42241 -18168
rect 42305 -18232 42540 -18168
rect 42000 -18460 42540 -18232
rect 49460 -11768 50000 -11540
rect 49460 -11832 49695 -11768
rect 49759 -11832 50000 -11768
rect 49460 -12088 50000 -11832
rect 49460 -12152 49695 -12088
rect 49759 -12152 50000 -12088
rect 49460 -12408 50000 -12152
rect 49460 -12472 49695 -12408
rect 49759 -12472 50000 -12408
rect 49460 -12728 50000 -12472
rect 49460 -12792 49695 -12728
rect 49759 -12792 50000 -12728
rect 49460 -13048 50000 -12792
rect 49460 -13112 49695 -13048
rect 49759 -13112 50000 -13048
rect 49460 -13368 50000 -13112
rect 49460 -13432 49695 -13368
rect 49759 -13432 50000 -13368
rect 49460 -13688 50000 -13432
rect 49460 -13752 49695 -13688
rect 49759 -13752 50000 -13688
rect 49460 -14008 50000 -13752
rect 49460 -14072 49695 -14008
rect 49759 -14072 50000 -14008
rect 49460 -14328 50000 -14072
rect 49460 -14392 49695 -14328
rect 49759 -14392 50000 -14328
rect 49460 -14648 50000 -14392
rect 49460 -14712 49695 -14648
rect 49759 -14712 50000 -14648
rect 49460 -14968 50000 -14712
rect 49460 -15032 49695 -14968
rect 49759 -15032 50000 -14968
rect 49460 -15288 50000 -15032
rect 49460 -15352 49695 -15288
rect 49759 -15352 50000 -15288
rect 49460 -15608 50000 -15352
rect 49460 -15672 49695 -15608
rect 49759 -15672 50000 -15608
rect 49460 -15928 50000 -15672
rect 49460 -15992 49695 -15928
rect 49759 -15992 50000 -15928
rect 49460 -16248 50000 -15992
rect 49460 -16312 49695 -16248
rect 49759 -16312 50000 -16248
rect 49460 -16568 50000 -16312
rect 49460 -16632 49695 -16568
rect 49759 -16632 50000 -16568
rect 49460 -16888 50000 -16632
rect 49460 -16952 49695 -16888
rect 49759 -16952 50000 -16888
rect 49460 -17208 50000 -16952
rect 49460 -17272 49695 -17208
rect 49759 -17272 50000 -17208
rect 49460 -17528 50000 -17272
rect 49460 -17592 49695 -17528
rect 49759 -17592 50000 -17528
rect 49460 -17848 50000 -17592
rect 49460 -17912 49695 -17848
rect 49759 -17912 50000 -17848
rect 49460 -18168 50000 -17912
rect 49460 -18232 49695 -18168
rect 49759 -18232 50000 -18168
rect 49460 -18460 50000 -18232
rect 42000 -18488 50000 -18460
rect 42000 -18552 42241 -18488
rect 42305 -18552 49695 -18488
rect 49759 -18552 50000 -18488
rect 42000 -18698 50000 -18552
rect 42000 -18762 42608 -18698
rect 42672 -18762 42928 -18698
rect 42992 -18762 43248 -18698
rect 43312 -18762 43568 -18698
rect 43632 -18762 43888 -18698
rect 43952 -18762 44208 -18698
rect 44272 -18762 44528 -18698
rect 44592 -18762 44848 -18698
rect 44912 -18762 45168 -18698
rect 45232 -18762 45488 -18698
rect 45552 -18762 45808 -18698
rect 45872 -18762 46128 -18698
rect 46192 -18762 46448 -18698
rect 46512 -18762 46768 -18698
rect 46832 -18762 47088 -18698
rect 47152 -18762 47408 -18698
rect 47472 -18762 47728 -18698
rect 47792 -18762 48048 -18698
rect 48112 -18762 48368 -18698
rect 48432 -18762 48688 -18698
rect 48752 -18762 49008 -18698
rect 49072 -18762 49328 -18698
rect 49392 -18762 50000 -18698
rect 42000 -19000 50000 -18762
rect 14200 -19700 14300 -19400
rect 14900 -19700 15000 -19400
rect 14200 -21800 15000 -19700
<< via3 >>
rect 13960 3480 14060 3720
rect 20080 3140 20480 3280
rect 15180 2680 15360 2940
rect 20020 1460 20260 1760
rect 14940 -580 15140 -200
rect 14120 -1620 14260 -1100
rect 20380 -2200 20620 -1680
rect 21360 -9380 21840 -9260
rect 6608 -11246 6672 -11242
rect 6608 -11302 6612 -11246
rect 6612 -11302 6668 -11246
rect 6668 -11302 6672 -11246
rect 6608 -11306 6672 -11302
rect 6928 -11246 6992 -11242
rect 6928 -11302 6932 -11246
rect 6932 -11302 6988 -11246
rect 6988 -11302 6992 -11246
rect 6928 -11306 6992 -11302
rect 7248 -11246 7312 -11242
rect 7248 -11302 7252 -11246
rect 7252 -11302 7308 -11246
rect 7308 -11302 7312 -11246
rect 7248 -11306 7312 -11302
rect 7568 -11246 7632 -11242
rect 7568 -11302 7572 -11246
rect 7572 -11302 7628 -11246
rect 7628 -11302 7632 -11246
rect 7568 -11306 7632 -11302
rect 7888 -11246 7952 -11242
rect 7888 -11302 7892 -11246
rect 7892 -11302 7948 -11246
rect 7948 -11302 7952 -11246
rect 7888 -11306 7952 -11302
rect 8208 -11246 8272 -11242
rect 8208 -11302 8212 -11246
rect 8212 -11302 8268 -11246
rect 8268 -11302 8272 -11246
rect 8208 -11306 8272 -11302
rect 8528 -11246 8592 -11242
rect 8528 -11302 8532 -11246
rect 8532 -11302 8588 -11246
rect 8588 -11302 8592 -11246
rect 8528 -11306 8592 -11302
rect 8848 -11246 8912 -11242
rect 8848 -11302 8852 -11246
rect 8852 -11302 8908 -11246
rect 8908 -11302 8912 -11246
rect 8848 -11306 8912 -11302
rect 9168 -11246 9232 -11242
rect 9168 -11302 9172 -11246
rect 9172 -11302 9228 -11246
rect 9228 -11302 9232 -11246
rect 9168 -11306 9232 -11302
rect 9488 -11246 9552 -11242
rect 9488 -11302 9492 -11246
rect 9492 -11302 9548 -11246
rect 9548 -11302 9552 -11246
rect 9488 -11306 9552 -11302
rect 9808 -11246 9872 -11242
rect 9808 -11302 9812 -11246
rect 9812 -11302 9868 -11246
rect 9868 -11302 9872 -11246
rect 9808 -11306 9872 -11302
rect 10128 -11246 10192 -11242
rect 10128 -11302 10132 -11246
rect 10132 -11302 10188 -11246
rect 10188 -11302 10192 -11246
rect 10128 -11306 10192 -11302
rect 10448 -11246 10512 -11242
rect 10448 -11302 10452 -11246
rect 10452 -11302 10508 -11246
rect 10508 -11302 10512 -11246
rect 10448 -11306 10512 -11302
rect 10768 -11246 10832 -11242
rect 10768 -11302 10772 -11246
rect 10772 -11302 10828 -11246
rect 10828 -11302 10832 -11246
rect 10768 -11306 10832 -11302
rect 11088 -11246 11152 -11242
rect 11088 -11302 11092 -11246
rect 11092 -11302 11148 -11246
rect 11148 -11302 11152 -11246
rect 11088 -11306 11152 -11302
rect 11408 -11246 11472 -11242
rect 11408 -11302 11412 -11246
rect 11412 -11302 11468 -11246
rect 11468 -11302 11472 -11246
rect 11408 -11306 11472 -11302
rect 11728 -11246 11792 -11242
rect 11728 -11302 11732 -11246
rect 11732 -11302 11788 -11246
rect 11788 -11302 11792 -11246
rect 11728 -11306 11792 -11302
rect 12048 -11246 12112 -11242
rect 12048 -11302 12052 -11246
rect 12052 -11302 12108 -11246
rect 12108 -11302 12112 -11246
rect 12048 -11306 12112 -11302
rect 12368 -11246 12432 -11242
rect 12368 -11302 12372 -11246
rect 12372 -11302 12428 -11246
rect 12428 -11302 12432 -11246
rect 12368 -11306 12432 -11302
rect 12688 -11246 12752 -11242
rect 12688 -11302 12692 -11246
rect 12692 -11302 12748 -11246
rect 12748 -11302 12752 -11246
rect 12688 -11306 12752 -11302
rect 13008 -11246 13072 -11242
rect 13008 -11302 13012 -11246
rect 13012 -11302 13068 -11246
rect 13068 -11302 13072 -11246
rect 13008 -11306 13072 -11302
rect 13328 -11246 13392 -11242
rect 13328 -11302 13332 -11246
rect 13332 -11302 13388 -11246
rect 13388 -11302 13392 -11246
rect 13328 -11306 13392 -11302
rect 6238 -11452 6302 -11448
rect 6238 -11508 6242 -11452
rect 6242 -11508 6298 -11452
rect 6298 -11508 6302 -11452
rect 6238 -11512 6302 -11508
rect 13704 -11452 13768 -11448
rect 13704 -11508 13708 -11452
rect 13708 -11508 13764 -11452
rect 13764 -11508 13768 -11452
rect 13704 -11512 13768 -11508
rect 18608 -11246 18672 -11242
rect 18608 -11302 18612 -11246
rect 18612 -11302 18668 -11246
rect 18668 -11302 18672 -11246
rect 18608 -11306 18672 -11302
rect 18928 -11246 18992 -11242
rect 18928 -11302 18932 -11246
rect 18932 -11302 18988 -11246
rect 18988 -11302 18992 -11246
rect 18928 -11306 18992 -11302
rect 19248 -11246 19312 -11242
rect 19248 -11302 19252 -11246
rect 19252 -11302 19308 -11246
rect 19308 -11302 19312 -11246
rect 19248 -11306 19312 -11302
rect 19568 -11246 19632 -11242
rect 19568 -11302 19572 -11246
rect 19572 -11302 19628 -11246
rect 19628 -11302 19632 -11246
rect 19568 -11306 19632 -11302
rect 19888 -11246 19952 -11242
rect 19888 -11302 19892 -11246
rect 19892 -11302 19948 -11246
rect 19948 -11302 19952 -11246
rect 19888 -11306 19952 -11302
rect 20208 -11246 20272 -11242
rect 20208 -11302 20212 -11246
rect 20212 -11302 20268 -11246
rect 20268 -11302 20272 -11246
rect 20208 -11306 20272 -11302
rect 20528 -11246 20592 -11242
rect 20528 -11302 20532 -11246
rect 20532 -11302 20588 -11246
rect 20588 -11302 20592 -11246
rect 20528 -11306 20592 -11302
rect 20848 -11246 20912 -11242
rect 20848 -11302 20852 -11246
rect 20852 -11302 20908 -11246
rect 20908 -11302 20912 -11246
rect 20848 -11306 20912 -11302
rect 21168 -11246 21232 -11242
rect 21168 -11302 21172 -11246
rect 21172 -11302 21228 -11246
rect 21228 -11302 21232 -11246
rect 21168 -11306 21232 -11302
rect 21488 -11246 21552 -11242
rect 21488 -11302 21492 -11246
rect 21492 -11302 21548 -11246
rect 21548 -11302 21552 -11246
rect 21488 -11306 21552 -11302
rect 21808 -11246 21872 -11242
rect 21808 -11302 21812 -11246
rect 21812 -11302 21868 -11246
rect 21868 -11302 21872 -11246
rect 21808 -11306 21872 -11302
rect 22128 -11246 22192 -11242
rect 22128 -11302 22132 -11246
rect 22132 -11302 22188 -11246
rect 22188 -11302 22192 -11246
rect 22128 -11306 22192 -11302
rect 22448 -11246 22512 -11242
rect 22448 -11302 22452 -11246
rect 22452 -11302 22508 -11246
rect 22508 -11302 22512 -11246
rect 22448 -11306 22512 -11302
rect 22768 -11246 22832 -11242
rect 22768 -11302 22772 -11246
rect 22772 -11302 22828 -11246
rect 22828 -11302 22832 -11246
rect 22768 -11306 22832 -11302
rect 23088 -11246 23152 -11242
rect 23088 -11302 23092 -11246
rect 23092 -11302 23148 -11246
rect 23148 -11302 23152 -11246
rect 23088 -11306 23152 -11302
rect 23408 -11246 23472 -11242
rect 23408 -11302 23412 -11246
rect 23412 -11302 23468 -11246
rect 23468 -11302 23472 -11246
rect 23408 -11306 23472 -11302
rect 23728 -11246 23792 -11242
rect 23728 -11302 23732 -11246
rect 23732 -11302 23788 -11246
rect 23788 -11302 23792 -11246
rect 23728 -11306 23792 -11302
rect 24048 -11246 24112 -11242
rect 24048 -11302 24052 -11246
rect 24052 -11302 24108 -11246
rect 24108 -11302 24112 -11246
rect 24048 -11306 24112 -11302
rect 24368 -11246 24432 -11242
rect 24368 -11302 24372 -11246
rect 24372 -11302 24428 -11246
rect 24428 -11302 24432 -11246
rect 24368 -11306 24432 -11302
rect 24688 -11246 24752 -11242
rect 24688 -11302 24692 -11246
rect 24692 -11302 24748 -11246
rect 24748 -11302 24752 -11246
rect 24688 -11306 24752 -11302
rect 25008 -11246 25072 -11242
rect 25008 -11302 25012 -11246
rect 25012 -11302 25068 -11246
rect 25068 -11302 25072 -11246
rect 25008 -11306 25072 -11302
rect 25328 -11246 25392 -11242
rect 25328 -11302 25332 -11246
rect 25332 -11302 25388 -11246
rect 25388 -11302 25392 -11246
rect 25328 -11306 25392 -11302
rect 18238 -11452 18302 -11448
rect 18238 -11508 18242 -11452
rect 18242 -11508 18298 -11452
rect 18298 -11508 18302 -11452
rect 18238 -11512 18302 -11508
rect 25704 -11452 25768 -11448
rect 25704 -11508 25708 -11452
rect 25708 -11508 25764 -11452
rect 25764 -11508 25768 -11452
rect 25704 -11512 25768 -11508
rect 6238 -11772 6302 -11768
rect 6238 -11828 6242 -11772
rect 6242 -11828 6298 -11772
rect 6298 -11828 6302 -11772
rect 6238 -11832 6302 -11828
rect 6238 -12092 6302 -12088
rect 6238 -12148 6242 -12092
rect 6242 -12148 6298 -12092
rect 6298 -12148 6302 -12092
rect 6238 -12152 6302 -12148
rect 6238 -12412 6302 -12408
rect 6238 -12468 6242 -12412
rect 6242 -12468 6298 -12412
rect 6298 -12468 6302 -12412
rect 6238 -12472 6302 -12468
rect 6238 -12732 6302 -12728
rect 6238 -12788 6242 -12732
rect 6242 -12788 6298 -12732
rect 6298 -12788 6302 -12732
rect 6238 -12792 6302 -12788
rect 6238 -13052 6302 -13048
rect 6238 -13108 6242 -13052
rect 6242 -13108 6298 -13052
rect 6298 -13108 6302 -13052
rect 6238 -13112 6302 -13108
rect 6238 -13372 6302 -13368
rect 6238 -13428 6242 -13372
rect 6242 -13428 6298 -13372
rect 6298 -13428 6302 -13372
rect 6238 -13432 6302 -13428
rect 6238 -13692 6302 -13688
rect 6238 -13748 6242 -13692
rect 6242 -13748 6298 -13692
rect 6298 -13748 6302 -13692
rect 6238 -13752 6302 -13748
rect 6238 -14012 6302 -14008
rect 6238 -14068 6242 -14012
rect 6242 -14068 6298 -14012
rect 6298 -14068 6302 -14012
rect 6238 -14072 6302 -14068
rect 6238 -14332 6302 -14328
rect 6238 -14388 6242 -14332
rect 6242 -14388 6298 -14332
rect 6298 -14388 6302 -14332
rect 6238 -14392 6302 -14388
rect 6238 -14652 6302 -14648
rect 6238 -14708 6242 -14652
rect 6242 -14708 6298 -14652
rect 6298 -14708 6302 -14652
rect 6238 -14712 6302 -14708
rect 6238 -14972 6302 -14968
rect 6238 -15028 6242 -14972
rect 6242 -15028 6298 -14972
rect 6298 -15028 6302 -14972
rect 6238 -15032 6302 -15028
rect 6238 -15292 6302 -15288
rect 6238 -15348 6242 -15292
rect 6242 -15348 6298 -15292
rect 6298 -15348 6302 -15292
rect 6238 -15352 6302 -15348
rect 6238 -15612 6302 -15608
rect 6238 -15668 6242 -15612
rect 6242 -15668 6298 -15612
rect 6298 -15668 6302 -15612
rect 6238 -15672 6302 -15668
rect 6238 -15932 6302 -15928
rect 6238 -15988 6242 -15932
rect 6242 -15988 6298 -15932
rect 6298 -15988 6302 -15932
rect 6238 -15992 6302 -15988
rect 6238 -16252 6302 -16248
rect 6238 -16308 6242 -16252
rect 6242 -16308 6298 -16252
rect 6298 -16308 6302 -16252
rect 6238 -16312 6302 -16308
rect 6238 -16572 6302 -16568
rect 6238 -16628 6242 -16572
rect 6242 -16628 6298 -16572
rect 6298 -16628 6302 -16572
rect 6238 -16632 6302 -16628
rect 6238 -16892 6302 -16888
rect 6238 -16948 6242 -16892
rect 6242 -16948 6298 -16892
rect 6298 -16948 6302 -16892
rect 6238 -16952 6302 -16948
rect 6238 -17212 6302 -17208
rect 6238 -17268 6242 -17212
rect 6242 -17268 6298 -17212
rect 6298 -17268 6302 -17212
rect 6238 -17272 6302 -17268
rect 6238 -17532 6302 -17528
rect 6238 -17588 6242 -17532
rect 6242 -17588 6298 -17532
rect 6298 -17588 6302 -17532
rect 6238 -17592 6302 -17588
rect 6238 -17852 6302 -17848
rect 6238 -17908 6242 -17852
rect 6242 -17908 6298 -17852
rect 6298 -17908 6302 -17852
rect 6238 -17912 6302 -17908
rect 6238 -18172 6302 -18168
rect 6238 -18228 6242 -18172
rect 6242 -18228 6298 -18172
rect 6298 -18228 6302 -18172
rect 6238 -18232 6302 -18228
rect 13704 -11772 13768 -11768
rect 13704 -11828 13708 -11772
rect 13708 -11828 13764 -11772
rect 13764 -11828 13768 -11772
rect 13704 -11832 13768 -11828
rect 13704 -12092 13768 -12088
rect 13704 -12148 13708 -12092
rect 13708 -12148 13764 -12092
rect 13764 -12148 13768 -12092
rect 13704 -12152 13768 -12148
rect 13704 -12412 13768 -12408
rect 13704 -12468 13708 -12412
rect 13708 -12468 13764 -12412
rect 13764 -12468 13768 -12412
rect 13704 -12472 13768 -12468
rect 13704 -12732 13768 -12728
rect 13704 -12788 13708 -12732
rect 13708 -12788 13764 -12732
rect 13764 -12788 13768 -12732
rect 13704 -12792 13768 -12788
rect 13704 -13052 13768 -13048
rect 13704 -13108 13708 -13052
rect 13708 -13108 13764 -13052
rect 13764 -13108 13768 -13052
rect 13704 -13112 13768 -13108
rect 13704 -13372 13768 -13368
rect 13704 -13428 13708 -13372
rect 13708 -13428 13764 -13372
rect 13764 -13428 13768 -13372
rect 13704 -13432 13768 -13428
rect 13704 -13692 13768 -13688
rect 13704 -13748 13708 -13692
rect 13708 -13748 13764 -13692
rect 13764 -13748 13768 -13692
rect 13704 -13752 13768 -13748
rect 13704 -14012 13768 -14008
rect 13704 -14068 13708 -14012
rect 13708 -14068 13764 -14012
rect 13764 -14068 13768 -14012
rect 13704 -14072 13768 -14068
rect 13704 -14332 13768 -14328
rect 13704 -14388 13708 -14332
rect 13708 -14388 13764 -14332
rect 13764 -14388 13768 -14332
rect 13704 -14392 13768 -14388
rect 13704 -14652 13768 -14648
rect 13704 -14708 13708 -14652
rect 13708 -14708 13764 -14652
rect 13764 -14708 13768 -14652
rect 13704 -14712 13768 -14708
rect 13704 -14972 13768 -14968
rect 13704 -15028 13708 -14972
rect 13708 -15028 13764 -14972
rect 13764 -15028 13768 -14972
rect 13704 -15032 13768 -15028
rect 13704 -15292 13768 -15288
rect 13704 -15348 13708 -15292
rect 13708 -15348 13764 -15292
rect 13764 -15348 13768 -15292
rect 13704 -15352 13768 -15348
rect 13704 -15612 13768 -15608
rect 13704 -15668 13708 -15612
rect 13708 -15668 13764 -15612
rect 13764 -15668 13768 -15612
rect 13704 -15672 13768 -15668
rect 13704 -15932 13768 -15928
rect 13704 -15988 13708 -15932
rect 13708 -15988 13764 -15932
rect 13764 -15988 13768 -15932
rect 13704 -15992 13768 -15988
rect 13704 -16252 13768 -16248
rect 13704 -16308 13708 -16252
rect 13708 -16308 13764 -16252
rect 13764 -16308 13768 -16252
rect 13704 -16312 13768 -16308
rect 13704 -16572 13768 -16568
rect 13704 -16628 13708 -16572
rect 13708 -16628 13764 -16572
rect 13764 -16628 13768 -16572
rect 13704 -16632 13768 -16628
rect 13704 -16892 13768 -16888
rect 13704 -16948 13708 -16892
rect 13708 -16948 13764 -16892
rect 13764 -16948 13768 -16892
rect 13704 -16952 13768 -16948
rect 13704 -17212 13768 -17208
rect 13704 -17268 13708 -17212
rect 13708 -17268 13764 -17212
rect 13764 -17268 13768 -17212
rect 13704 -17272 13768 -17268
rect 13704 -17532 13768 -17528
rect 13704 -17588 13708 -17532
rect 13708 -17588 13764 -17532
rect 13764 -17588 13768 -17532
rect 13704 -17592 13768 -17588
rect 13704 -17852 13768 -17848
rect 13704 -17908 13708 -17852
rect 13708 -17908 13764 -17852
rect 13764 -17908 13768 -17852
rect 13704 -17912 13768 -17908
rect 13704 -18172 13768 -18168
rect 13704 -18228 13708 -18172
rect 13708 -18228 13764 -18172
rect 13764 -18228 13768 -18172
rect 13704 -18232 13768 -18228
rect 6238 -18492 6302 -18488
rect 6238 -18548 6242 -18492
rect 6242 -18548 6298 -18492
rect 6298 -18548 6302 -18492
rect 6238 -18552 6302 -18548
rect 13704 -18492 13768 -18488
rect 13704 -18548 13708 -18492
rect 13708 -18548 13764 -18492
rect 13764 -18548 13768 -18492
rect 13704 -18552 13768 -18548
rect 6608 -18702 6672 -18698
rect 6608 -18758 6612 -18702
rect 6612 -18758 6668 -18702
rect 6668 -18758 6672 -18702
rect 6608 -18762 6672 -18758
rect 6928 -18702 6992 -18698
rect 6928 -18758 6932 -18702
rect 6932 -18758 6988 -18702
rect 6988 -18758 6992 -18702
rect 6928 -18762 6992 -18758
rect 7248 -18702 7312 -18698
rect 7248 -18758 7252 -18702
rect 7252 -18758 7308 -18702
rect 7308 -18758 7312 -18702
rect 7248 -18762 7312 -18758
rect 7568 -18702 7632 -18698
rect 7568 -18758 7572 -18702
rect 7572 -18758 7628 -18702
rect 7628 -18758 7632 -18702
rect 7568 -18762 7632 -18758
rect 7888 -18702 7952 -18698
rect 7888 -18758 7892 -18702
rect 7892 -18758 7948 -18702
rect 7948 -18758 7952 -18702
rect 7888 -18762 7952 -18758
rect 8208 -18702 8272 -18698
rect 8208 -18758 8212 -18702
rect 8212 -18758 8268 -18702
rect 8268 -18758 8272 -18702
rect 8208 -18762 8272 -18758
rect 8528 -18702 8592 -18698
rect 8528 -18758 8532 -18702
rect 8532 -18758 8588 -18702
rect 8588 -18758 8592 -18702
rect 8528 -18762 8592 -18758
rect 8848 -18702 8912 -18698
rect 8848 -18758 8852 -18702
rect 8852 -18758 8908 -18702
rect 8908 -18758 8912 -18702
rect 8848 -18762 8912 -18758
rect 9168 -18702 9232 -18698
rect 9168 -18758 9172 -18702
rect 9172 -18758 9228 -18702
rect 9228 -18758 9232 -18702
rect 9168 -18762 9232 -18758
rect 9488 -18702 9552 -18698
rect 9488 -18758 9492 -18702
rect 9492 -18758 9548 -18702
rect 9548 -18758 9552 -18702
rect 9488 -18762 9552 -18758
rect 9808 -18702 9872 -18698
rect 9808 -18758 9812 -18702
rect 9812 -18758 9868 -18702
rect 9868 -18758 9872 -18702
rect 9808 -18762 9872 -18758
rect 10128 -18702 10192 -18698
rect 10128 -18758 10132 -18702
rect 10132 -18758 10188 -18702
rect 10188 -18758 10192 -18702
rect 10128 -18762 10192 -18758
rect 10448 -18702 10512 -18698
rect 10448 -18758 10452 -18702
rect 10452 -18758 10508 -18702
rect 10508 -18758 10512 -18702
rect 10448 -18762 10512 -18758
rect 10768 -18702 10832 -18698
rect 10768 -18758 10772 -18702
rect 10772 -18758 10828 -18702
rect 10828 -18758 10832 -18702
rect 10768 -18762 10832 -18758
rect 11088 -18702 11152 -18698
rect 11088 -18758 11092 -18702
rect 11092 -18758 11148 -18702
rect 11148 -18758 11152 -18702
rect 11088 -18762 11152 -18758
rect 11408 -18702 11472 -18698
rect 11408 -18758 11412 -18702
rect 11412 -18758 11468 -18702
rect 11468 -18758 11472 -18702
rect 11408 -18762 11472 -18758
rect 11728 -18702 11792 -18698
rect 11728 -18758 11732 -18702
rect 11732 -18758 11788 -18702
rect 11788 -18758 11792 -18702
rect 11728 -18762 11792 -18758
rect 12048 -18702 12112 -18698
rect 12048 -18758 12052 -18702
rect 12052 -18758 12108 -18702
rect 12108 -18758 12112 -18702
rect 12048 -18762 12112 -18758
rect 12368 -18702 12432 -18698
rect 12368 -18758 12372 -18702
rect 12372 -18758 12428 -18702
rect 12428 -18758 12432 -18702
rect 12368 -18762 12432 -18758
rect 12688 -18702 12752 -18698
rect 12688 -18758 12692 -18702
rect 12692 -18758 12748 -18702
rect 12748 -18758 12752 -18702
rect 12688 -18762 12752 -18758
rect 13008 -18702 13072 -18698
rect 13008 -18758 13012 -18702
rect 13012 -18758 13068 -18702
rect 13068 -18758 13072 -18702
rect 13008 -18762 13072 -18758
rect 13328 -18702 13392 -18698
rect 13328 -18758 13332 -18702
rect 13332 -18758 13388 -18702
rect 13388 -18758 13392 -18702
rect 13328 -18762 13392 -18758
rect 18238 -11772 18302 -11768
rect 18238 -11828 18242 -11772
rect 18242 -11828 18298 -11772
rect 18298 -11828 18302 -11772
rect 18238 -11832 18302 -11828
rect 18238 -12092 18302 -12088
rect 18238 -12148 18242 -12092
rect 18242 -12148 18298 -12092
rect 18298 -12148 18302 -12092
rect 18238 -12152 18302 -12148
rect 18238 -12412 18302 -12408
rect 18238 -12468 18242 -12412
rect 18242 -12468 18298 -12412
rect 18298 -12468 18302 -12412
rect 18238 -12472 18302 -12468
rect 18238 -12732 18302 -12728
rect 18238 -12788 18242 -12732
rect 18242 -12788 18298 -12732
rect 18298 -12788 18302 -12732
rect 18238 -12792 18302 -12788
rect 18238 -13052 18302 -13048
rect 18238 -13108 18242 -13052
rect 18242 -13108 18298 -13052
rect 18298 -13108 18302 -13052
rect 18238 -13112 18302 -13108
rect 18238 -13372 18302 -13368
rect 18238 -13428 18242 -13372
rect 18242 -13428 18298 -13372
rect 18298 -13428 18302 -13372
rect 18238 -13432 18302 -13428
rect 18238 -13692 18302 -13688
rect 18238 -13748 18242 -13692
rect 18242 -13748 18298 -13692
rect 18298 -13748 18302 -13692
rect 18238 -13752 18302 -13748
rect 18238 -14012 18302 -14008
rect 18238 -14068 18242 -14012
rect 18242 -14068 18298 -14012
rect 18298 -14068 18302 -14012
rect 18238 -14072 18302 -14068
rect 18238 -14332 18302 -14328
rect 18238 -14388 18242 -14332
rect 18242 -14388 18298 -14332
rect 18298 -14388 18302 -14332
rect 18238 -14392 18302 -14388
rect 18238 -14652 18302 -14648
rect 18238 -14708 18242 -14652
rect 18242 -14708 18298 -14652
rect 18298 -14708 18302 -14652
rect 18238 -14712 18302 -14708
rect 18238 -14972 18302 -14968
rect 18238 -15028 18242 -14972
rect 18242 -15028 18298 -14972
rect 18298 -15028 18302 -14972
rect 18238 -15032 18302 -15028
rect 18238 -15292 18302 -15288
rect 18238 -15348 18242 -15292
rect 18242 -15348 18298 -15292
rect 18298 -15348 18302 -15292
rect 18238 -15352 18302 -15348
rect 18238 -15612 18302 -15608
rect 18238 -15668 18242 -15612
rect 18242 -15668 18298 -15612
rect 18298 -15668 18302 -15612
rect 18238 -15672 18302 -15668
rect 18238 -15932 18302 -15928
rect 18238 -15988 18242 -15932
rect 18242 -15988 18298 -15932
rect 18298 -15988 18302 -15932
rect 18238 -15992 18302 -15988
rect 18238 -16252 18302 -16248
rect 18238 -16308 18242 -16252
rect 18242 -16308 18298 -16252
rect 18298 -16308 18302 -16252
rect 18238 -16312 18302 -16308
rect 18238 -16572 18302 -16568
rect 18238 -16628 18242 -16572
rect 18242 -16628 18298 -16572
rect 18298 -16628 18302 -16572
rect 18238 -16632 18302 -16628
rect 18238 -16892 18302 -16888
rect 18238 -16948 18242 -16892
rect 18242 -16948 18298 -16892
rect 18298 -16948 18302 -16892
rect 18238 -16952 18302 -16948
rect 18238 -17212 18302 -17208
rect 18238 -17268 18242 -17212
rect 18242 -17268 18298 -17212
rect 18298 -17268 18302 -17212
rect 18238 -17272 18302 -17268
rect 18238 -17532 18302 -17528
rect 18238 -17588 18242 -17532
rect 18242 -17588 18298 -17532
rect 18298 -17588 18302 -17532
rect 18238 -17592 18302 -17588
rect 18238 -17852 18302 -17848
rect 18238 -17908 18242 -17852
rect 18242 -17908 18298 -17852
rect 18298 -17908 18302 -17852
rect 18238 -17912 18302 -17908
rect 18238 -18172 18302 -18168
rect 18238 -18228 18242 -18172
rect 18242 -18228 18298 -18172
rect 18298 -18228 18302 -18172
rect 18238 -18232 18302 -18228
rect 25704 -11772 25768 -11768
rect 25704 -11828 25708 -11772
rect 25708 -11828 25764 -11772
rect 25764 -11828 25768 -11772
rect 25704 -11832 25768 -11828
rect 25704 -12092 25768 -12088
rect 25704 -12148 25708 -12092
rect 25708 -12148 25764 -12092
rect 25764 -12148 25768 -12092
rect 25704 -12152 25768 -12148
rect 25704 -12412 25768 -12408
rect 25704 -12468 25708 -12412
rect 25708 -12468 25764 -12412
rect 25764 -12468 25768 -12412
rect 25704 -12472 25768 -12468
rect 25704 -12732 25768 -12728
rect 25704 -12788 25708 -12732
rect 25708 -12788 25764 -12732
rect 25764 -12788 25768 -12732
rect 25704 -12792 25768 -12788
rect 25704 -13052 25768 -13048
rect 25704 -13108 25708 -13052
rect 25708 -13108 25764 -13052
rect 25764 -13108 25768 -13052
rect 25704 -13112 25768 -13108
rect 25704 -13372 25768 -13368
rect 25704 -13428 25708 -13372
rect 25708 -13428 25764 -13372
rect 25764 -13428 25768 -13372
rect 25704 -13432 25768 -13428
rect 25704 -13692 25768 -13688
rect 25704 -13748 25708 -13692
rect 25708 -13748 25764 -13692
rect 25764 -13748 25768 -13692
rect 25704 -13752 25768 -13748
rect 25704 -14012 25768 -14008
rect 25704 -14068 25708 -14012
rect 25708 -14068 25764 -14012
rect 25764 -14068 25768 -14012
rect 25704 -14072 25768 -14068
rect 25704 -14332 25768 -14328
rect 25704 -14388 25708 -14332
rect 25708 -14388 25764 -14332
rect 25764 -14388 25768 -14332
rect 25704 -14392 25768 -14388
rect 25704 -14652 25768 -14648
rect 25704 -14708 25708 -14652
rect 25708 -14708 25764 -14652
rect 25764 -14708 25768 -14652
rect 25704 -14712 25768 -14708
rect 25704 -14972 25768 -14968
rect 25704 -15028 25708 -14972
rect 25708 -15028 25764 -14972
rect 25764 -15028 25768 -14972
rect 25704 -15032 25768 -15028
rect 25704 -15292 25768 -15288
rect 25704 -15348 25708 -15292
rect 25708 -15348 25764 -15292
rect 25764 -15348 25768 -15292
rect 25704 -15352 25768 -15348
rect 25704 -15612 25768 -15608
rect 25704 -15668 25708 -15612
rect 25708 -15668 25764 -15612
rect 25764 -15668 25768 -15612
rect 25704 -15672 25768 -15668
rect 25704 -15932 25768 -15928
rect 25704 -15988 25708 -15932
rect 25708 -15988 25764 -15932
rect 25764 -15988 25768 -15932
rect 25704 -15992 25768 -15988
rect 25704 -16252 25768 -16248
rect 25704 -16308 25708 -16252
rect 25708 -16308 25764 -16252
rect 25764 -16308 25768 -16252
rect 25704 -16312 25768 -16308
rect 25704 -16572 25768 -16568
rect 25704 -16628 25708 -16572
rect 25708 -16628 25764 -16572
rect 25764 -16628 25768 -16572
rect 25704 -16632 25768 -16628
rect 25704 -16892 25768 -16888
rect 25704 -16948 25708 -16892
rect 25708 -16948 25764 -16892
rect 25764 -16948 25768 -16892
rect 25704 -16952 25768 -16948
rect 25704 -17212 25768 -17208
rect 25704 -17268 25708 -17212
rect 25708 -17268 25764 -17212
rect 25764 -17268 25768 -17212
rect 25704 -17272 25768 -17268
rect 25704 -17532 25768 -17528
rect 25704 -17588 25708 -17532
rect 25708 -17588 25764 -17532
rect 25764 -17588 25768 -17532
rect 25704 -17592 25768 -17588
rect 25704 -17852 25768 -17848
rect 25704 -17908 25708 -17852
rect 25708 -17908 25764 -17852
rect 25764 -17908 25768 -17852
rect 25704 -17912 25768 -17908
rect 25704 -18172 25768 -18168
rect 25704 -18228 25708 -18172
rect 25708 -18228 25764 -18172
rect 25764 -18228 25768 -18172
rect 25704 -18232 25768 -18228
rect 18238 -18492 18302 -18488
rect 18238 -18548 18242 -18492
rect 18242 -18548 18298 -18492
rect 18298 -18548 18302 -18492
rect 18238 -18552 18302 -18548
rect 25704 -18492 25768 -18488
rect 25704 -18548 25708 -18492
rect 25708 -18548 25764 -18492
rect 25764 -18548 25768 -18492
rect 25704 -18552 25768 -18548
rect 18608 -18702 18672 -18698
rect 18608 -18758 18612 -18702
rect 18612 -18758 18668 -18702
rect 18668 -18758 18672 -18702
rect 18608 -18762 18672 -18758
rect 18928 -18702 18992 -18698
rect 18928 -18758 18932 -18702
rect 18932 -18758 18988 -18702
rect 18988 -18758 18992 -18702
rect 18928 -18762 18992 -18758
rect 19248 -18702 19312 -18698
rect 19248 -18758 19252 -18702
rect 19252 -18758 19308 -18702
rect 19308 -18758 19312 -18702
rect 19248 -18762 19312 -18758
rect 19568 -18702 19632 -18698
rect 19568 -18758 19572 -18702
rect 19572 -18758 19628 -18702
rect 19628 -18758 19632 -18702
rect 19568 -18762 19632 -18758
rect 19888 -18702 19952 -18698
rect 19888 -18758 19892 -18702
rect 19892 -18758 19948 -18702
rect 19948 -18758 19952 -18702
rect 19888 -18762 19952 -18758
rect 20208 -18702 20272 -18698
rect 20208 -18758 20212 -18702
rect 20212 -18758 20268 -18702
rect 20268 -18758 20272 -18702
rect 20208 -18762 20272 -18758
rect 20528 -18702 20592 -18698
rect 20528 -18758 20532 -18702
rect 20532 -18758 20588 -18702
rect 20588 -18758 20592 -18702
rect 20528 -18762 20592 -18758
rect 20848 -18702 20912 -18698
rect 20848 -18758 20852 -18702
rect 20852 -18758 20908 -18702
rect 20908 -18758 20912 -18702
rect 20848 -18762 20912 -18758
rect 21168 -18702 21232 -18698
rect 21168 -18758 21172 -18702
rect 21172 -18758 21228 -18702
rect 21228 -18758 21232 -18702
rect 21168 -18762 21232 -18758
rect 21488 -18702 21552 -18698
rect 21488 -18758 21492 -18702
rect 21492 -18758 21548 -18702
rect 21548 -18758 21552 -18702
rect 21488 -18762 21552 -18758
rect 21808 -18702 21872 -18698
rect 21808 -18758 21812 -18702
rect 21812 -18758 21868 -18702
rect 21868 -18758 21872 -18702
rect 21808 -18762 21872 -18758
rect 22128 -18702 22192 -18698
rect 22128 -18758 22132 -18702
rect 22132 -18758 22188 -18702
rect 22188 -18758 22192 -18702
rect 22128 -18762 22192 -18758
rect 22448 -18702 22512 -18698
rect 22448 -18758 22452 -18702
rect 22452 -18758 22508 -18702
rect 22508 -18758 22512 -18702
rect 22448 -18762 22512 -18758
rect 22768 -18702 22832 -18698
rect 22768 -18758 22772 -18702
rect 22772 -18758 22828 -18702
rect 22828 -18758 22832 -18702
rect 22768 -18762 22832 -18758
rect 23088 -18702 23152 -18698
rect 23088 -18758 23092 -18702
rect 23092 -18758 23148 -18702
rect 23148 -18758 23152 -18702
rect 23088 -18762 23152 -18758
rect 23408 -18702 23472 -18698
rect 23408 -18758 23412 -18702
rect 23412 -18758 23468 -18702
rect 23468 -18758 23472 -18702
rect 23408 -18762 23472 -18758
rect 23728 -18702 23792 -18698
rect 23728 -18758 23732 -18702
rect 23732 -18758 23788 -18702
rect 23788 -18758 23792 -18702
rect 23728 -18762 23792 -18758
rect 24048 -18702 24112 -18698
rect 24048 -18758 24052 -18702
rect 24052 -18758 24108 -18702
rect 24108 -18758 24112 -18702
rect 24048 -18762 24112 -18758
rect 24368 -18702 24432 -18698
rect 24368 -18758 24372 -18702
rect 24372 -18758 24428 -18702
rect 24428 -18758 24432 -18702
rect 24368 -18762 24432 -18758
rect 24688 -18702 24752 -18698
rect 24688 -18758 24692 -18702
rect 24692 -18758 24748 -18702
rect 24748 -18758 24752 -18702
rect 24688 -18762 24752 -18758
rect 25008 -18702 25072 -18698
rect 25008 -18758 25012 -18702
rect 25012 -18758 25068 -18702
rect 25068 -18758 25072 -18702
rect 25008 -18762 25072 -18758
rect 25328 -18702 25392 -18698
rect 25328 -18758 25332 -18702
rect 25332 -18758 25388 -18702
rect 25388 -18758 25392 -18702
rect 25328 -18762 25392 -18758
rect 30608 -11246 30672 -11242
rect 30608 -11302 30612 -11246
rect 30612 -11302 30668 -11246
rect 30668 -11302 30672 -11246
rect 30608 -11306 30672 -11302
rect 30928 -11246 30992 -11242
rect 30928 -11302 30932 -11246
rect 30932 -11302 30988 -11246
rect 30988 -11302 30992 -11246
rect 30928 -11306 30992 -11302
rect 31248 -11246 31312 -11242
rect 31248 -11302 31252 -11246
rect 31252 -11302 31308 -11246
rect 31308 -11302 31312 -11246
rect 31248 -11306 31312 -11302
rect 31568 -11246 31632 -11242
rect 31568 -11302 31572 -11246
rect 31572 -11302 31628 -11246
rect 31628 -11302 31632 -11246
rect 31568 -11306 31632 -11302
rect 31888 -11246 31952 -11242
rect 31888 -11302 31892 -11246
rect 31892 -11302 31948 -11246
rect 31948 -11302 31952 -11246
rect 31888 -11306 31952 -11302
rect 32208 -11246 32272 -11242
rect 32208 -11302 32212 -11246
rect 32212 -11302 32268 -11246
rect 32268 -11302 32272 -11246
rect 32208 -11306 32272 -11302
rect 32528 -11246 32592 -11242
rect 32528 -11302 32532 -11246
rect 32532 -11302 32588 -11246
rect 32588 -11302 32592 -11246
rect 32528 -11306 32592 -11302
rect 32848 -11246 32912 -11242
rect 32848 -11302 32852 -11246
rect 32852 -11302 32908 -11246
rect 32908 -11302 32912 -11246
rect 32848 -11306 32912 -11302
rect 33168 -11246 33232 -11242
rect 33168 -11302 33172 -11246
rect 33172 -11302 33228 -11246
rect 33228 -11302 33232 -11246
rect 33168 -11306 33232 -11302
rect 33488 -11246 33552 -11242
rect 33488 -11302 33492 -11246
rect 33492 -11302 33548 -11246
rect 33548 -11302 33552 -11246
rect 33488 -11306 33552 -11302
rect 33808 -11246 33872 -11242
rect 33808 -11302 33812 -11246
rect 33812 -11302 33868 -11246
rect 33868 -11302 33872 -11246
rect 33808 -11306 33872 -11302
rect 34128 -11246 34192 -11242
rect 34128 -11302 34132 -11246
rect 34132 -11302 34188 -11246
rect 34188 -11302 34192 -11246
rect 34128 -11306 34192 -11302
rect 34448 -11246 34512 -11242
rect 34448 -11302 34452 -11246
rect 34452 -11302 34508 -11246
rect 34508 -11302 34512 -11246
rect 34448 -11306 34512 -11302
rect 34768 -11246 34832 -11242
rect 34768 -11302 34772 -11246
rect 34772 -11302 34828 -11246
rect 34828 -11302 34832 -11246
rect 34768 -11306 34832 -11302
rect 35088 -11246 35152 -11242
rect 35088 -11302 35092 -11246
rect 35092 -11302 35148 -11246
rect 35148 -11302 35152 -11246
rect 35088 -11306 35152 -11302
rect 35408 -11246 35472 -11242
rect 35408 -11302 35412 -11246
rect 35412 -11302 35468 -11246
rect 35468 -11302 35472 -11246
rect 35408 -11306 35472 -11302
rect 35728 -11246 35792 -11242
rect 35728 -11302 35732 -11246
rect 35732 -11302 35788 -11246
rect 35788 -11302 35792 -11246
rect 35728 -11306 35792 -11302
rect 36048 -11246 36112 -11242
rect 36048 -11302 36052 -11246
rect 36052 -11302 36108 -11246
rect 36108 -11302 36112 -11246
rect 36048 -11306 36112 -11302
rect 36368 -11246 36432 -11242
rect 36368 -11302 36372 -11246
rect 36372 -11302 36428 -11246
rect 36428 -11302 36432 -11246
rect 36368 -11306 36432 -11302
rect 36688 -11246 36752 -11242
rect 36688 -11302 36692 -11246
rect 36692 -11302 36748 -11246
rect 36748 -11302 36752 -11246
rect 36688 -11306 36752 -11302
rect 37008 -11246 37072 -11242
rect 37008 -11302 37012 -11246
rect 37012 -11302 37068 -11246
rect 37068 -11302 37072 -11246
rect 37008 -11306 37072 -11302
rect 37328 -11246 37392 -11242
rect 37328 -11302 37332 -11246
rect 37332 -11302 37388 -11246
rect 37388 -11302 37392 -11246
rect 37328 -11306 37392 -11302
rect 30238 -11452 30302 -11448
rect 30238 -11508 30242 -11452
rect 30242 -11508 30298 -11452
rect 30298 -11508 30302 -11452
rect 30238 -11512 30302 -11508
rect 37704 -11452 37768 -11448
rect 37704 -11508 37708 -11452
rect 37708 -11508 37764 -11452
rect 37764 -11508 37768 -11452
rect 37704 -11512 37768 -11508
rect 30238 -11772 30302 -11768
rect 30238 -11828 30242 -11772
rect 30242 -11828 30298 -11772
rect 30298 -11828 30302 -11772
rect 30238 -11832 30302 -11828
rect 30238 -12092 30302 -12088
rect 30238 -12148 30242 -12092
rect 30242 -12148 30298 -12092
rect 30298 -12148 30302 -12092
rect 30238 -12152 30302 -12148
rect 30238 -12412 30302 -12408
rect 30238 -12468 30242 -12412
rect 30242 -12468 30298 -12412
rect 30298 -12468 30302 -12412
rect 30238 -12472 30302 -12468
rect 30238 -12732 30302 -12728
rect 30238 -12788 30242 -12732
rect 30242 -12788 30298 -12732
rect 30298 -12788 30302 -12732
rect 30238 -12792 30302 -12788
rect 30238 -13052 30302 -13048
rect 30238 -13108 30242 -13052
rect 30242 -13108 30298 -13052
rect 30298 -13108 30302 -13052
rect 30238 -13112 30302 -13108
rect 30238 -13372 30302 -13368
rect 30238 -13428 30242 -13372
rect 30242 -13428 30298 -13372
rect 30298 -13428 30302 -13372
rect 30238 -13432 30302 -13428
rect 30238 -13692 30302 -13688
rect 30238 -13748 30242 -13692
rect 30242 -13748 30298 -13692
rect 30298 -13748 30302 -13692
rect 30238 -13752 30302 -13748
rect 30238 -14012 30302 -14008
rect 30238 -14068 30242 -14012
rect 30242 -14068 30298 -14012
rect 30298 -14068 30302 -14012
rect 30238 -14072 30302 -14068
rect 30238 -14332 30302 -14328
rect 30238 -14388 30242 -14332
rect 30242 -14388 30298 -14332
rect 30298 -14388 30302 -14332
rect 30238 -14392 30302 -14388
rect 30238 -14652 30302 -14648
rect 30238 -14708 30242 -14652
rect 30242 -14708 30298 -14652
rect 30298 -14708 30302 -14652
rect 30238 -14712 30302 -14708
rect 30238 -14972 30302 -14968
rect 30238 -15028 30242 -14972
rect 30242 -15028 30298 -14972
rect 30298 -15028 30302 -14972
rect 30238 -15032 30302 -15028
rect 30238 -15292 30302 -15288
rect 30238 -15348 30242 -15292
rect 30242 -15348 30298 -15292
rect 30298 -15348 30302 -15292
rect 30238 -15352 30302 -15348
rect 30238 -15612 30302 -15608
rect 30238 -15668 30242 -15612
rect 30242 -15668 30298 -15612
rect 30298 -15668 30302 -15612
rect 30238 -15672 30302 -15668
rect 30238 -15932 30302 -15928
rect 30238 -15988 30242 -15932
rect 30242 -15988 30298 -15932
rect 30298 -15988 30302 -15932
rect 30238 -15992 30302 -15988
rect 30238 -16252 30302 -16248
rect 30238 -16308 30242 -16252
rect 30242 -16308 30298 -16252
rect 30298 -16308 30302 -16252
rect 30238 -16312 30302 -16308
rect 30238 -16572 30302 -16568
rect 30238 -16628 30242 -16572
rect 30242 -16628 30298 -16572
rect 30298 -16628 30302 -16572
rect 30238 -16632 30302 -16628
rect 30238 -16892 30302 -16888
rect 30238 -16948 30242 -16892
rect 30242 -16948 30298 -16892
rect 30298 -16948 30302 -16892
rect 30238 -16952 30302 -16948
rect 30238 -17212 30302 -17208
rect 30238 -17268 30242 -17212
rect 30242 -17268 30298 -17212
rect 30298 -17268 30302 -17212
rect 30238 -17272 30302 -17268
rect 30238 -17532 30302 -17528
rect 30238 -17588 30242 -17532
rect 30242 -17588 30298 -17532
rect 30298 -17588 30302 -17532
rect 30238 -17592 30302 -17588
rect 30238 -17852 30302 -17848
rect 30238 -17908 30242 -17852
rect 30242 -17908 30298 -17852
rect 30298 -17908 30302 -17852
rect 30238 -17912 30302 -17908
rect 30238 -18172 30302 -18168
rect 30238 -18228 30242 -18172
rect 30242 -18228 30298 -18172
rect 30298 -18228 30302 -18172
rect 30238 -18232 30302 -18228
rect 37704 -11772 37768 -11768
rect 37704 -11828 37708 -11772
rect 37708 -11828 37764 -11772
rect 37764 -11828 37768 -11772
rect 37704 -11832 37768 -11828
rect 37704 -12092 37768 -12088
rect 37704 -12148 37708 -12092
rect 37708 -12148 37764 -12092
rect 37764 -12148 37768 -12092
rect 37704 -12152 37768 -12148
rect 37704 -12412 37768 -12408
rect 37704 -12468 37708 -12412
rect 37708 -12468 37764 -12412
rect 37764 -12468 37768 -12412
rect 37704 -12472 37768 -12468
rect 37704 -12732 37768 -12728
rect 37704 -12788 37708 -12732
rect 37708 -12788 37764 -12732
rect 37764 -12788 37768 -12732
rect 37704 -12792 37768 -12788
rect 37704 -13052 37768 -13048
rect 37704 -13108 37708 -13052
rect 37708 -13108 37764 -13052
rect 37764 -13108 37768 -13052
rect 37704 -13112 37768 -13108
rect 37704 -13372 37768 -13368
rect 37704 -13428 37708 -13372
rect 37708 -13428 37764 -13372
rect 37764 -13428 37768 -13372
rect 37704 -13432 37768 -13428
rect 37704 -13692 37768 -13688
rect 37704 -13748 37708 -13692
rect 37708 -13748 37764 -13692
rect 37764 -13748 37768 -13692
rect 37704 -13752 37768 -13748
rect 37704 -14012 37768 -14008
rect 37704 -14068 37708 -14012
rect 37708 -14068 37764 -14012
rect 37764 -14068 37768 -14012
rect 37704 -14072 37768 -14068
rect 37704 -14332 37768 -14328
rect 37704 -14388 37708 -14332
rect 37708 -14388 37764 -14332
rect 37764 -14388 37768 -14332
rect 37704 -14392 37768 -14388
rect 37704 -14652 37768 -14648
rect 37704 -14708 37708 -14652
rect 37708 -14708 37764 -14652
rect 37764 -14708 37768 -14652
rect 37704 -14712 37768 -14708
rect 37704 -14972 37768 -14968
rect 37704 -15028 37708 -14972
rect 37708 -15028 37764 -14972
rect 37764 -15028 37768 -14972
rect 37704 -15032 37768 -15028
rect 37704 -15292 37768 -15288
rect 37704 -15348 37708 -15292
rect 37708 -15348 37764 -15292
rect 37764 -15348 37768 -15292
rect 37704 -15352 37768 -15348
rect 37704 -15612 37768 -15608
rect 37704 -15668 37708 -15612
rect 37708 -15668 37764 -15612
rect 37764 -15668 37768 -15612
rect 37704 -15672 37768 -15668
rect 37704 -15932 37768 -15928
rect 37704 -15988 37708 -15932
rect 37708 -15988 37764 -15932
rect 37764 -15988 37768 -15932
rect 37704 -15992 37768 -15988
rect 37704 -16252 37768 -16248
rect 37704 -16308 37708 -16252
rect 37708 -16308 37764 -16252
rect 37764 -16308 37768 -16252
rect 37704 -16312 37768 -16308
rect 37704 -16572 37768 -16568
rect 37704 -16628 37708 -16572
rect 37708 -16628 37764 -16572
rect 37764 -16628 37768 -16572
rect 37704 -16632 37768 -16628
rect 37704 -16892 37768 -16888
rect 37704 -16948 37708 -16892
rect 37708 -16948 37764 -16892
rect 37764 -16948 37768 -16892
rect 37704 -16952 37768 -16948
rect 37704 -17212 37768 -17208
rect 37704 -17268 37708 -17212
rect 37708 -17268 37764 -17212
rect 37764 -17268 37768 -17212
rect 37704 -17272 37768 -17268
rect 37704 -17532 37768 -17528
rect 37704 -17588 37708 -17532
rect 37708 -17588 37764 -17532
rect 37764 -17588 37768 -17532
rect 37704 -17592 37768 -17588
rect 37704 -17852 37768 -17848
rect 37704 -17908 37708 -17852
rect 37708 -17908 37764 -17852
rect 37764 -17908 37768 -17852
rect 37704 -17912 37768 -17908
rect 37704 -18172 37768 -18168
rect 37704 -18228 37708 -18172
rect 37708 -18228 37764 -18172
rect 37764 -18228 37768 -18172
rect 37704 -18232 37768 -18228
rect 30238 -18492 30302 -18488
rect 30238 -18548 30242 -18492
rect 30242 -18548 30298 -18492
rect 30298 -18548 30302 -18492
rect 30238 -18552 30302 -18548
rect 37704 -18492 37768 -18488
rect 37704 -18548 37708 -18492
rect 37708 -18548 37764 -18492
rect 37764 -18548 37768 -18492
rect 37704 -18552 37768 -18548
rect 30608 -18702 30672 -18698
rect 30608 -18758 30612 -18702
rect 30612 -18758 30668 -18702
rect 30668 -18758 30672 -18702
rect 30608 -18762 30672 -18758
rect 30928 -18702 30992 -18698
rect 30928 -18758 30932 -18702
rect 30932 -18758 30988 -18702
rect 30988 -18758 30992 -18702
rect 30928 -18762 30992 -18758
rect 31248 -18702 31312 -18698
rect 31248 -18758 31252 -18702
rect 31252 -18758 31308 -18702
rect 31308 -18758 31312 -18702
rect 31248 -18762 31312 -18758
rect 31568 -18702 31632 -18698
rect 31568 -18758 31572 -18702
rect 31572 -18758 31628 -18702
rect 31628 -18758 31632 -18702
rect 31568 -18762 31632 -18758
rect 31888 -18702 31952 -18698
rect 31888 -18758 31892 -18702
rect 31892 -18758 31948 -18702
rect 31948 -18758 31952 -18702
rect 31888 -18762 31952 -18758
rect 32208 -18702 32272 -18698
rect 32208 -18758 32212 -18702
rect 32212 -18758 32268 -18702
rect 32268 -18758 32272 -18702
rect 32208 -18762 32272 -18758
rect 32528 -18702 32592 -18698
rect 32528 -18758 32532 -18702
rect 32532 -18758 32588 -18702
rect 32588 -18758 32592 -18702
rect 32528 -18762 32592 -18758
rect 32848 -18702 32912 -18698
rect 32848 -18758 32852 -18702
rect 32852 -18758 32908 -18702
rect 32908 -18758 32912 -18702
rect 32848 -18762 32912 -18758
rect 33168 -18702 33232 -18698
rect 33168 -18758 33172 -18702
rect 33172 -18758 33228 -18702
rect 33228 -18758 33232 -18702
rect 33168 -18762 33232 -18758
rect 33488 -18702 33552 -18698
rect 33488 -18758 33492 -18702
rect 33492 -18758 33548 -18702
rect 33548 -18758 33552 -18702
rect 33488 -18762 33552 -18758
rect 33808 -18702 33872 -18698
rect 33808 -18758 33812 -18702
rect 33812 -18758 33868 -18702
rect 33868 -18758 33872 -18702
rect 33808 -18762 33872 -18758
rect 34128 -18702 34192 -18698
rect 34128 -18758 34132 -18702
rect 34132 -18758 34188 -18702
rect 34188 -18758 34192 -18702
rect 34128 -18762 34192 -18758
rect 34448 -18702 34512 -18698
rect 34448 -18758 34452 -18702
rect 34452 -18758 34508 -18702
rect 34508 -18758 34512 -18702
rect 34448 -18762 34512 -18758
rect 34768 -18702 34832 -18698
rect 34768 -18758 34772 -18702
rect 34772 -18758 34828 -18702
rect 34828 -18758 34832 -18702
rect 34768 -18762 34832 -18758
rect 35088 -18702 35152 -18698
rect 35088 -18758 35092 -18702
rect 35092 -18758 35148 -18702
rect 35148 -18758 35152 -18702
rect 35088 -18762 35152 -18758
rect 35408 -18702 35472 -18698
rect 35408 -18758 35412 -18702
rect 35412 -18758 35468 -18702
rect 35468 -18758 35472 -18702
rect 35408 -18762 35472 -18758
rect 35728 -18702 35792 -18698
rect 35728 -18758 35732 -18702
rect 35732 -18758 35788 -18702
rect 35788 -18758 35792 -18702
rect 35728 -18762 35792 -18758
rect 36048 -18702 36112 -18698
rect 36048 -18758 36052 -18702
rect 36052 -18758 36108 -18702
rect 36108 -18758 36112 -18702
rect 36048 -18762 36112 -18758
rect 36368 -18702 36432 -18698
rect 36368 -18758 36372 -18702
rect 36372 -18758 36428 -18702
rect 36428 -18758 36432 -18702
rect 36368 -18762 36432 -18758
rect 36688 -18702 36752 -18698
rect 36688 -18758 36692 -18702
rect 36692 -18758 36748 -18702
rect 36748 -18758 36752 -18702
rect 36688 -18762 36752 -18758
rect 37008 -18702 37072 -18698
rect 37008 -18758 37012 -18702
rect 37012 -18758 37068 -18702
rect 37068 -18758 37072 -18702
rect 37008 -18762 37072 -18758
rect 37328 -18702 37392 -18698
rect 37328 -18758 37332 -18702
rect 37332 -18758 37388 -18702
rect 37388 -18758 37392 -18702
rect 37328 -18762 37392 -18758
rect 42608 -11246 42672 -11242
rect 42608 -11302 42612 -11246
rect 42612 -11302 42668 -11246
rect 42668 -11302 42672 -11246
rect 42608 -11306 42672 -11302
rect 42928 -11246 42992 -11242
rect 42928 -11302 42932 -11246
rect 42932 -11302 42988 -11246
rect 42988 -11302 42992 -11246
rect 42928 -11306 42992 -11302
rect 43248 -11246 43312 -11242
rect 43248 -11302 43252 -11246
rect 43252 -11302 43308 -11246
rect 43308 -11302 43312 -11246
rect 43248 -11306 43312 -11302
rect 43568 -11246 43632 -11242
rect 43568 -11302 43572 -11246
rect 43572 -11302 43628 -11246
rect 43628 -11302 43632 -11246
rect 43568 -11306 43632 -11302
rect 43888 -11246 43952 -11242
rect 43888 -11302 43892 -11246
rect 43892 -11302 43948 -11246
rect 43948 -11302 43952 -11246
rect 43888 -11306 43952 -11302
rect 44208 -11246 44272 -11242
rect 44208 -11302 44212 -11246
rect 44212 -11302 44268 -11246
rect 44268 -11302 44272 -11246
rect 44208 -11306 44272 -11302
rect 44528 -11246 44592 -11242
rect 44528 -11302 44532 -11246
rect 44532 -11302 44588 -11246
rect 44588 -11302 44592 -11246
rect 44528 -11306 44592 -11302
rect 44848 -11246 44912 -11242
rect 44848 -11302 44852 -11246
rect 44852 -11302 44908 -11246
rect 44908 -11302 44912 -11246
rect 44848 -11306 44912 -11302
rect 45168 -11246 45232 -11242
rect 45168 -11302 45172 -11246
rect 45172 -11302 45228 -11246
rect 45228 -11302 45232 -11246
rect 45168 -11306 45232 -11302
rect 45488 -11246 45552 -11242
rect 45488 -11302 45492 -11246
rect 45492 -11302 45548 -11246
rect 45548 -11302 45552 -11246
rect 45488 -11306 45552 -11302
rect 45808 -11246 45872 -11242
rect 45808 -11302 45812 -11246
rect 45812 -11302 45868 -11246
rect 45868 -11302 45872 -11246
rect 45808 -11306 45872 -11302
rect 46128 -11246 46192 -11242
rect 46128 -11302 46132 -11246
rect 46132 -11302 46188 -11246
rect 46188 -11302 46192 -11246
rect 46128 -11306 46192 -11302
rect 46448 -11246 46512 -11242
rect 46448 -11302 46452 -11246
rect 46452 -11302 46508 -11246
rect 46508 -11302 46512 -11246
rect 46448 -11306 46512 -11302
rect 46768 -11246 46832 -11242
rect 46768 -11302 46772 -11246
rect 46772 -11302 46828 -11246
rect 46828 -11302 46832 -11246
rect 46768 -11306 46832 -11302
rect 47088 -11246 47152 -11242
rect 47088 -11302 47092 -11246
rect 47092 -11302 47148 -11246
rect 47148 -11302 47152 -11246
rect 47088 -11306 47152 -11302
rect 47408 -11246 47472 -11242
rect 47408 -11302 47412 -11246
rect 47412 -11302 47468 -11246
rect 47468 -11302 47472 -11246
rect 47408 -11306 47472 -11302
rect 47728 -11246 47792 -11242
rect 47728 -11302 47732 -11246
rect 47732 -11302 47788 -11246
rect 47788 -11302 47792 -11246
rect 47728 -11306 47792 -11302
rect 48048 -11246 48112 -11242
rect 48048 -11302 48052 -11246
rect 48052 -11302 48108 -11246
rect 48108 -11302 48112 -11246
rect 48048 -11306 48112 -11302
rect 48368 -11246 48432 -11242
rect 48368 -11302 48372 -11246
rect 48372 -11302 48428 -11246
rect 48428 -11302 48432 -11246
rect 48368 -11306 48432 -11302
rect 48688 -11246 48752 -11242
rect 48688 -11302 48692 -11246
rect 48692 -11302 48748 -11246
rect 48748 -11302 48752 -11246
rect 48688 -11306 48752 -11302
rect 49008 -11246 49072 -11242
rect 49008 -11302 49012 -11246
rect 49012 -11302 49068 -11246
rect 49068 -11302 49072 -11246
rect 49008 -11306 49072 -11302
rect 49328 -11246 49392 -11242
rect 49328 -11302 49332 -11246
rect 49332 -11302 49388 -11246
rect 49388 -11302 49392 -11246
rect 49328 -11306 49392 -11302
rect 42241 -11452 42305 -11448
rect 42241 -11508 42245 -11452
rect 42245 -11508 42301 -11452
rect 42301 -11508 42305 -11452
rect 42241 -11512 42305 -11508
rect 49695 -11452 49759 -11448
rect 49695 -11508 49699 -11452
rect 49699 -11508 49755 -11452
rect 49755 -11508 49759 -11452
rect 49695 -11512 49759 -11508
rect 42241 -11772 42305 -11768
rect 42241 -11828 42245 -11772
rect 42245 -11828 42301 -11772
rect 42301 -11828 42305 -11772
rect 42241 -11832 42305 -11828
rect 42241 -12092 42305 -12088
rect 42241 -12148 42245 -12092
rect 42245 -12148 42301 -12092
rect 42301 -12148 42305 -12092
rect 42241 -12152 42305 -12148
rect 42241 -12412 42305 -12408
rect 42241 -12468 42245 -12412
rect 42245 -12468 42301 -12412
rect 42301 -12468 42305 -12412
rect 42241 -12472 42305 -12468
rect 42241 -12732 42305 -12728
rect 42241 -12788 42245 -12732
rect 42245 -12788 42301 -12732
rect 42301 -12788 42305 -12732
rect 42241 -12792 42305 -12788
rect 42241 -13052 42305 -13048
rect 42241 -13108 42245 -13052
rect 42245 -13108 42301 -13052
rect 42301 -13108 42305 -13052
rect 42241 -13112 42305 -13108
rect 42241 -13372 42305 -13368
rect 42241 -13428 42245 -13372
rect 42245 -13428 42301 -13372
rect 42301 -13428 42305 -13372
rect 42241 -13432 42305 -13428
rect 42241 -13692 42305 -13688
rect 42241 -13748 42245 -13692
rect 42245 -13748 42301 -13692
rect 42301 -13748 42305 -13692
rect 42241 -13752 42305 -13748
rect 42241 -14012 42305 -14008
rect 42241 -14068 42245 -14012
rect 42245 -14068 42301 -14012
rect 42301 -14068 42305 -14012
rect 42241 -14072 42305 -14068
rect 42241 -14332 42305 -14328
rect 42241 -14388 42245 -14332
rect 42245 -14388 42301 -14332
rect 42301 -14388 42305 -14332
rect 42241 -14392 42305 -14388
rect 42241 -14652 42305 -14648
rect 42241 -14708 42245 -14652
rect 42245 -14708 42301 -14652
rect 42301 -14708 42305 -14652
rect 42241 -14712 42305 -14708
rect 42241 -14972 42305 -14968
rect 42241 -15028 42245 -14972
rect 42245 -15028 42301 -14972
rect 42301 -15028 42305 -14972
rect 42241 -15032 42305 -15028
rect 42241 -15292 42305 -15288
rect 42241 -15348 42245 -15292
rect 42245 -15348 42301 -15292
rect 42301 -15348 42305 -15292
rect 42241 -15352 42305 -15348
rect 42241 -15612 42305 -15608
rect 42241 -15668 42245 -15612
rect 42245 -15668 42301 -15612
rect 42301 -15668 42305 -15612
rect 42241 -15672 42305 -15668
rect 42241 -15932 42305 -15928
rect 42241 -15988 42245 -15932
rect 42245 -15988 42301 -15932
rect 42301 -15988 42305 -15932
rect 42241 -15992 42305 -15988
rect 42241 -16252 42305 -16248
rect 42241 -16308 42245 -16252
rect 42245 -16308 42301 -16252
rect 42301 -16308 42305 -16252
rect 42241 -16312 42305 -16308
rect 42241 -16572 42305 -16568
rect 42241 -16628 42245 -16572
rect 42245 -16628 42301 -16572
rect 42301 -16628 42305 -16572
rect 42241 -16632 42305 -16628
rect 42241 -16892 42305 -16888
rect 42241 -16948 42245 -16892
rect 42245 -16948 42301 -16892
rect 42301 -16948 42305 -16892
rect 42241 -16952 42305 -16948
rect 42241 -17212 42305 -17208
rect 42241 -17268 42245 -17212
rect 42245 -17268 42301 -17212
rect 42301 -17268 42305 -17212
rect 42241 -17272 42305 -17268
rect 42241 -17532 42305 -17528
rect 42241 -17588 42245 -17532
rect 42245 -17588 42301 -17532
rect 42301 -17588 42305 -17532
rect 42241 -17592 42305 -17588
rect 42241 -17852 42305 -17848
rect 42241 -17908 42245 -17852
rect 42245 -17908 42301 -17852
rect 42301 -17908 42305 -17852
rect 42241 -17912 42305 -17908
rect 42241 -18172 42305 -18168
rect 42241 -18228 42245 -18172
rect 42245 -18228 42301 -18172
rect 42301 -18228 42305 -18172
rect 42241 -18232 42305 -18228
rect 49695 -11772 49759 -11768
rect 49695 -11828 49699 -11772
rect 49699 -11828 49755 -11772
rect 49755 -11828 49759 -11772
rect 49695 -11832 49759 -11828
rect 49695 -12092 49759 -12088
rect 49695 -12148 49699 -12092
rect 49699 -12148 49755 -12092
rect 49755 -12148 49759 -12092
rect 49695 -12152 49759 -12148
rect 49695 -12412 49759 -12408
rect 49695 -12468 49699 -12412
rect 49699 -12468 49755 -12412
rect 49755 -12468 49759 -12412
rect 49695 -12472 49759 -12468
rect 49695 -12732 49759 -12728
rect 49695 -12788 49699 -12732
rect 49699 -12788 49755 -12732
rect 49755 -12788 49759 -12732
rect 49695 -12792 49759 -12788
rect 49695 -13052 49759 -13048
rect 49695 -13108 49699 -13052
rect 49699 -13108 49755 -13052
rect 49755 -13108 49759 -13052
rect 49695 -13112 49759 -13108
rect 49695 -13372 49759 -13368
rect 49695 -13428 49699 -13372
rect 49699 -13428 49755 -13372
rect 49755 -13428 49759 -13372
rect 49695 -13432 49759 -13428
rect 49695 -13692 49759 -13688
rect 49695 -13748 49699 -13692
rect 49699 -13748 49755 -13692
rect 49755 -13748 49759 -13692
rect 49695 -13752 49759 -13748
rect 49695 -14012 49759 -14008
rect 49695 -14068 49699 -14012
rect 49699 -14068 49755 -14012
rect 49755 -14068 49759 -14012
rect 49695 -14072 49759 -14068
rect 49695 -14332 49759 -14328
rect 49695 -14388 49699 -14332
rect 49699 -14388 49755 -14332
rect 49755 -14388 49759 -14332
rect 49695 -14392 49759 -14388
rect 49695 -14652 49759 -14648
rect 49695 -14708 49699 -14652
rect 49699 -14708 49755 -14652
rect 49755 -14708 49759 -14652
rect 49695 -14712 49759 -14708
rect 49695 -14972 49759 -14968
rect 49695 -15028 49699 -14972
rect 49699 -15028 49755 -14972
rect 49755 -15028 49759 -14972
rect 49695 -15032 49759 -15028
rect 49695 -15292 49759 -15288
rect 49695 -15348 49699 -15292
rect 49699 -15348 49755 -15292
rect 49755 -15348 49759 -15292
rect 49695 -15352 49759 -15348
rect 49695 -15612 49759 -15608
rect 49695 -15668 49699 -15612
rect 49699 -15668 49755 -15612
rect 49755 -15668 49759 -15612
rect 49695 -15672 49759 -15668
rect 49695 -15932 49759 -15928
rect 49695 -15988 49699 -15932
rect 49699 -15988 49755 -15932
rect 49755 -15988 49759 -15932
rect 49695 -15992 49759 -15988
rect 49695 -16252 49759 -16248
rect 49695 -16308 49699 -16252
rect 49699 -16308 49755 -16252
rect 49755 -16308 49759 -16252
rect 49695 -16312 49759 -16308
rect 49695 -16572 49759 -16568
rect 49695 -16628 49699 -16572
rect 49699 -16628 49755 -16572
rect 49755 -16628 49759 -16572
rect 49695 -16632 49759 -16628
rect 49695 -16892 49759 -16888
rect 49695 -16948 49699 -16892
rect 49699 -16948 49755 -16892
rect 49755 -16948 49759 -16892
rect 49695 -16952 49759 -16948
rect 49695 -17212 49759 -17208
rect 49695 -17268 49699 -17212
rect 49699 -17268 49755 -17212
rect 49755 -17268 49759 -17212
rect 49695 -17272 49759 -17268
rect 49695 -17532 49759 -17528
rect 49695 -17588 49699 -17532
rect 49699 -17588 49755 -17532
rect 49755 -17588 49759 -17532
rect 49695 -17592 49759 -17588
rect 49695 -17852 49759 -17848
rect 49695 -17908 49699 -17852
rect 49699 -17908 49755 -17852
rect 49755 -17908 49759 -17852
rect 49695 -17912 49759 -17908
rect 49695 -18172 49759 -18168
rect 49695 -18228 49699 -18172
rect 49699 -18228 49755 -18172
rect 49755 -18228 49759 -18172
rect 49695 -18232 49759 -18228
rect 42241 -18492 42305 -18488
rect 42241 -18548 42245 -18492
rect 42245 -18548 42301 -18492
rect 42301 -18548 42305 -18492
rect 42241 -18552 42305 -18548
rect 49695 -18492 49759 -18488
rect 49695 -18548 49699 -18492
rect 49699 -18548 49755 -18492
rect 49755 -18548 49759 -18492
rect 49695 -18552 49759 -18548
rect 42608 -18702 42672 -18698
rect 42608 -18758 42612 -18702
rect 42612 -18758 42668 -18702
rect 42668 -18758 42672 -18702
rect 42608 -18762 42672 -18758
rect 42928 -18702 42992 -18698
rect 42928 -18758 42932 -18702
rect 42932 -18758 42988 -18702
rect 42988 -18758 42992 -18702
rect 42928 -18762 42992 -18758
rect 43248 -18702 43312 -18698
rect 43248 -18758 43252 -18702
rect 43252 -18758 43308 -18702
rect 43308 -18758 43312 -18702
rect 43248 -18762 43312 -18758
rect 43568 -18702 43632 -18698
rect 43568 -18758 43572 -18702
rect 43572 -18758 43628 -18702
rect 43628 -18758 43632 -18702
rect 43568 -18762 43632 -18758
rect 43888 -18702 43952 -18698
rect 43888 -18758 43892 -18702
rect 43892 -18758 43948 -18702
rect 43948 -18758 43952 -18702
rect 43888 -18762 43952 -18758
rect 44208 -18702 44272 -18698
rect 44208 -18758 44212 -18702
rect 44212 -18758 44268 -18702
rect 44268 -18758 44272 -18702
rect 44208 -18762 44272 -18758
rect 44528 -18702 44592 -18698
rect 44528 -18758 44532 -18702
rect 44532 -18758 44588 -18702
rect 44588 -18758 44592 -18702
rect 44528 -18762 44592 -18758
rect 44848 -18702 44912 -18698
rect 44848 -18758 44852 -18702
rect 44852 -18758 44908 -18702
rect 44908 -18758 44912 -18702
rect 44848 -18762 44912 -18758
rect 45168 -18702 45232 -18698
rect 45168 -18758 45172 -18702
rect 45172 -18758 45228 -18702
rect 45228 -18758 45232 -18702
rect 45168 -18762 45232 -18758
rect 45488 -18702 45552 -18698
rect 45488 -18758 45492 -18702
rect 45492 -18758 45548 -18702
rect 45548 -18758 45552 -18702
rect 45488 -18762 45552 -18758
rect 45808 -18702 45872 -18698
rect 45808 -18758 45812 -18702
rect 45812 -18758 45868 -18702
rect 45868 -18758 45872 -18702
rect 45808 -18762 45872 -18758
rect 46128 -18702 46192 -18698
rect 46128 -18758 46132 -18702
rect 46132 -18758 46188 -18702
rect 46188 -18758 46192 -18702
rect 46128 -18762 46192 -18758
rect 46448 -18702 46512 -18698
rect 46448 -18758 46452 -18702
rect 46452 -18758 46508 -18702
rect 46508 -18758 46512 -18702
rect 46448 -18762 46512 -18758
rect 46768 -18702 46832 -18698
rect 46768 -18758 46772 -18702
rect 46772 -18758 46828 -18702
rect 46828 -18758 46832 -18702
rect 46768 -18762 46832 -18758
rect 47088 -18702 47152 -18698
rect 47088 -18758 47092 -18702
rect 47092 -18758 47148 -18702
rect 47148 -18758 47152 -18702
rect 47088 -18762 47152 -18758
rect 47408 -18702 47472 -18698
rect 47408 -18758 47412 -18702
rect 47412 -18758 47468 -18702
rect 47468 -18758 47472 -18702
rect 47408 -18762 47472 -18758
rect 47728 -18702 47792 -18698
rect 47728 -18758 47732 -18702
rect 47732 -18758 47788 -18702
rect 47788 -18758 47792 -18702
rect 47728 -18762 47792 -18758
rect 48048 -18702 48112 -18698
rect 48048 -18758 48052 -18702
rect 48052 -18758 48108 -18702
rect 48108 -18758 48112 -18702
rect 48048 -18762 48112 -18758
rect 48368 -18702 48432 -18698
rect 48368 -18758 48372 -18702
rect 48372 -18758 48428 -18702
rect 48428 -18758 48432 -18702
rect 48368 -18762 48432 -18758
rect 48688 -18702 48752 -18698
rect 48688 -18758 48692 -18702
rect 48692 -18758 48748 -18702
rect 48748 -18758 48752 -18702
rect 48688 -18762 48752 -18758
rect 49008 -18702 49072 -18698
rect 49008 -18758 49012 -18702
rect 49012 -18758 49068 -18702
rect 49068 -18758 49072 -18702
rect 49008 -18762 49072 -18758
rect 49328 -18702 49392 -18698
rect 49328 -18758 49332 -18702
rect 49332 -18758 49388 -18702
rect 49388 -18758 49392 -18702
rect 49328 -18762 49392 -18758
<< mimcap >>
rect 22840 1740 24400 1760
rect 22840 -540 22860 1740
rect 24380 -540 24400 1740
rect 22840 -560 24400 -540
rect 21300 -5560 21660 -5540
rect 21300 -8720 21320 -5560
rect 21640 -8720 21660 -5560
rect 21300 -8740 21660 -8720
<< mimcapcontact >>
rect 22860 -540 24380 1740
rect 21320 -8720 21640 -5560
<< metal4 >>
rect 3000 3720 51000 3740
rect 3000 3480 13960 3720
rect 14060 3480 51000 3720
rect 3000 3460 51000 3480
rect 20060 3360 20500 3400
rect 20060 3060 20080 3360
rect 20480 3060 20500 3360
rect 20060 3020 20500 3060
rect 3000 2940 51000 2960
rect 3000 2680 15180 2940
rect 15360 2680 51000 2940
rect 3000 2660 51000 2680
rect 3000 1880 51000 2160
rect 3000 1860 20840 1880
rect 24520 1860 51000 1880
rect 19980 1760 24440 1800
rect 11200 1600 12400 1700
rect 11200 1000 11400 1600
rect 12200 1000 12400 1600
rect 11200 -800 12400 1000
rect 15600 1600 16800 1700
rect 15600 1000 15800 1600
rect 16600 1000 16800 1600
rect 19980 1460 20020 1760
rect 20260 1740 24440 1760
rect 20260 1460 22860 1740
rect 19980 1420 22860 1460
rect 20000 1400 22860 1420
rect 14920 360 15220 400
rect 14920 -580 14940 360
rect 15200 -560 15220 360
rect 15140 -580 15220 -560
rect 14920 -600 15220 -580
rect 15600 -800 16800 1000
rect 22800 -540 22860 1400
rect 24380 -540 24440 1740
rect 22800 -600 24440 -540
rect 33000 1500 34700 1700
rect 33000 1000 33200 1500
rect 34500 1000 34700 1500
rect 33000 -700 34700 1000
rect 11200 -1100 20200 -800
rect 11200 -1200 14120 -1100
rect 12400 -1400 14120 -1200
rect 14260 -1400 20200 -1100
rect 20340 -1680 20660 -1640
rect 20340 -2200 20380 -1680
rect 20620 -2200 20660 -1680
rect 20340 -2240 20660 -2200
rect 21260 -5560 21860 -5500
rect 21260 -8720 21320 -5560
rect 21640 -8720 21860 -5560
rect 21260 -8840 21860 -8720
rect 19600 -9120 21860 -8840
rect 33000 -8400 33700 -700
rect 34000 -8400 34700 -700
rect 21340 -9260 21860 -9240
rect 21340 -9380 21360 -9260
rect 21840 -9380 21860 -9260
rect 21340 -9500 21380 -9380
rect 21820 -9500 21860 -9380
rect 21340 -9540 21860 -9500
rect 33000 -10100 43700 -8400
rect 42000 -11000 42700 -10100
rect 43000 -11000 43700 -10100
rect 6000 -11156 14000 -11000
rect 6000 -11362 6522 -11156
rect 6000 -11598 6152 -11362
rect 6388 -11392 6522 -11362
rect 6758 -11392 6842 -11156
rect 7078 -11392 7162 -11156
rect 7398 -11392 7482 -11156
rect 7718 -11392 7802 -11156
rect 8038 -11392 8122 -11156
rect 8358 -11392 8442 -11156
rect 8678 -11392 8762 -11156
rect 8998 -11392 9082 -11156
rect 9318 -11392 9402 -11156
rect 9638 -11392 9722 -11156
rect 9958 -11392 10042 -11156
rect 10278 -11392 10362 -11156
rect 10598 -11392 10682 -11156
rect 10918 -11392 11002 -11156
rect 11238 -11392 11322 -11156
rect 11558 -11392 11642 -11156
rect 11878 -11392 11962 -11156
rect 12198 -11392 12282 -11156
rect 12518 -11392 12602 -11156
rect 12838 -11392 12922 -11156
rect 13158 -11392 13242 -11156
rect 13478 -11362 14000 -11156
rect 13478 -11392 13618 -11362
rect 6388 -11540 13618 -11392
rect 6388 -11598 6540 -11540
rect 6000 -11682 6540 -11598
rect 6000 -11918 6152 -11682
rect 6388 -11918 6540 -11682
rect 6000 -12002 6540 -11918
rect 6000 -12238 6152 -12002
rect 6388 -12238 6540 -12002
rect 6000 -12322 6540 -12238
rect 6000 -12558 6152 -12322
rect 6388 -12558 6540 -12322
rect 6000 -12642 6540 -12558
rect 6000 -12878 6152 -12642
rect 6388 -12878 6540 -12642
rect 6000 -12962 6540 -12878
rect 6000 -13198 6152 -12962
rect 6388 -13198 6540 -12962
rect 6000 -13282 6540 -13198
rect 6000 -13518 6152 -13282
rect 6388 -13518 6540 -13282
rect 6000 -13602 6540 -13518
rect 6000 -13838 6152 -13602
rect 6388 -13838 6540 -13602
rect 6000 -13922 6540 -13838
rect 6000 -14158 6152 -13922
rect 6388 -14158 6540 -13922
rect 6000 -14242 6540 -14158
rect 6000 -14478 6152 -14242
rect 6388 -14478 6540 -14242
rect 6000 -14562 6540 -14478
rect 6000 -14798 6152 -14562
rect 6388 -14798 6540 -14562
rect 6000 -14882 6540 -14798
rect 6000 -15118 6152 -14882
rect 6388 -15118 6540 -14882
rect 6000 -15202 6540 -15118
rect 6000 -15438 6152 -15202
rect 6388 -15438 6540 -15202
rect 6000 -15522 6540 -15438
rect 6000 -15758 6152 -15522
rect 6388 -15758 6540 -15522
rect 6000 -15842 6540 -15758
rect 6000 -16078 6152 -15842
rect 6388 -16078 6540 -15842
rect 6000 -16162 6540 -16078
rect 6000 -16398 6152 -16162
rect 6388 -16398 6540 -16162
rect 6000 -16482 6540 -16398
rect 6000 -16718 6152 -16482
rect 6388 -16718 6540 -16482
rect 6000 -16802 6540 -16718
rect 6000 -17038 6152 -16802
rect 6388 -17038 6540 -16802
rect 6000 -17122 6540 -17038
rect 6000 -17358 6152 -17122
rect 6388 -17358 6540 -17122
rect 6000 -17442 6540 -17358
rect 6000 -17678 6152 -17442
rect 6388 -17678 6540 -17442
rect 6000 -17762 6540 -17678
rect 6000 -17998 6152 -17762
rect 6388 -17998 6540 -17762
rect 6000 -18082 6540 -17998
rect 6000 -18318 6152 -18082
rect 6388 -18318 6540 -18082
rect 6000 -18402 6540 -18318
rect 6000 -18638 6152 -18402
rect 6388 -18460 6540 -18402
rect 13460 -11598 13618 -11540
rect 13854 -11598 14000 -11362
rect 13460 -11682 14000 -11598
rect 13460 -11918 13618 -11682
rect 13854 -11918 14000 -11682
rect 13460 -12002 14000 -11918
rect 13460 -12238 13618 -12002
rect 13854 -12238 14000 -12002
rect 13460 -12322 14000 -12238
rect 13460 -12558 13618 -12322
rect 13854 -12558 14000 -12322
rect 13460 -12642 14000 -12558
rect 13460 -12878 13618 -12642
rect 13854 -12878 14000 -12642
rect 13460 -12962 14000 -12878
rect 13460 -13198 13618 -12962
rect 13854 -13198 14000 -12962
rect 13460 -13282 14000 -13198
rect 13460 -13518 13618 -13282
rect 13854 -13518 14000 -13282
rect 13460 -13602 14000 -13518
rect 13460 -13838 13618 -13602
rect 13854 -13838 14000 -13602
rect 13460 -13922 14000 -13838
rect 13460 -14158 13618 -13922
rect 13854 -14158 14000 -13922
rect 13460 -14242 14000 -14158
rect 13460 -14478 13618 -14242
rect 13854 -14478 14000 -14242
rect 13460 -14562 14000 -14478
rect 13460 -14798 13618 -14562
rect 13854 -14798 14000 -14562
rect 13460 -14882 14000 -14798
rect 13460 -15118 13618 -14882
rect 13854 -15118 14000 -14882
rect 13460 -15202 14000 -15118
rect 13460 -15438 13618 -15202
rect 13854 -15438 14000 -15202
rect 13460 -15522 14000 -15438
rect 13460 -15758 13618 -15522
rect 13854 -15758 14000 -15522
rect 13460 -15842 14000 -15758
rect 13460 -16078 13618 -15842
rect 13854 -16078 14000 -15842
rect 13460 -16162 14000 -16078
rect 13460 -16398 13618 -16162
rect 13854 -16398 14000 -16162
rect 13460 -16482 14000 -16398
rect 13460 -16718 13618 -16482
rect 13854 -16718 14000 -16482
rect 13460 -16802 14000 -16718
rect 13460 -17038 13618 -16802
rect 13854 -17038 14000 -16802
rect 13460 -17122 14000 -17038
rect 13460 -17358 13618 -17122
rect 13854 -17358 14000 -17122
rect 13460 -17442 14000 -17358
rect 13460 -17678 13618 -17442
rect 13854 -17678 14000 -17442
rect 13460 -17762 14000 -17678
rect 13460 -17998 13618 -17762
rect 13854 -17998 14000 -17762
rect 13460 -18082 14000 -17998
rect 13460 -18318 13618 -18082
rect 13854 -18318 14000 -18082
rect 13460 -18402 14000 -18318
rect 13460 -18460 13618 -18402
rect 6388 -18612 13618 -18460
rect 6388 -18638 6522 -18612
rect 6000 -18848 6522 -18638
rect 6758 -18848 6842 -18612
rect 7078 -18848 7162 -18612
rect 7398 -18848 7482 -18612
rect 7718 -18848 7802 -18612
rect 8038 -18848 8122 -18612
rect 8358 -18848 8442 -18612
rect 8678 -18848 8762 -18612
rect 8998 -18848 9082 -18612
rect 9318 -18848 9402 -18612
rect 9638 -18848 9722 -18612
rect 9958 -18848 10042 -18612
rect 10278 -18848 10362 -18612
rect 10598 -18848 10682 -18612
rect 10918 -18848 11002 -18612
rect 11238 -18848 11322 -18612
rect 11558 -18848 11642 -18612
rect 11878 -18848 11962 -18612
rect 12198 -18848 12282 -18612
rect 12518 -18848 12602 -18612
rect 12838 -18848 12922 -18612
rect 13158 -18848 13242 -18612
rect 13478 -18638 13618 -18612
rect 13854 -18638 14000 -18402
rect 13478 -18848 14000 -18638
rect 6000 -19000 14000 -18848
rect 18000 -11156 26000 -11000
rect 18000 -11362 18522 -11156
rect 18000 -11598 18152 -11362
rect 18388 -11392 18522 -11362
rect 18758 -11392 18842 -11156
rect 19078 -11392 19162 -11156
rect 19398 -11392 19482 -11156
rect 19718 -11392 19802 -11156
rect 20038 -11392 20122 -11156
rect 20358 -11392 20442 -11156
rect 20678 -11392 20762 -11156
rect 20998 -11392 21082 -11156
rect 21318 -11392 21402 -11156
rect 21638 -11392 21722 -11156
rect 21958 -11392 22042 -11156
rect 22278 -11392 22362 -11156
rect 22598 -11392 22682 -11156
rect 22918 -11392 23002 -11156
rect 23238 -11392 23322 -11156
rect 23558 -11392 23642 -11156
rect 23878 -11392 23962 -11156
rect 24198 -11392 24282 -11156
rect 24518 -11392 24602 -11156
rect 24838 -11392 24922 -11156
rect 25158 -11392 25242 -11156
rect 25478 -11362 26000 -11156
rect 25478 -11392 25618 -11362
rect 18388 -11540 25618 -11392
rect 18388 -11598 18540 -11540
rect 18000 -11682 18540 -11598
rect 18000 -11918 18152 -11682
rect 18388 -11918 18540 -11682
rect 18000 -12002 18540 -11918
rect 18000 -12238 18152 -12002
rect 18388 -12238 18540 -12002
rect 18000 -12322 18540 -12238
rect 18000 -12558 18152 -12322
rect 18388 -12558 18540 -12322
rect 18000 -12642 18540 -12558
rect 18000 -12878 18152 -12642
rect 18388 -12878 18540 -12642
rect 18000 -12962 18540 -12878
rect 18000 -13198 18152 -12962
rect 18388 -13198 18540 -12962
rect 18000 -13282 18540 -13198
rect 18000 -13518 18152 -13282
rect 18388 -13518 18540 -13282
rect 18000 -13602 18540 -13518
rect 18000 -13838 18152 -13602
rect 18388 -13838 18540 -13602
rect 18000 -13922 18540 -13838
rect 18000 -14158 18152 -13922
rect 18388 -14158 18540 -13922
rect 18000 -14242 18540 -14158
rect 18000 -14478 18152 -14242
rect 18388 -14478 18540 -14242
rect 18000 -14562 18540 -14478
rect 18000 -14798 18152 -14562
rect 18388 -14798 18540 -14562
rect 18000 -14882 18540 -14798
rect 18000 -15118 18152 -14882
rect 18388 -15118 18540 -14882
rect 18000 -15202 18540 -15118
rect 18000 -15438 18152 -15202
rect 18388 -15438 18540 -15202
rect 18000 -15522 18540 -15438
rect 18000 -15758 18152 -15522
rect 18388 -15758 18540 -15522
rect 18000 -15842 18540 -15758
rect 18000 -16078 18152 -15842
rect 18388 -16078 18540 -15842
rect 18000 -16162 18540 -16078
rect 18000 -16398 18152 -16162
rect 18388 -16398 18540 -16162
rect 18000 -16482 18540 -16398
rect 18000 -16718 18152 -16482
rect 18388 -16718 18540 -16482
rect 18000 -16802 18540 -16718
rect 18000 -17038 18152 -16802
rect 18388 -17038 18540 -16802
rect 18000 -17122 18540 -17038
rect 18000 -17358 18152 -17122
rect 18388 -17358 18540 -17122
rect 18000 -17442 18540 -17358
rect 18000 -17678 18152 -17442
rect 18388 -17678 18540 -17442
rect 18000 -17762 18540 -17678
rect 18000 -17998 18152 -17762
rect 18388 -17998 18540 -17762
rect 18000 -18082 18540 -17998
rect 18000 -18318 18152 -18082
rect 18388 -18318 18540 -18082
rect 18000 -18402 18540 -18318
rect 18000 -18638 18152 -18402
rect 18388 -18460 18540 -18402
rect 25460 -11598 25618 -11540
rect 25854 -11598 26000 -11362
rect 25460 -11682 26000 -11598
rect 25460 -11918 25618 -11682
rect 25854 -11918 26000 -11682
rect 25460 -12002 26000 -11918
rect 25460 -12238 25618 -12002
rect 25854 -12238 26000 -12002
rect 25460 -12322 26000 -12238
rect 25460 -12558 25618 -12322
rect 25854 -12558 26000 -12322
rect 25460 -12642 26000 -12558
rect 25460 -12878 25618 -12642
rect 25854 -12878 26000 -12642
rect 25460 -12962 26000 -12878
rect 25460 -13198 25618 -12962
rect 25854 -13198 26000 -12962
rect 25460 -13282 26000 -13198
rect 25460 -13518 25618 -13282
rect 25854 -13518 26000 -13282
rect 25460 -13602 26000 -13518
rect 25460 -13838 25618 -13602
rect 25854 -13838 26000 -13602
rect 25460 -13922 26000 -13838
rect 25460 -14158 25618 -13922
rect 25854 -14158 26000 -13922
rect 25460 -14242 26000 -14158
rect 25460 -14478 25618 -14242
rect 25854 -14478 26000 -14242
rect 25460 -14562 26000 -14478
rect 25460 -14798 25618 -14562
rect 25854 -14798 26000 -14562
rect 25460 -14882 26000 -14798
rect 25460 -15118 25618 -14882
rect 25854 -15118 26000 -14882
rect 25460 -15202 26000 -15118
rect 25460 -15438 25618 -15202
rect 25854 -15438 26000 -15202
rect 25460 -15522 26000 -15438
rect 25460 -15758 25618 -15522
rect 25854 -15758 26000 -15522
rect 25460 -15842 26000 -15758
rect 25460 -16078 25618 -15842
rect 25854 -16078 26000 -15842
rect 25460 -16162 26000 -16078
rect 25460 -16398 25618 -16162
rect 25854 -16398 26000 -16162
rect 25460 -16482 26000 -16398
rect 25460 -16718 25618 -16482
rect 25854 -16718 26000 -16482
rect 25460 -16802 26000 -16718
rect 25460 -17038 25618 -16802
rect 25854 -17038 26000 -16802
rect 25460 -17122 26000 -17038
rect 25460 -17358 25618 -17122
rect 25854 -17358 26000 -17122
rect 25460 -17442 26000 -17358
rect 25460 -17678 25618 -17442
rect 25854 -17678 26000 -17442
rect 25460 -17762 26000 -17678
rect 25460 -17998 25618 -17762
rect 25854 -17998 26000 -17762
rect 25460 -18082 26000 -17998
rect 25460 -18318 25618 -18082
rect 25854 -18318 26000 -18082
rect 25460 -18402 26000 -18318
rect 25460 -18460 25618 -18402
rect 18388 -18612 25618 -18460
rect 18388 -18638 18522 -18612
rect 18000 -18848 18522 -18638
rect 18758 -18848 18842 -18612
rect 19078 -18848 19162 -18612
rect 19398 -18848 19482 -18612
rect 19718 -18848 19802 -18612
rect 20038 -18848 20122 -18612
rect 20358 -18848 20442 -18612
rect 20678 -18848 20762 -18612
rect 20998 -18848 21082 -18612
rect 21318 -18848 21402 -18612
rect 21638 -18848 21722 -18612
rect 21958 -18848 22042 -18612
rect 22278 -18848 22362 -18612
rect 22598 -18848 22682 -18612
rect 22918 -18848 23002 -18612
rect 23238 -18848 23322 -18612
rect 23558 -18848 23642 -18612
rect 23878 -18848 23962 -18612
rect 24198 -18848 24282 -18612
rect 24518 -18848 24602 -18612
rect 24838 -18848 24922 -18612
rect 25158 -18848 25242 -18612
rect 25478 -18638 25618 -18612
rect 25854 -18638 26000 -18402
rect 25478 -18848 26000 -18638
rect 18000 -19000 26000 -18848
rect 30000 -11156 38000 -11000
rect 30000 -11362 30522 -11156
rect 30000 -11598 30152 -11362
rect 30388 -11392 30522 -11362
rect 30758 -11392 30842 -11156
rect 31078 -11392 31162 -11156
rect 31398 -11392 31482 -11156
rect 31718 -11392 31802 -11156
rect 32038 -11392 32122 -11156
rect 32358 -11392 32442 -11156
rect 32678 -11392 32762 -11156
rect 32998 -11392 33082 -11156
rect 33318 -11392 33402 -11156
rect 33638 -11392 33722 -11156
rect 33958 -11392 34042 -11156
rect 34278 -11392 34362 -11156
rect 34598 -11392 34682 -11156
rect 34918 -11392 35002 -11156
rect 35238 -11392 35322 -11156
rect 35558 -11392 35642 -11156
rect 35878 -11392 35962 -11156
rect 36198 -11392 36282 -11156
rect 36518 -11392 36602 -11156
rect 36838 -11392 36922 -11156
rect 37158 -11392 37242 -11156
rect 37478 -11362 38000 -11156
rect 37478 -11392 37618 -11362
rect 30388 -11540 37618 -11392
rect 30388 -11598 30540 -11540
rect 30000 -11682 30540 -11598
rect 30000 -11918 30152 -11682
rect 30388 -11918 30540 -11682
rect 30000 -12002 30540 -11918
rect 30000 -12238 30152 -12002
rect 30388 -12238 30540 -12002
rect 30000 -12322 30540 -12238
rect 30000 -12558 30152 -12322
rect 30388 -12558 30540 -12322
rect 30000 -12642 30540 -12558
rect 30000 -12878 30152 -12642
rect 30388 -12878 30540 -12642
rect 30000 -12962 30540 -12878
rect 30000 -13198 30152 -12962
rect 30388 -13198 30540 -12962
rect 30000 -13282 30540 -13198
rect 30000 -13518 30152 -13282
rect 30388 -13518 30540 -13282
rect 30000 -13602 30540 -13518
rect 30000 -13838 30152 -13602
rect 30388 -13838 30540 -13602
rect 30000 -13922 30540 -13838
rect 30000 -14158 30152 -13922
rect 30388 -14158 30540 -13922
rect 30000 -14242 30540 -14158
rect 30000 -14478 30152 -14242
rect 30388 -14478 30540 -14242
rect 30000 -14562 30540 -14478
rect 30000 -14798 30152 -14562
rect 30388 -14798 30540 -14562
rect 30000 -14882 30540 -14798
rect 30000 -15118 30152 -14882
rect 30388 -15118 30540 -14882
rect 30000 -15202 30540 -15118
rect 30000 -15438 30152 -15202
rect 30388 -15438 30540 -15202
rect 30000 -15522 30540 -15438
rect 30000 -15758 30152 -15522
rect 30388 -15758 30540 -15522
rect 30000 -15842 30540 -15758
rect 30000 -16078 30152 -15842
rect 30388 -16078 30540 -15842
rect 30000 -16162 30540 -16078
rect 30000 -16398 30152 -16162
rect 30388 -16398 30540 -16162
rect 30000 -16482 30540 -16398
rect 30000 -16718 30152 -16482
rect 30388 -16718 30540 -16482
rect 30000 -16802 30540 -16718
rect 30000 -17038 30152 -16802
rect 30388 -17038 30540 -16802
rect 30000 -17122 30540 -17038
rect 30000 -17358 30152 -17122
rect 30388 -17358 30540 -17122
rect 30000 -17442 30540 -17358
rect 30000 -17678 30152 -17442
rect 30388 -17678 30540 -17442
rect 30000 -17762 30540 -17678
rect 30000 -17998 30152 -17762
rect 30388 -17998 30540 -17762
rect 30000 -18082 30540 -17998
rect 30000 -18318 30152 -18082
rect 30388 -18318 30540 -18082
rect 30000 -18402 30540 -18318
rect 30000 -18638 30152 -18402
rect 30388 -18460 30540 -18402
rect 37460 -11598 37618 -11540
rect 37854 -11598 38000 -11362
rect 37460 -11682 38000 -11598
rect 37460 -11918 37618 -11682
rect 37854 -11918 38000 -11682
rect 37460 -12002 38000 -11918
rect 37460 -12238 37618 -12002
rect 37854 -12238 38000 -12002
rect 37460 -12322 38000 -12238
rect 37460 -12558 37618 -12322
rect 37854 -12558 38000 -12322
rect 37460 -12642 38000 -12558
rect 37460 -12878 37618 -12642
rect 37854 -12878 38000 -12642
rect 37460 -12962 38000 -12878
rect 37460 -13198 37618 -12962
rect 37854 -13198 38000 -12962
rect 37460 -13282 38000 -13198
rect 37460 -13518 37618 -13282
rect 37854 -13518 38000 -13282
rect 37460 -13602 38000 -13518
rect 37460 -13838 37618 -13602
rect 37854 -13838 38000 -13602
rect 37460 -13922 38000 -13838
rect 37460 -14158 37618 -13922
rect 37854 -14158 38000 -13922
rect 37460 -14242 38000 -14158
rect 37460 -14478 37618 -14242
rect 37854 -14478 38000 -14242
rect 37460 -14562 38000 -14478
rect 37460 -14798 37618 -14562
rect 37854 -14798 38000 -14562
rect 37460 -14882 38000 -14798
rect 37460 -15118 37618 -14882
rect 37854 -15118 38000 -14882
rect 37460 -15202 38000 -15118
rect 37460 -15438 37618 -15202
rect 37854 -15438 38000 -15202
rect 37460 -15522 38000 -15438
rect 37460 -15758 37618 -15522
rect 37854 -15758 38000 -15522
rect 37460 -15842 38000 -15758
rect 37460 -16078 37618 -15842
rect 37854 -16078 38000 -15842
rect 37460 -16162 38000 -16078
rect 37460 -16398 37618 -16162
rect 37854 -16398 38000 -16162
rect 37460 -16482 38000 -16398
rect 37460 -16718 37618 -16482
rect 37854 -16718 38000 -16482
rect 37460 -16802 38000 -16718
rect 37460 -17038 37618 -16802
rect 37854 -17038 38000 -16802
rect 37460 -17122 38000 -17038
rect 37460 -17358 37618 -17122
rect 37854 -17358 38000 -17122
rect 37460 -17442 38000 -17358
rect 37460 -17678 37618 -17442
rect 37854 -17678 38000 -17442
rect 37460 -17762 38000 -17678
rect 37460 -17998 37618 -17762
rect 37854 -17998 38000 -17762
rect 37460 -18082 38000 -17998
rect 37460 -18318 37618 -18082
rect 37854 -18318 38000 -18082
rect 37460 -18402 38000 -18318
rect 37460 -18460 37618 -18402
rect 30388 -18612 37618 -18460
rect 30388 -18638 30522 -18612
rect 30000 -18848 30522 -18638
rect 30758 -18848 30842 -18612
rect 31078 -18848 31162 -18612
rect 31398 -18848 31482 -18612
rect 31718 -18848 31802 -18612
rect 32038 -18848 32122 -18612
rect 32358 -18848 32442 -18612
rect 32678 -18848 32762 -18612
rect 32998 -18848 33082 -18612
rect 33318 -18848 33402 -18612
rect 33638 -18848 33722 -18612
rect 33958 -18848 34042 -18612
rect 34278 -18848 34362 -18612
rect 34598 -18848 34682 -18612
rect 34918 -18848 35002 -18612
rect 35238 -18848 35322 -18612
rect 35558 -18848 35642 -18612
rect 35878 -18848 35962 -18612
rect 36198 -18848 36282 -18612
rect 36518 -18848 36602 -18612
rect 36838 -18848 36922 -18612
rect 37158 -18848 37242 -18612
rect 37478 -18638 37618 -18612
rect 37854 -18638 38000 -18402
rect 37478 -18848 38000 -18638
rect 30000 -19000 38000 -18848
rect 42000 -11156 50000 -11000
rect 42000 -11362 42522 -11156
rect 42000 -11598 42155 -11362
rect 42391 -11392 42522 -11362
rect 42758 -11392 42842 -11156
rect 43078 -11392 43162 -11156
rect 43398 -11392 43482 -11156
rect 43718 -11392 43802 -11156
rect 44038 -11392 44122 -11156
rect 44358 -11392 44442 -11156
rect 44678 -11392 44762 -11156
rect 44998 -11392 45082 -11156
rect 45318 -11392 45402 -11156
rect 45638 -11392 45722 -11156
rect 45958 -11392 46042 -11156
rect 46278 -11392 46362 -11156
rect 46598 -11392 46682 -11156
rect 46918 -11392 47002 -11156
rect 47238 -11392 47322 -11156
rect 47558 -11392 47642 -11156
rect 47878 -11392 47962 -11156
rect 48198 -11392 48282 -11156
rect 48518 -11392 48602 -11156
rect 48838 -11392 48922 -11156
rect 49158 -11392 49242 -11156
rect 49478 -11362 50000 -11156
rect 49478 -11392 49609 -11362
rect 42391 -11540 49609 -11392
rect 42391 -11598 42540 -11540
rect 42000 -11682 42540 -11598
rect 42000 -11918 42155 -11682
rect 42391 -11918 42540 -11682
rect 42000 -12002 42540 -11918
rect 42000 -12238 42155 -12002
rect 42391 -12238 42540 -12002
rect 42000 -12322 42540 -12238
rect 42000 -12558 42155 -12322
rect 42391 -12558 42540 -12322
rect 42000 -12642 42540 -12558
rect 42000 -12878 42155 -12642
rect 42391 -12878 42540 -12642
rect 42000 -12962 42540 -12878
rect 42000 -13198 42155 -12962
rect 42391 -13198 42540 -12962
rect 42000 -13282 42540 -13198
rect 42000 -13518 42155 -13282
rect 42391 -13518 42540 -13282
rect 42000 -13602 42540 -13518
rect 42000 -13838 42155 -13602
rect 42391 -13838 42540 -13602
rect 42000 -13922 42540 -13838
rect 42000 -14158 42155 -13922
rect 42391 -14158 42540 -13922
rect 42000 -14242 42540 -14158
rect 42000 -14478 42155 -14242
rect 42391 -14478 42540 -14242
rect 42000 -14562 42540 -14478
rect 42000 -14798 42155 -14562
rect 42391 -14798 42540 -14562
rect 42000 -14882 42540 -14798
rect 42000 -15118 42155 -14882
rect 42391 -15118 42540 -14882
rect 42000 -15202 42540 -15118
rect 42000 -15438 42155 -15202
rect 42391 -15438 42540 -15202
rect 42000 -15522 42540 -15438
rect 42000 -15758 42155 -15522
rect 42391 -15758 42540 -15522
rect 42000 -15842 42540 -15758
rect 42000 -16078 42155 -15842
rect 42391 -16078 42540 -15842
rect 42000 -16162 42540 -16078
rect 42000 -16398 42155 -16162
rect 42391 -16398 42540 -16162
rect 42000 -16482 42540 -16398
rect 42000 -16718 42155 -16482
rect 42391 -16718 42540 -16482
rect 42000 -16802 42540 -16718
rect 42000 -17038 42155 -16802
rect 42391 -17038 42540 -16802
rect 42000 -17122 42540 -17038
rect 42000 -17358 42155 -17122
rect 42391 -17358 42540 -17122
rect 42000 -17442 42540 -17358
rect 42000 -17678 42155 -17442
rect 42391 -17678 42540 -17442
rect 42000 -17762 42540 -17678
rect 42000 -17998 42155 -17762
rect 42391 -17998 42540 -17762
rect 42000 -18082 42540 -17998
rect 42000 -18318 42155 -18082
rect 42391 -18318 42540 -18082
rect 42000 -18402 42540 -18318
rect 42000 -18638 42155 -18402
rect 42391 -18460 42540 -18402
rect 49460 -11598 49609 -11540
rect 49845 -11598 50000 -11362
rect 49460 -11682 50000 -11598
rect 49460 -11918 49609 -11682
rect 49845 -11918 50000 -11682
rect 49460 -12002 50000 -11918
rect 49460 -12238 49609 -12002
rect 49845 -12238 50000 -12002
rect 49460 -12322 50000 -12238
rect 49460 -12558 49609 -12322
rect 49845 -12558 50000 -12322
rect 49460 -12642 50000 -12558
rect 49460 -12878 49609 -12642
rect 49845 -12878 50000 -12642
rect 49460 -12962 50000 -12878
rect 49460 -13198 49609 -12962
rect 49845 -13198 50000 -12962
rect 49460 -13282 50000 -13198
rect 49460 -13518 49609 -13282
rect 49845 -13518 50000 -13282
rect 49460 -13602 50000 -13518
rect 49460 -13838 49609 -13602
rect 49845 -13838 50000 -13602
rect 49460 -13922 50000 -13838
rect 49460 -14158 49609 -13922
rect 49845 -14158 50000 -13922
rect 49460 -14242 50000 -14158
rect 49460 -14478 49609 -14242
rect 49845 -14478 50000 -14242
rect 49460 -14562 50000 -14478
rect 49460 -14798 49609 -14562
rect 49845 -14798 50000 -14562
rect 49460 -14882 50000 -14798
rect 49460 -15118 49609 -14882
rect 49845 -15118 50000 -14882
rect 49460 -15202 50000 -15118
rect 49460 -15438 49609 -15202
rect 49845 -15438 50000 -15202
rect 49460 -15522 50000 -15438
rect 49460 -15758 49609 -15522
rect 49845 -15758 50000 -15522
rect 49460 -15842 50000 -15758
rect 49460 -16078 49609 -15842
rect 49845 -16078 50000 -15842
rect 49460 -16162 50000 -16078
rect 49460 -16398 49609 -16162
rect 49845 -16398 50000 -16162
rect 49460 -16482 50000 -16398
rect 49460 -16718 49609 -16482
rect 49845 -16718 50000 -16482
rect 49460 -16802 50000 -16718
rect 49460 -17038 49609 -16802
rect 49845 -17038 50000 -16802
rect 49460 -17122 50000 -17038
rect 49460 -17358 49609 -17122
rect 49845 -17358 50000 -17122
rect 49460 -17442 50000 -17358
rect 49460 -17678 49609 -17442
rect 49845 -17678 50000 -17442
rect 49460 -17762 50000 -17678
rect 49460 -17998 49609 -17762
rect 49845 -17998 50000 -17762
rect 49460 -18082 50000 -17998
rect 49460 -18318 49609 -18082
rect 49845 -18318 50000 -18082
rect 49460 -18402 50000 -18318
rect 49460 -18460 49609 -18402
rect 42391 -18612 49609 -18460
rect 42391 -18638 42522 -18612
rect 42000 -18848 42522 -18638
rect 42758 -18848 42842 -18612
rect 43078 -18848 43162 -18612
rect 43398 -18848 43482 -18612
rect 43718 -18848 43802 -18612
rect 44038 -18848 44122 -18612
rect 44358 -18848 44442 -18612
rect 44678 -18848 44762 -18612
rect 44998 -18848 45082 -18612
rect 45318 -18848 45402 -18612
rect 45638 -18848 45722 -18612
rect 45958 -18848 46042 -18612
rect 46278 -18848 46362 -18612
rect 46598 -18848 46682 -18612
rect 46918 -18848 47002 -18612
rect 47238 -18848 47322 -18612
rect 47558 -18848 47642 -18612
rect 47878 -18848 47962 -18612
rect 48198 -18848 48282 -18612
rect 48518 -18848 48602 -18612
rect 48838 -18848 48922 -18612
rect 49158 -18848 49242 -18612
rect 49478 -18638 49609 -18612
rect 49845 -18638 50000 -18402
rect 49478 -18848 50000 -18638
rect 42000 -19000 50000 -18848
<< via4 >>
rect 20080 3280 20480 3360
rect 20080 3140 20480 3280
rect 20080 3060 20480 3140
rect 11400 1000 12200 1600
rect 15800 1000 16600 1600
rect 20020 1460 20260 1760
rect 14940 -200 15200 360
rect 14940 -560 15140 -200
rect 15140 -560 15200 -200
rect 33200 1000 34500 1500
rect 20380 -2200 20620 -1680
rect 21380 -9380 21820 -9260
rect 21380 -9500 21820 -9380
rect 6522 -11242 6758 -11156
rect 6522 -11306 6608 -11242
rect 6608 -11306 6672 -11242
rect 6672 -11306 6758 -11242
rect 6152 -11448 6388 -11362
rect 6522 -11392 6758 -11306
rect 6842 -11242 7078 -11156
rect 6842 -11306 6928 -11242
rect 6928 -11306 6992 -11242
rect 6992 -11306 7078 -11242
rect 6842 -11392 7078 -11306
rect 7162 -11242 7398 -11156
rect 7162 -11306 7248 -11242
rect 7248 -11306 7312 -11242
rect 7312 -11306 7398 -11242
rect 7162 -11392 7398 -11306
rect 7482 -11242 7718 -11156
rect 7482 -11306 7568 -11242
rect 7568 -11306 7632 -11242
rect 7632 -11306 7718 -11242
rect 7482 -11392 7718 -11306
rect 7802 -11242 8038 -11156
rect 7802 -11306 7888 -11242
rect 7888 -11306 7952 -11242
rect 7952 -11306 8038 -11242
rect 7802 -11392 8038 -11306
rect 8122 -11242 8358 -11156
rect 8122 -11306 8208 -11242
rect 8208 -11306 8272 -11242
rect 8272 -11306 8358 -11242
rect 8122 -11392 8358 -11306
rect 8442 -11242 8678 -11156
rect 8442 -11306 8528 -11242
rect 8528 -11306 8592 -11242
rect 8592 -11306 8678 -11242
rect 8442 -11392 8678 -11306
rect 8762 -11242 8998 -11156
rect 8762 -11306 8848 -11242
rect 8848 -11306 8912 -11242
rect 8912 -11306 8998 -11242
rect 8762 -11392 8998 -11306
rect 9082 -11242 9318 -11156
rect 9082 -11306 9168 -11242
rect 9168 -11306 9232 -11242
rect 9232 -11306 9318 -11242
rect 9082 -11392 9318 -11306
rect 9402 -11242 9638 -11156
rect 9402 -11306 9488 -11242
rect 9488 -11306 9552 -11242
rect 9552 -11306 9638 -11242
rect 9402 -11392 9638 -11306
rect 9722 -11242 9958 -11156
rect 9722 -11306 9808 -11242
rect 9808 -11306 9872 -11242
rect 9872 -11306 9958 -11242
rect 9722 -11392 9958 -11306
rect 10042 -11242 10278 -11156
rect 10042 -11306 10128 -11242
rect 10128 -11306 10192 -11242
rect 10192 -11306 10278 -11242
rect 10042 -11392 10278 -11306
rect 10362 -11242 10598 -11156
rect 10362 -11306 10448 -11242
rect 10448 -11306 10512 -11242
rect 10512 -11306 10598 -11242
rect 10362 -11392 10598 -11306
rect 10682 -11242 10918 -11156
rect 10682 -11306 10768 -11242
rect 10768 -11306 10832 -11242
rect 10832 -11306 10918 -11242
rect 10682 -11392 10918 -11306
rect 11002 -11242 11238 -11156
rect 11002 -11306 11088 -11242
rect 11088 -11306 11152 -11242
rect 11152 -11306 11238 -11242
rect 11002 -11392 11238 -11306
rect 11322 -11242 11558 -11156
rect 11322 -11306 11408 -11242
rect 11408 -11306 11472 -11242
rect 11472 -11306 11558 -11242
rect 11322 -11392 11558 -11306
rect 11642 -11242 11878 -11156
rect 11642 -11306 11728 -11242
rect 11728 -11306 11792 -11242
rect 11792 -11306 11878 -11242
rect 11642 -11392 11878 -11306
rect 11962 -11242 12198 -11156
rect 11962 -11306 12048 -11242
rect 12048 -11306 12112 -11242
rect 12112 -11306 12198 -11242
rect 11962 -11392 12198 -11306
rect 12282 -11242 12518 -11156
rect 12282 -11306 12368 -11242
rect 12368 -11306 12432 -11242
rect 12432 -11306 12518 -11242
rect 12282 -11392 12518 -11306
rect 12602 -11242 12838 -11156
rect 12602 -11306 12688 -11242
rect 12688 -11306 12752 -11242
rect 12752 -11306 12838 -11242
rect 12602 -11392 12838 -11306
rect 12922 -11242 13158 -11156
rect 12922 -11306 13008 -11242
rect 13008 -11306 13072 -11242
rect 13072 -11306 13158 -11242
rect 12922 -11392 13158 -11306
rect 13242 -11242 13478 -11156
rect 13242 -11306 13328 -11242
rect 13328 -11306 13392 -11242
rect 13392 -11306 13478 -11242
rect 13242 -11392 13478 -11306
rect 6152 -11512 6238 -11448
rect 6238 -11512 6302 -11448
rect 6302 -11512 6388 -11448
rect 6152 -11598 6388 -11512
rect 13618 -11448 13854 -11362
rect 13618 -11512 13704 -11448
rect 13704 -11512 13768 -11448
rect 13768 -11512 13854 -11448
rect 6152 -11768 6388 -11682
rect 6152 -11832 6238 -11768
rect 6238 -11832 6302 -11768
rect 6302 -11832 6388 -11768
rect 6152 -11918 6388 -11832
rect 6152 -12088 6388 -12002
rect 6152 -12152 6238 -12088
rect 6238 -12152 6302 -12088
rect 6302 -12152 6388 -12088
rect 6152 -12238 6388 -12152
rect 6152 -12408 6388 -12322
rect 6152 -12472 6238 -12408
rect 6238 -12472 6302 -12408
rect 6302 -12472 6388 -12408
rect 6152 -12558 6388 -12472
rect 6152 -12728 6388 -12642
rect 6152 -12792 6238 -12728
rect 6238 -12792 6302 -12728
rect 6302 -12792 6388 -12728
rect 6152 -12878 6388 -12792
rect 6152 -13048 6388 -12962
rect 6152 -13112 6238 -13048
rect 6238 -13112 6302 -13048
rect 6302 -13112 6388 -13048
rect 6152 -13198 6388 -13112
rect 6152 -13368 6388 -13282
rect 6152 -13432 6238 -13368
rect 6238 -13432 6302 -13368
rect 6302 -13432 6388 -13368
rect 6152 -13518 6388 -13432
rect 6152 -13688 6388 -13602
rect 6152 -13752 6238 -13688
rect 6238 -13752 6302 -13688
rect 6302 -13752 6388 -13688
rect 6152 -13838 6388 -13752
rect 6152 -14008 6388 -13922
rect 6152 -14072 6238 -14008
rect 6238 -14072 6302 -14008
rect 6302 -14072 6388 -14008
rect 6152 -14158 6388 -14072
rect 6152 -14328 6388 -14242
rect 6152 -14392 6238 -14328
rect 6238 -14392 6302 -14328
rect 6302 -14392 6388 -14328
rect 6152 -14478 6388 -14392
rect 6152 -14648 6388 -14562
rect 6152 -14712 6238 -14648
rect 6238 -14712 6302 -14648
rect 6302 -14712 6388 -14648
rect 6152 -14798 6388 -14712
rect 6152 -14968 6388 -14882
rect 6152 -15032 6238 -14968
rect 6238 -15032 6302 -14968
rect 6302 -15032 6388 -14968
rect 6152 -15118 6388 -15032
rect 6152 -15288 6388 -15202
rect 6152 -15352 6238 -15288
rect 6238 -15352 6302 -15288
rect 6302 -15352 6388 -15288
rect 6152 -15438 6388 -15352
rect 6152 -15608 6388 -15522
rect 6152 -15672 6238 -15608
rect 6238 -15672 6302 -15608
rect 6302 -15672 6388 -15608
rect 6152 -15758 6388 -15672
rect 6152 -15928 6388 -15842
rect 6152 -15992 6238 -15928
rect 6238 -15992 6302 -15928
rect 6302 -15992 6388 -15928
rect 6152 -16078 6388 -15992
rect 6152 -16248 6388 -16162
rect 6152 -16312 6238 -16248
rect 6238 -16312 6302 -16248
rect 6302 -16312 6388 -16248
rect 6152 -16398 6388 -16312
rect 6152 -16568 6388 -16482
rect 6152 -16632 6238 -16568
rect 6238 -16632 6302 -16568
rect 6302 -16632 6388 -16568
rect 6152 -16718 6388 -16632
rect 6152 -16888 6388 -16802
rect 6152 -16952 6238 -16888
rect 6238 -16952 6302 -16888
rect 6302 -16952 6388 -16888
rect 6152 -17038 6388 -16952
rect 6152 -17208 6388 -17122
rect 6152 -17272 6238 -17208
rect 6238 -17272 6302 -17208
rect 6302 -17272 6388 -17208
rect 6152 -17358 6388 -17272
rect 6152 -17528 6388 -17442
rect 6152 -17592 6238 -17528
rect 6238 -17592 6302 -17528
rect 6302 -17592 6388 -17528
rect 6152 -17678 6388 -17592
rect 6152 -17848 6388 -17762
rect 6152 -17912 6238 -17848
rect 6238 -17912 6302 -17848
rect 6302 -17912 6388 -17848
rect 6152 -17998 6388 -17912
rect 6152 -18168 6388 -18082
rect 6152 -18232 6238 -18168
rect 6238 -18232 6302 -18168
rect 6302 -18232 6388 -18168
rect 6152 -18318 6388 -18232
rect 6152 -18488 6388 -18402
rect 13618 -11598 13854 -11512
rect 13618 -11768 13854 -11682
rect 13618 -11832 13704 -11768
rect 13704 -11832 13768 -11768
rect 13768 -11832 13854 -11768
rect 13618 -11918 13854 -11832
rect 13618 -12088 13854 -12002
rect 13618 -12152 13704 -12088
rect 13704 -12152 13768 -12088
rect 13768 -12152 13854 -12088
rect 13618 -12238 13854 -12152
rect 13618 -12408 13854 -12322
rect 13618 -12472 13704 -12408
rect 13704 -12472 13768 -12408
rect 13768 -12472 13854 -12408
rect 13618 -12558 13854 -12472
rect 13618 -12728 13854 -12642
rect 13618 -12792 13704 -12728
rect 13704 -12792 13768 -12728
rect 13768 -12792 13854 -12728
rect 13618 -12878 13854 -12792
rect 13618 -13048 13854 -12962
rect 13618 -13112 13704 -13048
rect 13704 -13112 13768 -13048
rect 13768 -13112 13854 -13048
rect 13618 -13198 13854 -13112
rect 13618 -13368 13854 -13282
rect 13618 -13432 13704 -13368
rect 13704 -13432 13768 -13368
rect 13768 -13432 13854 -13368
rect 13618 -13518 13854 -13432
rect 13618 -13688 13854 -13602
rect 13618 -13752 13704 -13688
rect 13704 -13752 13768 -13688
rect 13768 -13752 13854 -13688
rect 13618 -13838 13854 -13752
rect 13618 -14008 13854 -13922
rect 13618 -14072 13704 -14008
rect 13704 -14072 13768 -14008
rect 13768 -14072 13854 -14008
rect 13618 -14158 13854 -14072
rect 13618 -14328 13854 -14242
rect 13618 -14392 13704 -14328
rect 13704 -14392 13768 -14328
rect 13768 -14392 13854 -14328
rect 13618 -14478 13854 -14392
rect 13618 -14648 13854 -14562
rect 13618 -14712 13704 -14648
rect 13704 -14712 13768 -14648
rect 13768 -14712 13854 -14648
rect 13618 -14798 13854 -14712
rect 13618 -14968 13854 -14882
rect 13618 -15032 13704 -14968
rect 13704 -15032 13768 -14968
rect 13768 -15032 13854 -14968
rect 13618 -15118 13854 -15032
rect 13618 -15288 13854 -15202
rect 13618 -15352 13704 -15288
rect 13704 -15352 13768 -15288
rect 13768 -15352 13854 -15288
rect 13618 -15438 13854 -15352
rect 13618 -15608 13854 -15522
rect 13618 -15672 13704 -15608
rect 13704 -15672 13768 -15608
rect 13768 -15672 13854 -15608
rect 13618 -15758 13854 -15672
rect 13618 -15928 13854 -15842
rect 13618 -15992 13704 -15928
rect 13704 -15992 13768 -15928
rect 13768 -15992 13854 -15928
rect 13618 -16078 13854 -15992
rect 13618 -16248 13854 -16162
rect 13618 -16312 13704 -16248
rect 13704 -16312 13768 -16248
rect 13768 -16312 13854 -16248
rect 13618 -16398 13854 -16312
rect 13618 -16568 13854 -16482
rect 13618 -16632 13704 -16568
rect 13704 -16632 13768 -16568
rect 13768 -16632 13854 -16568
rect 13618 -16718 13854 -16632
rect 13618 -16888 13854 -16802
rect 13618 -16952 13704 -16888
rect 13704 -16952 13768 -16888
rect 13768 -16952 13854 -16888
rect 13618 -17038 13854 -16952
rect 13618 -17208 13854 -17122
rect 13618 -17272 13704 -17208
rect 13704 -17272 13768 -17208
rect 13768 -17272 13854 -17208
rect 13618 -17358 13854 -17272
rect 13618 -17528 13854 -17442
rect 13618 -17592 13704 -17528
rect 13704 -17592 13768 -17528
rect 13768 -17592 13854 -17528
rect 13618 -17678 13854 -17592
rect 13618 -17848 13854 -17762
rect 13618 -17912 13704 -17848
rect 13704 -17912 13768 -17848
rect 13768 -17912 13854 -17848
rect 13618 -17998 13854 -17912
rect 13618 -18168 13854 -18082
rect 13618 -18232 13704 -18168
rect 13704 -18232 13768 -18168
rect 13768 -18232 13854 -18168
rect 13618 -18318 13854 -18232
rect 6152 -18552 6238 -18488
rect 6238 -18552 6302 -18488
rect 6302 -18552 6388 -18488
rect 6152 -18638 6388 -18552
rect 13618 -18488 13854 -18402
rect 13618 -18552 13704 -18488
rect 13704 -18552 13768 -18488
rect 13768 -18552 13854 -18488
rect 6522 -18698 6758 -18612
rect 6522 -18762 6608 -18698
rect 6608 -18762 6672 -18698
rect 6672 -18762 6758 -18698
rect 6522 -18848 6758 -18762
rect 6842 -18698 7078 -18612
rect 6842 -18762 6928 -18698
rect 6928 -18762 6992 -18698
rect 6992 -18762 7078 -18698
rect 6842 -18848 7078 -18762
rect 7162 -18698 7398 -18612
rect 7162 -18762 7248 -18698
rect 7248 -18762 7312 -18698
rect 7312 -18762 7398 -18698
rect 7162 -18848 7398 -18762
rect 7482 -18698 7718 -18612
rect 7482 -18762 7568 -18698
rect 7568 -18762 7632 -18698
rect 7632 -18762 7718 -18698
rect 7482 -18848 7718 -18762
rect 7802 -18698 8038 -18612
rect 7802 -18762 7888 -18698
rect 7888 -18762 7952 -18698
rect 7952 -18762 8038 -18698
rect 7802 -18848 8038 -18762
rect 8122 -18698 8358 -18612
rect 8122 -18762 8208 -18698
rect 8208 -18762 8272 -18698
rect 8272 -18762 8358 -18698
rect 8122 -18848 8358 -18762
rect 8442 -18698 8678 -18612
rect 8442 -18762 8528 -18698
rect 8528 -18762 8592 -18698
rect 8592 -18762 8678 -18698
rect 8442 -18848 8678 -18762
rect 8762 -18698 8998 -18612
rect 8762 -18762 8848 -18698
rect 8848 -18762 8912 -18698
rect 8912 -18762 8998 -18698
rect 8762 -18848 8998 -18762
rect 9082 -18698 9318 -18612
rect 9082 -18762 9168 -18698
rect 9168 -18762 9232 -18698
rect 9232 -18762 9318 -18698
rect 9082 -18848 9318 -18762
rect 9402 -18698 9638 -18612
rect 9402 -18762 9488 -18698
rect 9488 -18762 9552 -18698
rect 9552 -18762 9638 -18698
rect 9402 -18848 9638 -18762
rect 9722 -18698 9958 -18612
rect 9722 -18762 9808 -18698
rect 9808 -18762 9872 -18698
rect 9872 -18762 9958 -18698
rect 9722 -18848 9958 -18762
rect 10042 -18698 10278 -18612
rect 10042 -18762 10128 -18698
rect 10128 -18762 10192 -18698
rect 10192 -18762 10278 -18698
rect 10042 -18848 10278 -18762
rect 10362 -18698 10598 -18612
rect 10362 -18762 10448 -18698
rect 10448 -18762 10512 -18698
rect 10512 -18762 10598 -18698
rect 10362 -18848 10598 -18762
rect 10682 -18698 10918 -18612
rect 10682 -18762 10768 -18698
rect 10768 -18762 10832 -18698
rect 10832 -18762 10918 -18698
rect 10682 -18848 10918 -18762
rect 11002 -18698 11238 -18612
rect 11002 -18762 11088 -18698
rect 11088 -18762 11152 -18698
rect 11152 -18762 11238 -18698
rect 11002 -18848 11238 -18762
rect 11322 -18698 11558 -18612
rect 11322 -18762 11408 -18698
rect 11408 -18762 11472 -18698
rect 11472 -18762 11558 -18698
rect 11322 -18848 11558 -18762
rect 11642 -18698 11878 -18612
rect 11642 -18762 11728 -18698
rect 11728 -18762 11792 -18698
rect 11792 -18762 11878 -18698
rect 11642 -18848 11878 -18762
rect 11962 -18698 12198 -18612
rect 11962 -18762 12048 -18698
rect 12048 -18762 12112 -18698
rect 12112 -18762 12198 -18698
rect 11962 -18848 12198 -18762
rect 12282 -18698 12518 -18612
rect 12282 -18762 12368 -18698
rect 12368 -18762 12432 -18698
rect 12432 -18762 12518 -18698
rect 12282 -18848 12518 -18762
rect 12602 -18698 12838 -18612
rect 12602 -18762 12688 -18698
rect 12688 -18762 12752 -18698
rect 12752 -18762 12838 -18698
rect 12602 -18848 12838 -18762
rect 12922 -18698 13158 -18612
rect 12922 -18762 13008 -18698
rect 13008 -18762 13072 -18698
rect 13072 -18762 13158 -18698
rect 12922 -18848 13158 -18762
rect 13242 -18698 13478 -18612
rect 13618 -18638 13854 -18552
rect 13242 -18762 13328 -18698
rect 13328 -18762 13392 -18698
rect 13392 -18762 13478 -18698
rect 13242 -18848 13478 -18762
rect 18522 -11242 18758 -11156
rect 18522 -11306 18608 -11242
rect 18608 -11306 18672 -11242
rect 18672 -11306 18758 -11242
rect 18152 -11448 18388 -11362
rect 18522 -11392 18758 -11306
rect 18842 -11242 19078 -11156
rect 18842 -11306 18928 -11242
rect 18928 -11306 18992 -11242
rect 18992 -11306 19078 -11242
rect 18842 -11392 19078 -11306
rect 19162 -11242 19398 -11156
rect 19162 -11306 19248 -11242
rect 19248 -11306 19312 -11242
rect 19312 -11306 19398 -11242
rect 19162 -11392 19398 -11306
rect 19482 -11242 19718 -11156
rect 19482 -11306 19568 -11242
rect 19568 -11306 19632 -11242
rect 19632 -11306 19718 -11242
rect 19482 -11392 19718 -11306
rect 19802 -11242 20038 -11156
rect 19802 -11306 19888 -11242
rect 19888 -11306 19952 -11242
rect 19952 -11306 20038 -11242
rect 19802 -11392 20038 -11306
rect 20122 -11242 20358 -11156
rect 20122 -11306 20208 -11242
rect 20208 -11306 20272 -11242
rect 20272 -11306 20358 -11242
rect 20122 -11392 20358 -11306
rect 20442 -11242 20678 -11156
rect 20442 -11306 20528 -11242
rect 20528 -11306 20592 -11242
rect 20592 -11306 20678 -11242
rect 20442 -11392 20678 -11306
rect 20762 -11242 20998 -11156
rect 20762 -11306 20848 -11242
rect 20848 -11306 20912 -11242
rect 20912 -11306 20998 -11242
rect 20762 -11392 20998 -11306
rect 21082 -11242 21318 -11156
rect 21082 -11306 21168 -11242
rect 21168 -11306 21232 -11242
rect 21232 -11306 21318 -11242
rect 21082 -11392 21318 -11306
rect 21402 -11242 21638 -11156
rect 21402 -11306 21488 -11242
rect 21488 -11306 21552 -11242
rect 21552 -11306 21638 -11242
rect 21402 -11392 21638 -11306
rect 21722 -11242 21958 -11156
rect 21722 -11306 21808 -11242
rect 21808 -11306 21872 -11242
rect 21872 -11306 21958 -11242
rect 21722 -11392 21958 -11306
rect 22042 -11242 22278 -11156
rect 22042 -11306 22128 -11242
rect 22128 -11306 22192 -11242
rect 22192 -11306 22278 -11242
rect 22042 -11392 22278 -11306
rect 22362 -11242 22598 -11156
rect 22362 -11306 22448 -11242
rect 22448 -11306 22512 -11242
rect 22512 -11306 22598 -11242
rect 22362 -11392 22598 -11306
rect 22682 -11242 22918 -11156
rect 22682 -11306 22768 -11242
rect 22768 -11306 22832 -11242
rect 22832 -11306 22918 -11242
rect 22682 -11392 22918 -11306
rect 23002 -11242 23238 -11156
rect 23002 -11306 23088 -11242
rect 23088 -11306 23152 -11242
rect 23152 -11306 23238 -11242
rect 23002 -11392 23238 -11306
rect 23322 -11242 23558 -11156
rect 23322 -11306 23408 -11242
rect 23408 -11306 23472 -11242
rect 23472 -11306 23558 -11242
rect 23322 -11392 23558 -11306
rect 23642 -11242 23878 -11156
rect 23642 -11306 23728 -11242
rect 23728 -11306 23792 -11242
rect 23792 -11306 23878 -11242
rect 23642 -11392 23878 -11306
rect 23962 -11242 24198 -11156
rect 23962 -11306 24048 -11242
rect 24048 -11306 24112 -11242
rect 24112 -11306 24198 -11242
rect 23962 -11392 24198 -11306
rect 24282 -11242 24518 -11156
rect 24282 -11306 24368 -11242
rect 24368 -11306 24432 -11242
rect 24432 -11306 24518 -11242
rect 24282 -11392 24518 -11306
rect 24602 -11242 24838 -11156
rect 24602 -11306 24688 -11242
rect 24688 -11306 24752 -11242
rect 24752 -11306 24838 -11242
rect 24602 -11392 24838 -11306
rect 24922 -11242 25158 -11156
rect 24922 -11306 25008 -11242
rect 25008 -11306 25072 -11242
rect 25072 -11306 25158 -11242
rect 24922 -11392 25158 -11306
rect 25242 -11242 25478 -11156
rect 25242 -11306 25328 -11242
rect 25328 -11306 25392 -11242
rect 25392 -11306 25478 -11242
rect 25242 -11392 25478 -11306
rect 18152 -11512 18238 -11448
rect 18238 -11512 18302 -11448
rect 18302 -11512 18388 -11448
rect 18152 -11598 18388 -11512
rect 25618 -11448 25854 -11362
rect 25618 -11512 25704 -11448
rect 25704 -11512 25768 -11448
rect 25768 -11512 25854 -11448
rect 18152 -11768 18388 -11682
rect 18152 -11832 18238 -11768
rect 18238 -11832 18302 -11768
rect 18302 -11832 18388 -11768
rect 18152 -11918 18388 -11832
rect 18152 -12088 18388 -12002
rect 18152 -12152 18238 -12088
rect 18238 -12152 18302 -12088
rect 18302 -12152 18388 -12088
rect 18152 -12238 18388 -12152
rect 18152 -12408 18388 -12322
rect 18152 -12472 18238 -12408
rect 18238 -12472 18302 -12408
rect 18302 -12472 18388 -12408
rect 18152 -12558 18388 -12472
rect 18152 -12728 18388 -12642
rect 18152 -12792 18238 -12728
rect 18238 -12792 18302 -12728
rect 18302 -12792 18388 -12728
rect 18152 -12878 18388 -12792
rect 18152 -13048 18388 -12962
rect 18152 -13112 18238 -13048
rect 18238 -13112 18302 -13048
rect 18302 -13112 18388 -13048
rect 18152 -13198 18388 -13112
rect 18152 -13368 18388 -13282
rect 18152 -13432 18238 -13368
rect 18238 -13432 18302 -13368
rect 18302 -13432 18388 -13368
rect 18152 -13518 18388 -13432
rect 18152 -13688 18388 -13602
rect 18152 -13752 18238 -13688
rect 18238 -13752 18302 -13688
rect 18302 -13752 18388 -13688
rect 18152 -13838 18388 -13752
rect 18152 -14008 18388 -13922
rect 18152 -14072 18238 -14008
rect 18238 -14072 18302 -14008
rect 18302 -14072 18388 -14008
rect 18152 -14158 18388 -14072
rect 18152 -14328 18388 -14242
rect 18152 -14392 18238 -14328
rect 18238 -14392 18302 -14328
rect 18302 -14392 18388 -14328
rect 18152 -14478 18388 -14392
rect 18152 -14648 18388 -14562
rect 18152 -14712 18238 -14648
rect 18238 -14712 18302 -14648
rect 18302 -14712 18388 -14648
rect 18152 -14798 18388 -14712
rect 18152 -14968 18388 -14882
rect 18152 -15032 18238 -14968
rect 18238 -15032 18302 -14968
rect 18302 -15032 18388 -14968
rect 18152 -15118 18388 -15032
rect 18152 -15288 18388 -15202
rect 18152 -15352 18238 -15288
rect 18238 -15352 18302 -15288
rect 18302 -15352 18388 -15288
rect 18152 -15438 18388 -15352
rect 18152 -15608 18388 -15522
rect 18152 -15672 18238 -15608
rect 18238 -15672 18302 -15608
rect 18302 -15672 18388 -15608
rect 18152 -15758 18388 -15672
rect 18152 -15928 18388 -15842
rect 18152 -15992 18238 -15928
rect 18238 -15992 18302 -15928
rect 18302 -15992 18388 -15928
rect 18152 -16078 18388 -15992
rect 18152 -16248 18388 -16162
rect 18152 -16312 18238 -16248
rect 18238 -16312 18302 -16248
rect 18302 -16312 18388 -16248
rect 18152 -16398 18388 -16312
rect 18152 -16568 18388 -16482
rect 18152 -16632 18238 -16568
rect 18238 -16632 18302 -16568
rect 18302 -16632 18388 -16568
rect 18152 -16718 18388 -16632
rect 18152 -16888 18388 -16802
rect 18152 -16952 18238 -16888
rect 18238 -16952 18302 -16888
rect 18302 -16952 18388 -16888
rect 18152 -17038 18388 -16952
rect 18152 -17208 18388 -17122
rect 18152 -17272 18238 -17208
rect 18238 -17272 18302 -17208
rect 18302 -17272 18388 -17208
rect 18152 -17358 18388 -17272
rect 18152 -17528 18388 -17442
rect 18152 -17592 18238 -17528
rect 18238 -17592 18302 -17528
rect 18302 -17592 18388 -17528
rect 18152 -17678 18388 -17592
rect 18152 -17848 18388 -17762
rect 18152 -17912 18238 -17848
rect 18238 -17912 18302 -17848
rect 18302 -17912 18388 -17848
rect 18152 -17998 18388 -17912
rect 18152 -18168 18388 -18082
rect 18152 -18232 18238 -18168
rect 18238 -18232 18302 -18168
rect 18302 -18232 18388 -18168
rect 18152 -18318 18388 -18232
rect 18152 -18488 18388 -18402
rect 25618 -11598 25854 -11512
rect 25618 -11768 25854 -11682
rect 25618 -11832 25704 -11768
rect 25704 -11832 25768 -11768
rect 25768 -11832 25854 -11768
rect 25618 -11918 25854 -11832
rect 25618 -12088 25854 -12002
rect 25618 -12152 25704 -12088
rect 25704 -12152 25768 -12088
rect 25768 -12152 25854 -12088
rect 25618 -12238 25854 -12152
rect 25618 -12408 25854 -12322
rect 25618 -12472 25704 -12408
rect 25704 -12472 25768 -12408
rect 25768 -12472 25854 -12408
rect 25618 -12558 25854 -12472
rect 25618 -12728 25854 -12642
rect 25618 -12792 25704 -12728
rect 25704 -12792 25768 -12728
rect 25768 -12792 25854 -12728
rect 25618 -12878 25854 -12792
rect 25618 -13048 25854 -12962
rect 25618 -13112 25704 -13048
rect 25704 -13112 25768 -13048
rect 25768 -13112 25854 -13048
rect 25618 -13198 25854 -13112
rect 25618 -13368 25854 -13282
rect 25618 -13432 25704 -13368
rect 25704 -13432 25768 -13368
rect 25768 -13432 25854 -13368
rect 25618 -13518 25854 -13432
rect 25618 -13688 25854 -13602
rect 25618 -13752 25704 -13688
rect 25704 -13752 25768 -13688
rect 25768 -13752 25854 -13688
rect 25618 -13838 25854 -13752
rect 25618 -14008 25854 -13922
rect 25618 -14072 25704 -14008
rect 25704 -14072 25768 -14008
rect 25768 -14072 25854 -14008
rect 25618 -14158 25854 -14072
rect 25618 -14328 25854 -14242
rect 25618 -14392 25704 -14328
rect 25704 -14392 25768 -14328
rect 25768 -14392 25854 -14328
rect 25618 -14478 25854 -14392
rect 25618 -14648 25854 -14562
rect 25618 -14712 25704 -14648
rect 25704 -14712 25768 -14648
rect 25768 -14712 25854 -14648
rect 25618 -14798 25854 -14712
rect 25618 -14968 25854 -14882
rect 25618 -15032 25704 -14968
rect 25704 -15032 25768 -14968
rect 25768 -15032 25854 -14968
rect 25618 -15118 25854 -15032
rect 25618 -15288 25854 -15202
rect 25618 -15352 25704 -15288
rect 25704 -15352 25768 -15288
rect 25768 -15352 25854 -15288
rect 25618 -15438 25854 -15352
rect 25618 -15608 25854 -15522
rect 25618 -15672 25704 -15608
rect 25704 -15672 25768 -15608
rect 25768 -15672 25854 -15608
rect 25618 -15758 25854 -15672
rect 25618 -15928 25854 -15842
rect 25618 -15992 25704 -15928
rect 25704 -15992 25768 -15928
rect 25768 -15992 25854 -15928
rect 25618 -16078 25854 -15992
rect 25618 -16248 25854 -16162
rect 25618 -16312 25704 -16248
rect 25704 -16312 25768 -16248
rect 25768 -16312 25854 -16248
rect 25618 -16398 25854 -16312
rect 25618 -16568 25854 -16482
rect 25618 -16632 25704 -16568
rect 25704 -16632 25768 -16568
rect 25768 -16632 25854 -16568
rect 25618 -16718 25854 -16632
rect 25618 -16888 25854 -16802
rect 25618 -16952 25704 -16888
rect 25704 -16952 25768 -16888
rect 25768 -16952 25854 -16888
rect 25618 -17038 25854 -16952
rect 25618 -17208 25854 -17122
rect 25618 -17272 25704 -17208
rect 25704 -17272 25768 -17208
rect 25768 -17272 25854 -17208
rect 25618 -17358 25854 -17272
rect 25618 -17528 25854 -17442
rect 25618 -17592 25704 -17528
rect 25704 -17592 25768 -17528
rect 25768 -17592 25854 -17528
rect 25618 -17678 25854 -17592
rect 25618 -17848 25854 -17762
rect 25618 -17912 25704 -17848
rect 25704 -17912 25768 -17848
rect 25768 -17912 25854 -17848
rect 25618 -17998 25854 -17912
rect 25618 -18168 25854 -18082
rect 25618 -18232 25704 -18168
rect 25704 -18232 25768 -18168
rect 25768 -18232 25854 -18168
rect 25618 -18318 25854 -18232
rect 18152 -18552 18238 -18488
rect 18238 -18552 18302 -18488
rect 18302 -18552 18388 -18488
rect 18152 -18638 18388 -18552
rect 25618 -18488 25854 -18402
rect 25618 -18552 25704 -18488
rect 25704 -18552 25768 -18488
rect 25768 -18552 25854 -18488
rect 18522 -18698 18758 -18612
rect 18522 -18762 18608 -18698
rect 18608 -18762 18672 -18698
rect 18672 -18762 18758 -18698
rect 18522 -18848 18758 -18762
rect 18842 -18698 19078 -18612
rect 18842 -18762 18928 -18698
rect 18928 -18762 18992 -18698
rect 18992 -18762 19078 -18698
rect 18842 -18848 19078 -18762
rect 19162 -18698 19398 -18612
rect 19162 -18762 19248 -18698
rect 19248 -18762 19312 -18698
rect 19312 -18762 19398 -18698
rect 19162 -18848 19398 -18762
rect 19482 -18698 19718 -18612
rect 19482 -18762 19568 -18698
rect 19568 -18762 19632 -18698
rect 19632 -18762 19718 -18698
rect 19482 -18848 19718 -18762
rect 19802 -18698 20038 -18612
rect 19802 -18762 19888 -18698
rect 19888 -18762 19952 -18698
rect 19952 -18762 20038 -18698
rect 19802 -18848 20038 -18762
rect 20122 -18698 20358 -18612
rect 20122 -18762 20208 -18698
rect 20208 -18762 20272 -18698
rect 20272 -18762 20358 -18698
rect 20122 -18848 20358 -18762
rect 20442 -18698 20678 -18612
rect 20442 -18762 20528 -18698
rect 20528 -18762 20592 -18698
rect 20592 -18762 20678 -18698
rect 20442 -18848 20678 -18762
rect 20762 -18698 20998 -18612
rect 20762 -18762 20848 -18698
rect 20848 -18762 20912 -18698
rect 20912 -18762 20998 -18698
rect 20762 -18848 20998 -18762
rect 21082 -18698 21318 -18612
rect 21082 -18762 21168 -18698
rect 21168 -18762 21232 -18698
rect 21232 -18762 21318 -18698
rect 21082 -18848 21318 -18762
rect 21402 -18698 21638 -18612
rect 21402 -18762 21488 -18698
rect 21488 -18762 21552 -18698
rect 21552 -18762 21638 -18698
rect 21402 -18848 21638 -18762
rect 21722 -18698 21958 -18612
rect 21722 -18762 21808 -18698
rect 21808 -18762 21872 -18698
rect 21872 -18762 21958 -18698
rect 21722 -18848 21958 -18762
rect 22042 -18698 22278 -18612
rect 22042 -18762 22128 -18698
rect 22128 -18762 22192 -18698
rect 22192 -18762 22278 -18698
rect 22042 -18848 22278 -18762
rect 22362 -18698 22598 -18612
rect 22362 -18762 22448 -18698
rect 22448 -18762 22512 -18698
rect 22512 -18762 22598 -18698
rect 22362 -18848 22598 -18762
rect 22682 -18698 22918 -18612
rect 22682 -18762 22768 -18698
rect 22768 -18762 22832 -18698
rect 22832 -18762 22918 -18698
rect 22682 -18848 22918 -18762
rect 23002 -18698 23238 -18612
rect 23002 -18762 23088 -18698
rect 23088 -18762 23152 -18698
rect 23152 -18762 23238 -18698
rect 23002 -18848 23238 -18762
rect 23322 -18698 23558 -18612
rect 23322 -18762 23408 -18698
rect 23408 -18762 23472 -18698
rect 23472 -18762 23558 -18698
rect 23322 -18848 23558 -18762
rect 23642 -18698 23878 -18612
rect 23642 -18762 23728 -18698
rect 23728 -18762 23792 -18698
rect 23792 -18762 23878 -18698
rect 23642 -18848 23878 -18762
rect 23962 -18698 24198 -18612
rect 23962 -18762 24048 -18698
rect 24048 -18762 24112 -18698
rect 24112 -18762 24198 -18698
rect 23962 -18848 24198 -18762
rect 24282 -18698 24518 -18612
rect 24282 -18762 24368 -18698
rect 24368 -18762 24432 -18698
rect 24432 -18762 24518 -18698
rect 24282 -18848 24518 -18762
rect 24602 -18698 24838 -18612
rect 24602 -18762 24688 -18698
rect 24688 -18762 24752 -18698
rect 24752 -18762 24838 -18698
rect 24602 -18848 24838 -18762
rect 24922 -18698 25158 -18612
rect 24922 -18762 25008 -18698
rect 25008 -18762 25072 -18698
rect 25072 -18762 25158 -18698
rect 24922 -18848 25158 -18762
rect 25242 -18698 25478 -18612
rect 25618 -18638 25854 -18552
rect 25242 -18762 25328 -18698
rect 25328 -18762 25392 -18698
rect 25392 -18762 25478 -18698
rect 25242 -18848 25478 -18762
rect 30522 -11242 30758 -11156
rect 30522 -11306 30608 -11242
rect 30608 -11306 30672 -11242
rect 30672 -11306 30758 -11242
rect 30152 -11448 30388 -11362
rect 30522 -11392 30758 -11306
rect 30842 -11242 31078 -11156
rect 30842 -11306 30928 -11242
rect 30928 -11306 30992 -11242
rect 30992 -11306 31078 -11242
rect 30842 -11392 31078 -11306
rect 31162 -11242 31398 -11156
rect 31162 -11306 31248 -11242
rect 31248 -11306 31312 -11242
rect 31312 -11306 31398 -11242
rect 31162 -11392 31398 -11306
rect 31482 -11242 31718 -11156
rect 31482 -11306 31568 -11242
rect 31568 -11306 31632 -11242
rect 31632 -11306 31718 -11242
rect 31482 -11392 31718 -11306
rect 31802 -11242 32038 -11156
rect 31802 -11306 31888 -11242
rect 31888 -11306 31952 -11242
rect 31952 -11306 32038 -11242
rect 31802 -11392 32038 -11306
rect 32122 -11242 32358 -11156
rect 32122 -11306 32208 -11242
rect 32208 -11306 32272 -11242
rect 32272 -11306 32358 -11242
rect 32122 -11392 32358 -11306
rect 32442 -11242 32678 -11156
rect 32442 -11306 32528 -11242
rect 32528 -11306 32592 -11242
rect 32592 -11306 32678 -11242
rect 32442 -11392 32678 -11306
rect 32762 -11242 32998 -11156
rect 32762 -11306 32848 -11242
rect 32848 -11306 32912 -11242
rect 32912 -11306 32998 -11242
rect 32762 -11392 32998 -11306
rect 33082 -11242 33318 -11156
rect 33082 -11306 33168 -11242
rect 33168 -11306 33232 -11242
rect 33232 -11306 33318 -11242
rect 33082 -11392 33318 -11306
rect 33402 -11242 33638 -11156
rect 33402 -11306 33488 -11242
rect 33488 -11306 33552 -11242
rect 33552 -11306 33638 -11242
rect 33402 -11392 33638 -11306
rect 33722 -11242 33958 -11156
rect 33722 -11306 33808 -11242
rect 33808 -11306 33872 -11242
rect 33872 -11306 33958 -11242
rect 33722 -11392 33958 -11306
rect 34042 -11242 34278 -11156
rect 34042 -11306 34128 -11242
rect 34128 -11306 34192 -11242
rect 34192 -11306 34278 -11242
rect 34042 -11392 34278 -11306
rect 34362 -11242 34598 -11156
rect 34362 -11306 34448 -11242
rect 34448 -11306 34512 -11242
rect 34512 -11306 34598 -11242
rect 34362 -11392 34598 -11306
rect 34682 -11242 34918 -11156
rect 34682 -11306 34768 -11242
rect 34768 -11306 34832 -11242
rect 34832 -11306 34918 -11242
rect 34682 -11392 34918 -11306
rect 35002 -11242 35238 -11156
rect 35002 -11306 35088 -11242
rect 35088 -11306 35152 -11242
rect 35152 -11306 35238 -11242
rect 35002 -11392 35238 -11306
rect 35322 -11242 35558 -11156
rect 35322 -11306 35408 -11242
rect 35408 -11306 35472 -11242
rect 35472 -11306 35558 -11242
rect 35322 -11392 35558 -11306
rect 35642 -11242 35878 -11156
rect 35642 -11306 35728 -11242
rect 35728 -11306 35792 -11242
rect 35792 -11306 35878 -11242
rect 35642 -11392 35878 -11306
rect 35962 -11242 36198 -11156
rect 35962 -11306 36048 -11242
rect 36048 -11306 36112 -11242
rect 36112 -11306 36198 -11242
rect 35962 -11392 36198 -11306
rect 36282 -11242 36518 -11156
rect 36282 -11306 36368 -11242
rect 36368 -11306 36432 -11242
rect 36432 -11306 36518 -11242
rect 36282 -11392 36518 -11306
rect 36602 -11242 36838 -11156
rect 36602 -11306 36688 -11242
rect 36688 -11306 36752 -11242
rect 36752 -11306 36838 -11242
rect 36602 -11392 36838 -11306
rect 36922 -11242 37158 -11156
rect 36922 -11306 37008 -11242
rect 37008 -11306 37072 -11242
rect 37072 -11306 37158 -11242
rect 36922 -11392 37158 -11306
rect 37242 -11242 37478 -11156
rect 37242 -11306 37328 -11242
rect 37328 -11306 37392 -11242
rect 37392 -11306 37478 -11242
rect 37242 -11392 37478 -11306
rect 30152 -11512 30238 -11448
rect 30238 -11512 30302 -11448
rect 30302 -11512 30388 -11448
rect 30152 -11598 30388 -11512
rect 37618 -11448 37854 -11362
rect 37618 -11512 37704 -11448
rect 37704 -11512 37768 -11448
rect 37768 -11512 37854 -11448
rect 30152 -11768 30388 -11682
rect 30152 -11832 30238 -11768
rect 30238 -11832 30302 -11768
rect 30302 -11832 30388 -11768
rect 30152 -11918 30388 -11832
rect 30152 -12088 30388 -12002
rect 30152 -12152 30238 -12088
rect 30238 -12152 30302 -12088
rect 30302 -12152 30388 -12088
rect 30152 -12238 30388 -12152
rect 30152 -12408 30388 -12322
rect 30152 -12472 30238 -12408
rect 30238 -12472 30302 -12408
rect 30302 -12472 30388 -12408
rect 30152 -12558 30388 -12472
rect 30152 -12728 30388 -12642
rect 30152 -12792 30238 -12728
rect 30238 -12792 30302 -12728
rect 30302 -12792 30388 -12728
rect 30152 -12878 30388 -12792
rect 30152 -13048 30388 -12962
rect 30152 -13112 30238 -13048
rect 30238 -13112 30302 -13048
rect 30302 -13112 30388 -13048
rect 30152 -13198 30388 -13112
rect 30152 -13368 30388 -13282
rect 30152 -13432 30238 -13368
rect 30238 -13432 30302 -13368
rect 30302 -13432 30388 -13368
rect 30152 -13518 30388 -13432
rect 30152 -13688 30388 -13602
rect 30152 -13752 30238 -13688
rect 30238 -13752 30302 -13688
rect 30302 -13752 30388 -13688
rect 30152 -13838 30388 -13752
rect 30152 -14008 30388 -13922
rect 30152 -14072 30238 -14008
rect 30238 -14072 30302 -14008
rect 30302 -14072 30388 -14008
rect 30152 -14158 30388 -14072
rect 30152 -14328 30388 -14242
rect 30152 -14392 30238 -14328
rect 30238 -14392 30302 -14328
rect 30302 -14392 30388 -14328
rect 30152 -14478 30388 -14392
rect 30152 -14648 30388 -14562
rect 30152 -14712 30238 -14648
rect 30238 -14712 30302 -14648
rect 30302 -14712 30388 -14648
rect 30152 -14798 30388 -14712
rect 30152 -14968 30388 -14882
rect 30152 -15032 30238 -14968
rect 30238 -15032 30302 -14968
rect 30302 -15032 30388 -14968
rect 30152 -15118 30388 -15032
rect 30152 -15288 30388 -15202
rect 30152 -15352 30238 -15288
rect 30238 -15352 30302 -15288
rect 30302 -15352 30388 -15288
rect 30152 -15438 30388 -15352
rect 30152 -15608 30388 -15522
rect 30152 -15672 30238 -15608
rect 30238 -15672 30302 -15608
rect 30302 -15672 30388 -15608
rect 30152 -15758 30388 -15672
rect 30152 -15928 30388 -15842
rect 30152 -15992 30238 -15928
rect 30238 -15992 30302 -15928
rect 30302 -15992 30388 -15928
rect 30152 -16078 30388 -15992
rect 30152 -16248 30388 -16162
rect 30152 -16312 30238 -16248
rect 30238 -16312 30302 -16248
rect 30302 -16312 30388 -16248
rect 30152 -16398 30388 -16312
rect 30152 -16568 30388 -16482
rect 30152 -16632 30238 -16568
rect 30238 -16632 30302 -16568
rect 30302 -16632 30388 -16568
rect 30152 -16718 30388 -16632
rect 30152 -16888 30388 -16802
rect 30152 -16952 30238 -16888
rect 30238 -16952 30302 -16888
rect 30302 -16952 30388 -16888
rect 30152 -17038 30388 -16952
rect 30152 -17208 30388 -17122
rect 30152 -17272 30238 -17208
rect 30238 -17272 30302 -17208
rect 30302 -17272 30388 -17208
rect 30152 -17358 30388 -17272
rect 30152 -17528 30388 -17442
rect 30152 -17592 30238 -17528
rect 30238 -17592 30302 -17528
rect 30302 -17592 30388 -17528
rect 30152 -17678 30388 -17592
rect 30152 -17848 30388 -17762
rect 30152 -17912 30238 -17848
rect 30238 -17912 30302 -17848
rect 30302 -17912 30388 -17848
rect 30152 -17998 30388 -17912
rect 30152 -18168 30388 -18082
rect 30152 -18232 30238 -18168
rect 30238 -18232 30302 -18168
rect 30302 -18232 30388 -18168
rect 30152 -18318 30388 -18232
rect 30152 -18488 30388 -18402
rect 37618 -11598 37854 -11512
rect 37618 -11768 37854 -11682
rect 37618 -11832 37704 -11768
rect 37704 -11832 37768 -11768
rect 37768 -11832 37854 -11768
rect 37618 -11918 37854 -11832
rect 37618 -12088 37854 -12002
rect 37618 -12152 37704 -12088
rect 37704 -12152 37768 -12088
rect 37768 -12152 37854 -12088
rect 37618 -12238 37854 -12152
rect 37618 -12408 37854 -12322
rect 37618 -12472 37704 -12408
rect 37704 -12472 37768 -12408
rect 37768 -12472 37854 -12408
rect 37618 -12558 37854 -12472
rect 37618 -12728 37854 -12642
rect 37618 -12792 37704 -12728
rect 37704 -12792 37768 -12728
rect 37768 -12792 37854 -12728
rect 37618 -12878 37854 -12792
rect 37618 -13048 37854 -12962
rect 37618 -13112 37704 -13048
rect 37704 -13112 37768 -13048
rect 37768 -13112 37854 -13048
rect 37618 -13198 37854 -13112
rect 37618 -13368 37854 -13282
rect 37618 -13432 37704 -13368
rect 37704 -13432 37768 -13368
rect 37768 -13432 37854 -13368
rect 37618 -13518 37854 -13432
rect 37618 -13688 37854 -13602
rect 37618 -13752 37704 -13688
rect 37704 -13752 37768 -13688
rect 37768 -13752 37854 -13688
rect 37618 -13838 37854 -13752
rect 37618 -14008 37854 -13922
rect 37618 -14072 37704 -14008
rect 37704 -14072 37768 -14008
rect 37768 -14072 37854 -14008
rect 37618 -14158 37854 -14072
rect 37618 -14328 37854 -14242
rect 37618 -14392 37704 -14328
rect 37704 -14392 37768 -14328
rect 37768 -14392 37854 -14328
rect 37618 -14478 37854 -14392
rect 37618 -14648 37854 -14562
rect 37618 -14712 37704 -14648
rect 37704 -14712 37768 -14648
rect 37768 -14712 37854 -14648
rect 37618 -14798 37854 -14712
rect 37618 -14968 37854 -14882
rect 37618 -15032 37704 -14968
rect 37704 -15032 37768 -14968
rect 37768 -15032 37854 -14968
rect 37618 -15118 37854 -15032
rect 37618 -15288 37854 -15202
rect 37618 -15352 37704 -15288
rect 37704 -15352 37768 -15288
rect 37768 -15352 37854 -15288
rect 37618 -15438 37854 -15352
rect 37618 -15608 37854 -15522
rect 37618 -15672 37704 -15608
rect 37704 -15672 37768 -15608
rect 37768 -15672 37854 -15608
rect 37618 -15758 37854 -15672
rect 37618 -15928 37854 -15842
rect 37618 -15992 37704 -15928
rect 37704 -15992 37768 -15928
rect 37768 -15992 37854 -15928
rect 37618 -16078 37854 -15992
rect 37618 -16248 37854 -16162
rect 37618 -16312 37704 -16248
rect 37704 -16312 37768 -16248
rect 37768 -16312 37854 -16248
rect 37618 -16398 37854 -16312
rect 37618 -16568 37854 -16482
rect 37618 -16632 37704 -16568
rect 37704 -16632 37768 -16568
rect 37768 -16632 37854 -16568
rect 37618 -16718 37854 -16632
rect 37618 -16888 37854 -16802
rect 37618 -16952 37704 -16888
rect 37704 -16952 37768 -16888
rect 37768 -16952 37854 -16888
rect 37618 -17038 37854 -16952
rect 37618 -17208 37854 -17122
rect 37618 -17272 37704 -17208
rect 37704 -17272 37768 -17208
rect 37768 -17272 37854 -17208
rect 37618 -17358 37854 -17272
rect 37618 -17528 37854 -17442
rect 37618 -17592 37704 -17528
rect 37704 -17592 37768 -17528
rect 37768 -17592 37854 -17528
rect 37618 -17678 37854 -17592
rect 37618 -17848 37854 -17762
rect 37618 -17912 37704 -17848
rect 37704 -17912 37768 -17848
rect 37768 -17912 37854 -17848
rect 37618 -17998 37854 -17912
rect 37618 -18168 37854 -18082
rect 37618 -18232 37704 -18168
rect 37704 -18232 37768 -18168
rect 37768 -18232 37854 -18168
rect 37618 -18318 37854 -18232
rect 30152 -18552 30238 -18488
rect 30238 -18552 30302 -18488
rect 30302 -18552 30388 -18488
rect 30152 -18638 30388 -18552
rect 37618 -18488 37854 -18402
rect 37618 -18552 37704 -18488
rect 37704 -18552 37768 -18488
rect 37768 -18552 37854 -18488
rect 30522 -18698 30758 -18612
rect 30522 -18762 30608 -18698
rect 30608 -18762 30672 -18698
rect 30672 -18762 30758 -18698
rect 30522 -18848 30758 -18762
rect 30842 -18698 31078 -18612
rect 30842 -18762 30928 -18698
rect 30928 -18762 30992 -18698
rect 30992 -18762 31078 -18698
rect 30842 -18848 31078 -18762
rect 31162 -18698 31398 -18612
rect 31162 -18762 31248 -18698
rect 31248 -18762 31312 -18698
rect 31312 -18762 31398 -18698
rect 31162 -18848 31398 -18762
rect 31482 -18698 31718 -18612
rect 31482 -18762 31568 -18698
rect 31568 -18762 31632 -18698
rect 31632 -18762 31718 -18698
rect 31482 -18848 31718 -18762
rect 31802 -18698 32038 -18612
rect 31802 -18762 31888 -18698
rect 31888 -18762 31952 -18698
rect 31952 -18762 32038 -18698
rect 31802 -18848 32038 -18762
rect 32122 -18698 32358 -18612
rect 32122 -18762 32208 -18698
rect 32208 -18762 32272 -18698
rect 32272 -18762 32358 -18698
rect 32122 -18848 32358 -18762
rect 32442 -18698 32678 -18612
rect 32442 -18762 32528 -18698
rect 32528 -18762 32592 -18698
rect 32592 -18762 32678 -18698
rect 32442 -18848 32678 -18762
rect 32762 -18698 32998 -18612
rect 32762 -18762 32848 -18698
rect 32848 -18762 32912 -18698
rect 32912 -18762 32998 -18698
rect 32762 -18848 32998 -18762
rect 33082 -18698 33318 -18612
rect 33082 -18762 33168 -18698
rect 33168 -18762 33232 -18698
rect 33232 -18762 33318 -18698
rect 33082 -18848 33318 -18762
rect 33402 -18698 33638 -18612
rect 33402 -18762 33488 -18698
rect 33488 -18762 33552 -18698
rect 33552 -18762 33638 -18698
rect 33402 -18848 33638 -18762
rect 33722 -18698 33958 -18612
rect 33722 -18762 33808 -18698
rect 33808 -18762 33872 -18698
rect 33872 -18762 33958 -18698
rect 33722 -18848 33958 -18762
rect 34042 -18698 34278 -18612
rect 34042 -18762 34128 -18698
rect 34128 -18762 34192 -18698
rect 34192 -18762 34278 -18698
rect 34042 -18848 34278 -18762
rect 34362 -18698 34598 -18612
rect 34362 -18762 34448 -18698
rect 34448 -18762 34512 -18698
rect 34512 -18762 34598 -18698
rect 34362 -18848 34598 -18762
rect 34682 -18698 34918 -18612
rect 34682 -18762 34768 -18698
rect 34768 -18762 34832 -18698
rect 34832 -18762 34918 -18698
rect 34682 -18848 34918 -18762
rect 35002 -18698 35238 -18612
rect 35002 -18762 35088 -18698
rect 35088 -18762 35152 -18698
rect 35152 -18762 35238 -18698
rect 35002 -18848 35238 -18762
rect 35322 -18698 35558 -18612
rect 35322 -18762 35408 -18698
rect 35408 -18762 35472 -18698
rect 35472 -18762 35558 -18698
rect 35322 -18848 35558 -18762
rect 35642 -18698 35878 -18612
rect 35642 -18762 35728 -18698
rect 35728 -18762 35792 -18698
rect 35792 -18762 35878 -18698
rect 35642 -18848 35878 -18762
rect 35962 -18698 36198 -18612
rect 35962 -18762 36048 -18698
rect 36048 -18762 36112 -18698
rect 36112 -18762 36198 -18698
rect 35962 -18848 36198 -18762
rect 36282 -18698 36518 -18612
rect 36282 -18762 36368 -18698
rect 36368 -18762 36432 -18698
rect 36432 -18762 36518 -18698
rect 36282 -18848 36518 -18762
rect 36602 -18698 36838 -18612
rect 36602 -18762 36688 -18698
rect 36688 -18762 36752 -18698
rect 36752 -18762 36838 -18698
rect 36602 -18848 36838 -18762
rect 36922 -18698 37158 -18612
rect 36922 -18762 37008 -18698
rect 37008 -18762 37072 -18698
rect 37072 -18762 37158 -18698
rect 36922 -18848 37158 -18762
rect 37242 -18698 37478 -18612
rect 37618 -18638 37854 -18552
rect 37242 -18762 37328 -18698
rect 37328 -18762 37392 -18698
rect 37392 -18762 37478 -18698
rect 37242 -18848 37478 -18762
rect 42522 -11242 42758 -11156
rect 42522 -11306 42608 -11242
rect 42608 -11306 42672 -11242
rect 42672 -11306 42758 -11242
rect 42155 -11448 42391 -11362
rect 42522 -11392 42758 -11306
rect 42842 -11242 43078 -11156
rect 42842 -11306 42928 -11242
rect 42928 -11306 42992 -11242
rect 42992 -11306 43078 -11242
rect 42842 -11392 43078 -11306
rect 43162 -11242 43398 -11156
rect 43162 -11306 43248 -11242
rect 43248 -11306 43312 -11242
rect 43312 -11306 43398 -11242
rect 43162 -11392 43398 -11306
rect 43482 -11242 43718 -11156
rect 43482 -11306 43568 -11242
rect 43568 -11306 43632 -11242
rect 43632 -11306 43718 -11242
rect 43482 -11392 43718 -11306
rect 43802 -11242 44038 -11156
rect 43802 -11306 43888 -11242
rect 43888 -11306 43952 -11242
rect 43952 -11306 44038 -11242
rect 43802 -11392 44038 -11306
rect 44122 -11242 44358 -11156
rect 44122 -11306 44208 -11242
rect 44208 -11306 44272 -11242
rect 44272 -11306 44358 -11242
rect 44122 -11392 44358 -11306
rect 44442 -11242 44678 -11156
rect 44442 -11306 44528 -11242
rect 44528 -11306 44592 -11242
rect 44592 -11306 44678 -11242
rect 44442 -11392 44678 -11306
rect 44762 -11242 44998 -11156
rect 44762 -11306 44848 -11242
rect 44848 -11306 44912 -11242
rect 44912 -11306 44998 -11242
rect 44762 -11392 44998 -11306
rect 45082 -11242 45318 -11156
rect 45082 -11306 45168 -11242
rect 45168 -11306 45232 -11242
rect 45232 -11306 45318 -11242
rect 45082 -11392 45318 -11306
rect 45402 -11242 45638 -11156
rect 45402 -11306 45488 -11242
rect 45488 -11306 45552 -11242
rect 45552 -11306 45638 -11242
rect 45402 -11392 45638 -11306
rect 45722 -11242 45958 -11156
rect 45722 -11306 45808 -11242
rect 45808 -11306 45872 -11242
rect 45872 -11306 45958 -11242
rect 45722 -11392 45958 -11306
rect 46042 -11242 46278 -11156
rect 46042 -11306 46128 -11242
rect 46128 -11306 46192 -11242
rect 46192 -11306 46278 -11242
rect 46042 -11392 46278 -11306
rect 46362 -11242 46598 -11156
rect 46362 -11306 46448 -11242
rect 46448 -11306 46512 -11242
rect 46512 -11306 46598 -11242
rect 46362 -11392 46598 -11306
rect 46682 -11242 46918 -11156
rect 46682 -11306 46768 -11242
rect 46768 -11306 46832 -11242
rect 46832 -11306 46918 -11242
rect 46682 -11392 46918 -11306
rect 47002 -11242 47238 -11156
rect 47002 -11306 47088 -11242
rect 47088 -11306 47152 -11242
rect 47152 -11306 47238 -11242
rect 47002 -11392 47238 -11306
rect 47322 -11242 47558 -11156
rect 47322 -11306 47408 -11242
rect 47408 -11306 47472 -11242
rect 47472 -11306 47558 -11242
rect 47322 -11392 47558 -11306
rect 47642 -11242 47878 -11156
rect 47642 -11306 47728 -11242
rect 47728 -11306 47792 -11242
rect 47792 -11306 47878 -11242
rect 47642 -11392 47878 -11306
rect 47962 -11242 48198 -11156
rect 47962 -11306 48048 -11242
rect 48048 -11306 48112 -11242
rect 48112 -11306 48198 -11242
rect 47962 -11392 48198 -11306
rect 48282 -11242 48518 -11156
rect 48282 -11306 48368 -11242
rect 48368 -11306 48432 -11242
rect 48432 -11306 48518 -11242
rect 48282 -11392 48518 -11306
rect 48602 -11242 48838 -11156
rect 48602 -11306 48688 -11242
rect 48688 -11306 48752 -11242
rect 48752 -11306 48838 -11242
rect 48602 -11392 48838 -11306
rect 48922 -11242 49158 -11156
rect 48922 -11306 49008 -11242
rect 49008 -11306 49072 -11242
rect 49072 -11306 49158 -11242
rect 48922 -11392 49158 -11306
rect 49242 -11242 49478 -11156
rect 49242 -11306 49328 -11242
rect 49328 -11306 49392 -11242
rect 49392 -11306 49478 -11242
rect 49242 -11392 49478 -11306
rect 42155 -11512 42241 -11448
rect 42241 -11512 42305 -11448
rect 42305 -11512 42391 -11448
rect 42155 -11598 42391 -11512
rect 49609 -11448 49845 -11362
rect 49609 -11512 49695 -11448
rect 49695 -11512 49759 -11448
rect 49759 -11512 49845 -11448
rect 42155 -11768 42391 -11682
rect 42155 -11832 42241 -11768
rect 42241 -11832 42305 -11768
rect 42305 -11832 42391 -11768
rect 42155 -11918 42391 -11832
rect 42155 -12088 42391 -12002
rect 42155 -12152 42241 -12088
rect 42241 -12152 42305 -12088
rect 42305 -12152 42391 -12088
rect 42155 -12238 42391 -12152
rect 42155 -12408 42391 -12322
rect 42155 -12472 42241 -12408
rect 42241 -12472 42305 -12408
rect 42305 -12472 42391 -12408
rect 42155 -12558 42391 -12472
rect 42155 -12728 42391 -12642
rect 42155 -12792 42241 -12728
rect 42241 -12792 42305 -12728
rect 42305 -12792 42391 -12728
rect 42155 -12878 42391 -12792
rect 42155 -13048 42391 -12962
rect 42155 -13112 42241 -13048
rect 42241 -13112 42305 -13048
rect 42305 -13112 42391 -13048
rect 42155 -13198 42391 -13112
rect 42155 -13368 42391 -13282
rect 42155 -13432 42241 -13368
rect 42241 -13432 42305 -13368
rect 42305 -13432 42391 -13368
rect 42155 -13518 42391 -13432
rect 42155 -13688 42391 -13602
rect 42155 -13752 42241 -13688
rect 42241 -13752 42305 -13688
rect 42305 -13752 42391 -13688
rect 42155 -13838 42391 -13752
rect 42155 -14008 42391 -13922
rect 42155 -14072 42241 -14008
rect 42241 -14072 42305 -14008
rect 42305 -14072 42391 -14008
rect 42155 -14158 42391 -14072
rect 42155 -14328 42391 -14242
rect 42155 -14392 42241 -14328
rect 42241 -14392 42305 -14328
rect 42305 -14392 42391 -14328
rect 42155 -14478 42391 -14392
rect 42155 -14648 42391 -14562
rect 42155 -14712 42241 -14648
rect 42241 -14712 42305 -14648
rect 42305 -14712 42391 -14648
rect 42155 -14798 42391 -14712
rect 42155 -14968 42391 -14882
rect 42155 -15032 42241 -14968
rect 42241 -15032 42305 -14968
rect 42305 -15032 42391 -14968
rect 42155 -15118 42391 -15032
rect 42155 -15288 42391 -15202
rect 42155 -15352 42241 -15288
rect 42241 -15352 42305 -15288
rect 42305 -15352 42391 -15288
rect 42155 -15438 42391 -15352
rect 42155 -15608 42391 -15522
rect 42155 -15672 42241 -15608
rect 42241 -15672 42305 -15608
rect 42305 -15672 42391 -15608
rect 42155 -15758 42391 -15672
rect 42155 -15928 42391 -15842
rect 42155 -15992 42241 -15928
rect 42241 -15992 42305 -15928
rect 42305 -15992 42391 -15928
rect 42155 -16078 42391 -15992
rect 42155 -16248 42391 -16162
rect 42155 -16312 42241 -16248
rect 42241 -16312 42305 -16248
rect 42305 -16312 42391 -16248
rect 42155 -16398 42391 -16312
rect 42155 -16568 42391 -16482
rect 42155 -16632 42241 -16568
rect 42241 -16632 42305 -16568
rect 42305 -16632 42391 -16568
rect 42155 -16718 42391 -16632
rect 42155 -16888 42391 -16802
rect 42155 -16952 42241 -16888
rect 42241 -16952 42305 -16888
rect 42305 -16952 42391 -16888
rect 42155 -17038 42391 -16952
rect 42155 -17208 42391 -17122
rect 42155 -17272 42241 -17208
rect 42241 -17272 42305 -17208
rect 42305 -17272 42391 -17208
rect 42155 -17358 42391 -17272
rect 42155 -17528 42391 -17442
rect 42155 -17592 42241 -17528
rect 42241 -17592 42305 -17528
rect 42305 -17592 42391 -17528
rect 42155 -17678 42391 -17592
rect 42155 -17848 42391 -17762
rect 42155 -17912 42241 -17848
rect 42241 -17912 42305 -17848
rect 42305 -17912 42391 -17848
rect 42155 -17998 42391 -17912
rect 42155 -18168 42391 -18082
rect 42155 -18232 42241 -18168
rect 42241 -18232 42305 -18168
rect 42305 -18232 42391 -18168
rect 42155 -18318 42391 -18232
rect 42155 -18488 42391 -18402
rect 49609 -11598 49845 -11512
rect 49609 -11768 49845 -11682
rect 49609 -11832 49695 -11768
rect 49695 -11832 49759 -11768
rect 49759 -11832 49845 -11768
rect 49609 -11918 49845 -11832
rect 49609 -12088 49845 -12002
rect 49609 -12152 49695 -12088
rect 49695 -12152 49759 -12088
rect 49759 -12152 49845 -12088
rect 49609 -12238 49845 -12152
rect 49609 -12408 49845 -12322
rect 49609 -12472 49695 -12408
rect 49695 -12472 49759 -12408
rect 49759 -12472 49845 -12408
rect 49609 -12558 49845 -12472
rect 49609 -12728 49845 -12642
rect 49609 -12792 49695 -12728
rect 49695 -12792 49759 -12728
rect 49759 -12792 49845 -12728
rect 49609 -12878 49845 -12792
rect 49609 -13048 49845 -12962
rect 49609 -13112 49695 -13048
rect 49695 -13112 49759 -13048
rect 49759 -13112 49845 -13048
rect 49609 -13198 49845 -13112
rect 49609 -13368 49845 -13282
rect 49609 -13432 49695 -13368
rect 49695 -13432 49759 -13368
rect 49759 -13432 49845 -13368
rect 49609 -13518 49845 -13432
rect 49609 -13688 49845 -13602
rect 49609 -13752 49695 -13688
rect 49695 -13752 49759 -13688
rect 49759 -13752 49845 -13688
rect 49609 -13838 49845 -13752
rect 49609 -14008 49845 -13922
rect 49609 -14072 49695 -14008
rect 49695 -14072 49759 -14008
rect 49759 -14072 49845 -14008
rect 49609 -14158 49845 -14072
rect 49609 -14328 49845 -14242
rect 49609 -14392 49695 -14328
rect 49695 -14392 49759 -14328
rect 49759 -14392 49845 -14328
rect 49609 -14478 49845 -14392
rect 49609 -14648 49845 -14562
rect 49609 -14712 49695 -14648
rect 49695 -14712 49759 -14648
rect 49759 -14712 49845 -14648
rect 49609 -14798 49845 -14712
rect 49609 -14968 49845 -14882
rect 49609 -15032 49695 -14968
rect 49695 -15032 49759 -14968
rect 49759 -15032 49845 -14968
rect 49609 -15118 49845 -15032
rect 49609 -15288 49845 -15202
rect 49609 -15352 49695 -15288
rect 49695 -15352 49759 -15288
rect 49759 -15352 49845 -15288
rect 49609 -15438 49845 -15352
rect 49609 -15608 49845 -15522
rect 49609 -15672 49695 -15608
rect 49695 -15672 49759 -15608
rect 49759 -15672 49845 -15608
rect 49609 -15758 49845 -15672
rect 49609 -15928 49845 -15842
rect 49609 -15992 49695 -15928
rect 49695 -15992 49759 -15928
rect 49759 -15992 49845 -15928
rect 49609 -16078 49845 -15992
rect 49609 -16248 49845 -16162
rect 49609 -16312 49695 -16248
rect 49695 -16312 49759 -16248
rect 49759 -16312 49845 -16248
rect 49609 -16398 49845 -16312
rect 49609 -16568 49845 -16482
rect 49609 -16632 49695 -16568
rect 49695 -16632 49759 -16568
rect 49759 -16632 49845 -16568
rect 49609 -16718 49845 -16632
rect 49609 -16888 49845 -16802
rect 49609 -16952 49695 -16888
rect 49695 -16952 49759 -16888
rect 49759 -16952 49845 -16888
rect 49609 -17038 49845 -16952
rect 49609 -17208 49845 -17122
rect 49609 -17272 49695 -17208
rect 49695 -17272 49759 -17208
rect 49759 -17272 49845 -17208
rect 49609 -17358 49845 -17272
rect 49609 -17528 49845 -17442
rect 49609 -17592 49695 -17528
rect 49695 -17592 49759 -17528
rect 49759 -17592 49845 -17528
rect 49609 -17678 49845 -17592
rect 49609 -17848 49845 -17762
rect 49609 -17912 49695 -17848
rect 49695 -17912 49759 -17848
rect 49759 -17912 49845 -17848
rect 49609 -17998 49845 -17912
rect 49609 -18168 49845 -18082
rect 49609 -18232 49695 -18168
rect 49695 -18232 49759 -18168
rect 49759 -18232 49845 -18168
rect 49609 -18318 49845 -18232
rect 42155 -18552 42241 -18488
rect 42241 -18552 42305 -18488
rect 42305 -18552 42391 -18488
rect 42155 -18638 42391 -18552
rect 49609 -18488 49845 -18402
rect 49609 -18552 49695 -18488
rect 49695 -18552 49759 -18488
rect 49759 -18552 49845 -18488
rect 42522 -18698 42758 -18612
rect 42522 -18762 42608 -18698
rect 42608 -18762 42672 -18698
rect 42672 -18762 42758 -18698
rect 42522 -18848 42758 -18762
rect 42842 -18698 43078 -18612
rect 42842 -18762 42928 -18698
rect 42928 -18762 42992 -18698
rect 42992 -18762 43078 -18698
rect 42842 -18848 43078 -18762
rect 43162 -18698 43398 -18612
rect 43162 -18762 43248 -18698
rect 43248 -18762 43312 -18698
rect 43312 -18762 43398 -18698
rect 43162 -18848 43398 -18762
rect 43482 -18698 43718 -18612
rect 43482 -18762 43568 -18698
rect 43568 -18762 43632 -18698
rect 43632 -18762 43718 -18698
rect 43482 -18848 43718 -18762
rect 43802 -18698 44038 -18612
rect 43802 -18762 43888 -18698
rect 43888 -18762 43952 -18698
rect 43952 -18762 44038 -18698
rect 43802 -18848 44038 -18762
rect 44122 -18698 44358 -18612
rect 44122 -18762 44208 -18698
rect 44208 -18762 44272 -18698
rect 44272 -18762 44358 -18698
rect 44122 -18848 44358 -18762
rect 44442 -18698 44678 -18612
rect 44442 -18762 44528 -18698
rect 44528 -18762 44592 -18698
rect 44592 -18762 44678 -18698
rect 44442 -18848 44678 -18762
rect 44762 -18698 44998 -18612
rect 44762 -18762 44848 -18698
rect 44848 -18762 44912 -18698
rect 44912 -18762 44998 -18698
rect 44762 -18848 44998 -18762
rect 45082 -18698 45318 -18612
rect 45082 -18762 45168 -18698
rect 45168 -18762 45232 -18698
rect 45232 -18762 45318 -18698
rect 45082 -18848 45318 -18762
rect 45402 -18698 45638 -18612
rect 45402 -18762 45488 -18698
rect 45488 -18762 45552 -18698
rect 45552 -18762 45638 -18698
rect 45402 -18848 45638 -18762
rect 45722 -18698 45958 -18612
rect 45722 -18762 45808 -18698
rect 45808 -18762 45872 -18698
rect 45872 -18762 45958 -18698
rect 45722 -18848 45958 -18762
rect 46042 -18698 46278 -18612
rect 46042 -18762 46128 -18698
rect 46128 -18762 46192 -18698
rect 46192 -18762 46278 -18698
rect 46042 -18848 46278 -18762
rect 46362 -18698 46598 -18612
rect 46362 -18762 46448 -18698
rect 46448 -18762 46512 -18698
rect 46512 -18762 46598 -18698
rect 46362 -18848 46598 -18762
rect 46682 -18698 46918 -18612
rect 46682 -18762 46768 -18698
rect 46768 -18762 46832 -18698
rect 46832 -18762 46918 -18698
rect 46682 -18848 46918 -18762
rect 47002 -18698 47238 -18612
rect 47002 -18762 47088 -18698
rect 47088 -18762 47152 -18698
rect 47152 -18762 47238 -18698
rect 47002 -18848 47238 -18762
rect 47322 -18698 47558 -18612
rect 47322 -18762 47408 -18698
rect 47408 -18762 47472 -18698
rect 47472 -18762 47558 -18698
rect 47322 -18848 47558 -18762
rect 47642 -18698 47878 -18612
rect 47642 -18762 47728 -18698
rect 47728 -18762 47792 -18698
rect 47792 -18762 47878 -18698
rect 47642 -18848 47878 -18762
rect 47962 -18698 48198 -18612
rect 47962 -18762 48048 -18698
rect 48048 -18762 48112 -18698
rect 48112 -18762 48198 -18698
rect 47962 -18848 48198 -18762
rect 48282 -18698 48518 -18612
rect 48282 -18762 48368 -18698
rect 48368 -18762 48432 -18698
rect 48432 -18762 48518 -18698
rect 48282 -18848 48518 -18762
rect 48602 -18698 48838 -18612
rect 48602 -18762 48688 -18698
rect 48688 -18762 48752 -18698
rect 48752 -18762 48838 -18698
rect 48602 -18848 48838 -18762
rect 48922 -18698 49158 -18612
rect 48922 -18762 49008 -18698
rect 49008 -18762 49072 -18698
rect 49072 -18762 49158 -18698
rect 48922 -18848 49158 -18762
rect 49242 -18698 49478 -18612
rect 49609 -18638 49845 -18552
rect 49242 -18762 49328 -18698
rect 49328 -18762 49392 -18698
rect 49392 -18762 49478 -18698
rect 49242 -18848 49478 -18762
<< mimcap2 >>
rect 21380 -5560 21820 -5540
rect 21380 -9060 21400 -5560
rect 21800 -9060 21820 -5560
rect 21380 -9080 21820 -9060
<< mimcap2contact >>
rect 21400 -9060 21800 -5560
<< metal5 >>
rect 3000 3360 51000 3400
rect 3000 3060 20080 3360
rect 20480 3060 51000 3360
rect 3000 3000 51000 3060
rect 3000 1760 51000 1800
rect 3000 1600 20020 1760
rect 3000 1000 11400 1600
rect 12200 1000 15800 1600
rect 16600 1460 20020 1600
rect 20260 1500 51000 1760
rect 20260 1460 33200 1500
rect 16600 1000 33200 1460
rect 34500 1000 51000 1500
rect 3000 800 51000 1000
rect 3000 360 51000 400
rect 3000 -560 14940 360
rect 15200 -560 51000 360
rect 3000 -600 51000 -560
rect 11200 -1200 12200 -600
rect 13000 -1200 14000 -600
rect 20340 -1680 20660 -600
rect 20340 -2200 20380 -1680
rect 20620 -2200 20660 -1680
rect 20340 -2240 20660 -2200
rect 21340 -5560 21860 -5500
rect 21340 -9060 21400 -5560
rect 21800 -9060 21860 -5560
rect 21340 -9260 21860 -9060
rect 21340 -9500 21380 -9260
rect 21820 -9500 21860 -9260
rect 21340 -9540 21860 -9500
rect 6000 -11156 14000 -11000
rect 6000 -11362 6522 -11156
rect 6000 -11598 6152 -11362
rect 6388 -11392 6522 -11362
rect 6758 -11392 6842 -11156
rect 7078 -11392 7162 -11156
rect 7398 -11392 7482 -11156
rect 7718 -11392 7802 -11156
rect 8038 -11392 8122 -11156
rect 8358 -11392 8442 -11156
rect 8678 -11392 8762 -11156
rect 8998 -11392 9082 -11156
rect 9318 -11392 9402 -11156
rect 9638 -11392 9722 -11156
rect 9958 -11392 10042 -11156
rect 10278 -11392 10362 -11156
rect 10598 -11392 10682 -11156
rect 10918 -11392 11002 -11156
rect 11238 -11392 11322 -11156
rect 11558 -11392 11642 -11156
rect 11878 -11392 11962 -11156
rect 12198 -11392 12282 -11156
rect 12518 -11392 12602 -11156
rect 12838 -11392 12922 -11156
rect 13158 -11392 13242 -11156
rect 13478 -11362 14000 -11156
rect 13478 -11392 13618 -11362
rect 6388 -11598 13618 -11392
rect 13854 -11598 14000 -11362
rect 6000 -11682 14000 -11598
rect 6000 -11918 6152 -11682
rect 6388 -11918 13618 -11682
rect 13854 -11918 14000 -11682
rect 6000 -12002 14000 -11918
rect 6000 -12238 6152 -12002
rect 6388 -12238 13618 -12002
rect 13854 -12238 14000 -12002
rect 6000 -12322 14000 -12238
rect 6000 -12558 6152 -12322
rect 6388 -12558 13618 -12322
rect 13854 -12558 14000 -12322
rect 6000 -12642 14000 -12558
rect 6000 -12878 6152 -12642
rect 6388 -12878 13618 -12642
rect 13854 -12878 14000 -12642
rect 6000 -12962 14000 -12878
rect 6000 -13198 6152 -12962
rect 6388 -13198 13618 -12962
rect 13854 -13198 14000 -12962
rect 6000 -13282 14000 -13198
rect 6000 -13518 6152 -13282
rect 6388 -13518 13618 -13282
rect 13854 -13518 14000 -13282
rect 6000 -13602 14000 -13518
rect 6000 -13838 6152 -13602
rect 6388 -13838 13618 -13602
rect 13854 -13838 14000 -13602
rect 6000 -13922 14000 -13838
rect 6000 -14158 6152 -13922
rect 6388 -14158 13618 -13922
rect 13854 -14158 14000 -13922
rect 6000 -14242 14000 -14158
rect 6000 -14478 6152 -14242
rect 6388 -14478 13618 -14242
rect 13854 -14478 14000 -14242
rect 6000 -14562 14000 -14478
rect 6000 -14798 6152 -14562
rect 6388 -14798 13618 -14562
rect 13854 -14798 14000 -14562
rect 6000 -14882 14000 -14798
rect 6000 -15118 6152 -14882
rect 6388 -15118 13618 -14882
rect 13854 -15118 14000 -14882
rect 6000 -15202 14000 -15118
rect 6000 -15438 6152 -15202
rect 6388 -15438 13618 -15202
rect 13854 -15438 14000 -15202
rect 6000 -15522 14000 -15438
rect 6000 -15758 6152 -15522
rect 6388 -15758 13618 -15522
rect 13854 -15758 14000 -15522
rect 6000 -15842 14000 -15758
rect 6000 -16078 6152 -15842
rect 6388 -16078 13618 -15842
rect 13854 -16078 14000 -15842
rect 6000 -16162 14000 -16078
rect 6000 -16398 6152 -16162
rect 6388 -16398 13618 -16162
rect 13854 -16398 14000 -16162
rect 6000 -16482 14000 -16398
rect 6000 -16718 6152 -16482
rect 6388 -16718 13618 -16482
rect 13854 -16718 14000 -16482
rect 6000 -16802 14000 -16718
rect 6000 -17038 6152 -16802
rect 6388 -17038 13618 -16802
rect 13854 -17038 14000 -16802
rect 6000 -17122 14000 -17038
rect 6000 -17358 6152 -17122
rect 6388 -17358 13618 -17122
rect 13854 -17358 14000 -17122
rect 6000 -17442 14000 -17358
rect 6000 -17678 6152 -17442
rect 6388 -17678 13618 -17442
rect 13854 -17678 14000 -17442
rect 6000 -17762 14000 -17678
rect 6000 -17998 6152 -17762
rect 6388 -17998 13618 -17762
rect 13854 -17998 14000 -17762
rect 6000 -18082 14000 -17998
rect 6000 -18318 6152 -18082
rect 6388 -18318 13618 -18082
rect 13854 -18318 14000 -18082
rect 6000 -18402 14000 -18318
rect 6000 -18638 6152 -18402
rect 6388 -18612 13618 -18402
rect 6388 -18638 6522 -18612
rect 6000 -18848 6522 -18638
rect 6758 -18848 6842 -18612
rect 7078 -18848 7162 -18612
rect 7398 -18848 7482 -18612
rect 7718 -18848 7802 -18612
rect 8038 -18848 8122 -18612
rect 8358 -18848 8442 -18612
rect 8678 -18848 8762 -18612
rect 8998 -18848 9082 -18612
rect 9318 -18848 9402 -18612
rect 9638 -18848 9722 -18612
rect 9958 -18848 10042 -18612
rect 10278 -18848 10362 -18612
rect 10598 -18848 10682 -18612
rect 10918 -18848 11002 -18612
rect 11238 -18848 11322 -18612
rect 11558 -18848 11642 -18612
rect 11878 -18848 11962 -18612
rect 12198 -18848 12282 -18612
rect 12518 -18848 12602 -18612
rect 12838 -18848 12922 -18612
rect 13158 -18848 13242 -18612
rect 13478 -18638 13618 -18612
rect 13854 -18638 14000 -18402
rect 13478 -18848 14000 -18638
rect 6000 -19000 14000 -18848
rect 18000 -11156 26000 -11000
rect 18000 -11362 18522 -11156
rect 18000 -11598 18152 -11362
rect 18388 -11392 18522 -11362
rect 18758 -11392 18842 -11156
rect 19078 -11392 19162 -11156
rect 19398 -11392 19482 -11156
rect 19718 -11392 19802 -11156
rect 20038 -11392 20122 -11156
rect 20358 -11392 20442 -11156
rect 20678 -11392 20762 -11156
rect 20998 -11392 21082 -11156
rect 21318 -11392 21402 -11156
rect 21638 -11392 21722 -11156
rect 21958 -11392 22042 -11156
rect 22278 -11392 22362 -11156
rect 22598 -11392 22682 -11156
rect 22918 -11392 23002 -11156
rect 23238 -11392 23322 -11156
rect 23558 -11392 23642 -11156
rect 23878 -11392 23962 -11156
rect 24198 -11392 24282 -11156
rect 24518 -11392 24602 -11156
rect 24838 -11392 24922 -11156
rect 25158 -11392 25242 -11156
rect 25478 -11362 26000 -11156
rect 25478 -11392 25618 -11362
rect 18388 -11598 25618 -11392
rect 25854 -11598 26000 -11362
rect 18000 -11682 26000 -11598
rect 18000 -11918 18152 -11682
rect 18388 -11918 25618 -11682
rect 25854 -11918 26000 -11682
rect 18000 -12002 26000 -11918
rect 18000 -12238 18152 -12002
rect 18388 -12238 25618 -12002
rect 25854 -12238 26000 -12002
rect 18000 -12322 26000 -12238
rect 18000 -12558 18152 -12322
rect 18388 -12558 25618 -12322
rect 25854 -12558 26000 -12322
rect 18000 -12642 26000 -12558
rect 18000 -12878 18152 -12642
rect 18388 -12878 25618 -12642
rect 25854 -12878 26000 -12642
rect 18000 -12962 26000 -12878
rect 18000 -13198 18152 -12962
rect 18388 -13198 25618 -12962
rect 25854 -13198 26000 -12962
rect 18000 -13282 26000 -13198
rect 18000 -13518 18152 -13282
rect 18388 -13518 25618 -13282
rect 25854 -13518 26000 -13282
rect 18000 -13602 26000 -13518
rect 18000 -13838 18152 -13602
rect 18388 -13838 25618 -13602
rect 25854 -13838 26000 -13602
rect 18000 -13922 26000 -13838
rect 18000 -14158 18152 -13922
rect 18388 -14158 25618 -13922
rect 25854 -14158 26000 -13922
rect 18000 -14242 26000 -14158
rect 18000 -14478 18152 -14242
rect 18388 -14478 25618 -14242
rect 25854 -14478 26000 -14242
rect 18000 -14562 26000 -14478
rect 18000 -14798 18152 -14562
rect 18388 -14798 25618 -14562
rect 25854 -14798 26000 -14562
rect 18000 -14882 26000 -14798
rect 18000 -15118 18152 -14882
rect 18388 -15118 25618 -14882
rect 25854 -15118 26000 -14882
rect 18000 -15202 26000 -15118
rect 18000 -15438 18152 -15202
rect 18388 -15438 25618 -15202
rect 25854 -15438 26000 -15202
rect 18000 -15522 26000 -15438
rect 18000 -15758 18152 -15522
rect 18388 -15758 25618 -15522
rect 25854 -15758 26000 -15522
rect 18000 -15842 26000 -15758
rect 18000 -16078 18152 -15842
rect 18388 -16078 25618 -15842
rect 25854 -16078 26000 -15842
rect 18000 -16162 26000 -16078
rect 18000 -16398 18152 -16162
rect 18388 -16398 25618 -16162
rect 25854 -16398 26000 -16162
rect 18000 -16482 26000 -16398
rect 18000 -16718 18152 -16482
rect 18388 -16718 25618 -16482
rect 25854 -16718 26000 -16482
rect 18000 -16802 26000 -16718
rect 18000 -17038 18152 -16802
rect 18388 -17038 25618 -16802
rect 25854 -17038 26000 -16802
rect 18000 -17122 26000 -17038
rect 18000 -17358 18152 -17122
rect 18388 -17358 25618 -17122
rect 25854 -17358 26000 -17122
rect 18000 -17442 26000 -17358
rect 18000 -17678 18152 -17442
rect 18388 -17678 25618 -17442
rect 25854 -17678 26000 -17442
rect 18000 -17762 26000 -17678
rect 18000 -17998 18152 -17762
rect 18388 -17998 25618 -17762
rect 25854 -17998 26000 -17762
rect 18000 -18082 26000 -17998
rect 18000 -18318 18152 -18082
rect 18388 -18318 25618 -18082
rect 25854 -18318 26000 -18082
rect 18000 -18402 26000 -18318
rect 18000 -18638 18152 -18402
rect 18388 -18612 25618 -18402
rect 18388 -18638 18522 -18612
rect 18000 -18848 18522 -18638
rect 18758 -18848 18842 -18612
rect 19078 -18848 19162 -18612
rect 19398 -18848 19482 -18612
rect 19718 -18848 19802 -18612
rect 20038 -18848 20122 -18612
rect 20358 -18848 20442 -18612
rect 20678 -18848 20762 -18612
rect 20998 -18848 21082 -18612
rect 21318 -18848 21402 -18612
rect 21638 -18848 21722 -18612
rect 21958 -18848 22042 -18612
rect 22278 -18848 22362 -18612
rect 22598 -18848 22682 -18612
rect 22918 -18848 23002 -18612
rect 23238 -18848 23322 -18612
rect 23558 -18848 23642 -18612
rect 23878 -18848 23962 -18612
rect 24198 -18848 24282 -18612
rect 24518 -18848 24602 -18612
rect 24838 -18848 24922 -18612
rect 25158 -18848 25242 -18612
rect 25478 -18638 25618 -18612
rect 25854 -18638 26000 -18402
rect 25478 -18848 26000 -18638
rect 18000 -19000 26000 -18848
rect 30000 -11156 38000 -11000
rect 30000 -11362 30522 -11156
rect 30000 -11598 30152 -11362
rect 30388 -11392 30522 -11362
rect 30758 -11392 30842 -11156
rect 31078 -11392 31162 -11156
rect 31398 -11392 31482 -11156
rect 31718 -11392 31802 -11156
rect 32038 -11392 32122 -11156
rect 32358 -11392 32442 -11156
rect 32678 -11392 32762 -11156
rect 32998 -11392 33082 -11156
rect 33318 -11392 33402 -11156
rect 33638 -11392 33722 -11156
rect 33958 -11392 34042 -11156
rect 34278 -11392 34362 -11156
rect 34598 -11392 34682 -11156
rect 34918 -11392 35002 -11156
rect 35238 -11392 35322 -11156
rect 35558 -11392 35642 -11156
rect 35878 -11392 35962 -11156
rect 36198 -11392 36282 -11156
rect 36518 -11392 36602 -11156
rect 36838 -11392 36922 -11156
rect 37158 -11392 37242 -11156
rect 37478 -11362 38000 -11156
rect 37478 -11392 37618 -11362
rect 30388 -11598 37618 -11392
rect 37854 -11598 38000 -11362
rect 30000 -11682 38000 -11598
rect 30000 -11918 30152 -11682
rect 30388 -11918 37618 -11682
rect 37854 -11918 38000 -11682
rect 30000 -12002 38000 -11918
rect 30000 -12238 30152 -12002
rect 30388 -12238 37618 -12002
rect 37854 -12238 38000 -12002
rect 30000 -12322 38000 -12238
rect 30000 -12558 30152 -12322
rect 30388 -12558 37618 -12322
rect 37854 -12558 38000 -12322
rect 30000 -12642 38000 -12558
rect 30000 -12878 30152 -12642
rect 30388 -12878 37618 -12642
rect 37854 -12878 38000 -12642
rect 30000 -12962 38000 -12878
rect 30000 -13198 30152 -12962
rect 30388 -13198 37618 -12962
rect 37854 -13198 38000 -12962
rect 30000 -13282 38000 -13198
rect 30000 -13518 30152 -13282
rect 30388 -13518 37618 -13282
rect 37854 -13518 38000 -13282
rect 30000 -13602 38000 -13518
rect 30000 -13838 30152 -13602
rect 30388 -13838 37618 -13602
rect 37854 -13838 38000 -13602
rect 30000 -13922 38000 -13838
rect 30000 -14158 30152 -13922
rect 30388 -14158 37618 -13922
rect 37854 -14158 38000 -13922
rect 30000 -14242 38000 -14158
rect 30000 -14478 30152 -14242
rect 30388 -14478 37618 -14242
rect 37854 -14478 38000 -14242
rect 30000 -14562 38000 -14478
rect 30000 -14798 30152 -14562
rect 30388 -14798 37618 -14562
rect 37854 -14798 38000 -14562
rect 30000 -14882 38000 -14798
rect 30000 -15118 30152 -14882
rect 30388 -15118 37618 -14882
rect 37854 -15118 38000 -14882
rect 30000 -15202 38000 -15118
rect 30000 -15438 30152 -15202
rect 30388 -15438 37618 -15202
rect 37854 -15438 38000 -15202
rect 30000 -15522 38000 -15438
rect 30000 -15758 30152 -15522
rect 30388 -15758 37618 -15522
rect 37854 -15758 38000 -15522
rect 30000 -15842 38000 -15758
rect 30000 -16078 30152 -15842
rect 30388 -16078 37618 -15842
rect 37854 -16078 38000 -15842
rect 30000 -16162 38000 -16078
rect 30000 -16398 30152 -16162
rect 30388 -16398 37618 -16162
rect 37854 -16398 38000 -16162
rect 30000 -16482 38000 -16398
rect 30000 -16718 30152 -16482
rect 30388 -16718 37618 -16482
rect 37854 -16718 38000 -16482
rect 30000 -16802 38000 -16718
rect 30000 -17038 30152 -16802
rect 30388 -17038 37618 -16802
rect 37854 -17038 38000 -16802
rect 30000 -17122 38000 -17038
rect 30000 -17358 30152 -17122
rect 30388 -17358 37618 -17122
rect 37854 -17358 38000 -17122
rect 30000 -17442 38000 -17358
rect 30000 -17678 30152 -17442
rect 30388 -17678 37618 -17442
rect 37854 -17678 38000 -17442
rect 30000 -17762 38000 -17678
rect 30000 -17998 30152 -17762
rect 30388 -17998 37618 -17762
rect 37854 -17998 38000 -17762
rect 30000 -18082 38000 -17998
rect 30000 -18318 30152 -18082
rect 30388 -18318 37618 -18082
rect 37854 -18318 38000 -18082
rect 30000 -18402 38000 -18318
rect 30000 -18638 30152 -18402
rect 30388 -18612 37618 -18402
rect 30388 -18638 30522 -18612
rect 30000 -18848 30522 -18638
rect 30758 -18848 30842 -18612
rect 31078 -18848 31162 -18612
rect 31398 -18848 31482 -18612
rect 31718 -18848 31802 -18612
rect 32038 -18848 32122 -18612
rect 32358 -18848 32442 -18612
rect 32678 -18848 32762 -18612
rect 32998 -18848 33082 -18612
rect 33318 -18848 33402 -18612
rect 33638 -18848 33722 -18612
rect 33958 -18848 34042 -18612
rect 34278 -18848 34362 -18612
rect 34598 -18848 34682 -18612
rect 34918 -18848 35002 -18612
rect 35238 -18848 35322 -18612
rect 35558 -18848 35642 -18612
rect 35878 -18848 35962 -18612
rect 36198 -18848 36282 -18612
rect 36518 -18848 36602 -18612
rect 36838 -18848 36922 -18612
rect 37158 -18848 37242 -18612
rect 37478 -18638 37618 -18612
rect 37854 -18638 38000 -18402
rect 37478 -18848 38000 -18638
rect 30000 -19000 38000 -18848
rect 42000 -11156 50000 -11000
rect 42000 -11362 42522 -11156
rect 42000 -11598 42155 -11362
rect 42391 -11392 42522 -11362
rect 42758 -11392 42842 -11156
rect 43078 -11392 43162 -11156
rect 43398 -11392 43482 -11156
rect 43718 -11392 43802 -11156
rect 44038 -11392 44122 -11156
rect 44358 -11392 44442 -11156
rect 44678 -11392 44762 -11156
rect 44998 -11392 45082 -11156
rect 45318 -11392 45402 -11156
rect 45638 -11392 45722 -11156
rect 45958 -11392 46042 -11156
rect 46278 -11392 46362 -11156
rect 46598 -11392 46682 -11156
rect 46918 -11392 47002 -11156
rect 47238 -11392 47322 -11156
rect 47558 -11392 47642 -11156
rect 47878 -11392 47962 -11156
rect 48198 -11392 48282 -11156
rect 48518 -11392 48602 -11156
rect 48838 -11392 48922 -11156
rect 49158 -11392 49242 -11156
rect 49478 -11362 50000 -11156
rect 49478 -11392 49609 -11362
rect 42391 -11598 49609 -11392
rect 49845 -11598 50000 -11362
rect 42000 -11682 50000 -11598
rect 42000 -11918 42155 -11682
rect 42391 -11918 49609 -11682
rect 49845 -11918 50000 -11682
rect 42000 -12002 50000 -11918
rect 42000 -12238 42155 -12002
rect 42391 -12238 49609 -12002
rect 49845 -12238 50000 -12002
rect 42000 -12322 50000 -12238
rect 42000 -12558 42155 -12322
rect 42391 -12558 49609 -12322
rect 49845 -12558 50000 -12322
rect 42000 -12642 50000 -12558
rect 42000 -12878 42155 -12642
rect 42391 -12878 49609 -12642
rect 49845 -12878 50000 -12642
rect 42000 -12962 50000 -12878
rect 42000 -13198 42155 -12962
rect 42391 -13198 49609 -12962
rect 49845 -13198 50000 -12962
rect 42000 -13282 50000 -13198
rect 42000 -13518 42155 -13282
rect 42391 -13518 49609 -13282
rect 49845 -13518 50000 -13282
rect 42000 -13602 50000 -13518
rect 42000 -13838 42155 -13602
rect 42391 -13838 49609 -13602
rect 49845 -13838 50000 -13602
rect 42000 -13922 50000 -13838
rect 42000 -14158 42155 -13922
rect 42391 -14158 49609 -13922
rect 49845 -14158 50000 -13922
rect 42000 -14242 50000 -14158
rect 42000 -14478 42155 -14242
rect 42391 -14478 49609 -14242
rect 49845 -14478 50000 -14242
rect 42000 -14562 50000 -14478
rect 42000 -14798 42155 -14562
rect 42391 -14798 49609 -14562
rect 49845 -14798 50000 -14562
rect 42000 -14882 50000 -14798
rect 42000 -15118 42155 -14882
rect 42391 -15118 49609 -14882
rect 49845 -15118 50000 -14882
rect 42000 -15202 50000 -15118
rect 42000 -15438 42155 -15202
rect 42391 -15438 49609 -15202
rect 49845 -15438 50000 -15202
rect 42000 -15522 50000 -15438
rect 42000 -15758 42155 -15522
rect 42391 -15758 49609 -15522
rect 49845 -15758 50000 -15522
rect 42000 -15842 50000 -15758
rect 42000 -16078 42155 -15842
rect 42391 -16078 49609 -15842
rect 49845 -16078 50000 -15842
rect 42000 -16162 50000 -16078
rect 42000 -16398 42155 -16162
rect 42391 -16398 49609 -16162
rect 49845 -16398 50000 -16162
rect 42000 -16482 50000 -16398
rect 42000 -16718 42155 -16482
rect 42391 -16718 49609 -16482
rect 49845 -16718 50000 -16482
rect 42000 -16802 50000 -16718
rect 42000 -17038 42155 -16802
rect 42391 -17038 49609 -16802
rect 49845 -17038 50000 -16802
rect 42000 -17122 50000 -17038
rect 42000 -17358 42155 -17122
rect 42391 -17358 49609 -17122
rect 49845 -17358 50000 -17122
rect 42000 -17442 50000 -17358
rect 42000 -17678 42155 -17442
rect 42391 -17678 49609 -17442
rect 49845 -17678 50000 -17442
rect 42000 -17762 50000 -17678
rect 42000 -17998 42155 -17762
rect 42391 -17998 49609 -17762
rect 49845 -17998 50000 -17762
rect 42000 -18082 50000 -17998
rect 42000 -18318 42155 -18082
rect 42391 -18318 49609 -18082
rect 49845 -18318 50000 -18082
rect 42000 -18402 50000 -18318
rect 42000 -18638 42155 -18402
rect 42391 -18612 49609 -18402
rect 42391 -18638 42522 -18612
rect 42000 -18848 42522 -18638
rect 42758 -18848 42842 -18612
rect 43078 -18848 43162 -18612
rect 43398 -18848 43482 -18612
rect 43718 -18848 43802 -18612
rect 44038 -18848 44122 -18612
rect 44358 -18848 44442 -18612
rect 44678 -18848 44762 -18612
rect 44998 -18848 45082 -18612
rect 45318 -18848 45402 -18612
rect 45638 -18848 45722 -18612
rect 45958 -18848 46042 -18612
rect 46278 -18848 46362 -18612
rect 46598 -18848 46682 -18612
rect 46918 -18848 47002 -18612
rect 47238 -18848 47322 -18612
rect 47558 -18848 47642 -18612
rect 47878 -18848 47962 -18612
rect 48198 -18848 48282 -18612
rect 48518 -18848 48602 -18612
rect 48838 -18848 48922 -18612
rect 49158 -18848 49242 -18612
rect 49478 -18638 49609 -18612
rect 49845 -18638 50000 -18402
rect 49478 -18848 50000 -18638
rect 42000 -19000 50000 -18848
<< glass >>
rect 6600 -18400 13400 -11600
rect 18600 -18400 25400 -11600
rect 30600 -18400 37400 -11600
rect 42600 -18400 49400 -11600
<< fillblock >>
rect 21220 -3180 22140 -2260
<< comment >>
rect 1800 -19000 2000 -10600
<< res0p35 >>
rect 20503 3171 20907 3245
use QCS_unit1_flat_dnw  QCS_unit1_flat_dnw_0
timestamp 1668748373
transform 1 0 19080 0 1 -3120
box 1520 -680 3680 1480
use cellselect  cellselect_1
timestamp 1671823942
transform 0 1 14297 -1 0 -72
box 96 -97 1708 667
use cmota_gb_rp_gp  cmota_gb_rp_gp_1
timestamp 1671855392
transform 1 0 18200 0 -1 -9000
box -7000 -7800 2802 600
use sky130_fd_pr__res_xhigh_po_0p35_EP3CBP  sky130_fd_pr__res_xhigh_po_0p35_EP3CBP_0
timestamp 1671678338
transform 1 0 21304 0 -1 -4668
box -284 -748 284 748
<< labels >>
rlabel metal5 3000 3000 3440 3400 1 VMID
rlabel metal5 3000 800 3440 1800 1 VLO
rlabel metal5 3000 -600 3440 400 1 VHI
rlabel metal4 3000 1860 3440 2160 1 VTW
rlabel metal4 3000 3460 3440 3740 1 ROWSEL
rlabel metal4 3000 2660 3440 2960 1 VREF
rlabel metal3 21001 -2570 21044 -2510 1 TW
rlabel metal3 14200 -21800 15000 -21260 1 COLSEL
<< end >>
