* NGSPICE file created from twcon.ext - technology: sky130A

X0 tcap_50f_0/a_173_157# tcap_50f_0/C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=7.85e+06u
X1 tcap_50f_0/a_173_157# C100 VLO VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X2 tcap_50f_0/C tcap_50f_0/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=7.85e+06u
X3 tcap_50f_3/a_173_157# tcap_50f_3/C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=7.85e+06u
X4 tcap_50f_3/a_173_157# C100 VLO VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X5 tcap_50f_3/C tcap_50f_3/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=7.85e+06u
X6 tcap_50f_2/a_173_157# tcap_50f_2/C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=7.85e+06u
X7 tcap_50f_2/a_173_157# C50 VLO VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X8 tcap_50f_2/C tcap_50f_2/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=7.85e+06u
X9 tcap_100f_0/a_173_157# tcap_50f_0/C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=1.57e+07u
X10 tcap_100f_0/a_173_157# C50 VLO VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X11 tcap_50f_0/C tcap_100f_0/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=1.57e+07u
X12 tcap_100f_2/a_173_157# tcap_50f_2/C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=1.57e+07u
X13 tcap_100f_2/a_173_157# C100 VLO VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X14 tcap_50f_2/C tcap_100f_2/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=1.57e+07u
X15 tcap_100f_3/a_173_157# tcap_50f_3/C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=1.57e+07u
X16 tcap_100f_3/a_173_157# C50 VLO VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X17 tcap_50f_3/C tcap_100f_3/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=1.57e+07u
X18 twcon_tdly_0/sky130_fd_sc_hs__inv_1_0/Y tcap_50f_2/C VLO sky130_fd_pr__res_xhigh_po_1p41 l=500000u
X19 twcon_tdly_1/sky130_fd_sc_hs__inv_1_0/Y tcap_50f_0/C VLO sky130_fd_pr__res_xhigh_po_1p41 l=500000u
X20 twcon_tdly_2/sky130_fd_sc_hs__inv_1_0/Y tcap_50f_3/C VLO sky130_fd_pr__res_xhigh_po_1p41 l=500000u
C0 tcap_100f_3/a_173_157# tcap_50f_3/C 5.51fF
C1 sky130_fd_sc_hs__fill_4_0/VPB VHI 2.43fF
C2 sky130_fd_sc_hs__mux2_1_1/S VHI 2.13fF
C3 tcap_50f_3/C tcap_50f_3/a_173_157# 2.93fF
C4 tcap_50f_2/a_173_157# tcap_50f_2/C 3.17fF
C5 tcap_50f_2/C tcap_100f_2/a_173_157# 5.34fF
C6 tcap_50f_0/C tcap_100f_0/a_173_157# 5.48fF
C7 VHI sky130_fd_sc_hs__inv_2_1/VPB 3.40fF
C8 tcap_50f_0/C tcap_50f_0/a_173_157# 2.92fF
Xsky130_fd_sc_hs__decap_8_0 VLO VHI sky130_fd_sc_hs__decap_8
Xsky130_fd_sc_hs__decap_8_2 VLO VHI sky130_fd_sc_hs__decap_8
Xsky130_fd_sc_hs__decap_8_3 VLO VHI sky130_fd_sc_hs__decap_8
Xsky130_fd_sc_hs__decap_8_4 VLO VHI sky130_fd_sc_hs__decap_8
Xsky130_fd_sc_hs__decap_8_5 VLO VHI sky130_fd_sc_hs__decap_8
Xsky130_fd_sc_hs__mux2_1_1 VHI VLO sky130_fd_sc_hs__mux2_1_1/X sky130_fd_sc_hs__mux2_1_1/S
+ twcon_tdly_1/Y twcon_tdly_2/Y sky130_fd_sc_hs__mux2_1
Xsky130_fd_sc_hs__decap_8_6 VLO VHI sky130_fd_sc_hs__decap_8
Xsky130_fd_sc_hs__decap_4_0 VLO VHI sky130_fd_sc_hs__decap_4
Xsky130_fd_sc_hs__decap_8_7 VLO VHI sky130_fd_sc_hs__decap_8
Xsky130_fd_sc_hs__fill_1_0 VLO sky130_fd_sc_hs__fill_4_0/VPB VHI VLO sky130_fd_sc_hs__fill_1
Xsky130_fd_sc_hs__fill_1_1 VLO sky130_fd_sc_hs__fill_4_0/VPB VHI VLO sky130_fd_sc_hs__fill_1
Xsky130_fd_sc_hs__tapmet1_2_0 VLO sky130_fd_sc_hs__inv_2_1/VPB VHI VLO sky130_fd_sc_hs__tapmet1_2
Xsky130_fd_sc_hs__tapmet1_2_1 VLO sky130_fd_sc_hs__inv_2_1/VPB VHI VLO sky130_fd_sc_hs__tapmet1_2
Xsky130_fd_sc_hs__tapmet1_2_2 VLO sky130_fd_sc_hs__fill_4_0/VPB VHI VLO sky130_fd_sc_hs__tapmet1_2
Xsky130_fd_sc_hs__sdfbbn_2_0 VHI VHI VLO VLO VLO VHI sky130_fd_sc_hs__inv_2_1/Y sky130_fd_sc_hs__sdfbbn_2_0/Q_N
+ VHI sky130_fd_sc_hs__mux2_1_1/X sky130_fd_sc_hs__sdfbbn_2
Xsky130_fd_sc_hs__fill_4_0 VLO sky130_fd_sc_hs__fill_4_0/VPB VHI VLO sky130_fd_sc_hs__fill_4
Xsky130_fd_sc_hs__sdfbbn_2_1 VHI VHI VLO VLO VLO sky130_fd_sc_hs__mux2_1_1/S twcon_tdly_0/Y
+ sky130_fd_sc_hs__mux2_1_1/S UPDN RSTB sky130_fd_sc_hs__sdfbbn_2
Xsky130_fd_sc_hs__nand2_4_0 VHI VLO GN sky130_fd_sc_hs__mux2_1_1/S VHI sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__fill_2_0 VLO sky130_fd_sc_hs__fill_4_0/VPB VHI VLO sky130_fd_sc_hs__fill_2
Xtwcon_tdly_0/sky130_fd_sc_hs__inv_1_0 VHI VLO twcon_tdly_0/sky130_fd_sc_hs__inv_1_0/Y
+ CLKIN sky130_fd_sc_hs__inv_1
Xtwcon_tdly_0/sky130_fd_sc_hs__nand2_1_2 VHI VLO tcap_50f_2/C twcon_tdly_0/Y CLKIN
+ sky130_fd_sc_hs__nand2_1
Xtwcon_tdly_0/sky130_fd_sc_hs__fill_8_0 VLO sky130_fd_sc_hs__inv_2_1/VPB VHI VLO sky130_fd_sc_hs__fill_8
Xtwcon_tdly_0/sky130_fd_sc_hs__fill_4_0 VLO sky130_fd_sc_hs__inv_2_1/VPB VHI VLO sky130_fd_sc_hs__fill_4
Xtwcon_tdly_1/sky130_fd_sc_hs__inv_1_0 VHI VLO twcon_tdly_1/sky130_fd_sc_hs__inv_1_0/Y
+ A0 sky130_fd_sc_hs__inv_1
Xtwcon_tdly_1/sky130_fd_sc_hs__nand2_1_2 VHI VLO tcap_50f_0/C twcon_tdly_1/Y A0 sky130_fd_sc_hs__nand2_1
Xtwcon_tdly_1/sky130_fd_sc_hs__fill_8_0 VLO sky130_fd_sc_hs__inv_2_1/VPB VHI VLO sky130_fd_sc_hs__fill_8
Xtwcon_tdly_1/sky130_fd_sc_hs__fill_4_0 VLO sky130_fd_sc_hs__inv_2_1/VPB VHI VLO sky130_fd_sc_hs__fill_4
Xtwcon_tdly_2/sky130_fd_sc_hs__inv_1_0 VHI VLO twcon_tdly_2/sky130_fd_sc_hs__inv_1_0/Y
+ A1 sky130_fd_sc_hs__inv_1
Xtwcon_tdly_2/sky130_fd_sc_hs__nand2_1_2 VHI VLO tcap_50f_3/C twcon_tdly_2/Y A1 sky130_fd_sc_hs__nand2_1
Xtwcon_tdly_2/sky130_fd_sc_hs__fill_8_0 VLO sky130_fd_sc_hs__fill_4_0/VPB VHI VLO
+ sky130_fd_sc_hs__fill_8
Xtwcon_tdly_2/sky130_fd_sc_hs__fill_4_0 VLO sky130_fd_sc_hs__fill_4_0/VPB VHI VLO
+ sky130_fd_sc_hs__fill_4
Xsky130_fd_sc_hs__nand2_4_3 VHI VLO GP UPDN VHI sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__inv_2_1 VHI VLO CLKIN sky130_fd_sc_hs__inv_2_1/Y sky130_fd_sc_hs__inv_2
Xsky130_fd_sc_hs__fill_diode_2_1 VLO sky130_fd_sc_hs__inv_2_1/VPB VHI VLO sky130_fd_sc_hs__fill_diode_2
Xsky130_fd_sc_hs__fill_diode_2_3 VLO sky130_fd_sc_hs__inv_2_1/VPB VHI VLO sky130_fd_sc_hs__fill_diode_2
C9 sky130_fd_sc_hs__fill_4_0/VPB VLO 10.38fF
C10 tcap_50f_3/C VLO 2.47fF
C11 tcap_50f_0/C VLO 2.67fF
C12 VHI VLO 20.82fF
C13 sky130_fd_sc_hs__inv_2_1/VPB VLO 17.09fF
C14 tcap_50f_2/C VLO 3.19fF
C15 tcap_100f_3/a_173_157# VLO 5.80fF $ **FLOATING
C16 tcap_100f_2/a_173_157# VLO 5.37fF $ **FLOATING
C17 C100 VLO 3.36fF $ **FLOATING
C18 tcap_100f_0/a_173_157# VLO 5.04fF $ **FLOATING
C19 sky130_fd_sc_hs__mux2_1_1/S VLO 2.20fF
C20 tcap_50f_2/a_173_157# VLO 4.49fF $ **FLOATING
C21 C50 VLO 2.80fF $ **FLOATING
C22 tcap_50f_3/a_173_157# VLO 3.62fF $ **FLOATING
C23 tcap_50f_0/a_173_157# VLO 3.59fF $ **FLOATING
