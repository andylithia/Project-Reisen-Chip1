** sch_path: /home/andylithia/openmpw/Project-Reisen-Chip1/xschem/idrive_hs_PEX.sch
**.subckt idrive_hs_PEX
V1 vmid GND 0.9
.save i(v1)
V2 vdd GND 1.8
.save i(v2)
V5 net2 GND 1.1
.save i(v5)
V6 net1 GND 0.7
.save i(v6)
V7 clkin GND PULSE(1.8 0 0 1n 1n 200n 400n)
.save i(v7)
x5 vdd vout_amp net4 net3 GND i_type_ota_model
XR4 net3 vout_amp GND sky130_fd_pr__res_xhigh_po_0p35 L=2 mult=1 m=1
XR5 vmid net3 GND sky130_fd_pr__res_xhigh_po_0p35 L=1 mult=1 m=1
x16 vdd vdd vdd vdd vdd GND GND GND vout GND swcap_array_PEX
x17 gp vdd gn GND UPDN clkin limn_pulse udclk ulim enclk llim vdd vdd vdd twcon_PEX
x1 vdd GND vrefp vrefn vout net5 gp gn isrc_PEX
I2 vdd vrefn 10u
x2 vdd ulim net2 vout vrefn vdd GND GND i_type_ota_gb_rp_gp_PEX
x3 vdd llim vout net1 vrefn vdd GND GND i_type_ota_gb_rp_gp_PEX
x4 vdd vout_buf vout_buf net6 vrefn vdd GND GND i_type_ota_gb_rp_gp_PEX
R2 net6 vout 10k m=1
**** begin user architecture code
.lib /home/andylithia/openmpw/pdk_1/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.include /home/andylithia/openmpw/pdk_1/sky130A/libs.ref/sky130_fd_sc_hs/spice/sky130_fd_sc_hs.spice


*.ac dec 100 1e3 1e12
.ic v(vout)=0
.tran 1ns 2500ns
.save all
.control
run
display
plot vout gn gp
.endc


**** end user architecture code
**.ends

* expanding   symbol:  i_type_ota_model.sym # of pins=5
** sym_path: /home/andylithia/openmpw/Project-Reisen-Chip1/xschem/i_type_ota_model.sym
** sch_path: /home/andylithia/openmpw/Project-Reisen-Chip1/xschem/i_type_ota_model.sch
.subckt i_type_ota_model vhi vop vip vin vlo
*.ipin vip
*.ipin vin
*.opin vop
*.iopin vhi
*.iopin vlo
XM2 vmid net1 vlo vlo sky130_fd_pr__nfet_01v8 L=2 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=8 m=8
XM6 net1 net1 vlo vlo sky130_fd_pr__nfet_01v8 L=2 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
I1 vhi net1 20u
XM4 net2 vin vmid vlo sky130_fd_pr__nfet_01v8_lvt L=0.15 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2
XM1 net3 vip vmid vlo sky130_fd_pr__nfet_01v8_lvt L=0.15 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2
XM3 net2 net2 vhi vhi sky130_fd_pr__pfet_01v8 L=0.3 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2
XM5 net3 net3 vhi vhi sky130_fd_pr__pfet_01v8 L=0.3 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2
XM7 vop net3 vhi vhi sky130_fd_pr__pfet_01v8 L=0.3 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=8 m=8
XM8 net4 net2 vhi vhi sky130_fd_pr__pfet_01v8 L=0.3 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=8 m=8
XM9 net4 net4 vlo vlo sky130_fd_pr__nfet_01v8 L=0.3 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4
XM10 vop net4 vlo vlo sky130_fd_pr__nfet_01v8 L=0.3 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4
C1 vop net5 500f m=1
R2 net5 net4 2k m=1
.ends


* expanding   symbol:  swcap_array_PEX.sym # of pins=10
** sym_path: /home/andylithia/openmpw/Project-Reisen-Chip1/xschem/swcap_array_PEX.sym
** sch_path: /home/andylithia/openmpw/Project-Reisen-Chip1/xschem/swcap_array_PEX.sch
.subckt swcap_array_PEX b0 b1 b2 b3 b4 b5 b6 b7 c vsub
*.ipin b0
*.ipin b1
*.ipin b2
*.ipin b3
*.ipin b4
*.ipin b5
*.ipin b6
*.ipin b7
*.iopin c
*.iopin vsub
**** begin user architecture code

.subckt swcap_array C VSUB B0 B1 B2 B3 B4 B5 B6 B7

* NGSPICE file created from swcap_array_1.ext - technology: sky130A

X0 tcap_200f_60/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X1 tcap_200f_60/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X3 tcap_200f_50/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X4 tcap_200f_50/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X5 C tcap_200f_50/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X6 tcap_200f_61/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X7 tcap_200f_61/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X8 C tcap_200f_61/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X9 tcap_200f_40/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X10 tcap_200f_40/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X11 C tcap_200f_40/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X12 tcap_200f_51/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X13 tcap_200f_51/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X14 C tcap_200f_51/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X15 tcap_200f_62/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X16 tcap_200f_62/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X17 C tcap_200f_62/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X18 tcap_200f_30/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X19 tcap_200f_30/a_173_157# B6 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X20 C tcap_200f_30/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X21 tcap_200f_41/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X22 tcap_200f_41/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X23 C tcap_200f_41/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X24 tcap_200f_52/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X25 tcap_200f_52/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X26 C tcap_200f_52/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X27 tcap_200f_63/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X28 tcap_200f_63/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X29 C tcap_200f_63/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X30 tcap_50f_0/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=7.85e+06u
X31 tcap_50f_0/a_173_157# B0 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X32 C tcap_50f_0/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=7.85e+06u
X33 tcap_200f_31/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X34 tcap_200f_31/a_173_157# B6 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X35 C tcap_200f_31/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X36 tcap_200f_42/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X37 tcap_200f_42/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X38 C tcap_200f_42/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X39 tcap_200f_20/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X40 tcap_200f_20/a_173_157# B6 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X41 C tcap_200f_20/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X42 tcap_200f_53/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X43 tcap_200f_53/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X44 C tcap_200f_53/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X45 tcap_200f_64/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X46 tcap_200f_64/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X47 C tcap_200f_64/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X48 tcap_200f_32/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X49 tcap_200f_32/a_173_157# B6 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X50 C tcap_200f_32/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X51 tcap_200f_33/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X52 tcap_200f_33/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X53 C tcap_200f_33/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X54 tcap_200f_43/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X55 tcap_200f_43/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X56 C tcap_200f_43/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X57 tcap_200f_22/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X58 tcap_200f_22/a_173_157# B6 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X59 C tcap_200f_22/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X60 tcap_200f_44/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X61 tcap_200f_44/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X62 C tcap_200f_44/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X63 tcap_200f_21/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X64 tcap_200f_21/a_173_157# B6 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X65 C tcap_200f_21/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X66 tcap_200f_10/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X67 tcap_200f_10/a_173_157# B5 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X68 C tcap_200f_10/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X69 tcap_200f_54/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X70 tcap_200f_54/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X71 C tcap_200f_54/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X72 tcap_200f_11/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X73 tcap_200f_11/a_173_157# B5 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X74 C tcap_200f_11/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X75 tcap_200f_55/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X76 tcap_200f_55/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X77 C tcap_200f_55/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X78 tcap_200f_65/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X79 tcap_200f_65/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X80 C tcap_200f_65/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X81 tcap_200f_34/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X82 tcap_200f_34/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X83 C tcap_200f_34/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X84 tcap_200f_23/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X85 tcap_200f_23/a_173_157# B6 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X86 C tcap_200f_23/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X87 tcap_200f_45/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X88 tcap_200f_45/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X89 C tcap_200f_45/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X90 tcap_200f_12/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X91 tcap_200f_12/a_173_157# B5 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X92 C tcap_200f_12/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X93 tcap_200f_0/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X94 tcap_200f_0/a_173_157# B5 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X95 C tcap_200f_0/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X96 tcap_200f_56/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X97 tcap_200f_56/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X98 C tcap_200f_56/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X99 tcap_200f_35/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X100 tcap_200f_35/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X101 C tcap_200f_35/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X102 tcap_200f_24/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X103 tcap_200f_24/a_173_157# B6 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X104 C tcap_200f_24/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X105 tcap_200f_46/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X106 tcap_200f_46/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X107 C tcap_200f_46/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X108 tcap_200f_13/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X109 tcap_200f_13/a_173_157# B5 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X110 C tcap_200f_13/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X111 tcap_200f_57/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X112 tcap_200f_57/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X113 C tcap_200f_57/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X114 tcap_200f_36/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X115 tcap_200f_36/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X116 C tcap_200f_36/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X117 tcap_200f_25/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X118 tcap_200f_25/a_173_157# B6 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X119 C tcap_200f_25/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X120 tcap_200f_47/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X121 tcap_200f_47/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X122 C tcap_200f_47/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X123 tcap_200f_14/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X124 tcap_200f_14/a_173_157# B5 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X125 C tcap_200f_14/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X126 tcap_200f_58/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X127 tcap_200f_58/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X128 C tcap_200f_58/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X129 tcap_200f_37/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X130 tcap_200f_37/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X131 C tcap_200f_37/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X132 tcap_200f_26/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X133 tcap_200f_26/a_173_157# B6 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X134 C tcap_200f_26/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X135 tcap_200f_15/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X136 tcap_200f_15/a_173_157# B6 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X137 C tcap_200f_15/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X138 tcap_200f_48/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X139 tcap_200f_48/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X140 C tcap_200f_48/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X141 tcap_200f_59/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X142 tcap_200f_59/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X143 C tcap_200f_59/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X144 tcap_200f_3/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X145 tcap_200f_3/a_173_157# B2 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X146 C tcap_200f_3/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X147 tcap_200f_38/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X148 tcap_200f_38/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X149 C tcap_200f_38/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X150 tcap_200f_27/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X151 tcap_200f_27/a_173_157# B6 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X152 C tcap_200f_27/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X153 tcap_200f_16/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X154 tcap_200f_16/a_173_157# B5 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X155 C tcap_200f_16/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X156 tcap_200f_49/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X157 tcap_200f_49/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X158 C tcap_200f_49/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X159 tcap_200f_4/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X160 tcap_200f_4/a_173_157# B3 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X161 C tcap_200f_4/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X162 tcap_200f_28/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X163 tcap_200f_28/a_173_157# B6 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X164 C tcap_200f_28/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X165 tcap_200f_39/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X166 tcap_200f_39/a_173_157# B7 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X167 C tcap_200f_39/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X168 tcap_200f_17/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X169 tcap_200f_17/a_173_157# B5 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X170 C tcap_200f_17/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X171 tcap_200f_5/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X172 tcap_200f_5/a_173_157# B3 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X173 C tcap_200f_5/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X174 tcap_200f_29/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X175 tcap_200f_29/a_173_157# B6 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X176 C tcap_200f_29/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X177 tcap_200f_18/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X178 tcap_200f_18/a_173_157# B6 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X179 C tcap_200f_18/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X180 tcap_200f_6/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X181 tcap_200f_6/a_173_157# B4 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X182 C tcap_200f_6/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X183 tcap_200f_19/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X184 tcap_200f_19/a_173_157# B6 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X185 C tcap_200f_19/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X186 tcap_200f_8/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X187 tcap_200f_8/a_173_157# B4 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X188 C tcap_200f_8/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X189 tcap_200f_7/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X190 tcap_200f_7/a_173_157# B4 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X191 C tcap_200f_7/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X192 tcap_200f_9/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=3.14e+07u
X193 tcap_200f_9/a_173_157# B4 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X194 C tcap_200f_9/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=3.14e+07u
X195 tcap_100f_0/a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=1.57e+07u
X196 tcap_100f_0/a_173_157# B1 VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u
+ l=150000u
X197 C tcap_100f_0/a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=1.57e+07u
C0 C tcap_100f_0/a_173_157# 5.85fF
C1 tcap_200f_36/a_173_157# tcap_200f_37/a_173_157# 4.48fF
C2 tcap_200f_38/a_173_157# tcap_200f_37/a_173_157# 4.48fF
C3 tcap_200f_28/a_173_157# tcap_200f_31/a_173_157# 4.47fF
C4 tcap_200f_10/a_173_157# tcap_200f_13/a_173_157# 4.47fF
C5 tcap_200f_45/a_173_157# C 12.05fF
C6 tcap_200f_44/a_173_157# C 12.05fF
C7 tcap_200f_16/a_173_157# tcap_200f_14/a_173_157# 4.47fF
C8 C tcap_200f_52/a_173_157# 12.05fF
C9 tcap_200f_57/a_173_157# tcap_200f_58/a_173_157# 4.48fF
C10 tcap_200f_17/a_173_157# tcap_200f_16/a_173_157# 4.47fF
C11 tcap_200f_18/a_173_157# C 12.05fF
C12 tcap_200f_12/a_173_157# C 12.05fF
C13 tcap_200f_47/a_173_157# tcap_200f_46/a_173_157# 4.48fF
C14 tcap_200f_49/a_173_157# tcap_200f_50/a_173_157# 4.48fF
C15 tcap_200f_56/a_173_157# C 12.05fF
C16 tcap_200f_54/a_173_157# tcap_200f_53/a_173_157# 4.48fF
C17 tcap_200f_41/a_173_157# tcap_200f_40/a_173_157# 4.48fF
C18 tcap_200f_15/a_173_157# C 12.05fF
C19 C tcap_200f_7/a_173_157# 12.05fF
C20 tcap_200f_15/a_173_157# tcap_200f_25/a_173_157# 4.47fF
C21 tcap_200f_36/a_173_157# C 12.05fF
C22 tcap_200f_38/a_173_157# C 12.05fF
C23 tcap_200f_5/a_173_157# C 12.05fF
C24 tcap_200f_22/a_173_157# C 12.05fF
C25 tcap_200f_42/a_173_157# C 12.05fF
C26 tcap_200f_48/a_173_157# tcap_200f_47/a_173_157# 4.48fF
C27 tcap_200f_34/a_173_157# C 11.79fF
C28 tcap_200f_52/a_173_157# tcap_200f_53/a_173_157# 4.48fF
C29 C tcap_200f_6/a_173_157# 12.05fF
C30 tcap_200f_44/a_173_157# tcap_200f_43/a_173_157# 4.48fF
C31 tcap_200f_31/a_173_157# tcap_200f_30/a_173_157# 4.47fF
C32 tcap_200f_36/a_173_157# tcap_200f_35/a_173_157# 4.48fF
C33 tcap_200f_39/a_173_157# C 12.05fF
C34 tcap_200f_45/a_173_157# tcap_200f_46/a_173_157# 4.48fF
C35 tcap_200f_4/a_173_157# tcap_200f_3/a_173_157# 4.47fF
C36 tcap_200f_16/a_173_157# C 12.05fF
C37 tcap_200f_59/a_173_157# C 12.05fF
C38 tcap_200f_14/a_173_157# C 12.05fF
C39 tcap_200f_23/a_173_157# tcap_200f_22/a_173_157# 4.47fF
C40 tcap_200f_34/a_173_157# tcap_200f_35/a_173_157# 4.48fF
C41 tcap_200f_61/a_173_157# tcap_200f_62/a_173_157# 4.48fF
C42 tcap_200f_55/a_173_157# tcap_200f_54/a_173_157# 4.48fF
C43 C tcap_200f_37/a_173_157# 12.05fF
C44 tcap_200f_15/a_173_157# tcap_200f_27/a_173_157# 4.47fF
C45 tcap_200f_51/a_173_157# tcap_200f_50/a_173_157# 4.48fF
C46 tcap_200f_63/a_173_157# tcap_200f_62/a_173_157# 4.48fF
C47 tcap_200f_57/a_173_157# tcap_200f_56/a_173_157# 4.48fF
C48 tcap_200f_17/a_173_157# C 12.05fF
C49 tcap_200f_11/a_173_157# tcap_200f_0/a_173_157# 4.47fF
C50 tcap_50f_0/a_173_157# C 3.01fF
C51 tcap_200f_8/a_173_157# tcap_200f_7/a_173_157# 4.47fF
C52 tcap_200f_11/a_173_157# C 12.05fF
C53 tcap_200f_42/a_173_157# tcap_200f_43/a_173_157# 4.48fF
C54 tcap_200f_60/a_173_157# tcap_200f_61/a_173_157# 4.48fF
C55 tcap_200f_3/a_173_157# tcap_100f_0/a_173_157# 2.53fF
C56 tcap_200f_21/a_173_157# tcap_200f_22/a_173_157# 4.47fF
C57 tcap_200f_0/a_173_157# C 12.05fF
C58 tcap_200f_24/a_173_157# C 12.05fF
C59 tcap_200f_52/a_173_157# tcap_200f_51/a_173_157# 4.48fF
C60 tcap_200f_55/a_173_157# tcap_200f_56/a_173_157# 4.48fF
C61 tcap_200f_24/a_173_157# tcap_200f_25/a_173_157# 4.47fF
C62 tcap_200f_64/a_173_157# C 11.71fF
C63 tcap_200f_29/a_173_157# C 12.05fF
C64 B4 B5 3.35fF
C65 tcap_200f_20/a_173_157# C 12.05fF
C66 tcap_200f_42/a_173_157# tcap_200f_41/a_173_157# 4.48fF
C67 tcap_200f_25/a_173_157# C 12.05fF
C68 tcap_200f_18/a_173_157# tcap_200f_19/a_173_157# 4.47fF
C69 tcap_200f_23/a_173_157# tcap_200f_24/a_173_157# 4.47fF
C70 tcap_200f_10/a_173_157# tcap_200f_11/a_173_157# 4.47fF
C71 tcap_200f_12/a_173_157# tcap_200f_13/a_173_157# 4.47fF
C72 C tcap_200f_35/a_173_157# 12.05fF
C73 tcap_200f_5/a_173_157# tcap_200f_4/a_173_157# 4.47fF
C74 B5 B6 6.53fF
C75 tcap_200f_29/a_173_157# tcap_200f_28/a_173_157# 4.47fF
C76 tcap_200f_23/a_173_157# C 12.05fF
C77 tcap_200f_26/a_173_157# tcap_200f_29/a_173_157# 4.47fF
C78 tcap_200f_28/a_173_157# C 12.05fF
C79 tcap_200f_44/a_173_157# tcap_200f_45/a_173_157# 4.48fF
C80 tcap_200f_26/a_173_157# C 12.05fF
C81 tcap_200f_9/a_173_157# tcap_200f_0/a_173_157# 4.47fF
C82 tcap_200f_32/a_173_157# C 11.60fF
C83 tcap_200f_10/a_173_157# C 12.05fF
C84 tcap_200f_27/a_173_157# C 12.05fF
C85 tcap_200f_39/a_173_157# tcap_200f_40/a_173_157# 4.48fF
C86 tcap_200f_34/a_173_157# tcap_200f_33/a_173_157# 4.48fF
C87 C tcap_200f_53/a_173_157# 12.05fF
C88 tcap_200f_57/a_173_157# C 12.05fF
C89 tcap_200f_43/a_173_157# C 12.05fF
C90 tcap_200f_9/a_173_157# C 12.05fF
C91 tcap_200f_49/a_173_157# C 12.05fF
C92 C tcap_200f_8/a_173_157# 12.05fF
C93 C tcap_200f_46/a_173_157# 12.05fF
C94 tcap_200f_21/a_173_157# C 12.05fF
C95 tcap_200f_21/a_173_157# tcap_200f_20/a_173_157# 4.47fF
C96 tcap_200f_59/a_173_157# tcap_200f_58/a_173_157# 4.48fF
C97 tcap_200f_64/a_173_157# tcap_200f_65/a_173_157# 4.48fF
C98 C tcap_200f_65/a_173_157# 10.91fF
C99 tcap_200f_41/a_173_157# C 12.05fF
C100 tcap_200f_26/a_173_157# tcap_200f_27/a_173_157# 4.47fF
C101 tcap_200f_48/a_173_157# C 12.05fF
C102 tcap_200f_55/a_173_157# C 12.05fF
C103 tcap_200f_59/a_173_157# tcap_200f_60/a_173_157# 4.48fF
C104 C tcap_200f_30/a_173_157# 11.79fF
C105 tcap_200f_4/a_173_157# C 11.89fF
C106 B7 B6 9.55fF
C107 C tcap_200f_62/a_173_157# 12.05fF
C108 C tcap_200f_51/a_173_157# 12.05fF
C109 tcap_200f_19/a_173_157# C 12.05fF
C110 tcap_200f_19/a_173_157# tcap_200f_20/a_173_157# 4.47fF
C111 tcap_200f_9/a_173_157# tcap_200f_8/a_173_157# 4.47fF
C112 C tcap_200f_40/a_173_157# 12.05fF
C113 C tcap_200f_13/a_173_157# 12.05fF
C114 tcap_200f_6/a_173_157# tcap_200f_7/a_173_157# 4.47fF
C115 C tcap_200f_3/a_173_157# 11.41fF
C116 tcap_200f_33/a_173_157# C 11.60fF
C117 tcap_200f_61/a_173_157# C 12.05fF
C118 tcap_200f_14/a_173_157# tcap_200f_12/a_173_157# 4.47fF
C119 tcap_200f_47/a_173_157# C 12.05fF
C120 tcap_200f_58/a_173_157# C 12.05fF
C121 C tcap_200f_31/a_173_157# 12.05fF
C122 tcap_200f_64/a_173_157# tcap_200f_63/a_173_157# 4.48fF
C123 tcap_200f_5/a_173_157# tcap_200f_6/a_173_157# 4.47fF
C124 tcap_200f_32/a_173_157# tcap_200f_30/a_173_157# 4.47fF
C125 C tcap_200f_50/a_173_157# 12.05fF
C126 tcap_200f_39/a_173_157# tcap_200f_38/a_173_157# 4.48fF
C127 C tcap_200f_63/a_173_157# 12.04fF
C128 tcap_200f_18/a_173_157# tcap_200f_17/a_173_157# 4.47fF
C129 tcap_200f_48/a_173_157# tcap_200f_49/a_173_157# 4.48fF
C130 tcap_200f_60/a_173_157# C 12.05fF
C131 tcap_200f_54/a_173_157# C 12.05fF
C132 tcap_100f_0/a_173_157# VSUB 4.99fF $ **FLOATING
C133 tcap_200f_9/a_173_157# VSUB 7.94fF $ **FLOATING
C134 tcap_200f_7/a_173_157# VSUB 7.94fF $ **FLOATING
C135 tcap_200f_8/a_173_157# VSUB 7.94fF $ **FLOATING
C136 tcap_200f_19/a_173_157# VSUB 7.94fF $ **FLOATING
C137 tcap_200f_6/a_173_157# VSUB 7.94fF $ **FLOATING
C138 B4 VSUB 5.01fF $ **FLOATING
C139 tcap_200f_18/a_173_157# VSUB 7.94fF $ **FLOATING
C140 B6 VSUB 22.15fF $ **FLOATING
C141 tcap_200f_29/a_173_157# VSUB 7.94fF $ **FLOATING
C142 tcap_200f_5/a_173_157# VSUB 7.94fF $ **FLOATING
C143 tcap_200f_17/a_173_157# VSUB 7.94fF $ **FLOATING
C144 tcap_200f_39/a_173_157# VSUB 7.96fF $ **FLOATING
C145 tcap_200f_28/a_173_157# VSUB 7.94fF $ **FLOATING
C146 tcap_200f_4/a_173_157# VSUB 7.94fF $ **FLOATING
C147 B3 VSUB 2.41fF $ **FLOATING
C148 tcap_200f_49/a_173_157# VSUB 7.96fF $ **FLOATING
C149 tcap_200f_16/a_173_157# VSUB 7.94fF $ **FLOATING
C150 tcap_200f_27/a_173_157# VSUB 7.94fF $ **FLOATING
C151 tcap_200f_38/a_173_157# VSUB 7.96fF $ **FLOATING
C152 tcap_200f_3/a_173_157# VSUB 7.94fF $ **FLOATING
C153 tcap_200f_59/a_173_157# VSUB 7.95fF $ **FLOATING
C154 tcap_200f_48/a_173_157# VSUB 7.96fF $ **FLOATING
C155 tcap_200f_15/a_173_157# VSUB 7.94fF $ **FLOATING
C156 tcap_200f_26/a_173_157# VSUB 7.94fF $ **FLOATING
C157 tcap_200f_37/a_173_157# VSUB 7.96fF $ **FLOATING
C158 tcap_200f_58/a_173_157# VSUB 7.95fF $ **FLOATING
C159 tcap_200f_14/a_173_157# VSUB 7.94fF $ **FLOATING
C160 tcap_200f_47/a_173_157# VSUB 7.96fF $ **FLOATING
C161 tcap_200f_25/a_173_157# VSUB 7.94fF $ **FLOATING
C162 tcap_200f_36/a_173_157# VSUB 7.96fF $ **FLOATING
C163 tcap_200f_57/a_173_157# VSUB 7.95fF $ **FLOATING
C164 tcap_200f_13/a_173_157# VSUB 7.94fF $ **FLOATING
C165 tcap_200f_46/a_173_157# VSUB 7.96fF $ **FLOATING
C166 tcap_200f_24/a_173_157# VSUB 7.94fF $ **FLOATING
C167 tcap_200f_35/a_173_157# VSUB 7.96fF $ **FLOATING
C168 tcap_200f_56/a_173_157# VSUB 7.95fF $ **FLOATING
C169 tcap_200f_0/a_173_157# VSUB 7.94fF $ **FLOATING
C170 B5 VSUB 10.51fF $ **FLOATING
C171 tcap_200f_12/a_173_157# VSUB 7.94fF $ **FLOATING
C172 tcap_200f_45/a_173_157# VSUB 7.96fF $ **FLOATING
C173 tcap_200f_23/a_173_157# VSUB 7.94fF $ **FLOATING
C174 tcap_200f_34/a_173_157# VSUB 7.95fF $ **FLOATING
C175 C VSUB 71.74fF $ **FLOATING
C176 tcap_200f_65/a_173_157# VSUB 7.92fF $ **FLOATING
C177 B7 VSUB 28.92fF $ **FLOATING
C178 tcap_200f_55/a_173_157# VSUB 7.95fF $ **FLOATING
C179 tcap_200f_11/a_173_157# VSUB 7.94fF $ **FLOATING
C180 tcap_200f_54/a_173_157# VSUB 7.95fF $ **FLOATING
C181 tcap_200f_10/a_173_157# VSUB 7.94fF $ **FLOATING
C182 tcap_200f_21/a_173_157# VSUB 7.94fF $ **FLOATING
C183 tcap_200f_44/a_173_157# VSUB 7.96fF $ **FLOATING
C184 tcap_200f_22/a_173_157# VSUB 7.94fF $ **FLOATING
C185 tcap_200f_43/a_173_157# VSUB 7.96fF $ **FLOATING
C186 tcap_200f_33/a_173_157# VSUB 7.96fF $ **FLOATING
C187 tcap_200f_32/a_173_157# VSUB 7.96fF $ **FLOATING
C188 tcap_200f_64/a_173_157# VSUB 7.93fF $ **FLOATING
C189 tcap_200f_53/a_173_157# VSUB 7.95fF $ **FLOATING
C190 tcap_200f_20/a_173_157# VSUB 7.94fF $ **FLOATING
C191 tcap_200f_42/a_173_157# VSUB 7.96fF $ **FLOATING
C192 tcap_200f_31/a_173_157# VSUB 7.94fF $ **FLOATING
C193 tcap_50f_0/a_173_157# VSUB 3.60fF $ **FLOATING
C194 tcap_200f_63/a_173_157# VSUB 7.94fF $ **FLOATING
C195 tcap_200f_52/a_173_157# VSUB 7.95fF $ **FLOATING
C196 tcap_200f_41/a_173_157# VSUB 7.96fF $ **FLOATING
C197 tcap_200f_30/a_173_157# VSUB 7.94fF $ **FLOATING
C198 tcap_200f_62/a_173_157# VSUB 7.94fF $ **FLOATING
C199 tcap_200f_51/a_173_157# VSUB 7.95fF $ **FLOATING
C200 tcap_200f_40/a_173_157# VSUB 7.96fF $ **FLOATING
C201 tcap_200f_61/a_173_157# VSUB 7.95fF $ **FLOATING
C202 tcap_200f_50/a_173_157# VSUB 7.95fF $ **FLOATING
C203 tcap_200f_60/a_173_157# VSUB 7.95fF $ **FLOATING



.ends
XDUT c vsub b0 b1 b2 b3 b4 b5 b6 b7 swcap_array



**** end user architecture code
.ends


* expanding   symbol:  twcon_PEX.sym # of pins=14
** sym_path: /home/andylithia/openmpw/Project-Reisen-Chip1/xschem/twcon_PEX.sym
** sch_path: /home/andylithia/openmpw/Project-Reisen-Chip1/xschem/twcon_PEX.sch
.subckt twcon_PEX GP VHI GN VLO UPDN CLKIN MUX_OUT UDCLK A0 ENCLK A1 RSTB C100 C50
*.iopin VHI
*.iopin VLO
*.opin UPDN
*.ipin CLKIN
*.ipin A0
*.ipin A1
*.ipin RSTB
*.ipin C100
*.ipin C50
*.opin GP
*.opin GN
*.opin MUX_OUT
*.opin UDCLK
*.opin ENCLK
**** begin user architecture code

* NGSPICE file created from twcon.ext - technology: sky130A

* NGSPICE file created from twcon.ext - technology: sky130A

.subckt sky130_fd_sc_hs__decap_8 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8 ad=8.35e+11p pd=7.67e+06u as=0p ps=0u w=1e+06u
+ l=1e+06u
X1 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X2 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=3.465e+11p pd=4.17e+06u as=0p ps=0u w=420000u
+ l=1e+06u
X3 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=1e+06u
.ends

.subckt tcap_50f C S VLO
X0 a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=7.85e+06u
X1 a_173_157# S VLO VLO sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u
+ w=2e+06u l=150000u
X2 C a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=7.85e+06u
.ends

.subckt sky130_fd_sc_hs__mux2_1 A0 A1 S VGND VPWR X VNB VPB
X0 VGND a_27_112# a_443_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=7.0725e+11p pd=4.91e+06u
+ as=5.994e+11p ps=3.1e+06u w=740000u l=150000u
X1 VPWR S a_27_112# VPB sky130_fd_pr__pfet_01v8 ad=8.82e+11p pd=5.95e+06u as=2.478e+11p ps=2.27e+06u
+ w=840000u l=150000u
X2 X a_304_74# VPWR VPB sky130_fd_pr__pfet_01v8 ad=3.304e+11p pd=2.83e+06u as=0p ps=0u w=1.12e+06u
+ l=150000u
X3 VPWR a_27_112# a_524_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.2e+11p ps=2.84e+06u
+ w=1e+06u l=150000u
X4 a_304_74# A1 a_226_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=4.033e+11p pd=2.57e+06u as=1.776e+11p
+ ps=1.96e+06u w=740000u l=150000u
X5 X a_304_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=2.109e+11p pd=2.05e+06u as=0p ps=0u w=740000u
+ l=150000u
X6 a_223_368# S VPWR VPB sky130_fd_pr__pfet_01v8 ad=8.15e+11p pd=3.63e+06u as=0p ps=0u w=1e+06u
+ l=150000u
X7 a_304_74# A0 a_223_368# VPB sky130_fd_pr__pfet_01v8 ad=3.9e+11p pd=2.78e+06u as=0p ps=0u w=1e+06u
+ l=150000u
X8 a_443_74# A0 a_304_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u
+ l=150000u
X9 a_524_368# A1 a_304_74# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_226_74# S VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X11 VGND S a_27_112# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
+ w=550000u l=150000u
.ends

.subckt sky130_fd_sc_hs__decap_4 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8 ad=5.6e+11p pd=5.12e+06u as=0p ps=0u w=1e+06u l=1e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=2.31e+11p pd=2.78e+06u as=0p ps=0u w=420000u
+ l=1e+06u
.ends

.subckt tcap_100f C S VLO
X0 a_173_157# C sky130_fd_pr__cap_mim_m3_2 l=1.6e+06u w=1.57e+07u
X1 a_173_157# S VLO VLO sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u
+ w=2e+06u l=150000u
X2 C a_173_157# sky130_fd_pr__cap_mim_m3_1 l=1.6e+06u w=1.57e+07u
.ends

.subckt sky130_fd_sc_hs__sdfbbn_2 CLK_N D RESET_B SCD SCE SET_B VGND VPWR Q Q_N VNB  VPB
X0 a_1997_82# a_868_368# a_1986_424# VPB sky130_fd_pr__pfet_01v8 ad=2.856e+11p pd=2.45e+06u
+ as=2.016e+11p ps=2.16e+06u w=840000u l=150000u
X1 a_1185_125# a_1007_366# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=8.82e+10p pd=1.26e+06u
+ as=2.86405e+12p ps=2.37e+07u w=420000u l=150000u
X2 a_2452_74# SET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=5.7435e+11p pd=4.64e+06u as=0p ps=0u
+ w=740000u l=150000u
X3 a_1070_464# a_1007_366# VPWR VPB sky130_fd_pr__pfet_01v8 ad=1.134e+11p pd=1.38e+06u
+ as=4.12873e+12p ps=3.022e+07u w=420000u l=150000u
X4 a_363_119# D a_197_119# VNB sky130_fd_pr__nfet_01v8_lvt ad=1.008e+11p pd=1.32e+06u as=4.347e+11p
+ ps=3.75e+06u w=420000u l=150000u
X5 VGND a_2216_410# Q_N VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.072e+11p ps=2.04e+06u
+ w=740000u l=150000u
X6 VGND a_2216_410# a_3272_94# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.824e+11p
+ ps=1.85e+06u w=640000u l=150000u
X7 a_119_119# SCD VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
+ w=420000u l=150000u
X8 VGND SET_B a_1473_73# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=6.0335e+11p ps=4.55e+06u
+ w=550000u l=150000u
X9 a_2247_82# a_868_368# a_1997_82# VNB sky130_fd_pr__nfet_01v8_lvt ad=1.008e+11p pd=1.32e+06u
+ as=4.945e+11p ps=3.3e+06u w=420000u l=150000u
X10 VGND CLK_N a_688_98# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
+ w=740000u l=150000u
X11 a_868_368# a_688_98# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
+ w=740000u l=150000u
X12 VPWR a_3272_94# Q VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.36e+11p ps=2.84e+06u w=1.12e+06u
+ l=150000u
X13 a_2452_74# a_1997_82# a_2216_410# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.072e+11p
+ ps=2.04e+06u w=740000u l=150000u
X14 VPWR SCD a_27_464# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.776e+11p ps=3.74e+06u w=640000u
+ l=150000u
X15 Q a_3272_94# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X16 a_1986_424# a_1007_366# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u
+ l=150000u
X17 VPWR a_2216_410# a_2171_508# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
+ w=420000u l=150000u
X18 a_2216_410# a_1997_82# a_2556_392# VPB sky130_fd_pr__pfet_01v8 ad=5.9e+11p pd=5.18e+06u
+ as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X19 a_341_410# SCE VPWR VPB sky130_fd_pr__pfet_01v8 ad=1.888e+11p pd=1.87e+06u as=0p ps=0u w=640000u
+ l=150000u
X20 a_1007_366# a_1154_464# a_1473_73# VNB sky130_fd_pr__nfet_01v8_lvt ad=1.54e+11p pd=1.66e+06u
+ as=0p ps=0u w=550000u l=150000u
X21 VPWR SET_B a_2216_410# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VGND a_3272_94# Q VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.072e+11p ps=2.04e+06u
+ w=740000u l=150000u
X23 VPWR a_1643_257# a_1592_424# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.268e+11p ps=2.22e+06u
+ w=840000u l=150000u
X24 a_2171_508# a_688_98# a_1997_82# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u
+ l=150000u
X25 a_1997_82# a_688_98# a_1902_125# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.16375e+11p
+ ps=2.18e+06u w=550000u l=150000u
X26 a_2556_392# a_1643_257# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u
+ l=150000u
X27 a_1592_424# a_1154_464# a_1007_366# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=9.954e+11p
+ ps=5.73e+06u w=840000u l=150000u
X28 a_1007_366# SET_B VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X29 VPWR RESET_B a_1643_257# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.888e+11p ps=1.87e+06u
+ w=640000u l=150000u
X30 VPWR a_2216_410# Q_N VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.36e+11p ps=2.84e+06u
+ w=1.12e+06u l=150000u
X31 a_2216_410# a_1643_257# a_2452_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u
+ w=740000u l=150000u
X32 a_197_119# SCE a_119_119# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u
+ l=150000u
X33 Q_N a_2216_410# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X34 VGND a_2216_410# a_2247_82# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u
+ l=150000u
X35 a_27_464# a_341_410# a_197_119# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.128e+11p
+ ps=3.85e+06u w=640000u l=150000u
X36 a_1473_73# a_1643_257# a_1007_366# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u
+ w=550000u l=150000u
X37 a_197_119# D a_206_464# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.536e+11p ps=1.76e+06u
+ w=640000u l=150000u
X38 a_1154_464# a_688_98# a_1185_125# VNB sky130_fd_pr__nfet_01v8_lvt ad=1.281e+11p pd=1.45e+06u
+ as=0p ps=0u w=420000u l=150000u
X39 a_1902_125# a_1007_366# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=550000u
+ l=150000u
X40 Q a_3272_94# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X41 a_197_119# a_688_98# a_1154_464# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.266e+11p
+ ps=2.05e+06u w=640000u l=150000u
X42 VPWR a_2216_410# a_3272_94# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
+ w=1e+06u l=150000u
X43 VGND RESET_B a_1643_257# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
+ w=420000u l=150000u
X44 a_868_368# a_688_98# VPWR VPB sky130_fd_pr__pfet_01v8 ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
+ w=1.12e+06u l=150000u
X45 a_197_119# a_868_368# a_1154_464# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u
+ w=420000u l=150000u
X46 a_206_464# SCE VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X47 VPWR CLK_N a_688_98# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.304e+11p ps=2.83e+06u
+ w=1.12e+06u l=150000u
X48 a_1154_464# a_868_368# a_1070_464# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u
+ l=150000u
X49 VGND a_341_410# a_363_119# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u
+ l=150000u
X50 a_341_410# SCE VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
+ w=420000u l=150000u
X51 Q_N a_2216_410# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
.ends

.subckt sky130_fd_sc_hs__inv_1 A VGND VPWR Y VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8 ad=3.304e+11p pd=2.83e+06u as=3.864e+11p ps=2.93e+06u
+ w=1.12e+06u l=150000u
X1 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=2.109e+11p pd=2.05e+06u as=2.627e+11p ps=2.19e+06u
+ w=740000u l=150000u
.ends

.subckt sky130_fd_sc_hs__nand2_1 A B VGND VPWR Y VNB VPB
X0 a_117_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=1.776e+11p pd=1.96e+06u as=2.109e+11p
+ ps=2.05e+06u w=740000u l=150000u
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8 ad=6.384e+11p pd=5.62e+06u as=3.36e+11p ps=2.84e+06u
+ w=1.12e+06u l=150000u
X2 Y A a_117_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=2.109e+11p pd=2.05e+06u as=0p ps=0u w=740000u
+ l=150000u
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_GKKP9B a_n141_n482# a_n141_50# VSUBS
X0 a_n141_n482# a_n141_50# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=500000u
.ends

.subckt twcon_tdly C A Y sky130_fd_sc_hs__inv_1_0/VGND VSUBS sky130_fd_sc_hs__inv_1_0/VPWR
+  sky130_fd_sc_hs__inv_1_0/VPB
Xsky130_fd_sc_hs__inv_1_0 A sky130_fd_sc_hs__inv_1_0/VGND sky130_fd_sc_hs__inv_1_0/VPWR
+  sky130_fd_sc_hs__inv_1_0/Y VSUBS sky130_fd_sc_hs__inv_1_0/VPB sky130_fd_sc_hs__inv_1
Xsky130_fd_sc_hs__nand2_1_2 A C sky130_fd_sc_hs__inv_1_0/VGND sky130_fd_sc_hs__inv_1_0/VPWR  Y VSUBS
+ sky130_fd_sc_hs__inv_1_0/VPB sky130_fd_sc_hs__nand2_1
Xsky130_fd_pr__res_xhigh_po_1p41_GKKP9B_0 sky130_fd_sc_hs__inv_1_0/Y C VSUBS
+ sky130_fd_pr__res_xhigh_po_1p41_GKKP9B
.ends

.subckt sky130_fd_sc_hs__nand2_4 A B VGND VPWR Y VNB VPB
X0 Y A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=5.365e+11p pd=4.41e+06u as=1.1581e+12p
+ ps=1.053e+07u w=740000u l=150000u
X1 Y B VPWR VPB sky130_fd_pr__pfet_01v8 ad=2.7496e+12p pd=9.39e+06u as=1.1144e+12p ps=8.71e+06u
+ w=1.12e+06u l=150000u
X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X3 Y A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X4 Y A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X5 VGND B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=4.144e+11p pd=4.08e+06u as=0p ps=0u w=740000u
+ l=150000u
X6 a_27_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X7 VPWR B Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X8 a_27_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X9 a_27_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X10 a_27_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X11 VGND B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
.ends

.subckt sky130_fd_sc_hs__inv_2 A VGND VPWR Y VNB VPB
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=2.072e+11p pd=2.04e+06u as=4.218e+11p ps=4.1e+06u
+ w=740000u l=150000u
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8 ad=6.384e+11p pd=5.62e+06u as=3.36e+11p ps=2.84e+06u
+ w=1.12e+06u l=150000u
X2 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X3 Y A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
.ends

.subckt sky130_fd_sc_hs__and2_4 A B VGND VPWR X VNB VPB
X0 X a_83_269# VPWR VPB sky130_fd_pr__pfet_01v8 ad=6.944e+11p pd=5.72e+06u as=1.58705e+12p
+ ps=1.328e+07u w=1.12e+06u l=150000u
X1 a_83_269# B VPWR VPB sky130_fd_pr__pfet_01v8 ad=5.25e+11p pd=4.61e+06u as=0p ps=0u w=840000u
+ l=150000u
X2 a_83_269# A a_504_119# VNB sky130_fd_pr__nfet_01v8_lvt ad=2.08e+11p pd=1.93e+06u as=3.872e+11p
+ ps=3.77e+06u w=640000u l=150000u
X3 VPWR a_83_269# X VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X4 VGND a_83_269# X VNB sky130_fd_pr__nfet_01v8_lvt ad=8.594e+11p pd=8.14e+06u as=5.254e+11p
+ ps=4.38e+06u w=740000u l=150000u
X5 X a_83_269# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X6 X a_83_269# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X7 VPWR a_83_269# X VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X8 VPWR B a_83_269# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X9 a_83_269# A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X10 VGND a_83_269# X VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X11 VPWR A a_83_269# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X12 VGND B a_504_119# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X13 a_504_119# A a_83_269# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u
+ l=150000u
X14 X a_83_269# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X15 a_504_119# B VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
.ends

.subckt twcon UPDN CLKIN A0 A1 RSTB VHI VLO C100 C50 MUX_OUT ENCLK GN GP
Xsky130_fd_sc_hs__decap_8_0 VLO VHI VLO VHI sky130_fd_sc_hs__decap_8
Xtcap_50f_0 tcap_50f_0/C C100 VLO tcap_50f
Xsky130_fd_sc_hs__decap_8_2 VLO VHI VLO VHI sky130_fd_sc_hs__decap_8
Xsky130_fd_sc_hs__decap_8_3 VLO VHI VLO VHI sky130_fd_sc_hs__decap_8
Xtcap_50f_3 tcap_50f_3/C C100 VLO tcap_50f
Xsky130_fd_sc_hs__decap_8_4 VLO VHI VLO VHI sky130_fd_sc_hs__decap_8
Xtcap_50f_2 tcap_50f_2/C C50 VLO tcap_50f
Xsky130_fd_sc_hs__mux2_1_1 twcon_tdly_1/Y twcon_tdly_2/Y sky130_fd_sc_hs__mux2_1_1/S  VLO VHI
+ MUX_OUT VLO VHI sky130_fd_sc_hs__mux2_1
Xsky130_fd_sc_hs__decap_8_6 VLO VHI VLO VHI sky130_fd_sc_hs__decap_8
Xsky130_fd_sc_hs__decap_4_0 VLO VHI VLO VHI sky130_fd_sc_hs__decap_4
Xsky130_fd_sc_hs__decap_8_7 VLO VHI VLO VHI sky130_fd_sc_hs__decap_8
Xtcap_100f_0 tcap_50f_0/C C50 VLO tcap_100f
Xtcap_100f_2 tcap_50f_2/C C100 VLO tcap_100f
Xtcap_100f_3 tcap_50f_3/C C50 VLO tcap_100f
Xsky130_fd_sc_hs__sdfbbn_2_0 ENCLK VHI MUX_OUT VLO VLO VHI VLO VHI sky130_fd_sc_hs__and2_4_0/B
+  sky130_fd_sc_hs__sdfbbn_2_0/Q_N VLO VHI sky130_fd_sc_hs__sdfbbn_2
Xsky130_fd_sc_hs__sdfbbn_2_1 twcon_tdly_0/Y sky130_fd_sc_hs__mux2_1_1/S RSTB VLO VLO  VHI VLO VHI
+ UPDN sky130_fd_sc_hs__mux2_1_1/S VLO VHI sky130_fd_sc_hs__sdfbbn_2
Xtwcon_tdly_0 tcap_50f_2/C CLKIN twcon_tdly_0/Y VLO VLO VHI VHI twcon_tdly
Xtwcon_tdly_1 tcap_50f_0/C A0 twcon_tdly_1/Y VLO VLO VHI VHI twcon_tdly
Xtwcon_tdly_2 tcap_50f_3/C A1 twcon_tdly_2/Y VLO VLO VHI VHI twcon_tdly
Xsky130_fd_sc_hs__nand2_4_3 sky130_fd_sc_hs__and2_4_0/B UPDN VLO VHI GP VLO VHI
+ sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__inv_2_1 CLKIN VLO VHI ENCLK VLO VHI sky130_fd_sc_hs__inv_2
Xsky130_fd_sc_hs__and2_4_0 sky130_fd_sc_hs__mux2_1_1/S sky130_fd_sc_hs__and2_4_0/B  VLO VHI GN VLO
+ VHI sky130_fd_sc_hs__and2_4
.ends



XDUT UPDN CLKIN A0 A1 RSTB VHI VLO C100 C50 MUX_OUT ENCLK GN GP twcon


**** end user architecture code
.ends


* expanding   symbol:  isrc_PEX.sym # of pins=8
** sym_path: /home/andylithia/openmpw/Project-Reisen-Chip1/xschem/isrc_PEX.sym
** sch_path: /home/andylithia/openmpw/Project-Reisen-Chip1/xschem/isrc_PEX.sch
.subckt isrc_PEX VHI VLO VREFP VREFN IOUT IIN GP GN
*.iopin VHI
*.iopin VLO
*.iopin VREFP
*.iopin IOUT
*.iopin VREFN
*.iopin IIN
*.ipin GP
*.ipin GN
**** begin user architecture code

.subckt isrc VHI VLO IIN IOUT GN GP VREFP VREFN

X1 VHI GN IN VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X2 VHI VHI VREFP VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=2e+06u
X3 VLO GP IP VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4 VLO VLO a_314_3386# VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X5 a_314_3386# VREFP VLO sky130_fd_pr__res_xhigh_po w=350000u l=5.17e+06u
X7 VLO VLO VREFN VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X8 IP VREFP VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=2e+06u
X9 IN VREFN VLO VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X10 IOUT GP IP VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X11 VHI VHI IP VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=2e+06u
X12 VREFN VREFN VLO VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X13 IOUT GN IN VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X14 VLO VLO IN VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X15 VREFP VREFP VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=2e+06u
X16 a_314_3386# VREFN VLO VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
C0 VHI IN 2.47fF
C1 IOUT IP 2.22fF
C2 VHI IP 3.75fF
C3 VHI VREFP 6.31fF
C4 VREFN VLO 7.88fF $ **FLOATING
C5 IN VLO 2.16fF $ **FLOATING
C6 a_314_3386# VLO 2.09fF $ **FLOATING
C7 VHI VLO 30.82fF $ **FLOATING

.ends


XDUT VHI VLO IIN IOUT GN GP VREFP VREFN isrc


**** end user architecture code
.ends


* expanding   symbol:  i_type_ota_gb_rp_gp_PEX.sym # of pins=8
** sym_path: /home/andylithia/openmpw/Project-Reisen-Chip1/xschem/i_type_ota_gb_rp_gp_PEX.sym
** sch_path: /home/andylithia/openmpw/Project-Reisen-Chip1/xschem/i_type_ota_gb_rp_gp_PEX.sch
.subckt i_type_ota_gb_rp_gp_PEX vhi vop vin vip vref s sbar vlo
*.ipin vip
*.ipin vin
*.opin vop
*.iopin vhi
*.iopin vlo
*.ipin vref
*.ipin s
*.ipin sbar
*.iopin vlo
**** begin user architecture code

* NGSPICE file created from cmota_1_flat.ext - technology: sky130A
* NGSPICE file created from cmota_gb_rp_gp.ext - technology: sky130A
.subckt imirror2 OUT a_5468_1540# a_4094_1540# a_4493_207# VLO VHI a_5868_1637# IN  a_4036_1637#
X0 VHI a_4493_207# a_4493_207# VHI.t5 sky130_fd_pr__pfet_01v8 ad=2.9e+12p pd=2.058e+07u as=2.9e+12p
+ ps=2.058e+07u w=1e+07u l=2e+06u
X1 a_4493_207# VLO.t6 VLO.t8 VLO.t7 sky130_fd_pr__nfet_01v8 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u
+ w=5e+06u l=2e+06u
X2 VLO.t5 VLO.t3 OUT VLO.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.45e+12p ps=1.058e+07u w=5e+06u
+ l=2e+06u
X3 a_5868_1637# a_5468_1540# OUT VHI.t0 sky130_fd_pr__pfet_01v8 ad=2.9e+12p pd=2.058e+07u
+ as=2.9e+12p ps=2.058e+07u w=1e+07u l=2e+06u
X4 OUT OUT.t0 VLO VLO.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.35e+12p ps=3.174e+07u w=5e+06u
+ l=2e+06u
X5 VLO IN.t0 a_4493_207# VLO.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X6 a_4493_207# a_4094_1540# a_4036_1637# VHI.t1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.9e+12p
+ ps=2.058e+07u w=1e+07u l=2e+06u
X7 OUT a_4493_207# VHI VHI.t2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=2e+06u
R0 VHI.t2 VHI.t0 178.465
R1 VHI.t5 VHI.t1 178.465
R2 VHI.t0 VHI.n1 133.656
R3 VHI.t1 VHI.n3 133.656
R4 VHI.n6 VHI.t2 89.232
R5 VHI.n6 VHI.t5 89.232
R6 VHI.n9 VHI.n8 3.388
R7 VHI VHI.n9 1.702
R8 VHI.n5 VHI.n4 0.002
R9 VHI.n6 VHI.n5 0.002
R10 VHI.n8 VHI.n7 0.002
R11 VHI.n7 VHI.n6 0.002
R12 VHI.n3 VHI.n2 0.002
R13 VHI.n1 VHI.n0 0.002
R14 VLO.n4 VLO.t4 1062.83
R15 VLO.n7 VLO.t7 1062.83
R16 VLO.n15 VLO.t0 709.577
R17 VLO.n15 VLO.t9 709.577
R18 VLO.n13 VLO.n11 344.847
R19 VLO.n13 VLO.n12 344.847
R20 VLO.n6 VLO.n5 264.873
R21 VLO.n9 VLO.n8 264.496
R22 VLO.n21 VLO.n19 202.541
R23 VLO.n2 VLO.n0 202.541
R24 VLO.t6 VLO.n20 153.089
R25 VLO.n21 VLO.t6 153.089
R26 VLO.n2 VLO.t3 153.089
R27 VLO.t3 VLO.n1 153.089
R28 VLO.n22 VLO.n21 32.935
R29 VLO.n3 VLO.n2 32.935
R30 VLO.n24 VLO.n9 10.039
R31 VLO.n24 VLO.n6 10.037
R32 VLO.n24 VLO.n18 8.178
R33 VLO.n24 VLO.n23 8.178
R34 VLO.n23 VLO.n22 8.01
R35 VLO.n6 VLO.n3 6.032
R36 VLO.n24 VLO.n17 3.765
R37 VLO.n19 VLO.t8 3.48
R38 VLO.n0 VLO.t5 3.48
R39 VLO VLO.n24 1.562
R40 VLO.n17 VLO.n10 1.127
R41 VLO.n17 VLO.n16 0.014
R42 VLO.n16 VLO.n15 0.014
R43 VLO.n8 VLO.n7 0.012
R44 VLO.n5 VLO.n4 0.012
R45 VLO.n14 VLO.n13 0.007
R46 VLO.n15 VLO.n14 0.007
R47 OUT OUT.t0 68.216
R48 IN IN.t0 67.356
C0 a_4036_1637# VHI 0.68fF
C1 a_4493_207# VHI 3.25fF
C2 a_5468_1540# a_5868_1637# 0.15fF
C3 a_4094_1540# a_5868_1637# 0.01fF
C4 a_4493_207# a_4036_1637# 0.63fF
C5 IN OUT 0.22fF
C6 a_5468_1540# OUT 0.53fF
C7 a_4094_1540# OUT 0.10fF
C8 IN VHI 0.19fF
C9 a_5468_1540# VHI 0.99fF
C10 a_4036_1637# IN 0.03fF
C11 a_4094_1540# VHI 0.99fF
C12 a_4493_207# IN 0.46fF
C13 a_5468_1540# a_4036_1637# 0.01fF
C14 a_4493_207# a_5468_1540# 0.22fF
C15 a_4094_1540# a_4036_1637# 0.15fF
C16 a_4094_1540# a_4493_207# 0.44fF
C17 a_5868_1637# OUT 0.47fF
C18 a_5868_1637# VHI 0.45fF
C19 a_4493_207# a_5868_1637# 0.22fF
C20 a_4094_1540# IN 0.17fF
C21 a_4094_1540# a_5468_1540# 0.00fF
C22 VHI OUT 1.31fF
C23 a_4036_1637# OUT 0.03fF
C24 a_4493_207# OUT 0.88fF
C25 OUT VLO 5.14fF
C26 VHI VLO 19.08fF
C27 IN VLO 2.36fF
C28 a_5868_1637# VLO 0.34fF
C29 a_4036_1637# VLO 0.34fF
C30 a_5468_1540# VLO 0.34fF
C31 a_4493_207# VLO 1.55fF
C32 a_4094_1540# VLO 0.34fF
C33 OUT.t0 VLO 1.25fF
C34 VHI.n0 VLO 0.25fF $ **FLOATING
C35 VHI.n1 VLO 2.09fF $ **FLOATING
C36 VHI.t0 VLO 3.29fF
C37 VHI.t2 VLO 2.82fF
C38 VHI.n2 VLO 0.25fF $ **FLOATING
C39 VHI.n3 VLO 2.09fF $ **FLOATING
C40 VHI.t1 VLO 3.29fF
C41 VHI.t5 VLO 2.82fF
C42 VHI.n4 VLO 0.25fF $ **FLOATING
C43 VHI.n5 VLO 0.25fF $ **FLOATING
C44 VHI.n6 VLO 1.88fF $ **FLOATING
C45 VHI.n7 VLO 0.25fF $ **FLOATING
C46 VHI.n8 VLO 0.13fF $ **FLOATING
C47 VHI.n9 VLO 2.08fF $ **FLOATING
.ends

.subckt gated_iref_fix imirror2_0/a_5468_1540# imirror2_0/a_4094_1540# SBAR a_1444_106#
+  imirror2_0/OUT imirror2_0/a_5868_1637# VSUB imirror2_0/VHI imirror2_0/a_4493_207#  imirror2_0/a_4036_1637#
+ a_1712_150# S imirror2_0/IN
Ximirror2_0 imirror2_0/OUT imirror2_0/a_5468_1540# imirror2_0/a_4094_1540# imirror2_0/a_4493_207#
+  VSUB imirror2_0/VHI imirror2_0/a_5868_1637# imirror2_0/IN imirror2_0/a_4036_1637#  imirror2
X0 imirror2_0/OUT a_1444_106# VSUB sky130_fd_pr__res_xhigh_po w=350000u l=1.49e+06u
X1 VSUB SBAR a_1712_150# VSUB sky130_fd_pr__nfet_01v8 ad=5.95e+12p pd=4.302e+07u as=1.65e+12p
+ ps=1.132e+07u w=2.5e+06u l=150000u
X2 VSUB a_1712_150# sky130_fd_pr__cap_mim_m3_1 l=6.2e+06u w=2.76e+07u
X3 a_1712_150# VSUB sky130_fd_pr__cap_mim_m3_2 l=6.2e+06u w=2.76e+07u
X4 a_1712_150# S a_1444_106# VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.6e+12p ps=1.128e+07u
+ w=2.5e+06u l=150000u
X5 VSUB VSUB a_1444_106# VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X6 a_1712_150# SBAR VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X7 a_1444_106# S a_1712_150# VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.5e+06u
+ l=150000u
C0 a_1712_150# imirror2_0/a_5868_1637# 0.33fF
C1 imirror2_0/OUT S 0.13fF
C2 imirror2_0/VHI imirror2_0/OUT 0.03fF
C3 imirror2_0/OUT imirror2_0/a_4493_207# 0.00fF
C4 a_1444_106# a_1712_150# 0.93fF
C5 SBAR a_1444_106# 0.07fF
C6 S a_1712_150# 0.27fF
C7 S SBAR 0.71fF
C8 imirror2_0/OUT a_1712_150# 1.57fF
C9 imirror2_0/VHI a_1712_150# 0.88fF
C10 imirror2_0/OUT SBAR 0.14fF
C11 a_1444_106# imirror2_0/IN 0.00fF
C12 S imirror2_0/IN 0.01fF
C13 a_1712_150# imirror2_0/a_4493_207# 0.29fF
C14 imirror2_0/OUT imirror2_0/IN 0.07fF
C15 imirror2_0/VHI imirror2_0/IN 0.00fF
C16 imirror2_0/OUT imirror2_0/a_5468_1540# 0.00fF
C17 SBAR a_1712_150# 0.25fF
C18 imirror2_0/a_4493_207# imirror2_0/IN 0.12fF
C19 a_1712_150# imirror2_0/IN 0.12fF
C20 SBAR imirror2_0/IN 0.01fF
C21 a_1712_150# imirror2_0/a_5468_1540# 0.33fF
C22 imirror2_0/OUT imirror2_0/a_5868_1637# 0.00fF
C23 S a_1444_106# 0.03fF
C24 imirror2_0/OUT a_1444_106# 0.33fF
C25 a_1712_150# VSUB 39.40fF
C26 a_1444_106# VSUB 1.29fF
C27 SBAR VSUB 0.76fF
C28 S VSUB 0.77fF
C29 imirror2_0/OUT VSUB 6.83fF
C30 imirror2_0/VHI VSUB 19.56fF
C31 imirror2_0/IN VSUB 4.59fF
C32 imirror2_0/a_5868_1637# VSUB 0.44fF
C33 imirror2_0/a_4036_1637# VSUB 0.34fF
C34 imirror2_0/a_5468_1540# VSUB 0.49fF
C35 imirror2_0/a_4493_207# VSUB 1.64fF
C36 imirror2_0/a_4094_1540# VSUB 0.34fF
C37 imirror2_0/OUT.t0 VSUB 1.25fF $ **FLOATING
C38 imirror2_0/VHI.n0 VSUB 0.25fF $ **FLOATING
C39 imirror2_0/VHI.n1 VSUB 2.09fF $ **FLOATING
C40 imirror2_0/VHI.t0 VSUB 3.29fF $ **FLOATING
C41 imirror2_0/VHI.t2 VSUB 2.82fF $ **FLOATING
C42 imirror2_0/VHI.n2 VSUB 0.25fF $ **FLOATING
C43 imirror2_0/VHI.n3 VSUB 2.09fF $ **FLOATING
C44 imirror2_0/VHI.t1 VSUB 3.29fF $ **FLOATING
C45 imirror2_0/VHI.t5 VSUB 2.82fF $ **FLOATING
C46 imirror2_0/VHI.n4 VSUB 0.25fF $ **FLOATING
C47 imirror2_0/VHI.n5 VSUB 0.25fF $ **FLOATING
C48 imirror2_0/VHI.n6 VSUB 1.88fF $ **FLOATING
C49 imirror2_0/VHI.n7 VSUB 0.25fF $ **FLOATING
C50 imirror2_0/VHI.n8 VSUB 0.13fF $ **FLOATING
C51 imirror2_0/VHI.n9 VSUB 2.08fF $ **FLOATING
.ends

.subckt sky130_fd_pr__res_high_po_0p69_G8QCSG a_48_n518# a_n186_n518# a_n316_n648#
X0 a_n186_n518# a_48_n518# a_n316_n648# sky130_fd_pr__res_high_po w=690000u l=5.83e+06u
C0 a_n186_n518# a_48_n518# 0.18fF
C1 a_48_n518# a_n316_n648# 0.52fF
C2 a_n186_n518# a_n316_n648# 0.52fF
.ends

.subckt cmota_gb_rp VREF COM VIP VIN DP li_5300_n960# VLO a_2217_285# DN VOP VMN VHI  a_2925_285#
Xsky130_fd_pr__res_high_po_0p69_G8QCSG_0 li_5300_n960# VMN VLO sky130_fd_pr__res_high_po_0p69_G8QCSG
X0 VHI DN VMN VHI sky130_fd_pr__pfet_01v8 ad=4.93e+13p pd=3.4986e+08u as=1.16e+13p ps=8.232e+07u
+ w=1e+07u l=300000u
X1 VHI DN DN VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+12p ps=6.174e+07u w=1e+07u l=300000u
X2 VHI DP VOP VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.16e+13p ps=8.232e+07u w=1e+07u l=300000u
X3 DN VIN COM VLO sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.264e+07u as=1.3225e+13p ps=9.21e+07u
+ w=2.5e+06u l=150000u
X4 COM VIN DN VLO sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X5 DP VIP COM VLO sky130_fd_pr__nfet_01v8_lvt ad=3.3e+12p pd=2.264e+07u as=0p ps=0u w=2.5e+06u
+ l=150000u
X6 VMN DN VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X7 VMN DN VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X8 VHI VHI VOP VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X9 a_2925_285# DN VHI VHI sky130_fd_pr__pfet_01v8 ad=2.9e+12p pd=2.058e+07u as=0p ps=0u w=1e+07u
+ l=300000u
X10 DP VIP COM VLO sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X11 li_5300_n960# VOP sky130_fd_pr__cap_mim_m3_2 l=1.32e+07u w=3.7e+06u
X12 VOP DP VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X13 VOP DP VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X14 VOP DP VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X15 COM VLO VLO VLO sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.8e+13p ps=2.69525e+08u w=2.5e+06u
+ l=150000u
X16 VLO VMN VOP VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+12p ps=4.116e+07u w=1e+07u l=300000u
X17 VHI DN VMN VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X18 VLO VLO VLO VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X19 VHI DN DP VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+12p ps=6.174e+07u w=1e+07u l=300000u
X20 VHI DP DP VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X21 COM VIP DP VLO sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X22 VLO VREF COM VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=2e+06u
X23 VMN VHI VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X24 DN DN VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X25 VHI DP VOP VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X26 VLO VLO VLO VLO sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X27 VLO VREF COM VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=2e+06u
X28 COM VIN DN VLO sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X29 DN DN VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X30 DP DN VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X31 DN DP VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X32 DP DP VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X33 DN VIN COM VLO sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X34 VLO VLO VLO VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X35 COM VIP DP VLO sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X36 VHI DN DN VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X37 VOP DP VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X38 VMN VMN VLO VLO sky130_fd_pr__nfet_01v8 ad=5.8e+12p pd=4.116e+07u as=0p ps=0u w=1e+07u l=300000u
X39 VLO VMN VMN VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X40 VLO VLO VLO VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X41 VOP VMN VLO VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X42 VHI DP DN VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X43 VLO VMN VOP VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X44 VHI DN VMN VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X45 VLO VLO COM VLO sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X46 DN VIN COM VLO sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X47 VHI DP a_2217_285# VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.9e+12p ps=2.058e+07u w=1e+07u
+ l=300000u
X48 VHI DP DP VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X49 VLO VLO VLO VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X50 COM VREF VLO VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=2e+06u
X51 VLO VLO VLO VLO sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X52 COM VIN DN VLO sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X53 COM VREF VLO VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=2e+06u
X54 DP VIP COM VLO sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X55 COM VIN DN VLO sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X56 VMN DN VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X57 DP DP VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X58 DP VIP COM VLO sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X59 a_2217_285# DP VHI VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X60 VMN VMN VLO VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X61 COM VIP DP VLO sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X62 VLO VMN VMN VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X63 VOP VMN VLO VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X64 COM VIP DP VLO sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X65 VHI DN VMN VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X66 DN VIN COM VLO sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=150000u
X67 VOP li_5300_n960# sky130_fd_pr__cap_mim_m3_1 l=1.32e+07u w=3.7e+06u
X68 VHI DN a_2925_285# VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
X69 VHI DP VOP VHI sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=300000u
C0 VOP VREF 0.03fF
C1 DN COM 6.05fF
C2 VOP VIP 0.01fF
C3 VMN VREF 0.10fF
C4 li_5300_n960# DP 0.48fF
C5 VOP a_2217_285# 0.01fF
C6 VMN VIP 0.14fF
C7 VHI a_2925_285# 4.31fF
C8 DN DP 1.21fF
C9 VHI VIN 0.11fF
C10 VMN a_2217_285# 0.06fF
C11 COM a_2925_285# 0.01fF
C12 VIN COM 0.71fF
C13 VHI VREF 0.04fF
C14 COM VREF 2.35fF
C15 VHI VIP 0.10fF
C16 DP a_2925_285# 0.17fF
C17 VHI a_2217_285# 4.31fF
C18 COM VIP 0.71fF
C19 VIN DP 0.04fF
C20 a_2217_285# COM 0.01fF
C21 DP VREF 0.14fF
C22 VIP DP 0.53fF
C23 a_2217_285# DP 0.13fF
C24 DN a_2925_285# 0.13fF
C25 DN VIN 0.53fF
C26 DN VREF 0.14fF
C27 DN VIP 0.05fF
C28 VMN VOP 0.72fF
C29 DN a_2217_285# 0.17fF
C30 VREF a_2925_285# 0.00fF
C31 VIN VREF 0.36fF
C32 VIP a_2925_285# 0.00fF
C33 VIN VIP 0.11fF
C34 VHI VOP 18.23fF
C35 a_2217_285# a_2925_285# 0.02fF
C36 a_2217_285# VIN 0.00fF
C37 VOP COM 0.05fF
C38 VIP VREF 0.36fF
C39 VHI VMN 17.75fF
C40 a_2217_285# VREF 0.00fF
C41 VMN COM 0.33fF
C42 VOP DP 0.97fF
C43 VMN DP 0.34fF
C44 VHI COM 0.10fF
C45 li_5300_n960# VOP 9.33fF
C46 VHI DP 16.22fF
C47 VMN li_5300_n960# 1.12fF
C48 DN VOP 0.06fF
C49 COM DP 6.02fF
C50 DN VMN 1.12fF
C51 VHI li_5300_n960# 2.02fF
C52 VOP a_2925_285# 0.05fF
C53 VHI DN 16.22fF
C54 VMN a_2925_285# 0.01fF
C55 VMN VIN 0.15fF
C56 VREF VLO 7.20fF
C57 COM VLO 6.11fF
C58 VIP VLO 0.78fF
C59 VIN VLO 0.79fF
C60 VOP VLO 9.34fF
C61 a_2925_285# VLO -0.04fF
C62 a_2217_285# VLO -0.04fF
C63 DP VLO 1.36fF
C64 DN VLO 1.42fF
C65 VHI VLO 35.14fF
C66 li_5300_n960# VLO 3.02fF
C67 VMN VLO 13.45fF
.ends

.subckt cmota_gb_rp_gp VHI VLO VREF VIP VIN VOP S SBAR
Xgated_iref_fix_0 gated_iref_fix_0/imirror2_0/a_5468_1540# gated_iref_fix_0/imirror2_0/a_4094_1540#
+  SBAR gated_iref_fix_0/a_1444_106# gated_iref_fix_0/imirror2_0/OUT
+ gated_iref_fix_0/imirror2_0/a_5868_1637#  VLO VHI gated_iref_fix_0/imirror2_0/a_4493_207# gated_iref_fix_0/imirror2_0/a_4036_1637#
+  VREF_GATED S VREF gated_iref_fix
Xcmota_gb_rp_0 VREF_GATED cmota_gb_rp_0/COM VIP VIN cmota_gb_rp_0/DP cmota_gb_rp_0/li_5300_n960#
+  VLO cmota_gb_rp_0/a_2217_285# cmota_gb_rp_0/DN VOP cmota_gb_rp_0/VMN VHI cmota_gb_rp_0/a_2925_285#
+  cmota_gb_rp
X0 VLO VHI sky130_fd_pr__cap_mim_m3_2 l=3.1e+07u w=1.3e+07u
X1 VHI VLO sky130_fd_pr__cap_mim_m3_1 l=3.1e+07u w=1.3e+07u
C0 cmota_gb_rp_0/VMN VIN -0.00fF
C1 VREF_GATED cmota_gb_rp_0/VMN 1.54fF
C2 cmota_gb_rp_0/DN VHI 0.89fF
C3 VIN VIP 0.00fF
C4 VREF gated_iref_fix_0/a_1444_106# 0.00fF
C5 VREF S 0.03fF
C6 VREF gated_iref_fix_0/imirror2_0/OUT 0.00fF
C7 VREF_GATED VREF -0.04fF
C8 gated_iref_fix_0/imirror2_0/a_5868_1637# VHI 0.03fF
C9 VOP cmota_gb_rp_0/VMN 0.00fF
C10 VHI gated_iref_fix_0/a_1444_106# 0.00fF
C11 VREF_GATED gated_iref_fix_0/imirror2_0/a_5468_1540# -0.31fF
C12 cmota_gb_rp_0/a_2925_285# VHI 0.04fF
C13 VHI S 0.00fF
C14 cmota_gb_rp_0/DP VHI 0.81fF
C15 VIN cmota_gb_rp_0/COM -0.00fF
C16 VHI gated_iref_fix_0/imirror2_0/OUT 0.17fF
C17 VREF_GATED cmota_gb_rp_0/COM 0.17fF
C18 VREF_GATED cmota_gb_rp_0/DN 0.40fF
C19 VREF_GATED VHI 3.68fF
C20 VREF SBAR 0.02fF
C21 VOP cmota_gb_rp_0/li_5300_n960# 0.00fF
C22 VREF_GATED gated_iref_fix_0/imirror2_0/a_5868_1637# -0.07fF
C23 gated_iref_fix_0/imirror2_0/a_4036_1637# VHI 0.07fF
C24 VREF_GATED gated_iref_fix_0/a_1444_106# 0.00fF
C25 VOP VHI 0.11fF
C26 gated_iref_fix_0/imirror2_0/a_4493_207# VHI 0.19fF
C27 gated_iref_fix_0/imirror2_0/OUT S 0.00fF
C28 VHI SBAR 0.00fF
C29 cmota_gb_rp_0/VMN cmota_gb_rp_0/COM -0.00fF
C30 VREF_GATED S 0.00fF
C31 VHI cmota_gb_rp_0/VMN 0.15fF
C32 VREF_GATED gated_iref_fix_0/imirror2_0/OUT -0.37fF
C33 VREF_GATED VIN 0.00fF
C34 SBAR gated_iref_fix_0/a_1444_106# 0.00fF
C35 VREF VHI 0.16fF
C36 S SBAR 0.10fF
C37 cmota_gb_rp_0/DP VOP -0.00fF
C38 gated_iref_fix_0/imirror2_0/a_5468_1540# VHI 0.00fF
C39 gated_iref_fix_0/imirror2_0/OUT SBAR 0.00fF
C40 VHI cmota_gb_rp_0/li_5300_n960# 0.03fF
C41 VREF_GATED gated_iref_fix_0/imirror2_0/a_4493_207# -0.29fF
C42 VREF_GATED SBAR 0.02fF
C43 cmota_gb_rp_0/a_2217_285# VHI 0.04fF
C44 gated_iref_fix_0/imirror2_0/a_4094_1540# VHI 0.01fF
C45 VREF_GATED VLO 52.16fF
C46 cmota_gb_rp_0/COM VLO 6.15fF
C47 VIP VLO 0.78fF
C48 VIN VLO 0.79fF
C49 VOP VLO 9.31fF
C50 cmota_gb_rp_0/a_2925_285# VLO -0.04fF
C51 cmota_gb_rp_0/a_2217_285# VLO -0.04fF
C52 cmota_gb_rp_0/DP VLO 1.36fF
C53 cmota_gb_rp_0/DN VLO 1.55fF
C54 cmota_gb_rp_0/li_5300_n960# VLO 2.88fF
C55 cmota_gb_rp_0/VMN VLO 14.06fF
C56 gated_iref_fix_0/a_1444_106# VLO 1.29fF
C57 SBAR VLO 0.76fF
C58 S VLO 0.78fF
C59 gated_iref_fix_0/imirror2_0/OUT VLO 8.38fF
C60 VHI VLO 134.49fF
C61 VREF VLO 6.75fF
C62 gated_iref_fix_0/imirror2_0/a_5868_1637# VLO 0.48fF
C63 gated_iref_fix_0/imirror2_0/a_4036_1637# VLO 0.88fF
C64 gated_iref_fix_0/imirror2_0/a_5468_1540# VLO 0.63fF
C65 gated_iref_fix_0/imirror2_0/a_4493_207# VLO 4.55fF
C66 gated_iref_fix_0/imirror2_0/a_4094_1540# VLO 0.94fF
C67 gated_iref_fix_0/imirror2_0/OUT.t0 VLO 1.25fF $ **FLOATING
C68 gated_iref_fix_0/imirror2_0/VHI.n0 VLO 0.25fF $ **FLOATING
C69 gated_iref_fix_0/imirror2_0/VHI.n1 VLO 2.09fF $ **FLOATING
C70 gated_iref_fix_0/imirror2_0/VHI.t0 VLO 3.29fF $ **FLOATING
C71 gated_iref_fix_0/imirror2_0/VHI.t2 VLO 2.82fF $ **FLOATING
C72 gated_iref_fix_0/imirror2_0/VHI.n2 VLO 0.25fF $ **FLOATING
C73 gated_iref_fix_0/imirror2_0/VHI.n3 VLO 2.09fF $ **FLOATING
C74 gated_iref_fix_0/imirror2_0/VHI.t1 VLO 3.29fF $ **FLOATING
C75 gated_iref_fix_0/imirror2_0/VHI.t5 VLO 2.82fF $ **FLOATING
C76 gated_iref_fix_0/imirror2_0/VHI.n4 VLO 0.25fF $ **FLOATING
C77 gated_iref_fix_0/imirror2_0/VHI.n5 VLO 0.25fF $ **FLOATING
C78 gated_iref_fix_0/imirror2_0/VHI.n6 VLO 1.88fF $ **FLOATING
C79 gated_iref_fix_0/imirror2_0/VHI.n7 VLO 0.25fF $ **FLOATING
C80 gated_iref_fix_0/imirror2_0/VHI.n8 VLO 0.13fF $ **FLOATING
C81 gated_iref_fix_0/imirror2_0/VHI.n9 VLO 2.08fF $ **FLOATING
.ends



XDUT vhi vlo vref vip vin vop s sbar cmota_gb_rp_gp


**** end user architecture code
.ends

.GLOBAL GND
.end
