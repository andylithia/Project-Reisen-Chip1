magic
tech sky130B
magscale 1 2
timestamp 1668466684
<< pwell >>
rect 30 -6050 390 -5410
<< nmos >>
rect 100 -5920 130 -5520
rect 196 -5920 226 -5520
rect 292 -5920 322 -5520
<< ndiff >>
rect 38 -5532 100 -5520
rect 38 -5908 50 -5532
rect 84 -5908 100 -5532
rect 38 -5920 100 -5908
rect 130 -5532 196 -5520
rect 130 -5908 146 -5532
rect 180 -5908 196 -5532
rect 130 -5920 196 -5908
rect 226 -5532 292 -5520
rect 226 -5908 242 -5532
rect 276 -5908 292 -5532
rect 226 -5920 292 -5908
rect 322 -5532 388 -5520
rect 322 -5908 338 -5532
rect 372 -5908 388 -5532
rect 322 -5920 388 -5908
<< ndiffc >>
rect 50 -5908 84 -5532
rect 146 -5908 180 -5532
rect 242 -5908 276 -5532
rect 338 -5908 372 -5532
<< poly >>
rect 100 -5448 226 -5432
rect 100 -5482 110 -5448
rect 215 -5482 226 -5448
rect 100 -5498 226 -5482
rect 100 -5520 130 -5498
rect 196 -5520 226 -5498
rect 292 -5520 322 -5494
rect 100 -5946 130 -5920
rect 196 -5946 226 -5920
rect 292 -5942 322 -5920
rect 274 -6008 340 -5942
<< polycont >>
rect 110 -5482 215 -5448
<< locali >>
rect 87 -5482 110 -5448
rect 240 -5482 254 -5448
rect 50 -5532 84 -5516
rect 50 -5924 84 -5908
rect 146 -5532 180 -5516
rect 146 -5924 180 -5908
rect 242 -5532 276 -5516
rect 242 -5924 276 -5908
rect 338 -5532 372 -5516
rect 338 -5924 372 -5908
<< viali >>
rect 110 -5482 215 -5448
rect 215 -5482 240 -5448
rect 50 -5908 84 -5532
rect 146 -5908 180 -5532
rect 242 -5908 276 -5532
rect 338 -5908 372 -5532
<< metal1 >>
rect 87 -5448 254 -5442
rect 87 -5482 110 -5448
rect 240 -5482 254 -5448
rect 87 -5488 254 -5482
rect 44 -5532 90 -5520
rect 44 -5908 50 -5532
rect 84 -5908 90 -5532
rect 44 -5920 90 -5908
rect 137 -5532 189 -5516
rect 137 -5924 189 -5910
rect 236 -5532 282 -5520
rect 236 -5908 242 -5532
rect 276 -5908 282 -5532
rect 236 -5920 282 -5908
rect 332 -5532 378 -5520
rect 332 -5908 338 -5532
rect 372 -5908 378 -5532
rect 332 -5920 378 -5908
<< via1 >>
rect 137 -5908 146 -5532
rect 146 -5908 180 -5532
rect 180 -5908 189 -5532
rect 137 -5910 189 -5908
<< metal2 >>
rect 134 -5532 191 -5516
rect 134 -5924 191 -5910
<< via2 >>
rect 134 -5910 137 -5532
rect 137 -5910 189 -5532
rect 189 -5910 191 -5532
<< metal3 >>
rect 129 -5532 197 -5516
rect 129 -5910 134 -5532
rect 191 -5910 197 -5532
rect 129 -5924 197 -5910
<< end >>
