magic
tech sky130A
magscale 1 2
timestamp 1670863210
<< viali >>
rect 1685 7497 1719 7531
rect 4077 7497 4111 7531
rect 5733 7497 5767 7531
rect 7941 7497 7975 7531
rect 12449 7497 12483 7531
rect 14657 7497 14691 7531
rect 17049 7497 17083 7531
rect 18245 7497 18279 7531
rect 9597 7429 9631 7463
rect 10149 7429 10183 7463
rect 1869 7361 1903 7395
rect 4261 7361 4295 7395
rect 5917 7361 5951 7395
rect 8125 7361 8159 7395
rect 12265 7361 12299 7395
rect 14473 7361 14507 7395
rect 16865 7361 16899 7395
rect 18061 7361 18095 7395
rect 10333 7225 10367 7259
rect 8033 6273 8067 6307
rect 8217 6273 8251 6307
rect 8401 6069 8435 6103
rect 8309 5865 8343 5899
rect 7757 5729 7791 5763
rect 6929 5661 6963 5695
rect 7941 5593 7975 5627
rect 11529 5593 11563 5627
rect 11713 5593 11747 5627
rect 12817 5593 12851 5627
rect 13001 5593 13035 5627
rect 6745 5525 6779 5559
rect 7849 5525 7883 5559
rect 11897 5525 11931 5559
rect 13185 5525 13219 5559
rect 4537 5321 4571 5355
rect 7021 5321 7055 5355
rect 7113 5321 7147 5355
rect 10425 5321 10459 5355
rect 11713 5321 11747 5355
rect 12173 5321 12207 5355
rect 13185 5321 13219 5355
rect 10333 5253 10367 5287
rect 12081 5253 12115 5287
rect 13277 5185 13311 5219
rect 2789 5117 2823 5151
rect 3065 5117 3099 5151
rect 7205 5117 7239 5151
rect 7849 5117 7883 5151
rect 8125 5117 8159 5151
rect 10149 5117 10183 5151
rect 12265 5117 12299 5151
rect 13093 5117 13127 5151
rect 6653 4981 6687 5015
rect 9597 4981 9631 5015
rect 10793 4981 10827 5015
rect 13645 4981 13679 5015
rect 7205 4777 7239 4811
rect 12725 4777 12759 4811
rect 7849 4709 7883 4743
rect 11529 4709 11563 4743
rect 8401 4641 8435 4675
rect 12081 4641 12115 4675
rect 12265 4641 12299 4675
rect 3065 4573 3099 4607
rect 4905 4573 4939 4607
rect 6377 4573 6411 4607
rect 6837 4573 6871 4607
rect 8309 4573 8343 4607
rect 9965 4573 9999 4607
rect 10517 4573 10551 4607
rect 11345 4573 11379 4607
rect 13369 4573 13403 4607
rect 15209 4573 15243 4607
rect 16221 4573 16255 4607
rect 16865 4573 16899 4607
rect 4353 4505 4387 4539
rect 6193 4505 6227 4539
rect 7021 4505 7055 4539
rect 9137 4505 9171 4539
rect 9321 4505 9355 4539
rect 10701 4505 10735 4539
rect 15393 4505 15427 4539
rect 15577 4505 15611 4539
rect 2421 4437 2455 4471
rect 4077 4437 4111 4471
rect 6009 4437 6043 4471
rect 8217 4437 8251 4471
rect 9505 4437 9539 4471
rect 10885 4437 10919 4471
rect 12357 4437 12391 4471
rect 13185 4437 13219 4471
rect 16037 4437 16071 4471
rect 16681 4437 16715 4471
rect 2421 4233 2455 4267
rect 8033 4233 8067 4267
rect 8401 4233 8435 4267
rect 11713 4233 11747 4267
rect 8955 4165 8989 4199
rect 2237 4097 2271 4131
rect 6837 4097 6871 4131
rect 2881 4029 2915 4063
rect 3157 4029 3191 4063
rect 7757 4029 7791 4063
rect 7941 4029 7975 4063
rect 13185 4029 13219 4063
rect 13461 4029 13495 4063
rect 13921 4029 13955 4063
rect 14197 4029 14231 4063
rect 5089 3961 5123 3995
rect 6653 3961 6687 3995
rect 4629 3893 4663 3927
rect 10241 3893 10275 3927
rect 15669 3893 15703 3927
rect 1948 3689 1982 3723
rect 4997 3689 5031 3723
rect 8493 3621 8527 3655
rect 9321 3621 9355 3655
rect 11161 3621 11195 3655
rect 11989 3621 12023 3655
rect 1685 3553 1719 3587
rect 13737 3553 13771 3587
rect 6285 3485 6319 3519
rect 6745 3485 6779 3519
rect 9137 3485 9171 3519
rect 10241 3485 10275 3519
rect 10977 3485 11011 3519
rect 7021 3417 7055 3451
rect 13461 3417 13495 3451
rect 3433 3349 3467 3383
rect 10057 3349 10091 3383
rect 1961 3145 1995 3179
rect 7205 3145 7239 3179
rect 3433 3077 3467 3111
rect 8689 3077 8723 3111
rect 9413 3077 9447 3111
rect 13185 3077 13219 3111
rect 3709 3009 3743 3043
rect 4169 3009 4203 3043
rect 4537 3009 4571 3043
rect 13921 3009 13955 3043
rect 5963 2941 5997 2975
rect 8953 2941 8987 2975
rect 13461 2941 13495 2975
rect 10701 2873 10735 2907
rect 11713 2873 11747 2907
rect 14105 2805 14139 2839
rect 3433 2601 3467 2635
rect 6009 2601 6043 2635
rect 9137 2601 9171 2635
rect 14289 2601 14323 2635
rect 11989 2533 12023 2567
rect 1685 2465 1719 2499
rect 4261 2465 4295 2499
rect 4537 2465 4571 2499
rect 10609 2465 10643 2499
rect 13461 2465 13495 2499
rect 13737 2465 13771 2499
rect 16037 2465 16071 2499
rect 10885 2397 10919 2431
rect 17509 2397 17543 2431
rect 1961 2329 1995 2363
rect 15761 2329 15795 2363
rect 17693 2261 17727 2295
<< metal1 >>
rect 1104 7642 19019 7664
rect 1104 7590 5388 7642
rect 5440 7590 5452 7642
rect 5504 7590 5516 7642
rect 5568 7590 5580 7642
rect 5632 7590 5644 7642
rect 5696 7590 9827 7642
rect 9879 7590 9891 7642
rect 9943 7590 9955 7642
rect 10007 7590 10019 7642
rect 10071 7590 10083 7642
rect 10135 7590 14266 7642
rect 14318 7590 14330 7642
rect 14382 7590 14394 7642
rect 14446 7590 14458 7642
rect 14510 7590 14522 7642
rect 14574 7590 18705 7642
rect 18757 7590 18769 7642
rect 18821 7590 18833 7642
rect 18885 7590 18897 7642
rect 18949 7590 18961 7642
rect 19013 7590 19019 7642
rect 1104 7568 19019 7590
rect 1118 7488 1124 7540
rect 1176 7528 1182 7540
rect 1673 7531 1731 7537
rect 1673 7528 1685 7531
rect 1176 7500 1685 7528
rect 1176 7488 1182 7500
rect 1673 7497 1685 7500
rect 1719 7497 1731 7531
rect 1673 7491 1731 7497
rect 3326 7488 3332 7540
rect 3384 7528 3390 7540
rect 4065 7531 4123 7537
rect 4065 7528 4077 7531
rect 3384 7500 4077 7528
rect 3384 7488 3390 7500
rect 4065 7497 4077 7500
rect 4111 7497 4123 7531
rect 5718 7528 5724 7540
rect 5679 7500 5724 7528
rect 4065 7491 4123 7497
rect 5718 7488 5724 7500
rect 5776 7488 5782 7540
rect 7926 7528 7932 7540
rect 7887 7500 7932 7528
rect 7926 7488 7932 7500
rect 7984 7488 7990 7540
rect 12434 7528 12440 7540
rect 12395 7500 12440 7528
rect 12434 7488 12440 7500
rect 12492 7488 12498 7540
rect 14642 7528 14648 7540
rect 14603 7500 14648 7528
rect 14642 7488 14648 7500
rect 14700 7488 14706 7540
rect 16574 7488 16580 7540
rect 16632 7528 16638 7540
rect 17037 7531 17095 7537
rect 17037 7528 17049 7531
rect 16632 7500 17049 7528
rect 16632 7488 16638 7500
rect 17037 7497 17049 7500
rect 17083 7497 17095 7531
rect 17037 7491 17095 7497
rect 18233 7531 18291 7537
rect 18233 7497 18245 7531
rect 18279 7528 18291 7531
rect 18414 7528 18420 7540
rect 18279 7500 18420 7528
rect 18279 7497 18291 7500
rect 18233 7491 18291 7497
rect 18414 7488 18420 7500
rect 18472 7488 18478 7540
rect 7282 7420 7288 7472
rect 7340 7460 7346 7472
rect 9585 7463 9643 7469
rect 7340 7432 8248 7460
rect 7340 7420 7346 7432
rect 1857 7395 1915 7401
rect 1857 7361 1869 7395
rect 1903 7361 1915 7395
rect 1857 7355 1915 7361
rect 4249 7395 4307 7401
rect 4249 7361 4261 7395
rect 4295 7361 4307 7395
rect 4249 7355 4307 7361
rect 5905 7395 5963 7401
rect 5905 7361 5917 7395
rect 5951 7392 5963 7395
rect 7006 7392 7012 7404
rect 5951 7364 7012 7392
rect 5951 7361 5963 7364
rect 5905 7355 5963 7361
rect 1872 7324 1900 7355
rect 4264 7324 4292 7355
rect 7006 7352 7012 7364
rect 7064 7352 7070 7404
rect 7466 7352 7472 7404
rect 7524 7392 7530 7404
rect 8113 7395 8171 7401
rect 8113 7392 8125 7395
rect 7524 7364 8125 7392
rect 7524 7352 7530 7364
rect 8113 7361 8125 7364
rect 8159 7361 8171 7395
rect 8220 7392 8248 7432
rect 9585 7429 9597 7463
rect 9631 7460 9643 7463
rect 10137 7463 10195 7469
rect 10137 7460 10149 7463
rect 9631 7432 10149 7460
rect 9631 7429 9643 7432
rect 9585 7423 9643 7429
rect 10137 7429 10149 7432
rect 10183 7460 10195 7463
rect 10226 7460 10232 7472
rect 10183 7432 10232 7460
rect 10183 7429 10195 7432
rect 10137 7423 10195 7429
rect 10226 7420 10232 7432
rect 10284 7420 10290 7472
rect 12253 7395 12311 7401
rect 12253 7392 12265 7395
rect 8220 7364 12265 7392
rect 8113 7355 8171 7361
rect 12253 7361 12265 7364
rect 12299 7361 12311 7395
rect 12253 7355 12311 7361
rect 13814 7352 13820 7404
rect 13872 7392 13878 7404
rect 14461 7395 14519 7401
rect 14461 7392 14473 7395
rect 13872 7364 14473 7392
rect 13872 7352 13878 7364
rect 14461 7361 14473 7364
rect 14507 7361 14519 7395
rect 16850 7392 16856 7404
rect 16811 7364 16856 7392
rect 14461 7355 14519 7361
rect 16850 7352 16856 7364
rect 16908 7352 16914 7404
rect 18049 7395 18107 7401
rect 18049 7361 18061 7395
rect 18095 7361 18107 7395
rect 18049 7355 18107 7361
rect 7926 7324 7932 7336
rect 1872 7296 2774 7324
rect 4264 7296 7932 7324
rect 2746 7188 2774 7296
rect 7926 7284 7932 7296
rect 7984 7284 7990 7336
rect 13354 7284 13360 7336
rect 13412 7324 13418 7336
rect 18064 7324 18092 7355
rect 13412 7296 18092 7324
rect 13412 7284 13418 7296
rect 10318 7256 10324 7268
rect 10279 7228 10324 7256
rect 10318 7216 10324 7228
rect 10376 7216 10382 7268
rect 11054 7188 11060 7200
rect 2746 7160 11060 7188
rect 11054 7148 11060 7160
rect 11112 7148 11118 7200
rect 1104 7098 18860 7120
rect 1104 7046 3169 7098
rect 3221 7046 3233 7098
rect 3285 7046 3297 7098
rect 3349 7046 3361 7098
rect 3413 7046 3425 7098
rect 3477 7046 7608 7098
rect 7660 7046 7672 7098
rect 7724 7046 7736 7098
rect 7788 7046 7800 7098
rect 7852 7046 7864 7098
rect 7916 7046 12047 7098
rect 12099 7046 12111 7098
rect 12163 7046 12175 7098
rect 12227 7046 12239 7098
rect 12291 7046 12303 7098
rect 12355 7046 16486 7098
rect 16538 7046 16550 7098
rect 16602 7046 16614 7098
rect 16666 7046 16678 7098
rect 16730 7046 16742 7098
rect 16794 7046 18860 7098
rect 1104 7024 18860 7046
rect 1104 6554 19019 6576
rect 1104 6502 5388 6554
rect 5440 6502 5452 6554
rect 5504 6502 5516 6554
rect 5568 6502 5580 6554
rect 5632 6502 5644 6554
rect 5696 6502 9827 6554
rect 9879 6502 9891 6554
rect 9943 6502 9955 6554
rect 10007 6502 10019 6554
rect 10071 6502 10083 6554
rect 10135 6502 14266 6554
rect 14318 6502 14330 6554
rect 14382 6502 14394 6554
rect 14446 6502 14458 6554
rect 14510 6502 14522 6554
rect 14574 6502 18705 6554
rect 18757 6502 18769 6554
rect 18821 6502 18833 6554
rect 18885 6502 18897 6554
rect 18949 6502 18961 6554
rect 19013 6502 19019 6554
rect 1104 6480 19019 6502
rect 8018 6304 8024 6316
rect 7979 6276 8024 6304
rect 8018 6264 8024 6276
rect 8076 6264 8082 6316
rect 8202 6304 8208 6316
rect 8163 6276 8208 6304
rect 8202 6264 8208 6276
rect 8260 6264 8266 6316
rect 8389 6103 8447 6109
rect 8389 6069 8401 6103
rect 8435 6100 8447 6103
rect 10962 6100 10968 6112
rect 8435 6072 10968 6100
rect 8435 6069 8447 6072
rect 8389 6063 8447 6069
rect 10962 6060 10968 6072
rect 11020 6060 11026 6112
rect 1104 6010 18860 6032
rect 1104 5958 3169 6010
rect 3221 5958 3233 6010
rect 3285 5958 3297 6010
rect 3349 5958 3361 6010
rect 3413 5958 3425 6010
rect 3477 5958 7608 6010
rect 7660 5958 7672 6010
rect 7724 5958 7736 6010
rect 7788 5958 7800 6010
rect 7852 5958 7864 6010
rect 7916 5958 12047 6010
rect 12099 5958 12111 6010
rect 12163 5958 12175 6010
rect 12227 5958 12239 6010
rect 12291 5958 12303 6010
rect 12355 5958 16486 6010
rect 16538 5958 16550 6010
rect 16602 5958 16614 6010
rect 16666 5958 16678 6010
rect 16730 5958 16742 6010
rect 16794 5958 18860 6010
rect 1104 5936 18860 5958
rect 8018 5856 8024 5908
rect 8076 5896 8082 5908
rect 8297 5899 8355 5905
rect 8297 5896 8309 5899
rect 8076 5868 8309 5896
rect 8076 5856 8082 5868
rect 8297 5865 8309 5868
rect 8343 5865 8355 5899
rect 8297 5859 8355 5865
rect 7745 5763 7803 5769
rect 7745 5729 7757 5763
rect 7791 5760 7803 5763
rect 8110 5760 8116 5772
rect 7791 5732 8116 5760
rect 7791 5729 7803 5732
rect 7745 5723 7803 5729
rect 8110 5720 8116 5732
rect 8168 5720 8174 5772
rect 6914 5692 6920 5704
rect 6875 5664 6920 5692
rect 6914 5652 6920 5664
rect 6972 5652 6978 5704
rect 7466 5584 7472 5636
rect 7524 5624 7530 5636
rect 7929 5627 7987 5633
rect 7929 5624 7941 5627
rect 7524 5596 7941 5624
rect 7524 5584 7530 5596
rect 7929 5593 7941 5596
rect 7975 5593 7987 5627
rect 11514 5624 11520 5636
rect 11475 5596 11520 5624
rect 7929 5587 7987 5593
rect 11514 5584 11520 5596
rect 11572 5584 11578 5636
rect 11698 5624 11704 5636
rect 11659 5596 11704 5624
rect 11698 5584 11704 5596
rect 11756 5584 11762 5636
rect 12802 5624 12808 5636
rect 12763 5596 12808 5624
rect 12802 5584 12808 5596
rect 12860 5584 12866 5636
rect 12894 5584 12900 5636
rect 12952 5624 12958 5636
rect 12989 5627 13047 5633
rect 12989 5624 13001 5627
rect 12952 5596 13001 5624
rect 12952 5584 12958 5596
rect 12989 5593 13001 5596
rect 13035 5593 13047 5627
rect 12989 5587 13047 5593
rect 4614 5516 4620 5568
rect 4672 5556 4678 5568
rect 6733 5559 6791 5565
rect 6733 5556 6745 5559
rect 4672 5528 6745 5556
rect 4672 5516 4678 5528
rect 6733 5525 6745 5528
rect 6779 5525 6791 5559
rect 6733 5519 6791 5525
rect 7374 5516 7380 5568
rect 7432 5556 7438 5568
rect 7837 5559 7895 5565
rect 7837 5556 7849 5559
rect 7432 5528 7849 5556
rect 7432 5516 7438 5528
rect 7837 5525 7849 5528
rect 7883 5525 7895 5559
rect 7837 5519 7895 5525
rect 11885 5559 11943 5565
rect 11885 5525 11897 5559
rect 11931 5556 11943 5559
rect 13078 5556 13084 5568
rect 11931 5528 13084 5556
rect 11931 5525 11943 5528
rect 11885 5519 11943 5525
rect 13078 5516 13084 5528
rect 13136 5516 13142 5568
rect 13173 5559 13231 5565
rect 13173 5525 13185 5559
rect 13219 5556 13231 5559
rect 15102 5556 15108 5568
rect 13219 5528 15108 5556
rect 13219 5525 13231 5528
rect 13173 5519 13231 5525
rect 15102 5516 15108 5528
rect 15160 5516 15166 5568
rect 1104 5466 19019 5488
rect 1104 5414 5388 5466
rect 5440 5414 5452 5466
rect 5504 5414 5516 5466
rect 5568 5414 5580 5466
rect 5632 5414 5644 5466
rect 5696 5414 9827 5466
rect 9879 5414 9891 5466
rect 9943 5414 9955 5466
rect 10007 5414 10019 5466
rect 10071 5414 10083 5466
rect 10135 5414 14266 5466
rect 14318 5414 14330 5466
rect 14382 5414 14394 5466
rect 14446 5414 14458 5466
rect 14510 5414 14522 5466
rect 14574 5414 18705 5466
rect 18757 5414 18769 5466
rect 18821 5414 18833 5466
rect 18885 5414 18897 5466
rect 18949 5414 18961 5466
rect 19013 5414 19019 5466
rect 1104 5392 19019 5414
rect 4525 5355 4583 5361
rect 4525 5321 4537 5355
rect 4571 5321 4583 5355
rect 7006 5352 7012 5364
rect 6967 5324 7012 5352
rect 4525 5315 4583 5321
rect 4430 5284 4436 5296
rect 4278 5256 4436 5284
rect 4430 5244 4436 5256
rect 4488 5244 4494 5296
rect 4540 5284 4568 5315
rect 7006 5312 7012 5324
rect 7064 5312 7070 5364
rect 7101 5355 7159 5361
rect 7101 5321 7113 5355
rect 7147 5352 7159 5355
rect 7374 5352 7380 5364
rect 7147 5324 7380 5352
rect 7147 5321 7159 5324
rect 7101 5315 7159 5321
rect 7374 5312 7380 5324
rect 7432 5312 7438 5364
rect 10413 5355 10471 5361
rect 8496 5324 9720 5352
rect 8496 5284 8524 5324
rect 4540 5256 8524 5284
rect 6730 5176 6736 5228
rect 6788 5216 6794 5228
rect 6788 5188 7880 5216
rect 6788 5176 6794 5188
rect 2777 5151 2835 5157
rect 2777 5117 2789 5151
rect 2823 5148 2835 5151
rect 3050 5148 3056 5160
rect 2823 5120 2912 5148
rect 3011 5120 3056 5148
rect 2823 5117 2835 5120
rect 2777 5111 2835 5117
rect 2884 5012 2912 5120
rect 3050 5108 3056 5120
rect 3108 5108 3114 5160
rect 7852 5157 7880 5188
rect 9214 5176 9220 5228
rect 9272 5176 9278 5228
rect 9692 5216 9720 5324
rect 10413 5321 10425 5355
rect 10459 5352 10471 5355
rect 11054 5352 11060 5364
rect 10459 5324 11060 5352
rect 10459 5321 10471 5324
rect 10413 5315 10471 5321
rect 11054 5312 11060 5324
rect 11112 5312 11118 5364
rect 11514 5312 11520 5364
rect 11572 5352 11578 5364
rect 11701 5355 11759 5361
rect 11701 5352 11713 5355
rect 11572 5324 11713 5352
rect 11572 5312 11578 5324
rect 11701 5321 11713 5324
rect 11747 5321 11759 5355
rect 12161 5355 12219 5361
rect 12161 5352 12173 5355
rect 11701 5315 11759 5321
rect 11808 5324 12173 5352
rect 10318 5284 10324 5296
rect 10231 5256 10324 5284
rect 10318 5244 10324 5256
rect 10376 5284 10382 5296
rect 11808 5284 11836 5324
rect 12161 5321 12173 5324
rect 12207 5352 12219 5355
rect 12434 5352 12440 5364
rect 12207 5324 12440 5352
rect 12207 5321 12219 5324
rect 12161 5315 12219 5321
rect 12434 5312 12440 5324
rect 12492 5352 12498 5364
rect 13173 5355 13231 5361
rect 13173 5352 13185 5355
rect 12492 5324 13185 5352
rect 12492 5312 12498 5324
rect 13173 5321 13185 5324
rect 13219 5321 13231 5355
rect 13173 5315 13231 5321
rect 10376 5256 11836 5284
rect 12069 5287 12127 5293
rect 10376 5244 10382 5256
rect 12069 5253 12081 5287
rect 12115 5253 12127 5287
rect 13814 5284 13820 5296
rect 12069 5247 12127 5253
rect 12406 5256 13820 5284
rect 12084 5216 12112 5247
rect 12406 5216 12434 5256
rect 13814 5244 13820 5256
rect 13872 5244 13878 5296
rect 9692 5188 12434 5216
rect 12986 5176 12992 5228
rect 13044 5216 13050 5228
rect 13265 5219 13323 5225
rect 13265 5216 13277 5219
rect 13044 5188 13277 5216
rect 13044 5176 13050 5188
rect 13265 5185 13277 5188
rect 13311 5216 13323 5219
rect 13354 5216 13360 5228
rect 13311 5188 13360 5216
rect 13311 5185 13323 5188
rect 13265 5179 13323 5185
rect 13354 5176 13360 5188
rect 13412 5176 13418 5228
rect 7193 5151 7251 5157
rect 7193 5117 7205 5151
rect 7239 5117 7251 5151
rect 7193 5111 7251 5117
rect 7837 5151 7895 5157
rect 7837 5117 7849 5151
rect 7883 5117 7895 5151
rect 8110 5148 8116 5160
rect 8071 5120 8116 5148
rect 7837 5111 7895 5117
rect 4246 5040 4252 5092
rect 4304 5080 4310 5092
rect 7208 5080 7236 5111
rect 8110 5108 8116 5120
rect 8168 5108 8174 5160
rect 9674 5108 9680 5160
rect 9732 5148 9738 5160
rect 10137 5151 10195 5157
rect 10137 5148 10149 5151
rect 9732 5120 10149 5148
rect 9732 5108 9738 5120
rect 10137 5117 10149 5120
rect 10183 5117 10195 5151
rect 10137 5111 10195 5117
rect 4304 5052 7236 5080
rect 10152 5080 10180 5111
rect 11882 5108 11888 5160
rect 11940 5148 11946 5160
rect 12253 5151 12311 5157
rect 12253 5148 12265 5151
rect 11940 5120 12265 5148
rect 11940 5108 11946 5120
rect 12253 5117 12265 5120
rect 12299 5117 12311 5151
rect 12253 5111 12311 5117
rect 12894 5108 12900 5160
rect 12952 5148 12958 5160
rect 13081 5151 13139 5157
rect 13081 5148 13093 5151
rect 12952 5120 13093 5148
rect 12952 5108 12958 5120
rect 13081 5117 13093 5120
rect 13127 5117 13139 5151
rect 13081 5111 13139 5117
rect 13906 5080 13912 5092
rect 10152 5052 13912 5080
rect 4304 5040 4310 5052
rect 4154 5012 4160 5024
rect 2884 4984 4160 5012
rect 4154 4972 4160 4984
rect 4212 4972 4218 5024
rect 6641 5015 6699 5021
rect 6641 4981 6653 5015
rect 6687 5012 6699 5015
rect 6822 5012 6828 5024
rect 6687 4984 6828 5012
rect 6687 4981 6699 4984
rect 6641 4975 6699 4981
rect 6822 4972 6828 4984
rect 6880 4972 6886 5024
rect 7208 5012 7236 5052
rect 13906 5040 13912 5052
rect 13964 5040 13970 5092
rect 9306 5012 9312 5024
rect 7208 4984 9312 5012
rect 9306 4972 9312 4984
rect 9364 5012 9370 5024
rect 9585 5015 9643 5021
rect 9585 5012 9597 5015
rect 9364 4984 9597 5012
rect 9364 4972 9370 4984
rect 9585 4981 9597 4984
rect 9631 4981 9643 5015
rect 9585 4975 9643 4981
rect 10502 4972 10508 5024
rect 10560 5012 10566 5024
rect 10781 5015 10839 5021
rect 10781 5012 10793 5015
rect 10560 4984 10793 5012
rect 10560 4972 10566 4984
rect 10781 4981 10793 4984
rect 10827 4981 10839 5015
rect 10781 4975 10839 4981
rect 13633 5015 13691 5021
rect 13633 4981 13645 5015
rect 13679 5012 13691 5015
rect 15194 5012 15200 5024
rect 13679 4984 15200 5012
rect 13679 4981 13691 4984
rect 13633 4975 13691 4981
rect 15194 4972 15200 4984
rect 15252 4972 15258 5024
rect 1104 4922 18860 4944
rect 1104 4870 3169 4922
rect 3221 4870 3233 4922
rect 3285 4870 3297 4922
rect 3349 4870 3361 4922
rect 3413 4870 3425 4922
rect 3477 4870 7608 4922
rect 7660 4870 7672 4922
rect 7724 4870 7736 4922
rect 7788 4870 7800 4922
rect 7852 4870 7864 4922
rect 7916 4870 12047 4922
rect 12099 4870 12111 4922
rect 12163 4870 12175 4922
rect 12227 4870 12239 4922
rect 12291 4870 12303 4922
rect 12355 4870 16486 4922
rect 16538 4870 16550 4922
rect 16602 4870 16614 4922
rect 16666 4870 16678 4922
rect 16730 4870 16742 4922
rect 16794 4870 18860 4922
rect 1104 4848 18860 4870
rect 6914 4768 6920 4820
rect 6972 4808 6978 4820
rect 7193 4811 7251 4817
rect 7193 4808 7205 4811
rect 6972 4780 7205 4808
rect 6972 4768 6978 4780
rect 7193 4777 7205 4780
rect 7239 4777 7251 4811
rect 12713 4811 12771 4817
rect 7193 4771 7251 4777
rect 7760 4780 12204 4808
rect 3050 4700 3056 4752
rect 3108 4740 3114 4752
rect 7760 4740 7788 4780
rect 3108 4712 7788 4740
rect 7837 4743 7895 4749
rect 3108 4700 3114 4712
rect 7837 4709 7849 4743
rect 7883 4709 7895 4743
rect 7837 4703 7895 4709
rect 7852 4672 7880 4703
rect 8294 4700 8300 4752
rect 8352 4740 8358 4752
rect 11517 4743 11575 4749
rect 8352 4712 10824 4740
rect 8352 4700 8358 4712
rect 6380 4644 7880 4672
rect 2774 4564 2780 4616
rect 2832 4604 2838 4616
rect 6380 4613 6408 4644
rect 8018 4632 8024 4684
rect 8076 4672 8082 4684
rect 8202 4672 8208 4684
rect 8076 4644 8208 4672
rect 8076 4632 8082 4644
rect 8202 4632 8208 4644
rect 8260 4672 8266 4684
rect 8389 4675 8447 4681
rect 8389 4672 8401 4675
rect 8260 4644 8401 4672
rect 8260 4632 8266 4644
rect 8389 4641 8401 4644
rect 8435 4641 8447 4675
rect 10318 4672 10324 4684
rect 8389 4635 8447 4641
rect 8496 4644 10324 4672
rect 3053 4607 3111 4613
rect 3053 4604 3065 4607
rect 2832 4576 3065 4604
rect 2832 4564 2838 4576
rect 3053 4573 3065 4576
rect 3099 4604 3111 4607
rect 4893 4607 4951 4613
rect 4893 4604 4905 4607
rect 3099 4576 4905 4604
rect 3099 4573 3111 4576
rect 3053 4567 3111 4573
rect 4893 4573 4905 4576
rect 4939 4573 4951 4607
rect 4893 4567 4951 4573
rect 6365 4607 6423 4613
rect 6365 4573 6377 4607
rect 6411 4573 6423 4607
rect 6822 4604 6828 4616
rect 6783 4576 6828 4604
rect 6365 4567 6423 4573
rect 6822 4564 6828 4576
rect 6880 4564 6886 4616
rect 7374 4564 7380 4616
rect 7432 4604 7438 4616
rect 7834 4604 7840 4616
rect 7432 4576 7840 4604
rect 7432 4564 7438 4576
rect 7834 4564 7840 4576
rect 7892 4604 7898 4616
rect 8297 4607 8355 4613
rect 8297 4604 8309 4607
rect 7892 4576 8309 4604
rect 7892 4564 7898 4576
rect 8297 4573 8309 4576
rect 8343 4604 8355 4607
rect 8496 4604 8524 4644
rect 10318 4632 10324 4644
rect 10376 4632 10382 4684
rect 8343 4576 8524 4604
rect 8343 4573 8355 4576
rect 8297 4567 8355 4573
rect 9030 4564 9036 4616
rect 9088 4604 9094 4616
rect 9582 4604 9588 4616
rect 9088 4576 9588 4604
rect 9088 4564 9094 4576
rect 9582 4564 9588 4576
rect 9640 4604 9646 4616
rect 9953 4607 10011 4613
rect 9953 4604 9965 4607
rect 9640 4576 9965 4604
rect 9640 4564 9646 4576
rect 9953 4573 9965 4576
rect 9999 4573 10011 4607
rect 10502 4604 10508 4616
rect 10463 4576 10508 4604
rect 9953 4567 10011 4573
rect 10502 4564 10508 4576
rect 10560 4564 10566 4616
rect 4341 4539 4399 4545
rect 4341 4505 4353 4539
rect 4387 4536 4399 4539
rect 4982 4536 4988 4548
rect 4387 4508 4988 4536
rect 4387 4505 4399 4508
rect 4341 4499 4399 4505
rect 4982 4496 4988 4508
rect 5040 4496 5046 4548
rect 6178 4536 6184 4548
rect 6139 4508 6184 4536
rect 6178 4496 6184 4508
rect 6236 4496 6242 4548
rect 7009 4539 7067 4545
rect 7009 4505 7021 4539
rect 7055 4536 7067 4539
rect 8110 4536 8116 4548
rect 7055 4508 8116 4536
rect 7055 4505 7067 4508
rect 7009 4499 7067 4505
rect 8110 4496 8116 4508
rect 8168 4496 8174 4548
rect 8386 4496 8392 4548
rect 8444 4536 8450 4548
rect 9125 4539 9183 4545
rect 9125 4536 9137 4539
rect 8444 4508 9137 4536
rect 8444 4496 8450 4508
rect 9125 4505 9137 4508
rect 9171 4505 9183 4539
rect 9306 4536 9312 4548
rect 9267 4508 9312 4536
rect 9125 4499 9183 4505
rect 9306 4496 9312 4508
rect 9364 4496 9370 4548
rect 10686 4536 10692 4548
rect 10647 4508 10692 4536
rect 10686 4496 10692 4508
rect 10744 4496 10750 4548
rect 10796 4536 10824 4712
rect 11517 4709 11529 4743
rect 11563 4740 11575 4743
rect 11974 4740 11980 4752
rect 11563 4712 11980 4740
rect 11563 4709 11575 4712
rect 11517 4703 11575 4709
rect 11974 4700 11980 4712
rect 12032 4700 12038 4752
rect 11698 4632 11704 4684
rect 11756 4672 11762 4684
rect 12069 4675 12127 4681
rect 12069 4672 12081 4675
rect 11756 4644 12081 4672
rect 11756 4632 11762 4644
rect 12069 4641 12081 4644
rect 12115 4641 12127 4675
rect 12069 4635 12127 4641
rect 10962 4564 10968 4616
rect 11020 4604 11026 4616
rect 11333 4607 11391 4613
rect 11333 4604 11345 4607
rect 11020 4576 11345 4604
rect 11020 4564 11026 4576
rect 11333 4573 11345 4576
rect 11379 4573 11391 4607
rect 11333 4567 11391 4573
rect 11882 4536 11888 4548
rect 10796 4508 11888 4536
rect 11882 4496 11888 4508
rect 11940 4496 11946 4548
rect 12176 4536 12204 4780
rect 12713 4777 12725 4811
rect 12759 4808 12771 4811
rect 12802 4808 12808 4820
rect 12759 4780 12808 4808
rect 12759 4777 12771 4780
rect 12713 4771 12771 4777
rect 12802 4768 12808 4780
rect 12860 4768 12866 4820
rect 12342 4700 12348 4752
rect 12400 4740 12406 4752
rect 13722 4740 13728 4752
rect 12400 4712 13728 4740
rect 12400 4700 12406 4712
rect 13722 4700 13728 4712
rect 13780 4700 13786 4752
rect 16850 4740 16856 4752
rect 13832 4712 16856 4740
rect 12253 4675 12311 4681
rect 12253 4641 12265 4675
rect 12299 4672 12311 4675
rect 12434 4672 12440 4684
rect 12299 4644 12440 4672
rect 12299 4641 12311 4644
rect 12253 4635 12311 4641
rect 12434 4632 12440 4644
rect 12492 4632 12498 4684
rect 13832 4672 13860 4712
rect 16850 4700 16856 4712
rect 16908 4700 16914 4752
rect 13004 4644 13860 4672
rect 12342 4564 12348 4616
rect 12400 4604 12406 4616
rect 13004 4604 13032 4644
rect 15102 4632 15108 4684
rect 15160 4672 15166 4684
rect 15160 4644 16252 4672
rect 15160 4632 15166 4644
rect 12400 4576 13032 4604
rect 12400 4564 12406 4576
rect 13078 4564 13084 4616
rect 13136 4604 13142 4616
rect 13357 4607 13415 4613
rect 13357 4604 13369 4607
rect 13136 4576 13369 4604
rect 13136 4564 13142 4576
rect 13357 4573 13369 4576
rect 13403 4573 13415 4607
rect 15194 4604 15200 4616
rect 15155 4576 15200 4604
rect 13357 4567 13415 4573
rect 15194 4564 15200 4576
rect 15252 4564 15258 4616
rect 16224 4613 16252 4644
rect 16209 4607 16267 4613
rect 16209 4573 16221 4607
rect 16255 4573 16267 4607
rect 16853 4607 16911 4613
rect 16853 4604 16865 4607
rect 16209 4567 16267 4573
rect 16546 4576 16865 4604
rect 15378 4536 15384 4548
rect 12176 4508 13216 4536
rect 15339 4508 15384 4536
rect 2222 4428 2228 4480
rect 2280 4468 2286 4480
rect 2409 4471 2467 4477
rect 2409 4468 2421 4471
rect 2280 4440 2421 4468
rect 2280 4428 2286 4440
rect 2409 4437 2421 4440
rect 2455 4437 2467 4471
rect 2409 4431 2467 4437
rect 4065 4471 4123 4477
rect 4065 4437 4077 4471
rect 4111 4468 4123 4471
rect 4430 4468 4436 4480
rect 4111 4440 4436 4468
rect 4111 4437 4123 4440
rect 4065 4431 4123 4437
rect 4430 4428 4436 4440
rect 4488 4428 4494 4480
rect 5997 4471 6055 4477
rect 5997 4437 6009 4471
rect 6043 4468 6055 4471
rect 6822 4468 6828 4480
rect 6043 4440 6828 4468
rect 6043 4437 6055 4440
rect 5997 4431 6055 4437
rect 6822 4428 6828 4440
rect 6880 4428 6886 4480
rect 7282 4428 7288 4480
rect 7340 4468 7346 4480
rect 8205 4471 8263 4477
rect 8205 4468 8217 4471
rect 7340 4440 8217 4468
rect 7340 4428 7346 4440
rect 8205 4437 8217 4440
rect 8251 4437 8263 4471
rect 8205 4431 8263 4437
rect 8846 4428 8852 4480
rect 8904 4468 8910 4480
rect 9398 4468 9404 4480
rect 8904 4440 9404 4468
rect 8904 4428 8910 4440
rect 9398 4428 9404 4440
rect 9456 4428 9462 4480
rect 9493 4471 9551 4477
rect 9493 4437 9505 4471
rect 9539 4468 9551 4471
rect 10226 4468 10232 4480
rect 9539 4440 10232 4468
rect 9539 4437 9551 4440
rect 9493 4431 9551 4437
rect 10226 4428 10232 4440
rect 10284 4428 10290 4480
rect 10873 4471 10931 4477
rect 10873 4437 10885 4471
rect 10919 4468 10931 4471
rect 10962 4468 10968 4480
rect 10919 4440 10968 4468
rect 10919 4437 10931 4440
rect 10873 4431 10931 4437
rect 10962 4428 10968 4440
rect 11020 4428 11026 4480
rect 11054 4428 11060 4480
rect 11112 4468 11118 4480
rect 12342 4468 12348 4480
rect 11112 4440 12348 4468
rect 11112 4428 11118 4440
rect 12342 4428 12348 4440
rect 12400 4428 12406 4480
rect 13188 4477 13216 4508
rect 15378 4496 15384 4508
rect 15436 4496 15442 4548
rect 15565 4539 15623 4545
rect 15565 4505 15577 4539
rect 15611 4536 15623 4539
rect 16546 4536 16574 4576
rect 16853 4573 16865 4576
rect 16899 4573 16911 4607
rect 16853 4567 16911 4573
rect 15611 4508 16574 4536
rect 15611 4505 15623 4508
rect 15565 4499 15623 4505
rect 13173 4471 13231 4477
rect 13173 4437 13185 4471
rect 13219 4437 13231 4471
rect 16022 4468 16028 4480
rect 15983 4440 16028 4468
rect 13173 4431 13231 4437
rect 16022 4428 16028 4440
rect 16080 4428 16086 4480
rect 16669 4471 16727 4477
rect 16669 4437 16681 4471
rect 16715 4468 16727 4471
rect 16850 4468 16856 4480
rect 16715 4440 16856 4468
rect 16715 4437 16727 4440
rect 16669 4431 16727 4437
rect 16850 4428 16856 4440
rect 16908 4428 16914 4480
rect 1104 4378 19019 4400
rect 1104 4326 5388 4378
rect 5440 4326 5452 4378
rect 5504 4326 5516 4378
rect 5568 4326 5580 4378
rect 5632 4326 5644 4378
rect 5696 4326 9827 4378
rect 9879 4326 9891 4378
rect 9943 4326 9955 4378
rect 10007 4326 10019 4378
rect 10071 4326 10083 4378
rect 10135 4326 14266 4378
rect 14318 4326 14330 4378
rect 14382 4326 14394 4378
rect 14446 4326 14458 4378
rect 14510 4326 14522 4378
rect 14574 4326 18705 4378
rect 18757 4326 18769 4378
rect 18821 4326 18833 4378
rect 18885 4326 18897 4378
rect 18949 4326 18961 4378
rect 19013 4326 19019 4378
rect 1104 4304 19019 4326
rect 2409 4267 2467 4273
rect 2409 4233 2421 4267
rect 2455 4264 2467 4267
rect 4982 4264 4988 4276
rect 2455 4236 4988 4264
rect 2455 4233 2467 4236
rect 2409 4227 2467 4233
rect 4982 4224 4988 4236
rect 5040 4224 5046 4276
rect 6178 4224 6184 4276
rect 6236 4264 6242 4276
rect 6236 4236 7880 4264
rect 6236 4224 6242 4236
rect 4430 4196 4436 4208
rect 4343 4168 4436 4196
rect 4430 4156 4436 4168
rect 4488 4196 4494 4208
rect 5258 4196 5264 4208
rect 4488 4168 5264 4196
rect 4488 4156 4494 4168
rect 5258 4156 5264 4168
rect 5316 4156 5322 4208
rect 7282 4196 7288 4208
rect 6656 4168 7288 4196
rect 2222 4128 2228 4140
rect 2183 4100 2228 4128
rect 2222 4088 2228 4100
rect 2280 4088 2286 4140
rect 4706 4088 4712 4140
rect 4764 4128 4770 4140
rect 6656 4128 6684 4168
rect 7282 4156 7288 4168
rect 7340 4156 7346 4208
rect 7852 4196 7880 4236
rect 7926 4224 7932 4276
rect 7984 4264 7990 4276
rect 8021 4267 8079 4273
rect 8021 4264 8033 4267
rect 7984 4236 8033 4264
rect 7984 4224 7990 4236
rect 8021 4233 8033 4236
rect 8067 4233 8079 4267
rect 8386 4264 8392 4276
rect 8347 4236 8392 4264
rect 8021 4227 8079 4233
rect 8386 4224 8392 4236
rect 8444 4224 8450 4276
rect 9030 4264 9036 4276
rect 8956 4236 9036 4264
rect 8846 4196 8852 4208
rect 7852 4168 8852 4196
rect 8846 4156 8852 4168
rect 8904 4156 8910 4208
rect 8956 4205 8984 4236
rect 9030 4224 9036 4236
rect 9088 4224 9094 4276
rect 11146 4224 11152 4276
rect 11204 4264 11210 4276
rect 11701 4267 11759 4273
rect 11701 4264 11713 4267
rect 11204 4236 11713 4264
rect 11204 4224 11210 4236
rect 11701 4233 11713 4236
rect 11747 4233 11759 4267
rect 11701 4227 11759 4233
rect 11882 4224 11888 4276
rect 11940 4264 11946 4276
rect 11940 4236 12848 4264
rect 11940 4224 11946 4236
rect 8943 4199 9001 4205
rect 8943 4165 8955 4199
rect 8989 4165 9001 4199
rect 8943 4159 9001 4165
rect 9398 4156 9404 4208
rect 9456 4196 9462 4208
rect 11790 4196 11796 4208
rect 9456 4168 11796 4196
rect 9456 4156 9462 4168
rect 11790 4156 11796 4168
rect 11848 4156 11854 4208
rect 12820 4196 12848 4236
rect 12742 4168 14674 4196
rect 6822 4128 6828 4140
rect 4764 4100 6684 4128
rect 6783 4100 6828 4128
rect 4764 4088 4770 4100
rect 6822 4088 6828 4100
rect 6880 4088 6886 4140
rect 7466 4088 7472 4140
rect 7524 4128 7530 4140
rect 11882 4128 11888 4140
rect 7524 4100 11888 4128
rect 7524 4088 7530 4100
rect 11882 4088 11888 4100
rect 11940 4088 11946 4140
rect 2869 4063 2927 4069
rect 2869 4029 2881 4063
rect 2915 4029 2927 4063
rect 2869 4023 2927 4029
rect 3145 4063 3203 4069
rect 3145 4029 3157 4063
rect 3191 4060 3203 4063
rect 3191 4032 6684 4060
rect 3191 4029 3203 4032
rect 3145 4023 3203 4029
rect 2498 3884 2504 3936
rect 2556 3924 2562 3936
rect 2884 3924 2912 4023
rect 4522 3952 4528 4004
rect 4580 3992 4586 4004
rect 6656 4001 6684 4032
rect 7098 4020 7104 4072
rect 7156 4060 7162 4072
rect 7745 4063 7803 4069
rect 7745 4060 7757 4063
rect 7156 4032 7757 4060
rect 7156 4020 7162 4032
rect 7745 4029 7757 4032
rect 7791 4029 7803 4063
rect 7745 4023 7803 4029
rect 7834 4020 7840 4072
rect 7892 4060 7898 4072
rect 7929 4063 7987 4069
rect 7929 4060 7941 4063
rect 7892 4032 7941 4060
rect 7892 4020 7898 4032
rect 7929 4029 7941 4032
rect 7975 4029 7987 4063
rect 11054 4060 11060 4072
rect 7929 4023 7987 4029
rect 8404 4032 11060 4060
rect 5077 3995 5135 4001
rect 5077 3992 5089 3995
rect 4580 3964 5089 3992
rect 4580 3952 4586 3964
rect 5077 3961 5089 3964
rect 5123 3961 5135 3995
rect 5077 3955 5135 3961
rect 6641 3995 6699 4001
rect 6641 3961 6653 3995
rect 6687 3961 6699 3995
rect 6641 3955 6699 3961
rect 6914 3952 6920 4004
rect 6972 3992 6978 4004
rect 8404 3992 8432 4032
rect 11054 4020 11060 4032
rect 11112 4020 11118 4072
rect 11146 4020 11152 4072
rect 11204 4060 11210 4072
rect 13173 4063 13231 4069
rect 13173 4060 13185 4063
rect 11204 4032 13185 4060
rect 11204 4020 11210 4032
rect 13173 4029 13185 4032
rect 13219 4029 13231 4063
rect 13173 4023 13231 4029
rect 13449 4063 13507 4069
rect 13449 4029 13461 4063
rect 13495 4060 13507 4063
rect 13630 4060 13636 4072
rect 13495 4032 13636 4060
rect 13495 4029 13507 4032
rect 13449 4023 13507 4029
rect 13630 4020 13636 4032
rect 13688 4060 13694 4072
rect 13909 4063 13967 4069
rect 13909 4060 13921 4063
rect 13688 4032 13921 4060
rect 13688 4020 13694 4032
rect 13909 4029 13921 4032
rect 13955 4029 13967 4063
rect 14185 4063 14243 4069
rect 14185 4060 14197 4063
rect 13909 4023 13967 4029
rect 14016 4032 14197 4060
rect 6972 3964 8432 3992
rect 6972 3952 6978 3964
rect 8478 3952 8484 4004
rect 8536 3992 8542 4004
rect 8536 3964 11836 3992
rect 8536 3952 8542 3964
rect 4154 3924 4160 3936
rect 2556 3896 4160 3924
rect 2556 3884 2562 3896
rect 4154 3884 4160 3896
rect 4212 3884 4218 3936
rect 4617 3927 4675 3933
rect 4617 3893 4629 3927
rect 4663 3924 4675 3927
rect 4706 3924 4712 3936
rect 4663 3896 4712 3924
rect 4663 3893 4675 3896
rect 4617 3887 4675 3893
rect 4706 3884 4712 3896
rect 4764 3884 4770 3936
rect 4982 3884 4988 3936
rect 5040 3924 5046 3936
rect 9122 3924 9128 3936
rect 5040 3896 9128 3924
rect 5040 3884 5046 3896
rect 9122 3884 9128 3896
rect 9180 3884 9186 3936
rect 9398 3884 9404 3936
rect 9456 3924 9462 3936
rect 10229 3927 10287 3933
rect 10229 3924 10241 3927
rect 9456 3896 10241 3924
rect 9456 3884 9462 3896
rect 10229 3893 10241 3896
rect 10275 3893 10287 3927
rect 11808 3924 11836 3964
rect 13722 3952 13728 4004
rect 13780 3992 13786 4004
rect 14016 3992 14044 4032
rect 14185 4029 14197 4032
rect 14231 4029 14243 4063
rect 14185 4023 14243 4029
rect 13780 3964 14044 3992
rect 13780 3952 13786 3964
rect 12986 3924 12992 3936
rect 11808 3896 12992 3924
rect 10229 3887 10287 3893
rect 12986 3884 12992 3896
rect 13044 3884 13050 3936
rect 13078 3884 13084 3936
rect 13136 3924 13142 3936
rect 15657 3927 15715 3933
rect 15657 3924 15669 3927
rect 13136 3896 15669 3924
rect 13136 3884 13142 3896
rect 15657 3893 15669 3896
rect 15703 3893 15715 3927
rect 15657 3887 15715 3893
rect 1104 3834 18860 3856
rect 1104 3782 3169 3834
rect 3221 3782 3233 3834
rect 3285 3782 3297 3834
rect 3349 3782 3361 3834
rect 3413 3782 3425 3834
rect 3477 3782 7608 3834
rect 7660 3782 7672 3834
rect 7724 3782 7736 3834
rect 7788 3782 7800 3834
rect 7852 3782 7864 3834
rect 7916 3782 12047 3834
rect 12099 3782 12111 3834
rect 12163 3782 12175 3834
rect 12227 3782 12239 3834
rect 12291 3782 12303 3834
rect 12355 3782 16486 3834
rect 16538 3782 16550 3834
rect 16602 3782 16614 3834
rect 16666 3782 16678 3834
rect 16730 3782 16742 3834
rect 16794 3782 18860 3834
rect 1104 3760 18860 3782
rect 1936 3723 1994 3729
rect 1936 3689 1948 3723
rect 1982 3720 1994 3723
rect 1982 3692 4108 3720
rect 1982 3689 1994 3692
rect 1936 3683 1994 3689
rect 4080 3652 4108 3692
rect 4154 3680 4160 3732
rect 4212 3720 4218 3732
rect 4985 3723 5043 3729
rect 4985 3720 4997 3723
rect 4212 3692 4997 3720
rect 4212 3680 4218 3692
rect 4985 3689 4997 3692
rect 5031 3720 5043 3723
rect 6730 3720 6736 3732
rect 5031 3692 6736 3720
rect 5031 3689 5043 3692
rect 4985 3683 5043 3689
rect 6730 3680 6736 3692
rect 6788 3680 6794 3732
rect 16022 3720 16028 3732
rect 6840 3692 16028 3720
rect 6840 3652 6868 3692
rect 16022 3680 16028 3692
rect 16080 3680 16086 3732
rect 8478 3652 8484 3664
rect 4080 3624 6868 3652
rect 8439 3624 8484 3652
rect 8478 3612 8484 3624
rect 8536 3612 8542 3664
rect 9214 3612 9220 3664
rect 9272 3652 9278 3664
rect 9309 3655 9367 3661
rect 9309 3652 9321 3655
rect 9272 3624 9321 3652
rect 9272 3612 9278 3624
rect 9309 3621 9321 3624
rect 9355 3621 9367 3655
rect 11146 3652 11152 3664
rect 11107 3624 11152 3652
rect 9309 3615 9367 3621
rect 11146 3612 11152 3624
rect 11204 3612 11210 3664
rect 11790 3612 11796 3664
rect 11848 3652 11854 3664
rect 11977 3655 12035 3661
rect 11977 3652 11989 3655
rect 11848 3624 11989 3652
rect 11848 3612 11854 3624
rect 11977 3621 11989 3624
rect 12023 3621 12035 3655
rect 11977 3615 12035 3621
rect 1673 3587 1731 3593
rect 1673 3553 1685 3587
rect 1719 3584 1731 3587
rect 2498 3584 2504 3596
rect 1719 3556 2504 3584
rect 1719 3553 1731 3556
rect 1673 3547 1731 3553
rect 2498 3544 2504 3556
rect 2556 3544 2562 3596
rect 9398 3584 9404 3596
rect 6288 3556 9404 3584
rect 6288 3525 6316 3556
rect 9398 3544 9404 3556
rect 9456 3544 9462 3596
rect 13446 3584 13452 3596
rect 9692 3556 13452 3584
rect 6273 3519 6331 3525
rect 6273 3485 6285 3519
rect 6319 3485 6331 3519
rect 6730 3516 6736 3528
rect 6691 3488 6736 3516
rect 6273 3479 6331 3485
rect 6730 3476 6736 3488
rect 6788 3476 6794 3528
rect 8294 3516 8300 3528
rect 8142 3488 8300 3516
rect 8294 3476 8300 3488
rect 8352 3476 8358 3528
rect 9122 3516 9128 3528
rect 9083 3488 9128 3516
rect 9122 3476 9128 3488
rect 9180 3476 9186 3528
rect 4430 3448 4436 3460
rect 3174 3420 4436 3448
rect 2958 3340 2964 3392
rect 3016 3380 3022 3392
rect 3252 3380 3280 3420
rect 4430 3408 4436 3420
rect 4488 3408 4494 3460
rect 7009 3451 7067 3457
rect 7009 3417 7021 3451
rect 7055 3417 7067 3451
rect 9692 3448 9720 3556
rect 13446 3544 13452 3556
rect 13504 3544 13510 3596
rect 13722 3584 13728 3596
rect 13683 3556 13728 3584
rect 13722 3544 13728 3556
rect 13780 3544 13786 3596
rect 10226 3516 10232 3528
rect 10187 3488 10232 3516
rect 10226 3476 10232 3488
rect 10284 3476 10290 3528
rect 10962 3516 10968 3528
rect 10923 3488 10968 3516
rect 10962 3476 10968 3488
rect 11020 3476 11026 3528
rect 7009 3411 7067 3417
rect 8404 3420 9720 3448
rect 3016 3352 3280 3380
rect 3421 3383 3479 3389
rect 3016 3340 3022 3352
rect 3421 3349 3433 3383
rect 3467 3380 3479 3383
rect 6914 3380 6920 3392
rect 3467 3352 6920 3380
rect 3467 3349 3479 3352
rect 3421 3343 3479 3349
rect 6914 3340 6920 3352
rect 6972 3340 6978 3392
rect 7024 3380 7052 3411
rect 8404 3380 8432 3420
rect 11698 3408 11704 3460
rect 11756 3448 11762 3460
rect 11756 3420 12112 3448
rect 11756 3408 11762 3420
rect 7024 3352 8432 3380
rect 8662 3340 8668 3392
rect 8720 3380 8726 3392
rect 10045 3383 10103 3389
rect 10045 3380 10057 3383
rect 8720 3352 10057 3380
rect 8720 3340 8726 3352
rect 10045 3349 10057 3352
rect 10091 3349 10103 3383
rect 12084 3380 12112 3420
rect 12710 3408 12716 3460
rect 12768 3408 12774 3460
rect 13449 3451 13507 3457
rect 13449 3417 13461 3451
rect 13495 3417 13507 3451
rect 13449 3411 13507 3417
rect 13464 3380 13492 3411
rect 12084 3352 13492 3380
rect 10045 3343 10103 3349
rect 1104 3290 19019 3312
rect 1104 3238 5388 3290
rect 5440 3238 5452 3290
rect 5504 3238 5516 3290
rect 5568 3238 5580 3290
rect 5632 3238 5644 3290
rect 5696 3238 9827 3290
rect 9879 3238 9891 3290
rect 9943 3238 9955 3290
rect 10007 3238 10019 3290
rect 10071 3238 10083 3290
rect 10135 3238 14266 3290
rect 14318 3238 14330 3290
rect 14382 3238 14394 3290
rect 14446 3238 14458 3290
rect 14510 3238 14522 3290
rect 14574 3238 18705 3290
rect 18757 3238 18769 3290
rect 18821 3238 18833 3290
rect 18885 3238 18897 3290
rect 18949 3238 18961 3290
rect 19013 3238 19019 3290
rect 1104 3216 19019 3238
rect 1946 3176 1952 3188
rect 1859 3148 1952 3176
rect 1946 3136 1952 3148
rect 2004 3176 2010 3188
rect 7098 3176 7104 3188
rect 2004 3148 7104 3176
rect 2004 3136 2010 3148
rect 7098 3136 7104 3148
rect 7156 3136 7162 3188
rect 7193 3179 7251 3185
rect 7193 3145 7205 3179
rect 7239 3176 7251 3179
rect 7926 3176 7932 3188
rect 7239 3148 7932 3176
rect 7239 3145 7251 3148
rect 7193 3139 7251 3145
rect 7926 3136 7932 3148
rect 7984 3136 7990 3188
rect 9214 3176 9220 3188
rect 8588 3148 9220 3176
rect 2958 3068 2964 3120
rect 3016 3068 3022 3120
rect 3421 3111 3479 3117
rect 3421 3077 3433 3111
rect 3467 3108 3479 3111
rect 4246 3108 4252 3120
rect 3467 3080 4252 3108
rect 3467 3077 3479 3080
rect 3421 3071 3479 3077
rect 4246 3068 4252 3080
rect 4304 3068 4310 3120
rect 7374 3108 7380 3120
rect 5566 3094 7380 3108
rect 5552 3080 7380 3094
rect 3697 3043 3755 3049
rect 3697 3009 3709 3043
rect 3743 3040 3755 3043
rect 4154 3040 4160 3052
rect 3743 3012 4160 3040
rect 3743 3009 3755 3012
rect 3697 3003 3755 3009
rect 4154 3000 4160 3012
rect 4212 3000 4218 3052
rect 4522 3040 4528 3052
rect 4483 3012 4528 3040
rect 4522 3000 4528 3012
rect 4580 3000 4586 3052
rect 5258 2932 5264 2984
rect 5316 2972 5322 2984
rect 5552 2972 5580 3080
rect 7374 3068 7380 3080
rect 7432 3068 7438 3120
rect 8588 3108 8616 3148
rect 9214 3136 9220 3148
rect 9272 3136 9278 3188
rect 10870 3136 10876 3188
rect 10928 3176 10934 3188
rect 13722 3176 13728 3188
rect 10928 3148 13728 3176
rect 10928 3136 10934 3148
rect 13722 3136 13728 3148
rect 13780 3136 13786 3188
rect 8234 3080 8616 3108
rect 8662 3068 8668 3120
rect 8720 3117 8726 3120
rect 8720 3111 8735 3117
rect 8723 3077 8735 3111
rect 9398 3108 9404 3120
rect 9359 3080 9404 3108
rect 8720 3071 8735 3077
rect 8720 3068 8726 3071
rect 9398 3068 9404 3080
rect 9456 3068 9462 3120
rect 12710 3068 12716 3120
rect 12768 3068 12774 3120
rect 12894 3068 12900 3120
rect 12952 3108 12958 3120
rect 13173 3111 13231 3117
rect 13173 3108 13185 3111
rect 12952 3080 13185 3108
rect 12952 3068 12958 3080
rect 13173 3077 13185 3080
rect 13219 3077 13231 3111
rect 13173 3071 13231 3077
rect 13446 3068 13452 3120
rect 13504 3108 13510 3120
rect 13504 3080 16574 3108
rect 13504 3068 13510 3080
rect 9030 3000 9036 3052
rect 9088 3040 9094 3052
rect 10686 3040 10692 3052
rect 9088 3012 10692 3040
rect 9088 3000 9094 3012
rect 10686 3000 10692 3012
rect 10744 3000 10750 3052
rect 13906 3040 13912 3052
rect 13867 3012 13912 3040
rect 13906 3000 13912 3012
rect 13964 3000 13970 3052
rect 5316 2944 5580 2972
rect 5951 2975 6009 2981
rect 5316 2932 5322 2944
rect 5951 2941 5963 2975
rect 5997 2972 6009 2975
rect 8941 2975 8999 2981
rect 5997 2944 8892 2972
rect 5997 2941 6009 2944
rect 5951 2935 6009 2941
rect 8864 2904 8892 2944
rect 8941 2941 8953 2975
rect 8987 2972 8999 2975
rect 13449 2975 13507 2981
rect 8987 2944 10732 2972
rect 8987 2941 8999 2944
rect 8941 2935 8999 2941
rect 10704 2913 10732 2944
rect 10980 2944 13400 2972
rect 10689 2907 10747 2913
rect 8864 2876 10640 2904
rect 7466 2796 7472 2848
rect 7524 2836 7530 2848
rect 9582 2836 9588 2848
rect 7524 2808 9588 2836
rect 7524 2796 7530 2808
rect 9582 2796 9588 2808
rect 9640 2796 9646 2848
rect 10612 2836 10640 2876
rect 10689 2873 10701 2907
rect 10735 2904 10747 2907
rect 10870 2904 10876 2916
rect 10735 2876 10876 2904
rect 10735 2873 10747 2876
rect 10689 2867 10747 2873
rect 10870 2864 10876 2876
rect 10928 2864 10934 2916
rect 10980 2836 11008 2944
rect 11698 2904 11704 2916
rect 11659 2876 11704 2904
rect 11698 2864 11704 2876
rect 11756 2864 11762 2916
rect 13372 2904 13400 2944
rect 13449 2941 13461 2975
rect 13495 2972 13507 2975
rect 13722 2972 13728 2984
rect 13495 2944 13728 2972
rect 13495 2941 13507 2944
rect 13449 2935 13507 2941
rect 13722 2932 13728 2944
rect 13780 2932 13786 2984
rect 15378 2904 15384 2916
rect 13372 2876 15384 2904
rect 15378 2864 15384 2876
rect 15436 2904 15442 2916
rect 15746 2904 15752 2916
rect 15436 2876 15752 2904
rect 15436 2864 15442 2876
rect 15746 2864 15752 2876
rect 15804 2864 15810 2916
rect 16546 2904 16574 3080
rect 16850 2904 16856 2916
rect 16546 2876 16856 2904
rect 16850 2864 16856 2876
rect 16908 2864 16914 2916
rect 10612 2808 11008 2836
rect 12434 2796 12440 2848
rect 12492 2836 12498 2848
rect 14093 2839 14151 2845
rect 14093 2836 14105 2839
rect 12492 2808 14105 2836
rect 12492 2796 12498 2808
rect 14093 2805 14105 2808
rect 14139 2805 14151 2839
rect 14093 2799 14151 2805
rect 1104 2746 18860 2768
rect 1104 2694 3169 2746
rect 3221 2694 3233 2746
rect 3285 2694 3297 2746
rect 3349 2694 3361 2746
rect 3413 2694 3425 2746
rect 3477 2694 7608 2746
rect 7660 2694 7672 2746
rect 7724 2694 7736 2746
rect 7788 2694 7800 2746
rect 7852 2694 7864 2746
rect 7916 2694 12047 2746
rect 12099 2694 12111 2746
rect 12163 2694 12175 2746
rect 12227 2694 12239 2746
rect 12291 2694 12303 2746
rect 12355 2694 16486 2746
rect 16538 2694 16550 2746
rect 16602 2694 16614 2746
rect 16666 2694 16678 2746
rect 16730 2694 16742 2746
rect 16794 2694 18860 2746
rect 1104 2672 18860 2694
rect 3421 2635 3479 2641
rect 3421 2601 3433 2635
rect 3467 2632 3479 2635
rect 5997 2635 6055 2641
rect 3467 2604 5948 2632
rect 3467 2601 3479 2604
rect 3421 2595 3479 2601
rect 5920 2564 5948 2604
rect 5997 2601 6009 2635
rect 6043 2632 6055 2635
rect 7006 2632 7012 2644
rect 6043 2604 7012 2632
rect 6043 2601 6055 2604
rect 5997 2595 6055 2601
rect 7006 2592 7012 2604
rect 7064 2592 7070 2644
rect 8202 2592 8208 2644
rect 8260 2632 8266 2644
rect 9125 2635 9183 2641
rect 9125 2632 9137 2635
rect 8260 2604 9137 2632
rect 8260 2592 8266 2604
rect 9125 2601 9137 2604
rect 9171 2601 9183 2635
rect 9125 2595 9183 2601
rect 12894 2592 12900 2644
rect 12952 2632 12958 2644
rect 14277 2635 14335 2641
rect 14277 2632 14289 2635
rect 12952 2604 14289 2632
rect 12952 2592 12958 2604
rect 14277 2601 14289 2604
rect 14323 2601 14335 2635
rect 14277 2595 14335 2601
rect 9582 2564 9588 2576
rect 5920 2536 9588 2564
rect 9582 2524 9588 2536
rect 9640 2524 9646 2576
rect 11977 2567 12035 2573
rect 11977 2564 11989 2567
rect 10796 2536 11989 2564
rect 1673 2499 1731 2505
rect 1673 2465 1685 2499
rect 1719 2496 1731 2499
rect 2498 2496 2504 2508
rect 1719 2468 2504 2496
rect 1719 2465 1731 2468
rect 1673 2459 1731 2465
rect 2498 2456 2504 2468
rect 2556 2456 2562 2508
rect 4154 2456 4160 2508
rect 4212 2496 4218 2508
rect 4249 2499 4307 2505
rect 4249 2496 4261 2499
rect 4212 2468 4261 2496
rect 4212 2456 4218 2468
rect 4249 2465 4261 2468
rect 4295 2465 4307 2499
rect 4249 2459 4307 2465
rect 4525 2499 4583 2505
rect 4525 2465 4537 2499
rect 4571 2496 4583 2499
rect 4614 2496 4620 2508
rect 4571 2468 4620 2496
rect 4571 2465 4583 2468
rect 4525 2459 4583 2465
rect 4614 2456 4620 2468
rect 4672 2456 4678 2508
rect 8018 2456 8024 2508
rect 8076 2496 8082 2508
rect 10597 2499 10655 2505
rect 10597 2496 10609 2499
rect 8076 2468 10609 2496
rect 8076 2456 8082 2468
rect 10597 2465 10609 2468
rect 10643 2496 10655 2499
rect 10796 2496 10824 2536
rect 11977 2533 11989 2536
rect 12023 2533 12035 2567
rect 11977 2527 12035 2533
rect 10643 2468 10824 2496
rect 10643 2465 10655 2468
rect 10597 2459 10655 2465
rect 11698 2456 11704 2508
rect 11756 2496 11762 2508
rect 13449 2499 13507 2505
rect 13449 2496 13461 2499
rect 11756 2468 13461 2496
rect 11756 2456 11762 2468
rect 13449 2465 13461 2468
rect 13495 2465 13507 2499
rect 13722 2496 13728 2508
rect 13635 2468 13728 2496
rect 13449 2459 13507 2465
rect 13722 2456 13728 2468
rect 13780 2496 13786 2508
rect 16025 2499 16083 2505
rect 16025 2496 16037 2499
rect 13780 2468 16037 2496
rect 13780 2456 13786 2468
rect 16025 2465 16037 2468
rect 16071 2465 16083 2499
rect 16025 2459 16083 2465
rect 10870 2388 10876 2440
rect 10928 2428 10934 2440
rect 17494 2428 17500 2440
rect 10928 2400 10973 2428
rect 17455 2400 17500 2428
rect 10928 2388 10934 2400
rect 17494 2388 17500 2400
rect 17552 2388 17558 2440
rect 1946 2360 1952 2372
rect 1907 2332 1952 2360
rect 1946 2320 1952 2332
rect 2004 2320 2010 2372
rect 15746 2360 15752 2372
rect 3174 2332 5014 2360
rect 10166 2332 11836 2360
rect 13018 2332 14582 2360
rect 15707 2332 15752 2360
rect 4908 2292 4936 2332
rect 5258 2292 5264 2304
rect 4908 2264 5264 2292
rect 5258 2252 5264 2264
rect 5316 2252 5322 2304
rect 9306 2252 9312 2304
rect 9364 2292 9370 2304
rect 10244 2292 10272 2332
rect 9364 2264 10272 2292
rect 11808 2292 11836 2332
rect 12710 2292 12716 2304
rect 11808 2264 12716 2292
rect 9364 2252 9370 2264
rect 12710 2252 12716 2264
rect 12768 2292 12774 2304
rect 13096 2292 13124 2332
rect 15746 2320 15752 2332
rect 15804 2320 15810 2372
rect 12768 2264 13124 2292
rect 12768 2252 12774 2264
rect 17402 2252 17408 2304
rect 17460 2292 17466 2304
rect 17681 2295 17739 2301
rect 17681 2292 17693 2295
rect 17460 2264 17693 2292
rect 17460 2252 17466 2264
rect 17681 2261 17693 2264
rect 17727 2261 17739 2295
rect 17681 2255 17739 2261
rect 1104 2202 19019 2224
rect 1104 2150 5388 2202
rect 5440 2150 5452 2202
rect 5504 2150 5516 2202
rect 5568 2150 5580 2202
rect 5632 2150 5644 2202
rect 5696 2150 9827 2202
rect 9879 2150 9891 2202
rect 9943 2150 9955 2202
rect 10007 2150 10019 2202
rect 10071 2150 10083 2202
rect 10135 2150 14266 2202
rect 14318 2150 14330 2202
rect 14382 2150 14394 2202
rect 14446 2150 14458 2202
rect 14510 2150 14522 2202
rect 14574 2150 18705 2202
rect 18757 2150 18769 2202
rect 18821 2150 18833 2202
rect 18885 2150 18897 2202
rect 18949 2150 18961 2202
rect 19013 2150 19019 2202
rect 1104 2128 19019 2150
rect 10686 2048 10692 2100
rect 10744 2088 10750 2100
rect 17494 2088 17500 2100
rect 10744 2060 17500 2088
rect 10744 2048 10750 2060
rect 17494 2048 17500 2060
rect 17552 2048 17558 2100
<< via1 >>
rect 5388 7590 5440 7642
rect 5452 7590 5504 7642
rect 5516 7590 5568 7642
rect 5580 7590 5632 7642
rect 5644 7590 5696 7642
rect 9827 7590 9879 7642
rect 9891 7590 9943 7642
rect 9955 7590 10007 7642
rect 10019 7590 10071 7642
rect 10083 7590 10135 7642
rect 14266 7590 14318 7642
rect 14330 7590 14382 7642
rect 14394 7590 14446 7642
rect 14458 7590 14510 7642
rect 14522 7590 14574 7642
rect 18705 7590 18757 7642
rect 18769 7590 18821 7642
rect 18833 7590 18885 7642
rect 18897 7590 18949 7642
rect 18961 7590 19013 7642
rect 1124 7488 1176 7540
rect 3332 7488 3384 7540
rect 5724 7531 5776 7540
rect 5724 7497 5733 7531
rect 5733 7497 5767 7531
rect 5767 7497 5776 7531
rect 5724 7488 5776 7497
rect 7932 7531 7984 7540
rect 7932 7497 7941 7531
rect 7941 7497 7975 7531
rect 7975 7497 7984 7531
rect 7932 7488 7984 7497
rect 12440 7531 12492 7540
rect 12440 7497 12449 7531
rect 12449 7497 12483 7531
rect 12483 7497 12492 7531
rect 12440 7488 12492 7497
rect 14648 7531 14700 7540
rect 14648 7497 14657 7531
rect 14657 7497 14691 7531
rect 14691 7497 14700 7531
rect 14648 7488 14700 7497
rect 16580 7488 16632 7540
rect 18420 7488 18472 7540
rect 7288 7420 7340 7472
rect 7012 7352 7064 7404
rect 7472 7352 7524 7404
rect 10232 7420 10284 7472
rect 13820 7352 13872 7404
rect 16856 7395 16908 7404
rect 16856 7361 16865 7395
rect 16865 7361 16899 7395
rect 16899 7361 16908 7395
rect 16856 7352 16908 7361
rect 7932 7284 7984 7336
rect 13360 7284 13412 7336
rect 10324 7259 10376 7268
rect 10324 7225 10333 7259
rect 10333 7225 10367 7259
rect 10367 7225 10376 7259
rect 10324 7216 10376 7225
rect 11060 7148 11112 7200
rect 3169 7046 3221 7098
rect 3233 7046 3285 7098
rect 3297 7046 3349 7098
rect 3361 7046 3413 7098
rect 3425 7046 3477 7098
rect 7608 7046 7660 7098
rect 7672 7046 7724 7098
rect 7736 7046 7788 7098
rect 7800 7046 7852 7098
rect 7864 7046 7916 7098
rect 12047 7046 12099 7098
rect 12111 7046 12163 7098
rect 12175 7046 12227 7098
rect 12239 7046 12291 7098
rect 12303 7046 12355 7098
rect 16486 7046 16538 7098
rect 16550 7046 16602 7098
rect 16614 7046 16666 7098
rect 16678 7046 16730 7098
rect 16742 7046 16794 7098
rect 5388 6502 5440 6554
rect 5452 6502 5504 6554
rect 5516 6502 5568 6554
rect 5580 6502 5632 6554
rect 5644 6502 5696 6554
rect 9827 6502 9879 6554
rect 9891 6502 9943 6554
rect 9955 6502 10007 6554
rect 10019 6502 10071 6554
rect 10083 6502 10135 6554
rect 14266 6502 14318 6554
rect 14330 6502 14382 6554
rect 14394 6502 14446 6554
rect 14458 6502 14510 6554
rect 14522 6502 14574 6554
rect 18705 6502 18757 6554
rect 18769 6502 18821 6554
rect 18833 6502 18885 6554
rect 18897 6502 18949 6554
rect 18961 6502 19013 6554
rect 8024 6307 8076 6316
rect 8024 6273 8033 6307
rect 8033 6273 8067 6307
rect 8067 6273 8076 6307
rect 8024 6264 8076 6273
rect 8208 6307 8260 6316
rect 8208 6273 8217 6307
rect 8217 6273 8251 6307
rect 8251 6273 8260 6307
rect 8208 6264 8260 6273
rect 10968 6060 11020 6112
rect 3169 5958 3221 6010
rect 3233 5958 3285 6010
rect 3297 5958 3349 6010
rect 3361 5958 3413 6010
rect 3425 5958 3477 6010
rect 7608 5958 7660 6010
rect 7672 5958 7724 6010
rect 7736 5958 7788 6010
rect 7800 5958 7852 6010
rect 7864 5958 7916 6010
rect 12047 5958 12099 6010
rect 12111 5958 12163 6010
rect 12175 5958 12227 6010
rect 12239 5958 12291 6010
rect 12303 5958 12355 6010
rect 16486 5958 16538 6010
rect 16550 5958 16602 6010
rect 16614 5958 16666 6010
rect 16678 5958 16730 6010
rect 16742 5958 16794 6010
rect 8024 5856 8076 5908
rect 8116 5720 8168 5772
rect 6920 5695 6972 5704
rect 6920 5661 6929 5695
rect 6929 5661 6963 5695
rect 6963 5661 6972 5695
rect 6920 5652 6972 5661
rect 7472 5584 7524 5636
rect 11520 5627 11572 5636
rect 11520 5593 11529 5627
rect 11529 5593 11563 5627
rect 11563 5593 11572 5627
rect 11520 5584 11572 5593
rect 11704 5627 11756 5636
rect 11704 5593 11713 5627
rect 11713 5593 11747 5627
rect 11747 5593 11756 5627
rect 11704 5584 11756 5593
rect 12808 5627 12860 5636
rect 12808 5593 12817 5627
rect 12817 5593 12851 5627
rect 12851 5593 12860 5627
rect 12808 5584 12860 5593
rect 12900 5584 12952 5636
rect 4620 5516 4672 5568
rect 7380 5516 7432 5568
rect 13084 5516 13136 5568
rect 15108 5516 15160 5568
rect 5388 5414 5440 5466
rect 5452 5414 5504 5466
rect 5516 5414 5568 5466
rect 5580 5414 5632 5466
rect 5644 5414 5696 5466
rect 9827 5414 9879 5466
rect 9891 5414 9943 5466
rect 9955 5414 10007 5466
rect 10019 5414 10071 5466
rect 10083 5414 10135 5466
rect 14266 5414 14318 5466
rect 14330 5414 14382 5466
rect 14394 5414 14446 5466
rect 14458 5414 14510 5466
rect 14522 5414 14574 5466
rect 18705 5414 18757 5466
rect 18769 5414 18821 5466
rect 18833 5414 18885 5466
rect 18897 5414 18949 5466
rect 18961 5414 19013 5466
rect 7012 5355 7064 5364
rect 4436 5244 4488 5296
rect 7012 5321 7021 5355
rect 7021 5321 7055 5355
rect 7055 5321 7064 5355
rect 7012 5312 7064 5321
rect 7380 5312 7432 5364
rect 6736 5176 6788 5228
rect 3056 5151 3108 5160
rect 3056 5117 3065 5151
rect 3065 5117 3099 5151
rect 3099 5117 3108 5151
rect 3056 5108 3108 5117
rect 9220 5176 9272 5228
rect 11060 5312 11112 5364
rect 11520 5312 11572 5364
rect 10324 5287 10376 5296
rect 10324 5253 10333 5287
rect 10333 5253 10367 5287
rect 10367 5253 10376 5287
rect 12440 5312 12492 5364
rect 10324 5244 10376 5253
rect 13820 5244 13872 5296
rect 12992 5176 13044 5228
rect 13360 5176 13412 5228
rect 8116 5151 8168 5160
rect 4252 5040 4304 5092
rect 8116 5117 8125 5151
rect 8125 5117 8159 5151
rect 8159 5117 8168 5151
rect 8116 5108 8168 5117
rect 9680 5108 9732 5160
rect 11888 5108 11940 5160
rect 12900 5108 12952 5160
rect 4160 4972 4212 5024
rect 6828 4972 6880 5024
rect 13912 5040 13964 5092
rect 9312 4972 9364 5024
rect 10508 4972 10560 5024
rect 15200 4972 15252 5024
rect 3169 4870 3221 4922
rect 3233 4870 3285 4922
rect 3297 4870 3349 4922
rect 3361 4870 3413 4922
rect 3425 4870 3477 4922
rect 7608 4870 7660 4922
rect 7672 4870 7724 4922
rect 7736 4870 7788 4922
rect 7800 4870 7852 4922
rect 7864 4870 7916 4922
rect 12047 4870 12099 4922
rect 12111 4870 12163 4922
rect 12175 4870 12227 4922
rect 12239 4870 12291 4922
rect 12303 4870 12355 4922
rect 16486 4870 16538 4922
rect 16550 4870 16602 4922
rect 16614 4870 16666 4922
rect 16678 4870 16730 4922
rect 16742 4870 16794 4922
rect 6920 4768 6972 4820
rect 3056 4700 3108 4752
rect 8300 4700 8352 4752
rect 2780 4564 2832 4616
rect 8024 4632 8076 4684
rect 8208 4632 8260 4684
rect 6828 4607 6880 4616
rect 6828 4573 6837 4607
rect 6837 4573 6871 4607
rect 6871 4573 6880 4607
rect 6828 4564 6880 4573
rect 7380 4564 7432 4616
rect 7840 4564 7892 4616
rect 10324 4632 10376 4684
rect 9036 4564 9088 4616
rect 9588 4564 9640 4616
rect 10508 4607 10560 4616
rect 10508 4573 10517 4607
rect 10517 4573 10551 4607
rect 10551 4573 10560 4607
rect 10508 4564 10560 4573
rect 4988 4496 5040 4548
rect 6184 4539 6236 4548
rect 6184 4505 6193 4539
rect 6193 4505 6227 4539
rect 6227 4505 6236 4539
rect 6184 4496 6236 4505
rect 8116 4496 8168 4548
rect 8392 4496 8444 4548
rect 9312 4539 9364 4548
rect 9312 4505 9321 4539
rect 9321 4505 9355 4539
rect 9355 4505 9364 4539
rect 9312 4496 9364 4505
rect 10692 4539 10744 4548
rect 10692 4505 10701 4539
rect 10701 4505 10735 4539
rect 10735 4505 10744 4539
rect 10692 4496 10744 4505
rect 11980 4700 12032 4752
rect 11704 4632 11756 4684
rect 10968 4564 11020 4616
rect 11888 4496 11940 4548
rect 12808 4768 12860 4820
rect 12348 4700 12400 4752
rect 13728 4700 13780 4752
rect 12440 4632 12492 4684
rect 16856 4700 16908 4752
rect 12348 4564 12400 4616
rect 15108 4632 15160 4684
rect 13084 4564 13136 4616
rect 15200 4607 15252 4616
rect 15200 4573 15209 4607
rect 15209 4573 15243 4607
rect 15243 4573 15252 4607
rect 15200 4564 15252 4573
rect 15384 4539 15436 4548
rect 2228 4428 2280 4480
rect 4436 4428 4488 4480
rect 6828 4428 6880 4480
rect 7288 4428 7340 4480
rect 8852 4428 8904 4480
rect 9404 4428 9456 4480
rect 10232 4428 10284 4480
rect 10968 4428 11020 4480
rect 11060 4428 11112 4480
rect 12348 4471 12400 4480
rect 12348 4437 12357 4471
rect 12357 4437 12391 4471
rect 12391 4437 12400 4471
rect 12348 4428 12400 4437
rect 15384 4505 15393 4539
rect 15393 4505 15427 4539
rect 15427 4505 15436 4539
rect 15384 4496 15436 4505
rect 16028 4471 16080 4480
rect 16028 4437 16037 4471
rect 16037 4437 16071 4471
rect 16071 4437 16080 4471
rect 16028 4428 16080 4437
rect 16856 4428 16908 4480
rect 5388 4326 5440 4378
rect 5452 4326 5504 4378
rect 5516 4326 5568 4378
rect 5580 4326 5632 4378
rect 5644 4326 5696 4378
rect 9827 4326 9879 4378
rect 9891 4326 9943 4378
rect 9955 4326 10007 4378
rect 10019 4326 10071 4378
rect 10083 4326 10135 4378
rect 14266 4326 14318 4378
rect 14330 4326 14382 4378
rect 14394 4326 14446 4378
rect 14458 4326 14510 4378
rect 14522 4326 14574 4378
rect 18705 4326 18757 4378
rect 18769 4326 18821 4378
rect 18833 4326 18885 4378
rect 18897 4326 18949 4378
rect 18961 4326 19013 4378
rect 4988 4224 5040 4276
rect 6184 4224 6236 4276
rect 4436 4156 4488 4208
rect 5264 4156 5316 4208
rect 2228 4131 2280 4140
rect 2228 4097 2237 4131
rect 2237 4097 2271 4131
rect 2271 4097 2280 4131
rect 2228 4088 2280 4097
rect 4712 4088 4764 4140
rect 7288 4156 7340 4208
rect 7932 4224 7984 4276
rect 8392 4267 8444 4276
rect 8392 4233 8401 4267
rect 8401 4233 8435 4267
rect 8435 4233 8444 4267
rect 8392 4224 8444 4233
rect 8852 4156 8904 4208
rect 9036 4224 9088 4276
rect 11152 4224 11204 4276
rect 11888 4224 11940 4276
rect 9404 4156 9456 4208
rect 11796 4156 11848 4208
rect 6828 4131 6880 4140
rect 6828 4097 6837 4131
rect 6837 4097 6871 4131
rect 6871 4097 6880 4131
rect 6828 4088 6880 4097
rect 7472 4088 7524 4140
rect 11888 4088 11940 4140
rect 2504 3884 2556 3936
rect 4528 3952 4580 4004
rect 7104 4020 7156 4072
rect 7840 4020 7892 4072
rect 6920 3952 6972 4004
rect 11060 4020 11112 4072
rect 11152 4020 11204 4072
rect 13636 4020 13688 4072
rect 8484 3952 8536 4004
rect 4160 3884 4212 3936
rect 4712 3884 4764 3936
rect 4988 3884 5040 3936
rect 9128 3884 9180 3936
rect 9404 3884 9456 3936
rect 13728 3952 13780 4004
rect 12992 3884 13044 3936
rect 13084 3884 13136 3936
rect 3169 3782 3221 3834
rect 3233 3782 3285 3834
rect 3297 3782 3349 3834
rect 3361 3782 3413 3834
rect 3425 3782 3477 3834
rect 7608 3782 7660 3834
rect 7672 3782 7724 3834
rect 7736 3782 7788 3834
rect 7800 3782 7852 3834
rect 7864 3782 7916 3834
rect 12047 3782 12099 3834
rect 12111 3782 12163 3834
rect 12175 3782 12227 3834
rect 12239 3782 12291 3834
rect 12303 3782 12355 3834
rect 16486 3782 16538 3834
rect 16550 3782 16602 3834
rect 16614 3782 16666 3834
rect 16678 3782 16730 3834
rect 16742 3782 16794 3834
rect 4160 3680 4212 3732
rect 6736 3680 6788 3732
rect 16028 3680 16080 3732
rect 8484 3655 8536 3664
rect 8484 3621 8493 3655
rect 8493 3621 8527 3655
rect 8527 3621 8536 3655
rect 8484 3612 8536 3621
rect 9220 3612 9272 3664
rect 11152 3655 11204 3664
rect 11152 3621 11161 3655
rect 11161 3621 11195 3655
rect 11195 3621 11204 3655
rect 11152 3612 11204 3621
rect 11796 3612 11848 3664
rect 2504 3544 2556 3596
rect 9404 3544 9456 3596
rect 6736 3519 6788 3528
rect 6736 3485 6745 3519
rect 6745 3485 6779 3519
rect 6779 3485 6788 3519
rect 6736 3476 6788 3485
rect 8300 3476 8352 3528
rect 9128 3519 9180 3528
rect 9128 3485 9137 3519
rect 9137 3485 9171 3519
rect 9171 3485 9180 3519
rect 9128 3476 9180 3485
rect 2964 3340 3016 3392
rect 4436 3408 4488 3460
rect 13452 3544 13504 3596
rect 13728 3587 13780 3596
rect 13728 3553 13737 3587
rect 13737 3553 13771 3587
rect 13771 3553 13780 3587
rect 13728 3544 13780 3553
rect 10232 3519 10284 3528
rect 10232 3485 10241 3519
rect 10241 3485 10275 3519
rect 10275 3485 10284 3519
rect 10232 3476 10284 3485
rect 10968 3519 11020 3528
rect 10968 3485 10977 3519
rect 10977 3485 11011 3519
rect 11011 3485 11020 3519
rect 10968 3476 11020 3485
rect 6920 3340 6972 3392
rect 11704 3408 11756 3460
rect 8668 3340 8720 3392
rect 12716 3408 12768 3460
rect 5388 3238 5440 3290
rect 5452 3238 5504 3290
rect 5516 3238 5568 3290
rect 5580 3238 5632 3290
rect 5644 3238 5696 3290
rect 9827 3238 9879 3290
rect 9891 3238 9943 3290
rect 9955 3238 10007 3290
rect 10019 3238 10071 3290
rect 10083 3238 10135 3290
rect 14266 3238 14318 3290
rect 14330 3238 14382 3290
rect 14394 3238 14446 3290
rect 14458 3238 14510 3290
rect 14522 3238 14574 3290
rect 18705 3238 18757 3290
rect 18769 3238 18821 3290
rect 18833 3238 18885 3290
rect 18897 3238 18949 3290
rect 18961 3238 19013 3290
rect 1952 3179 2004 3188
rect 1952 3145 1961 3179
rect 1961 3145 1995 3179
rect 1995 3145 2004 3179
rect 1952 3136 2004 3145
rect 7104 3136 7156 3188
rect 7932 3136 7984 3188
rect 2964 3068 3016 3120
rect 4252 3068 4304 3120
rect 4160 3043 4212 3052
rect 4160 3009 4169 3043
rect 4169 3009 4203 3043
rect 4203 3009 4212 3043
rect 4160 3000 4212 3009
rect 4528 3043 4580 3052
rect 4528 3009 4537 3043
rect 4537 3009 4571 3043
rect 4571 3009 4580 3043
rect 4528 3000 4580 3009
rect 5264 2932 5316 2984
rect 7380 3068 7432 3120
rect 9220 3136 9272 3188
rect 10876 3136 10928 3188
rect 13728 3136 13780 3188
rect 8668 3111 8720 3120
rect 8668 3077 8689 3111
rect 8689 3077 8720 3111
rect 9404 3111 9456 3120
rect 8668 3068 8720 3077
rect 9404 3077 9413 3111
rect 9413 3077 9447 3111
rect 9447 3077 9456 3111
rect 9404 3068 9456 3077
rect 12716 3068 12768 3120
rect 12900 3068 12952 3120
rect 13452 3068 13504 3120
rect 9036 3000 9088 3052
rect 10692 3000 10744 3052
rect 13912 3043 13964 3052
rect 13912 3009 13921 3043
rect 13921 3009 13955 3043
rect 13955 3009 13964 3043
rect 13912 3000 13964 3009
rect 7472 2796 7524 2848
rect 9588 2796 9640 2848
rect 10876 2864 10928 2916
rect 11704 2907 11756 2916
rect 11704 2873 11713 2907
rect 11713 2873 11747 2907
rect 11747 2873 11756 2907
rect 11704 2864 11756 2873
rect 13728 2932 13780 2984
rect 15384 2864 15436 2916
rect 15752 2864 15804 2916
rect 16856 2864 16908 2916
rect 12440 2796 12492 2848
rect 3169 2694 3221 2746
rect 3233 2694 3285 2746
rect 3297 2694 3349 2746
rect 3361 2694 3413 2746
rect 3425 2694 3477 2746
rect 7608 2694 7660 2746
rect 7672 2694 7724 2746
rect 7736 2694 7788 2746
rect 7800 2694 7852 2746
rect 7864 2694 7916 2746
rect 12047 2694 12099 2746
rect 12111 2694 12163 2746
rect 12175 2694 12227 2746
rect 12239 2694 12291 2746
rect 12303 2694 12355 2746
rect 16486 2694 16538 2746
rect 16550 2694 16602 2746
rect 16614 2694 16666 2746
rect 16678 2694 16730 2746
rect 16742 2694 16794 2746
rect 7012 2592 7064 2644
rect 8208 2592 8260 2644
rect 12900 2592 12952 2644
rect 9588 2524 9640 2576
rect 2504 2456 2556 2508
rect 4160 2456 4212 2508
rect 4620 2456 4672 2508
rect 8024 2456 8076 2508
rect 11704 2456 11756 2508
rect 13728 2499 13780 2508
rect 13728 2465 13737 2499
rect 13737 2465 13771 2499
rect 13771 2465 13780 2499
rect 13728 2456 13780 2465
rect 10876 2431 10928 2440
rect 10876 2397 10885 2431
rect 10885 2397 10919 2431
rect 10919 2397 10928 2431
rect 17500 2431 17552 2440
rect 10876 2388 10928 2397
rect 17500 2397 17509 2431
rect 17509 2397 17543 2431
rect 17543 2397 17552 2431
rect 17500 2388 17552 2397
rect 1952 2363 2004 2372
rect 1952 2329 1961 2363
rect 1961 2329 1995 2363
rect 1995 2329 2004 2363
rect 1952 2320 2004 2329
rect 15752 2363 15804 2372
rect 5264 2252 5316 2304
rect 9312 2252 9364 2304
rect 12716 2252 12768 2304
rect 15752 2329 15761 2363
rect 15761 2329 15795 2363
rect 15795 2329 15804 2363
rect 15752 2320 15804 2329
rect 17408 2252 17460 2304
rect 5388 2150 5440 2202
rect 5452 2150 5504 2202
rect 5516 2150 5568 2202
rect 5580 2150 5632 2202
rect 5644 2150 5696 2202
rect 9827 2150 9879 2202
rect 9891 2150 9943 2202
rect 9955 2150 10007 2202
rect 10019 2150 10071 2202
rect 10083 2150 10135 2202
rect 14266 2150 14318 2202
rect 14330 2150 14382 2202
rect 14394 2150 14446 2202
rect 14458 2150 14510 2202
rect 14522 2150 14574 2202
rect 18705 2150 18757 2202
rect 18769 2150 18821 2202
rect 18833 2150 18885 2202
rect 18897 2150 18949 2202
rect 18961 2150 19013 2202
rect 10692 2048 10744 2100
rect 17500 2048 17552 2100
<< metal2 >>
rect 1122 9200 1178 10000
rect 3330 9200 3386 10000
rect 5538 9330 5594 10000
rect 7746 9330 7802 10000
rect 9954 9330 10010 10000
rect 12162 9330 12218 10000
rect 14370 9330 14426 10000
rect 5538 9302 5764 9330
rect 5538 9200 5594 9302
rect 1136 7546 1164 9200
rect 3344 7546 3372 9200
rect 5388 7644 5696 7653
rect 5388 7642 5394 7644
rect 5450 7642 5474 7644
rect 5530 7642 5554 7644
rect 5610 7642 5634 7644
rect 5690 7642 5696 7644
rect 5450 7590 5452 7642
rect 5632 7590 5634 7642
rect 5388 7588 5394 7590
rect 5450 7588 5474 7590
rect 5530 7588 5554 7590
rect 5610 7588 5634 7590
rect 5690 7588 5696 7590
rect 5388 7579 5696 7588
rect 5736 7546 5764 9302
rect 7746 9302 7972 9330
rect 7746 9200 7802 9302
rect 7944 7546 7972 9302
rect 9954 9302 10272 9330
rect 9954 9200 10010 9302
rect 9827 7644 10135 7653
rect 9827 7642 9833 7644
rect 9889 7642 9913 7644
rect 9969 7642 9993 7644
rect 10049 7642 10073 7644
rect 10129 7642 10135 7644
rect 9889 7590 9891 7642
rect 10071 7590 10073 7642
rect 9827 7588 9833 7590
rect 9889 7588 9913 7590
rect 9969 7588 9993 7590
rect 10049 7588 10073 7590
rect 10129 7588 10135 7590
rect 9827 7579 10135 7588
rect 1124 7540 1176 7546
rect 1124 7482 1176 7488
rect 3332 7540 3384 7546
rect 3332 7482 3384 7488
rect 5724 7540 5776 7546
rect 5724 7482 5776 7488
rect 7932 7540 7984 7546
rect 7932 7482 7984 7488
rect 10244 7478 10272 9302
rect 12162 9302 12388 9330
rect 12162 9200 12218 9302
rect 12360 7528 12388 9302
rect 14370 9302 14688 9330
rect 14370 9200 14426 9302
rect 14266 7644 14574 7653
rect 14266 7642 14272 7644
rect 14328 7642 14352 7644
rect 14408 7642 14432 7644
rect 14488 7642 14512 7644
rect 14568 7642 14574 7644
rect 14328 7590 14330 7642
rect 14510 7590 14512 7642
rect 14266 7588 14272 7590
rect 14328 7588 14352 7590
rect 14408 7588 14432 7590
rect 14488 7588 14512 7590
rect 14568 7588 14574 7590
rect 14266 7579 14574 7588
rect 14660 7546 14688 9302
rect 16578 9200 16634 10000
rect 18786 9330 18842 10000
rect 18432 9302 18842 9330
rect 16592 7546 16620 9200
rect 18432 7546 18460 9302
rect 18786 9200 18842 9302
rect 18705 7644 19013 7653
rect 18705 7642 18711 7644
rect 18767 7642 18791 7644
rect 18847 7642 18871 7644
rect 18927 7642 18951 7644
rect 19007 7642 19013 7644
rect 18767 7590 18769 7642
rect 18949 7590 18951 7642
rect 18705 7588 18711 7590
rect 18767 7588 18791 7590
rect 18847 7588 18871 7590
rect 18927 7588 18951 7590
rect 19007 7588 19013 7590
rect 18705 7579 19013 7588
rect 12440 7540 12492 7546
rect 12360 7500 12440 7528
rect 12440 7482 12492 7488
rect 14648 7540 14700 7546
rect 14648 7482 14700 7488
rect 16580 7540 16632 7546
rect 16580 7482 16632 7488
rect 18420 7540 18472 7546
rect 18420 7482 18472 7488
rect 7288 7472 7340 7478
rect 7288 7414 7340 7420
rect 10232 7472 10284 7478
rect 10232 7414 10284 7420
rect 7012 7404 7064 7410
rect 7012 7346 7064 7352
rect 3169 7100 3477 7109
rect 3169 7098 3175 7100
rect 3231 7098 3255 7100
rect 3311 7098 3335 7100
rect 3391 7098 3415 7100
rect 3471 7098 3477 7100
rect 3231 7046 3233 7098
rect 3413 7046 3415 7098
rect 3169 7044 3175 7046
rect 3231 7044 3255 7046
rect 3311 7044 3335 7046
rect 3391 7044 3415 7046
rect 3471 7044 3477 7046
rect 3169 7035 3477 7044
rect 5388 6556 5696 6565
rect 5388 6554 5394 6556
rect 5450 6554 5474 6556
rect 5530 6554 5554 6556
rect 5610 6554 5634 6556
rect 5690 6554 5696 6556
rect 5450 6502 5452 6554
rect 5632 6502 5634 6554
rect 5388 6500 5394 6502
rect 5450 6500 5474 6502
rect 5530 6500 5554 6502
rect 5610 6500 5634 6502
rect 5690 6500 5696 6502
rect 5388 6491 5696 6500
rect 3169 6012 3477 6021
rect 3169 6010 3175 6012
rect 3231 6010 3255 6012
rect 3311 6010 3335 6012
rect 3391 6010 3415 6012
rect 3471 6010 3477 6012
rect 3231 5958 3233 6010
rect 3413 5958 3415 6010
rect 3169 5956 3175 5958
rect 3231 5956 3255 5958
rect 3311 5956 3335 5958
rect 3391 5956 3415 5958
rect 3471 5956 3477 5958
rect 3169 5947 3477 5956
rect 6920 5704 6972 5710
rect 6920 5646 6972 5652
rect 4620 5568 4672 5574
rect 4620 5510 4672 5516
rect 4436 5296 4488 5302
rect 4436 5238 4488 5244
rect 3056 5160 3108 5166
rect 3056 5102 3108 5108
rect 3068 4758 3096 5102
rect 4252 5092 4304 5098
rect 4252 5034 4304 5040
rect 4160 5024 4212 5030
rect 4160 4966 4212 4972
rect 3169 4924 3477 4933
rect 3169 4922 3175 4924
rect 3231 4922 3255 4924
rect 3311 4922 3335 4924
rect 3391 4922 3415 4924
rect 3471 4922 3477 4924
rect 3231 4870 3233 4922
rect 3413 4870 3415 4922
rect 3169 4868 3175 4870
rect 3231 4868 3255 4870
rect 3311 4868 3335 4870
rect 3391 4868 3415 4870
rect 3471 4868 3477 4870
rect 3169 4859 3477 4868
rect 3056 4752 3108 4758
rect 3056 4694 3108 4700
rect 2780 4616 2832 4622
rect 2780 4558 2832 4564
rect 2228 4480 2280 4486
rect 2228 4422 2280 4428
rect 2240 4146 2268 4422
rect 2228 4140 2280 4146
rect 2228 4082 2280 4088
rect 2792 4060 2820 4558
rect 2700 4032 2820 4060
rect 2504 3936 2556 3942
rect 2504 3878 2556 3884
rect 2516 3602 2544 3878
rect 2504 3596 2556 3602
rect 2504 3538 2556 3544
rect 1952 3188 2004 3194
rect 1952 3130 2004 3136
rect 1964 2378 1992 3130
rect 2516 2514 2544 3538
rect 2504 2508 2556 2514
rect 2504 2450 2556 2456
rect 2700 2394 2728 4032
rect 4172 3942 4200 4966
rect 4160 3936 4212 3942
rect 4160 3878 4212 3884
rect 3169 3836 3477 3845
rect 3169 3834 3175 3836
rect 3231 3834 3255 3836
rect 3311 3834 3335 3836
rect 3391 3834 3415 3836
rect 3471 3834 3477 3836
rect 3231 3782 3233 3834
rect 3413 3782 3415 3834
rect 3169 3780 3175 3782
rect 3231 3780 3255 3782
rect 3311 3780 3335 3782
rect 3391 3780 3415 3782
rect 3471 3780 3477 3782
rect 3169 3771 3477 3780
rect 4172 3738 4200 3878
rect 4160 3732 4212 3738
rect 4160 3674 4212 3680
rect 2964 3392 3016 3398
rect 2964 3334 3016 3340
rect 2976 3126 3004 3334
rect 2964 3120 3016 3126
rect 2964 3062 3016 3068
rect 4172 3058 4200 3674
rect 4264 3126 4292 5034
rect 4448 4486 4476 5238
rect 4436 4480 4488 4486
rect 4436 4422 4488 4428
rect 4448 4214 4476 4422
rect 4436 4208 4488 4214
rect 4436 4150 4488 4156
rect 4448 3466 4476 4150
rect 4528 4004 4580 4010
rect 4528 3946 4580 3952
rect 4436 3460 4488 3466
rect 4436 3402 4488 3408
rect 4252 3120 4304 3126
rect 4252 3062 4304 3068
rect 4540 3058 4568 3946
rect 4160 3052 4212 3058
rect 4160 2994 4212 3000
rect 4528 3052 4580 3058
rect 4528 2994 4580 3000
rect 3169 2748 3477 2757
rect 3169 2746 3175 2748
rect 3231 2746 3255 2748
rect 3311 2746 3335 2748
rect 3391 2746 3415 2748
rect 3471 2746 3477 2748
rect 3231 2694 3233 2746
rect 3413 2694 3415 2746
rect 3169 2692 3175 2694
rect 3231 2692 3255 2694
rect 3311 2692 3335 2694
rect 3391 2692 3415 2694
rect 3471 2692 3477 2694
rect 3169 2683 3477 2692
rect 4172 2514 4200 2994
rect 4632 2514 4660 5510
rect 5388 5468 5696 5477
rect 5388 5466 5394 5468
rect 5450 5466 5474 5468
rect 5530 5466 5554 5468
rect 5610 5466 5634 5468
rect 5690 5466 5696 5468
rect 5450 5414 5452 5466
rect 5632 5414 5634 5466
rect 5388 5412 5394 5414
rect 5450 5412 5474 5414
rect 5530 5412 5554 5414
rect 5610 5412 5634 5414
rect 5690 5412 5696 5414
rect 5388 5403 5696 5412
rect 6736 5228 6788 5234
rect 6736 5170 6788 5176
rect 4988 4548 5040 4554
rect 4988 4490 5040 4496
rect 6184 4548 6236 4554
rect 6184 4490 6236 4496
rect 5000 4282 5028 4490
rect 5388 4380 5696 4389
rect 5388 4378 5394 4380
rect 5450 4378 5474 4380
rect 5530 4378 5554 4380
rect 5610 4378 5634 4380
rect 5690 4378 5696 4380
rect 5450 4326 5452 4378
rect 5632 4326 5634 4378
rect 5388 4324 5394 4326
rect 5450 4324 5474 4326
rect 5530 4324 5554 4326
rect 5610 4324 5634 4326
rect 5690 4324 5696 4326
rect 5388 4315 5696 4324
rect 6196 4282 6224 4490
rect 4988 4276 5040 4282
rect 4988 4218 5040 4224
rect 6184 4276 6236 4282
rect 6184 4218 6236 4224
rect 4712 4140 4764 4146
rect 4712 4082 4764 4088
rect 4724 3942 4752 4082
rect 5000 3942 5028 4218
rect 5264 4208 5316 4214
rect 5264 4150 5316 4156
rect 4712 3936 4764 3942
rect 4712 3878 4764 3884
rect 4988 3936 5040 3942
rect 4988 3878 5040 3884
rect 5276 2990 5304 4150
rect 6748 3738 6776 5170
rect 6828 5024 6880 5030
rect 6828 4966 6880 4972
rect 6840 4622 6868 4966
rect 6932 4826 6960 5646
rect 7024 5370 7052 7346
rect 7012 5364 7064 5370
rect 7012 5306 7064 5312
rect 6920 4820 6972 4826
rect 6920 4762 6972 4768
rect 6828 4616 6880 4622
rect 6828 4558 6880 4564
rect 6828 4480 6880 4486
rect 6828 4422 6880 4428
rect 6840 4146 6868 4422
rect 6828 4140 6880 4146
rect 6828 4082 6880 4088
rect 6920 4004 6972 4010
rect 6920 3946 6972 3952
rect 6736 3732 6788 3738
rect 6736 3674 6788 3680
rect 6748 3534 6776 3674
rect 6736 3528 6788 3534
rect 6736 3470 6788 3476
rect 6932 3398 6960 3946
rect 6920 3392 6972 3398
rect 6920 3334 6972 3340
rect 5388 3292 5696 3301
rect 5388 3290 5394 3292
rect 5450 3290 5474 3292
rect 5530 3290 5554 3292
rect 5610 3290 5634 3292
rect 5690 3290 5696 3292
rect 5450 3238 5452 3290
rect 5632 3238 5634 3290
rect 5388 3236 5394 3238
rect 5450 3236 5474 3238
rect 5530 3236 5554 3238
rect 5610 3236 5634 3238
rect 5690 3236 5696 3238
rect 5388 3227 5696 3236
rect 5264 2984 5316 2990
rect 5264 2926 5316 2932
rect 4160 2508 4212 2514
rect 4160 2450 4212 2456
rect 4620 2508 4672 2514
rect 4620 2450 4672 2456
rect 1952 2372 2004 2378
rect 1952 2314 2004 2320
rect 2516 2366 2728 2394
rect 2516 800 2544 2366
rect 5276 2310 5304 2926
rect 7024 2650 7052 5306
rect 7300 4486 7328 7414
rect 7472 7404 7524 7410
rect 7472 7346 7524 7352
rect 13820 7404 13872 7410
rect 13820 7346 13872 7352
rect 16856 7404 16908 7410
rect 16856 7346 16908 7352
rect 7484 5642 7512 7346
rect 7932 7336 7984 7342
rect 7932 7278 7984 7284
rect 13360 7336 13412 7342
rect 13360 7278 13412 7284
rect 7608 7100 7916 7109
rect 7608 7098 7614 7100
rect 7670 7098 7694 7100
rect 7750 7098 7774 7100
rect 7830 7098 7854 7100
rect 7910 7098 7916 7100
rect 7670 7046 7672 7098
rect 7852 7046 7854 7098
rect 7608 7044 7614 7046
rect 7670 7044 7694 7046
rect 7750 7044 7774 7046
rect 7830 7044 7854 7046
rect 7910 7044 7916 7046
rect 7608 7035 7916 7044
rect 7608 6012 7916 6021
rect 7608 6010 7614 6012
rect 7670 6010 7694 6012
rect 7750 6010 7774 6012
rect 7830 6010 7854 6012
rect 7910 6010 7916 6012
rect 7670 5958 7672 6010
rect 7852 5958 7854 6010
rect 7608 5956 7614 5958
rect 7670 5956 7694 5958
rect 7750 5956 7774 5958
rect 7830 5956 7854 5958
rect 7910 5956 7916 5958
rect 7608 5947 7916 5956
rect 7472 5636 7524 5642
rect 7472 5578 7524 5584
rect 7380 5568 7432 5574
rect 7380 5510 7432 5516
rect 7392 5370 7420 5510
rect 7380 5364 7432 5370
rect 7380 5306 7432 5312
rect 7392 4622 7420 5306
rect 7380 4616 7432 4622
rect 7380 4558 7432 4564
rect 7288 4480 7340 4486
rect 7288 4422 7340 4428
rect 7300 4214 7328 4422
rect 7288 4208 7340 4214
rect 7288 4150 7340 4156
rect 7484 4146 7512 5578
rect 7608 4924 7916 4933
rect 7608 4922 7614 4924
rect 7670 4922 7694 4924
rect 7750 4922 7774 4924
rect 7830 4922 7854 4924
rect 7910 4922 7916 4924
rect 7670 4870 7672 4922
rect 7852 4870 7854 4922
rect 7608 4868 7614 4870
rect 7670 4868 7694 4870
rect 7750 4868 7774 4870
rect 7830 4868 7854 4870
rect 7910 4868 7916 4870
rect 7608 4859 7916 4868
rect 7840 4616 7892 4622
rect 7840 4558 7892 4564
rect 7472 4140 7524 4146
rect 7472 4082 7524 4088
rect 7852 4078 7880 4558
rect 7944 4282 7972 7278
rect 10324 7268 10376 7274
rect 10324 7210 10376 7216
rect 9827 6556 10135 6565
rect 9827 6554 9833 6556
rect 9889 6554 9913 6556
rect 9969 6554 9993 6556
rect 10049 6554 10073 6556
rect 10129 6554 10135 6556
rect 9889 6502 9891 6554
rect 10071 6502 10073 6554
rect 9827 6500 9833 6502
rect 9889 6500 9913 6502
rect 9969 6500 9993 6502
rect 10049 6500 10073 6502
rect 10129 6500 10135 6502
rect 9827 6491 10135 6500
rect 8024 6316 8076 6322
rect 8024 6258 8076 6264
rect 8208 6316 8260 6322
rect 8208 6258 8260 6264
rect 8036 5914 8064 6258
rect 8024 5908 8076 5914
rect 8024 5850 8076 5856
rect 8116 5772 8168 5778
rect 8116 5714 8168 5720
rect 8128 5166 8156 5714
rect 8116 5160 8168 5166
rect 8116 5102 8168 5108
rect 8024 4684 8076 4690
rect 8024 4626 8076 4632
rect 7932 4276 7984 4282
rect 7932 4218 7984 4224
rect 7104 4072 7156 4078
rect 7104 4014 7156 4020
rect 7840 4072 7892 4078
rect 7840 4014 7892 4020
rect 7116 3194 7144 4014
rect 7608 3836 7916 3845
rect 7608 3834 7614 3836
rect 7670 3834 7694 3836
rect 7750 3834 7774 3836
rect 7830 3834 7854 3836
rect 7910 3834 7916 3836
rect 7670 3782 7672 3834
rect 7852 3782 7854 3834
rect 7608 3780 7614 3782
rect 7670 3780 7694 3782
rect 7750 3780 7774 3782
rect 7830 3780 7854 3782
rect 7910 3780 7916 3782
rect 7608 3771 7916 3780
rect 7378 3360 7434 3369
rect 7378 3295 7434 3304
rect 7104 3188 7156 3194
rect 7104 3130 7156 3136
rect 7116 3097 7144 3130
rect 7392 3126 7420 3295
rect 7944 3194 7972 4218
rect 7932 3188 7984 3194
rect 7932 3130 7984 3136
rect 7380 3120 7432 3126
rect 7102 3088 7158 3097
rect 7380 3062 7432 3068
rect 7102 3023 7158 3032
rect 7472 2848 7524 2854
rect 7472 2790 7524 2796
rect 7012 2644 7064 2650
rect 7012 2586 7064 2592
rect 5264 2304 5316 2310
rect 5264 2246 5316 2252
rect 5388 2204 5696 2213
rect 5388 2202 5394 2204
rect 5450 2202 5474 2204
rect 5530 2202 5554 2204
rect 5610 2202 5634 2204
rect 5690 2202 5696 2204
rect 5450 2150 5452 2202
rect 5632 2150 5634 2202
rect 5388 2148 5394 2150
rect 5450 2148 5474 2150
rect 5530 2148 5554 2150
rect 5610 2148 5634 2150
rect 5690 2148 5696 2150
rect 5388 2139 5696 2148
rect 7484 800 7512 2790
rect 7608 2748 7916 2757
rect 7608 2746 7614 2748
rect 7670 2746 7694 2748
rect 7750 2746 7774 2748
rect 7830 2746 7854 2748
rect 7910 2746 7916 2748
rect 7670 2694 7672 2746
rect 7852 2694 7854 2746
rect 7608 2692 7614 2694
rect 7670 2692 7694 2694
rect 7750 2692 7774 2694
rect 7830 2692 7854 2694
rect 7910 2692 7916 2694
rect 7608 2683 7916 2692
rect 8036 2514 8064 4626
rect 8128 4554 8156 5102
rect 8220 4690 8248 6258
rect 9827 5468 10135 5477
rect 9827 5466 9833 5468
rect 9889 5466 9913 5468
rect 9969 5466 9993 5468
rect 10049 5466 10073 5468
rect 10129 5466 10135 5468
rect 9889 5414 9891 5466
rect 10071 5414 10073 5466
rect 9827 5412 9833 5414
rect 9889 5412 9913 5414
rect 9969 5412 9993 5414
rect 10049 5412 10073 5414
rect 10129 5412 10135 5414
rect 9827 5403 10135 5412
rect 10336 5302 10364 7210
rect 11060 7200 11112 7206
rect 11060 7142 11112 7148
rect 10968 6112 11020 6118
rect 10968 6054 11020 6060
rect 10324 5296 10376 5302
rect 10324 5238 10376 5244
rect 9220 5228 9272 5234
rect 9220 5170 9272 5176
rect 8300 4752 8352 4758
rect 8300 4694 8352 4700
rect 8208 4684 8260 4690
rect 8208 4626 8260 4632
rect 8116 4548 8168 4554
rect 8116 4490 8168 4496
rect 8128 2774 8156 4490
rect 8312 3534 8340 4694
rect 9036 4616 9088 4622
rect 9036 4558 9088 4564
rect 8392 4548 8444 4554
rect 8392 4490 8444 4496
rect 8404 4282 8432 4490
rect 8852 4480 8904 4486
rect 8852 4422 8904 4428
rect 8392 4276 8444 4282
rect 8392 4218 8444 4224
rect 8864 4214 8892 4422
rect 9048 4282 9076 4558
rect 9036 4276 9088 4282
rect 9036 4218 9088 4224
rect 8852 4208 8904 4214
rect 8852 4150 8904 4156
rect 8484 4004 8536 4010
rect 8484 3946 8536 3952
rect 8496 3670 8524 3946
rect 9128 3936 9180 3942
rect 9128 3878 9180 3884
rect 8484 3664 8536 3670
rect 8484 3606 8536 3612
rect 9140 3534 9168 3878
rect 9232 3670 9260 5170
rect 9680 5160 9732 5166
rect 9680 5102 9732 5108
rect 9312 5024 9364 5030
rect 9312 4966 9364 4972
rect 9324 4554 9352 4966
rect 9588 4616 9640 4622
rect 9588 4558 9640 4564
rect 9312 4548 9364 4554
rect 9312 4490 9364 4496
rect 9404 4480 9456 4486
rect 9404 4422 9456 4428
rect 9416 4214 9444 4422
rect 9404 4208 9456 4214
rect 9404 4150 9456 4156
rect 9404 3936 9456 3942
rect 9404 3878 9456 3884
rect 9220 3664 9272 3670
rect 9220 3606 9272 3612
rect 8300 3528 8352 3534
rect 8300 3470 8352 3476
rect 9128 3528 9180 3534
rect 9128 3470 9180 3476
rect 8312 3369 8340 3470
rect 8668 3392 8720 3398
rect 8298 3360 8354 3369
rect 8668 3334 8720 3340
rect 8298 3295 8354 3304
rect 8680 3126 8708 3334
rect 9232 3194 9260 3606
rect 9416 3602 9444 3878
rect 9404 3596 9456 3602
rect 9404 3538 9456 3544
rect 9220 3188 9272 3194
rect 9220 3130 9272 3136
rect 8668 3120 8720 3126
rect 8668 3062 8720 3068
rect 9034 3088 9090 3097
rect 9034 3023 9036 3032
rect 9088 3023 9090 3032
rect 9036 2994 9088 3000
rect 9232 2774 9260 3130
rect 9416 3126 9444 3538
rect 9404 3120 9456 3126
rect 9404 3062 9456 3068
rect 9600 2854 9628 4558
rect 9588 2848 9640 2854
rect 9588 2790 9640 2796
rect 8128 2746 8248 2774
rect 9232 2746 9352 2774
rect 8220 2650 8248 2746
rect 8208 2644 8260 2650
rect 8208 2586 8260 2592
rect 8024 2508 8076 2514
rect 8024 2450 8076 2456
rect 9324 2310 9352 2746
rect 9692 2666 9720 5102
rect 10336 4690 10364 5238
rect 10508 5024 10560 5030
rect 10508 4966 10560 4972
rect 10324 4684 10376 4690
rect 10324 4626 10376 4632
rect 10520 4622 10548 4966
rect 10980 4622 11008 6054
rect 11072 5370 11100 7142
rect 12047 7100 12355 7109
rect 12047 7098 12053 7100
rect 12109 7098 12133 7100
rect 12189 7098 12213 7100
rect 12269 7098 12293 7100
rect 12349 7098 12355 7100
rect 12109 7046 12111 7098
rect 12291 7046 12293 7098
rect 12047 7044 12053 7046
rect 12109 7044 12133 7046
rect 12189 7044 12213 7046
rect 12269 7044 12293 7046
rect 12349 7044 12355 7046
rect 12047 7035 12355 7044
rect 12047 6012 12355 6021
rect 12047 6010 12053 6012
rect 12109 6010 12133 6012
rect 12189 6010 12213 6012
rect 12269 6010 12293 6012
rect 12349 6010 12355 6012
rect 12109 5958 12111 6010
rect 12291 5958 12293 6010
rect 12047 5956 12053 5958
rect 12109 5956 12133 5958
rect 12189 5956 12213 5958
rect 12269 5956 12293 5958
rect 12349 5956 12355 5958
rect 12047 5947 12355 5956
rect 11520 5636 11572 5642
rect 11520 5578 11572 5584
rect 11704 5636 11756 5642
rect 11704 5578 11756 5584
rect 12808 5636 12860 5642
rect 12808 5578 12860 5584
rect 12900 5636 12952 5642
rect 12900 5578 12952 5584
rect 11532 5370 11560 5578
rect 11060 5364 11112 5370
rect 11520 5364 11572 5370
rect 11112 5324 11192 5352
rect 11060 5306 11112 5312
rect 10508 4616 10560 4622
rect 10508 4558 10560 4564
rect 10968 4616 11020 4622
rect 10968 4558 11020 4564
rect 10692 4548 10744 4554
rect 10692 4490 10744 4496
rect 10232 4480 10284 4486
rect 10232 4422 10284 4428
rect 9827 4380 10135 4389
rect 9827 4378 9833 4380
rect 9889 4378 9913 4380
rect 9969 4378 9993 4380
rect 10049 4378 10073 4380
rect 10129 4378 10135 4380
rect 9889 4326 9891 4378
rect 10071 4326 10073 4378
rect 9827 4324 9833 4326
rect 9889 4324 9913 4326
rect 9969 4324 9993 4326
rect 10049 4324 10073 4326
rect 10129 4324 10135 4326
rect 9827 4315 10135 4324
rect 10244 3534 10272 4422
rect 10232 3528 10284 3534
rect 10232 3470 10284 3476
rect 9827 3292 10135 3301
rect 9827 3290 9833 3292
rect 9889 3290 9913 3292
rect 9969 3290 9993 3292
rect 10049 3290 10073 3292
rect 10129 3290 10135 3292
rect 9889 3238 9891 3290
rect 10071 3238 10073 3290
rect 9827 3236 9833 3238
rect 9889 3236 9913 3238
rect 9969 3236 9993 3238
rect 10049 3236 10073 3238
rect 10129 3236 10135 3238
rect 9827 3227 10135 3236
rect 10704 3058 10732 4490
rect 10968 4480 11020 4486
rect 10968 4422 11020 4428
rect 11060 4480 11112 4486
rect 11060 4422 11112 4428
rect 10980 3534 11008 4422
rect 11072 4078 11100 4422
rect 11164 4282 11192 5324
rect 11520 5306 11572 5312
rect 11716 4690 11744 5578
rect 12440 5364 12492 5370
rect 12440 5306 12492 5312
rect 11888 5160 11940 5166
rect 11808 5108 11888 5114
rect 11808 5102 11940 5108
rect 11808 5086 11928 5102
rect 11704 4684 11756 4690
rect 11704 4626 11756 4632
rect 11152 4276 11204 4282
rect 11152 4218 11204 4224
rect 11060 4072 11112 4078
rect 11060 4014 11112 4020
rect 11152 4072 11204 4078
rect 11152 4014 11204 4020
rect 11164 3670 11192 4014
rect 11152 3664 11204 3670
rect 11152 3606 11204 3612
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 11716 3466 11744 4626
rect 11808 4214 11836 5086
rect 12047 4924 12355 4933
rect 12047 4922 12053 4924
rect 12109 4922 12133 4924
rect 12189 4922 12213 4924
rect 12269 4922 12293 4924
rect 12349 4922 12355 4924
rect 12109 4870 12111 4922
rect 12291 4870 12293 4922
rect 12047 4868 12053 4870
rect 12109 4868 12133 4870
rect 12189 4868 12213 4870
rect 12269 4868 12293 4870
rect 12349 4868 12355 4870
rect 12047 4859 12355 4868
rect 11980 4752 12032 4758
rect 12348 4752 12400 4758
rect 12032 4700 12348 4706
rect 11980 4694 12400 4700
rect 11992 4678 12388 4694
rect 12452 4690 12480 5306
rect 12820 4826 12848 5578
rect 12912 5166 12940 5578
rect 13084 5568 13136 5574
rect 13084 5510 13136 5516
rect 12992 5228 13044 5234
rect 12992 5170 13044 5176
rect 12900 5160 12952 5166
rect 12900 5102 12952 5108
rect 12808 4820 12860 4826
rect 12808 4762 12860 4768
rect 12440 4684 12492 4690
rect 12440 4626 12492 4632
rect 12348 4616 12400 4622
rect 12348 4558 12400 4564
rect 11888 4548 11940 4554
rect 11888 4490 11940 4496
rect 11900 4282 11928 4490
rect 12360 4486 12388 4558
rect 12348 4480 12400 4486
rect 12348 4422 12400 4428
rect 11888 4276 11940 4282
rect 11888 4218 11940 4224
rect 11796 4208 11848 4214
rect 11796 4150 11848 4156
rect 11808 3670 11836 4150
rect 11888 4140 11940 4146
rect 11888 4082 11940 4088
rect 11900 4049 11928 4082
rect 11886 4040 11942 4049
rect 11886 3975 11942 3984
rect 12047 3836 12355 3845
rect 12047 3834 12053 3836
rect 12109 3834 12133 3836
rect 12189 3834 12213 3836
rect 12269 3834 12293 3836
rect 12349 3834 12355 3836
rect 12109 3782 12111 3834
rect 12291 3782 12293 3834
rect 12047 3780 12053 3782
rect 12109 3780 12133 3782
rect 12189 3780 12213 3782
rect 12269 3780 12293 3782
rect 12349 3780 12355 3782
rect 12047 3771 12355 3780
rect 11796 3664 11848 3670
rect 11796 3606 11848 3612
rect 11704 3460 11756 3466
rect 11704 3402 11756 3408
rect 10876 3188 10928 3194
rect 10876 3130 10928 3136
rect 10692 3052 10744 3058
rect 10692 2994 10744 3000
rect 9600 2638 9720 2666
rect 9600 2582 9628 2638
rect 9588 2576 9640 2582
rect 9588 2518 9640 2524
rect 9312 2304 9364 2310
rect 9312 2246 9364 2252
rect 9827 2204 10135 2213
rect 9827 2202 9833 2204
rect 9889 2202 9913 2204
rect 9969 2202 9993 2204
rect 10049 2202 10073 2204
rect 10129 2202 10135 2204
rect 9889 2150 9891 2202
rect 10071 2150 10073 2202
rect 9827 2148 9833 2150
rect 9889 2148 9913 2150
rect 9969 2148 9993 2150
rect 10049 2148 10073 2150
rect 10129 2148 10135 2150
rect 9827 2139 10135 2148
rect 10704 2106 10732 2994
rect 10888 2922 10916 3130
rect 11716 2922 11744 3402
rect 10876 2916 10928 2922
rect 10876 2858 10928 2864
rect 11704 2916 11756 2922
rect 11704 2858 11756 2864
rect 10888 2446 10916 2858
rect 11808 2774 11836 3606
rect 12716 3460 12768 3466
rect 12716 3402 12768 3408
rect 12728 3126 12756 3402
rect 12912 3126 12940 5102
rect 13004 3942 13032 5170
rect 13096 4622 13124 5510
rect 13372 5234 13400 7278
rect 13832 5302 13860 7346
rect 16486 7100 16794 7109
rect 16486 7098 16492 7100
rect 16548 7098 16572 7100
rect 16628 7098 16652 7100
rect 16708 7098 16732 7100
rect 16788 7098 16794 7100
rect 16548 7046 16550 7098
rect 16730 7046 16732 7098
rect 16486 7044 16492 7046
rect 16548 7044 16572 7046
rect 16628 7044 16652 7046
rect 16708 7044 16732 7046
rect 16788 7044 16794 7046
rect 16486 7035 16794 7044
rect 14266 6556 14574 6565
rect 14266 6554 14272 6556
rect 14328 6554 14352 6556
rect 14408 6554 14432 6556
rect 14488 6554 14512 6556
rect 14568 6554 14574 6556
rect 14328 6502 14330 6554
rect 14510 6502 14512 6554
rect 14266 6500 14272 6502
rect 14328 6500 14352 6502
rect 14408 6500 14432 6502
rect 14488 6500 14512 6502
rect 14568 6500 14574 6502
rect 14266 6491 14574 6500
rect 16486 6012 16794 6021
rect 16486 6010 16492 6012
rect 16548 6010 16572 6012
rect 16628 6010 16652 6012
rect 16708 6010 16732 6012
rect 16788 6010 16794 6012
rect 16548 5958 16550 6010
rect 16730 5958 16732 6010
rect 16486 5956 16492 5958
rect 16548 5956 16572 5958
rect 16628 5956 16652 5958
rect 16708 5956 16732 5958
rect 16788 5956 16794 5958
rect 16486 5947 16794 5956
rect 15108 5568 15160 5574
rect 15108 5510 15160 5516
rect 14266 5468 14574 5477
rect 14266 5466 14272 5468
rect 14328 5466 14352 5468
rect 14408 5466 14432 5468
rect 14488 5466 14512 5468
rect 14568 5466 14574 5468
rect 14328 5414 14330 5466
rect 14510 5414 14512 5466
rect 14266 5412 14272 5414
rect 14328 5412 14352 5414
rect 14408 5412 14432 5414
rect 14488 5412 14512 5414
rect 14568 5412 14574 5414
rect 14266 5403 14574 5412
rect 13820 5296 13872 5302
rect 13820 5238 13872 5244
rect 13360 5228 13412 5234
rect 13360 5170 13412 5176
rect 13912 5092 13964 5098
rect 13912 5034 13964 5040
rect 13728 4752 13780 4758
rect 13728 4694 13780 4700
rect 13084 4616 13136 4622
rect 13084 4558 13136 4564
rect 13636 4072 13688 4078
rect 13082 4040 13138 4049
rect 13636 4014 13688 4020
rect 13082 3975 13138 3984
rect 13096 3942 13124 3975
rect 12992 3936 13044 3942
rect 12992 3878 13044 3884
rect 13084 3936 13136 3942
rect 13084 3878 13136 3884
rect 13452 3596 13504 3602
rect 13648 3584 13676 4014
rect 13740 4010 13768 4694
rect 13728 4004 13780 4010
rect 13728 3946 13780 3952
rect 13728 3596 13780 3602
rect 13648 3556 13728 3584
rect 13452 3538 13504 3544
rect 13728 3538 13780 3544
rect 13464 3126 13492 3538
rect 13740 3194 13768 3538
rect 13728 3188 13780 3194
rect 13728 3130 13780 3136
rect 12716 3120 12768 3126
rect 12716 3062 12768 3068
rect 12900 3120 12952 3126
rect 12900 3062 12952 3068
rect 13452 3120 13504 3126
rect 13452 3062 13504 3068
rect 12440 2848 12492 2854
rect 12440 2790 12492 2796
rect 11716 2746 11836 2774
rect 12047 2748 12355 2757
rect 12047 2746 12053 2748
rect 12109 2746 12133 2748
rect 12189 2746 12213 2748
rect 12269 2746 12293 2748
rect 12349 2746 12355 2748
rect 11716 2514 11744 2746
rect 12109 2694 12111 2746
rect 12291 2694 12293 2746
rect 12047 2692 12053 2694
rect 12109 2692 12133 2694
rect 12189 2692 12213 2694
rect 12269 2692 12293 2694
rect 12349 2692 12355 2694
rect 12047 2683 12355 2692
rect 11704 2508 11756 2514
rect 11704 2450 11756 2456
rect 10876 2440 10928 2446
rect 10876 2382 10928 2388
rect 10692 2100 10744 2106
rect 10692 2042 10744 2048
rect 12452 800 12480 2790
rect 12728 2310 12756 3062
rect 12912 2650 12940 3062
rect 13740 2990 13768 3130
rect 13924 3058 13952 5034
rect 15120 4690 15148 5510
rect 15200 5024 15252 5030
rect 15200 4966 15252 4972
rect 15108 4684 15160 4690
rect 15108 4626 15160 4632
rect 15212 4622 15240 4966
rect 16486 4924 16794 4933
rect 16486 4922 16492 4924
rect 16548 4922 16572 4924
rect 16628 4922 16652 4924
rect 16708 4922 16732 4924
rect 16788 4922 16794 4924
rect 16548 4870 16550 4922
rect 16730 4870 16732 4922
rect 16486 4868 16492 4870
rect 16548 4868 16572 4870
rect 16628 4868 16652 4870
rect 16708 4868 16732 4870
rect 16788 4868 16794 4870
rect 16486 4859 16794 4868
rect 16868 4758 16896 7346
rect 18705 6556 19013 6565
rect 18705 6554 18711 6556
rect 18767 6554 18791 6556
rect 18847 6554 18871 6556
rect 18927 6554 18951 6556
rect 19007 6554 19013 6556
rect 18767 6502 18769 6554
rect 18949 6502 18951 6554
rect 18705 6500 18711 6502
rect 18767 6500 18791 6502
rect 18847 6500 18871 6502
rect 18927 6500 18951 6502
rect 19007 6500 19013 6502
rect 18705 6491 19013 6500
rect 18705 5468 19013 5477
rect 18705 5466 18711 5468
rect 18767 5466 18791 5468
rect 18847 5466 18871 5468
rect 18927 5466 18951 5468
rect 19007 5466 19013 5468
rect 18767 5414 18769 5466
rect 18949 5414 18951 5466
rect 18705 5412 18711 5414
rect 18767 5412 18791 5414
rect 18847 5412 18871 5414
rect 18927 5412 18951 5414
rect 19007 5412 19013 5414
rect 18705 5403 19013 5412
rect 16856 4752 16908 4758
rect 16856 4694 16908 4700
rect 15200 4616 15252 4622
rect 15200 4558 15252 4564
rect 15384 4548 15436 4554
rect 15384 4490 15436 4496
rect 14266 4380 14574 4389
rect 14266 4378 14272 4380
rect 14328 4378 14352 4380
rect 14408 4378 14432 4380
rect 14488 4378 14512 4380
rect 14568 4378 14574 4380
rect 14328 4326 14330 4378
rect 14510 4326 14512 4378
rect 14266 4324 14272 4326
rect 14328 4324 14352 4326
rect 14408 4324 14432 4326
rect 14488 4324 14512 4326
rect 14568 4324 14574 4326
rect 14266 4315 14574 4324
rect 14266 3292 14574 3301
rect 14266 3290 14272 3292
rect 14328 3290 14352 3292
rect 14408 3290 14432 3292
rect 14488 3290 14512 3292
rect 14568 3290 14574 3292
rect 14328 3238 14330 3290
rect 14510 3238 14512 3290
rect 14266 3236 14272 3238
rect 14328 3236 14352 3238
rect 14408 3236 14432 3238
rect 14488 3236 14512 3238
rect 14568 3236 14574 3238
rect 14266 3227 14574 3236
rect 13912 3052 13964 3058
rect 13912 2994 13964 3000
rect 13728 2984 13780 2990
rect 13728 2926 13780 2932
rect 12900 2644 12952 2650
rect 12900 2586 12952 2592
rect 13740 2514 13768 2926
rect 15396 2922 15424 4490
rect 16028 4480 16080 4486
rect 16028 4422 16080 4428
rect 16856 4480 16908 4486
rect 16856 4422 16908 4428
rect 16040 3738 16068 4422
rect 16486 3836 16794 3845
rect 16486 3834 16492 3836
rect 16548 3834 16572 3836
rect 16628 3834 16652 3836
rect 16708 3834 16732 3836
rect 16788 3834 16794 3836
rect 16548 3782 16550 3834
rect 16730 3782 16732 3834
rect 16486 3780 16492 3782
rect 16548 3780 16572 3782
rect 16628 3780 16652 3782
rect 16708 3780 16732 3782
rect 16788 3780 16794 3782
rect 16486 3771 16794 3780
rect 16028 3732 16080 3738
rect 16028 3674 16080 3680
rect 16868 2922 16896 4422
rect 18705 4380 19013 4389
rect 18705 4378 18711 4380
rect 18767 4378 18791 4380
rect 18847 4378 18871 4380
rect 18927 4378 18951 4380
rect 19007 4378 19013 4380
rect 18767 4326 18769 4378
rect 18949 4326 18951 4378
rect 18705 4324 18711 4326
rect 18767 4324 18791 4326
rect 18847 4324 18871 4326
rect 18927 4324 18951 4326
rect 19007 4324 19013 4326
rect 18705 4315 19013 4324
rect 18705 3292 19013 3301
rect 18705 3290 18711 3292
rect 18767 3290 18791 3292
rect 18847 3290 18871 3292
rect 18927 3290 18951 3292
rect 19007 3290 19013 3292
rect 18767 3238 18769 3290
rect 18949 3238 18951 3290
rect 18705 3236 18711 3238
rect 18767 3236 18791 3238
rect 18847 3236 18871 3238
rect 18927 3236 18951 3238
rect 19007 3236 19013 3238
rect 18705 3227 19013 3236
rect 15384 2916 15436 2922
rect 15384 2858 15436 2864
rect 15752 2916 15804 2922
rect 15752 2858 15804 2864
rect 16856 2916 16908 2922
rect 16856 2858 16908 2864
rect 13728 2508 13780 2514
rect 13728 2450 13780 2456
rect 15764 2378 15792 2858
rect 16486 2748 16794 2757
rect 16486 2746 16492 2748
rect 16548 2746 16572 2748
rect 16628 2746 16652 2748
rect 16708 2746 16732 2748
rect 16788 2746 16794 2748
rect 16548 2694 16550 2746
rect 16730 2694 16732 2746
rect 16486 2692 16492 2694
rect 16548 2692 16572 2694
rect 16628 2692 16652 2694
rect 16708 2692 16732 2694
rect 16788 2692 16794 2694
rect 16486 2683 16794 2692
rect 17500 2440 17552 2446
rect 17500 2382 17552 2388
rect 15752 2372 15804 2378
rect 15752 2314 15804 2320
rect 12716 2304 12768 2310
rect 12716 2246 12768 2252
rect 17408 2304 17460 2310
rect 17408 2246 17460 2252
rect 14266 2204 14574 2213
rect 14266 2202 14272 2204
rect 14328 2202 14352 2204
rect 14408 2202 14432 2204
rect 14488 2202 14512 2204
rect 14568 2202 14574 2204
rect 14328 2150 14330 2202
rect 14510 2150 14512 2202
rect 14266 2148 14272 2150
rect 14328 2148 14352 2150
rect 14408 2148 14432 2150
rect 14488 2148 14512 2150
rect 14568 2148 14574 2150
rect 14266 2139 14574 2148
rect 17420 800 17448 2246
rect 17512 2106 17540 2382
rect 18705 2204 19013 2213
rect 18705 2202 18711 2204
rect 18767 2202 18791 2204
rect 18847 2202 18871 2204
rect 18927 2202 18951 2204
rect 19007 2202 19013 2204
rect 18767 2150 18769 2202
rect 18949 2150 18951 2202
rect 18705 2148 18711 2150
rect 18767 2148 18791 2150
rect 18847 2148 18871 2150
rect 18927 2148 18951 2150
rect 19007 2148 19013 2150
rect 18705 2139 19013 2148
rect 17500 2100 17552 2106
rect 17500 2042 17552 2048
rect 2502 0 2558 800
rect 7470 0 7526 800
rect 12438 0 12494 800
rect 17406 0 17462 800
<< via2 >>
rect 5394 7642 5450 7644
rect 5474 7642 5530 7644
rect 5554 7642 5610 7644
rect 5634 7642 5690 7644
rect 5394 7590 5440 7642
rect 5440 7590 5450 7642
rect 5474 7590 5504 7642
rect 5504 7590 5516 7642
rect 5516 7590 5530 7642
rect 5554 7590 5568 7642
rect 5568 7590 5580 7642
rect 5580 7590 5610 7642
rect 5634 7590 5644 7642
rect 5644 7590 5690 7642
rect 5394 7588 5450 7590
rect 5474 7588 5530 7590
rect 5554 7588 5610 7590
rect 5634 7588 5690 7590
rect 9833 7642 9889 7644
rect 9913 7642 9969 7644
rect 9993 7642 10049 7644
rect 10073 7642 10129 7644
rect 9833 7590 9879 7642
rect 9879 7590 9889 7642
rect 9913 7590 9943 7642
rect 9943 7590 9955 7642
rect 9955 7590 9969 7642
rect 9993 7590 10007 7642
rect 10007 7590 10019 7642
rect 10019 7590 10049 7642
rect 10073 7590 10083 7642
rect 10083 7590 10129 7642
rect 9833 7588 9889 7590
rect 9913 7588 9969 7590
rect 9993 7588 10049 7590
rect 10073 7588 10129 7590
rect 14272 7642 14328 7644
rect 14352 7642 14408 7644
rect 14432 7642 14488 7644
rect 14512 7642 14568 7644
rect 14272 7590 14318 7642
rect 14318 7590 14328 7642
rect 14352 7590 14382 7642
rect 14382 7590 14394 7642
rect 14394 7590 14408 7642
rect 14432 7590 14446 7642
rect 14446 7590 14458 7642
rect 14458 7590 14488 7642
rect 14512 7590 14522 7642
rect 14522 7590 14568 7642
rect 14272 7588 14328 7590
rect 14352 7588 14408 7590
rect 14432 7588 14488 7590
rect 14512 7588 14568 7590
rect 18711 7642 18767 7644
rect 18791 7642 18847 7644
rect 18871 7642 18927 7644
rect 18951 7642 19007 7644
rect 18711 7590 18757 7642
rect 18757 7590 18767 7642
rect 18791 7590 18821 7642
rect 18821 7590 18833 7642
rect 18833 7590 18847 7642
rect 18871 7590 18885 7642
rect 18885 7590 18897 7642
rect 18897 7590 18927 7642
rect 18951 7590 18961 7642
rect 18961 7590 19007 7642
rect 18711 7588 18767 7590
rect 18791 7588 18847 7590
rect 18871 7588 18927 7590
rect 18951 7588 19007 7590
rect 3175 7098 3231 7100
rect 3255 7098 3311 7100
rect 3335 7098 3391 7100
rect 3415 7098 3471 7100
rect 3175 7046 3221 7098
rect 3221 7046 3231 7098
rect 3255 7046 3285 7098
rect 3285 7046 3297 7098
rect 3297 7046 3311 7098
rect 3335 7046 3349 7098
rect 3349 7046 3361 7098
rect 3361 7046 3391 7098
rect 3415 7046 3425 7098
rect 3425 7046 3471 7098
rect 3175 7044 3231 7046
rect 3255 7044 3311 7046
rect 3335 7044 3391 7046
rect 3415 7044 3471 7046
rect 5394 6554 5450 6556
rect 5474 6554 5530 6556
rect 5554 6554 5610 6556
rect 5634 6554 5690 6556
rect 5394 6502 5440 6554
rect 5440 6502 5450 6554
rect 5474 6502 5504 6554
rect 5504 6502 5516 6554
rect 5516 6502 5530 6554
rect 5554 6502 5568 6554
rect 5568 6502 5580 6554
rect 5580 6502 5610 6554
rect 5634 6502 5644 6554
rect 5644 6502 5690 6554
rect 5394 6500 5450 6502
rect 5474 6500 5530 6502
rect 5554 6500 5610 6502
rect 5634 6500 5690 6502
rect 3175 6010 3231 6012
rect 3255 6010 3311 6012
rect 3335 6010 3391 6012
rect 3415 6010 3471 6012
rect 3175 5958 3221 6010
rect 3221 5958 3231 6010
rect 3255 5958 3285 6010
rect 3285 5958 3297 6010
rect 3297 5958 3311 6010
rect 3335 5958 3349 6010
rect 3349 5958 3361 6010
rect 3361 5958 3391 6010
rect 3415 5958 3425 6010
rect 3425 5958 3471 6010
rect 3175 5956 3231 5958
rect 3255 5956 3311 5958
rect 3335 5956 3391 5958
rect 3415 5956 3471 5958
rect 3175 4922 3231 4924
rect 3255 4922 3311 4924
rect 3335 4922 3391 4924
rect 3415 4922 3471 4924
rect 3175 4870 3221 4922
rect 3221 4870 3231 4922
rect 3255 4870 3285 4922
rect 3285 4870 3297 4922
rect 3297 4870 3311 4922
rect 3335 4870 3349 4922
rect 3349 4870 3361 4922
rect 3361 4870 3391 4922
rect 3415 4870 3425 4922
rect 3425 4870 3471 4922
rect 3175 4868 3231 4870
rect 3255 4868 3311 4870
rect 3335 4868 3391 4870
rect 3415 4868 3471 4870
rect 3175 3834 3231 3836
rect 3255 3834 3311 3836
rect 3335 3834 3391 3836
rect 3415 3834 3471 3836
rect 3175 3782 3221 3834
rect 3221 3782 3231 3834
rect 3255 3782 3285 3834
rect 3285 3782 3297 3834
rect 3297 3782 3311 3834
rect 3335 3782 3349 3834
rect 3349 3782 3361 3834
rect 3361 3782 3391 3834
rect 3415 3782 3425 3834
rect 3425 3782 3471 3834
rect 3175 3780 3231 3782
rect 3255 3780 3311 3782
rect 3335 3780 3391 3782
rect 3415 3780 3471 3782
rect 3175 2746 3231 2748
rect 3255 2746 3311 2748
rect 3335 2746 3391 2748
rect 3415 2746 3471 2748
rect 3175 2694 3221 2746
rect 3221 2694 3231 2746
rect 3255 2694 3285 2746
rect 3285 2694 3297 2746
rect 3297 2694 3311 2746
rect 3335 2694 3349 2746
rect 3349 2694 3361 2746
rect 3361 2694 3391 2746
rect 3415 2694 3425 2746
rect 3425 2694 3471 2746
rect 3175 2692 3231 2694
rect 3255 2692 3311 2694
rect 3335 2692 3391 2694
rect 3415 2692 3471 2694
rect 5394 5466 5450 5468
rect 5474 5466 5530 5468
rect 5554 5466 5610 5468
rect 5634 5466 5690 5468
rect 5394 5414 5440 5466
rect 5440 5414 5450 5466
rect 5474 5414 5504 5466
rect 5504 5414 5516 5466
rect 5516 5414 5530 5466
rect 5554 5414 5568 5466
rect 5568 5414 5580 5466
rect 5580 5414 5610 5466
rect 5634 5414 5644 5466
rect 5644 5414 5690 5466
rect 5394 5412 5450 5414
rect 5474 5412 5530 5414
rect 5554 5412 5610 5414
rect 5634 5412 5690 5414
rect 5394 4378 5450 4380
rect 5474 4378 5530 4380
rect 5554 4378 5610 4380
rect 5634 4378 5690 4380
rect 5394 4326 5440 4378
rect 5440 4326 5450 4378
rect 5474 4326 5504 4378
rect 5504 4326 5516 4378
rect 5516 4326 5530 4378
rect 5554 4326 5568 4378
rect 5568 4326 5580 4378
rect 5580 4326 5610 4378
rect 5634 4326 5644 4378
rect 5644 4326 5690 4378
rect 5394 4324 5450 4326
rect 5474 4324 5530 4326
rect 5554 4324 5610 4326
rect 5634 4324 5690 4326
rect 5394 3290 5450 3292
rect 5474 3290 5530 3292
rect 5554 3290 5610 3292
rect 5634 3290 5690 3292
rect 5394 3238 5440 3290
rect 5440 3238 5450 3290
rect 5474 3238 5504 3290
rect 5504 3238 5516 3290
rect 5516 3238 5530 3290
rect 5554 3238 5568 3290
rect 5568 3238 5580 3290
rect 5580 3238 5610 3290
rect 5634 3238 5644 3290
rect 5644 3238 5690 3290
rect 5394 3236 5450 3238
rect 5474 3236 5530 3238
rect 5554 3236 5610 3238
rect 5634 3236 5690 3238
rect 7614 7098 7670 7100
rect 7694 7098 7750 7100
rect 7774 7098 7830 7100
rect 7854 7098 7910 7100
rect 7614 7046 7660 7098
rect 7660 7046 7670 7098
rect 7694 7046 7724 7098
rect 7724 7046 7736 7098
rect 7736 7046 7750 7098
rect 7774 7046 7788 7098
rect 7788 7046 7800 7098
rect 7800 7046 7830 7098
rect 7854 7046 7864 7098
rect 7864 7046 7910 7098
rect 7614 7044 7670 7046
rect 7694 7044 7750 7046
rect 7774 7044 7830 7046
rect 7854 7044 7910 7046
rect 7614 6010 7670 6012
rect 7694 6010 7750 6012
rect 7774 6010 7830 6012
rect 7854 6010 7910 6012
rect 7614 5958 7660 6010
rect 7660 5958 7670 6010
rect 7694 5958 7724 6010
rect 7724 5958 7736 6010
rect 7736 5958 7750 6010
rect 7774 5958 7788 6010
rect 7788 5958 7800 6010
rect 7800 5958 7830 6010
rect 7854 5958 7864 6010
rect 7864 5958 7910 6010
rect 7614 5956 7670 5958
rect 7694 5956 7750 5958
rect 7774 5956 7830 5958
rect 7854 5956 7910 5958
rect 7614 4922 7670 4924
rect 7694 4922 7750 4924
rect 7774 4922 7830 4924
rect 7854 4922 7910 4924
rect 7614 4870 7660 4922
rect 7660 4870 7670 4922
rect 7694 4870 7724 4922
rect 7724 4870 7736 4922
rect 7736 4870 7750 4922
rect 7774 4870 7788 4922
rect 7788 4870 7800 4922
rect 7800 4870 7830 4922
rect 7854 4870 7864 4922
rect 7864 4870 7910 4922
rect 7614 4868 7670 4870
rect 7694 4868 7750 4870
rect 7774 4868 7830 4870
rect 7854 4868 7910 4870
rect 9833 6554 9889 6556
rect 9913 6554 9969 6556
rect 9993 6554 10049 6556
rect 10073 6554 10129 6556
rect 9833 6502 9879 6554
rect 9879 6502 9889 6554
rect 9913 6502 9943 6554
rect 9943 6502 9955 6554
rect 9955 6502 9969 6554
rect 9993 6502 10007 6554
rect 10007 6502 10019 6554
rect 10019 6502 10049 6554
rect 10073 6502 10083 6554
rect 10083 6502 10129 6554
rect 9833 6500 9889 6502
rect 9913 6500 9969 6502
rect 9993 6500 10049 6502
rect 10073 6500 10129 6502
rect 7614 3834 7670 3836
rect 7694 3834 7750 3836
rect 7774 3834 7830 3836
rect 7854 3834 7910 3836
rect 7614 3782 7660 3834
rect 7660 3782 7670 3834
rect 7694 3782 7724 3834
rect 7724 3782 7736 3834
rect 7736 3782 7750 3834
rect 7774 3782 7788 3834
rect 7788 3782 7800 3834
rect 7800 3782 7830 3834
rect 7854 3782 7864 3834
rect 7864 3782 7910 3834
rect 7614 3780 7670 3782
rect 7694 3780 7750 3782
rect 7774 3780 7830 3782
rect 7854 3780 7910 3782
rect 7378 3304 7434 3360
rect 7102 3032 7158 3088
rect 5394 2202 5450 2204
rect 5474 2202 5530 2204
rect 5554 2202 5610 2204
rect 5634 2202 5690 2204
rect 5394 2150 5440 2202
rect 5440 2150 5450 2202
rect 5474 2150 5504 2202
rect 5504 2150 5516 2202
rect 5516 2150 5530 2202
rect 5554 2150 5568 2202
rect 5568 2150 5580 2202
rect 5580 2150 5610 2202
rect 5634 2150 5644 2202
rect 5644 2150 5690 2202
rect 5394 2148 5450 2150
rect 5474 2148 5530 2150
rect 5554 2148 5610 2150
rect 5634 2148 5690 2150
rect 7614 2746 7670 2748
rect 7694 2746 7750 2748
rect 7774 2746 7830 2748
rect 7854 2746 7910 2748
rect 7614 2694 7660 2746
rect 7660 2694 7670 2746
rect 7694 2694 7724 2746
rect 7724 2694 7736 2746
rect 7736 2694 7750 2746
rect 7774 2694 7788 2746
rect 7788 2694 7800 2746
rect 7800 2694 7830 2746
rect 7854 2694 7864 2746
rect 7864 2694 7910 2746
rect 7614 2692 7670 2694
rect 7694 2692 7750 2694
rect 7774 2692 7830 2694
rect 7854 2692 7910 2694
rect 9833 5466 9889 5468
rect 9913 5466 9969 5468
rect 9993 5466 10049 5468
rect 10073 5466 10129 5468
rect 9833 5414 9879 5466
rect 9879 5414 9889 5466
rect 9913 5414 9943 5466
rect 9943 5414 9955 5466
rect 9955 5414 9969 5466
rect 9993 5414 10007 5466
rect 10007 5414 10019 5466
rect 10019 5414 10049 5466
rect 10073 5414 10083 5466
rect 10083 5414 10129 5466
rect 9833 5412 9889 5414
rect 9913 5412 9969 5414
rect 9993 5412 10049 5414
rect 10073 5412 10129 5414
rect 8298 3304 8354 3360
rect 9034 3052 9090 3088
rect 9034 3032 9036 3052
rect 9036 3032 9088 3052
rect 9088 3032 9090 3052
rect 12053 7098 12109 7100
rect 12133 7098 12189 7100
rect 12213 7098 12269 7100
rect 12293 7098 12349 7100
rect 12053 7046 12099 7098
rect 12099 7046 12109 7098
rect 12133 7046 12163 7098
rect 12163 7046 12175 7098
rect 12175 7046 12189 7098
rect 12213 7046 12227 7098
rect 12227 7046 12239 7098
rect 12239 7046 12269 7098
rect 12293 7046 12303 7098
rect 12303 7046 12349 7098
rect 12053 7044 12109 7046
rect 12133 7044 12189 7046
rect 12213 7044 12269 7046
rect 12293 7044 12349 7046
rect 12053 6010 12109 6012
rect 12133 6010 12189 6012
rect 12213 6010 12269 6012
rect 12293 6010 12349 6012
rect 12053 5958 12099 6010
rect 12099 5958 12109 6010
rect 12133 5958 12163 6010
rect 12163 5958 12175 6010
rect 12175 5958 12189 6010
rect 12213 5958 12227 6010
rect 12227 5958 12239 6010
rect 12239 5958 12269 6010
rect 12293 5958 12303 6010
rect 12303 5958 12349 6010
rect 12053 5956 12109 5958
rect 12133 5956 12189 5958
rect 12213 5956 12269 5958
rect 12293 5956 12349 5958
rect 9833 4378 9889 4380
rect 9913 4378 9969 4380
rect 9993 4378 10049 4380
rect 10073 4378 10129 4380
rect 9833 4326 9879 4378
rect 9879 4326 9889 4378
rect 9913 4326 9943 4378
rect 9943 4326 9955 4378
rect 9955 4326 9969 4378
rect 9993 4326 10007 4378
rect 10007 4326 10019 4378
rect 10019 4326 10049 4378
rect 10073 4326 10083 4378
rect 10083 4326 10129 4378
rect 9833 4324 9889 4326
rect 9913 4324 9969 4326
rect 9993 4324 10049 4326
rect 10073 4324 10129 4326
rect 9833 3290 9889 3292
rect 9913 3290 9969 3292
rect 9993 3290 10049 3292
rect 10073 3290 10129 3292
rect 9833 3238 9879 3290
rect 9879 3238 9889 3290
rect 9913 3238 9943 3290
rect 9943 3238 9955 3290
rect 9955 3238 9969 3290
rect 9993 3238 10007 3290
rect 10007 3238 10019 3290
rect 10019 3238 10049 3290
rect 10073 3238 10083 3290
rect 10083 3238 10129 3290
rect 9833 3236 9889 3238
rect 9913 3236 9969 3238
rect 9993 3236 10049 3238
rect 10073 3236 10129 3238
rect 12053 4922 12109 4924
rect 12133 4922 12189 4924
rect 12213 4922 12269 4924
rect 12293 4922 12349 4924
rect 12053 4870 12099 4922
rect 12099 4870 12109 4922
rect 12133 4870 12163 4922
rect 12163 4870 12175 4922
rect 12175 4870 12189 4922
rect 12213 4870 12227 4922
rect 12227 4870 12239 4922
rect 12239 4870 12269 4922
rect 12293 4870 12303 4922
rect 12303 4870 12349 4922
rect 12053 4868 12109 4870
rect 12133 4868 12189 4870
rect 12213 4868 12269 4870
rect 12293 4868 12349 4870
rect 11886 3984 11942 4040
rect 12053 3834 12109 3836
rect 12133 3834 12189 3836
rect 12213 3834 12269 3836
rect 12293 3834 12349 3836
rect 12053 3782 12099 3834
rect 12099 3782 12109 3834
rect 12133 3782 12163 3834
rect 12163 3782 12175 3834
rect 12175 3782 12189 3834
rect 12213 3782 12227 3834
rect 12227 3782 12239 3834
rect 12239 3782 12269 3834
rect 12293 3782 12303 3834
rect 12303 3782 12349 3834
rect 12053 3780 12109 3782
rect 12133 3780 12189 3782
rect 12213 3780 12269 3782
rect 12293 3780 12349 3782
rect 9833 2202 9889 2204
rect 9913 2202 9969 2204
rect 9993 2202 10049 2204
rect 10073 2202 10129 2204
rect 9833 2150 9879 2202
rect 9879 2150 9889 2202
rect 9913 2150 9943 2202
rect 9943 2150 9955 2202
rect 9955 2150 9969 2202
rect 9993 2150 10007 2202
rect 10007 2150 10019 2202
rect 10019 2150 10049 2202
rect 10073 2150 10083 2202
rect 10083 2150 10129 2202
rect 9833 2148 9889 2150
rect 9913 2148 9969 2150
rect 9993 2148 10049 2150
rect 10073 2148 10129 2150
rect 16492 7098 16548 7100
rect 16572 7098 16628 7100
rect 16652 7098 16708 7100
rect 16732 7098 16788 7100
rect 16492 7046 16538 7098
rect 16538 7046 16548 7098
rect 16572 7046 16602 7098
rect 16602 7046 16614 7098
rect 16614 7046 16628 7098
rect 16652 7046 16666 7098
rect 16666 7046 16678 7098
rect 16678 7046 16708 7098
rect 16732 7046 16742 7098
rect 16742 7046 16788 7098
rect 16492 7044 16548 7046
rect 16572 7044 16628 7046
rect 16652 7044 16708 7046
rect 16732 7044 16788 7046
rect 14272 6554 14328 6556
rect 14352 6554 14408 6556
rect 14432 6554 14488 6556
rect 14512 6554 14568 6556
rect 14272 6502 14318 6554
rect 14318 6502 14328 6554
rect 14352 6502 14382 6554
rect 14382 6502 14394 6554
rect 14394 6502 14408 6554
rect 14432 6502 14446 6554
rect 14446 6502 14458 6554
rect 14458 6502 14488 6554
rect 14512 6502 14522 6554
rect 14522 6502 14568 6554
rect 14272 6500 14328 6502
rect 14352 6500 14408 6502
rect 14432 6500 14488 6502
rect 14512 6500 14568 6502
rect 16492 6010 16548 6012
rect 16572 6010 16628 6012
rect 16652 6010 16708 6012
rect 16732 6010 16788 6012
rect 16492 5958 16538 6010
rect 16538 5958 16548 6010
rect 16572 5958 16602 6010
rect 16602 5958 16614 6010
rect 16614 5958 16628 6010
rect 16652 5958 16666 6010
rect 16666 5958 16678 6010
rect 16678 5958 16708 6010
rect 16732 5958 16742 6010
rect 16742 5958 16788 6010
rect 16492 5956 16548 5958
rect 16572 5956 16628 5958
rect 16652 5956 16708 5958
rect 16732 5956 16788 5958
rect 14272 5466 14328 5468
rect 14352 5466 14408 5468
rect 14432 5466 14488 5468
rect 14512 5466 14568 5468
rect 14272 5414 14318 5466
rect 14318 5414 14328 5466
rect 14352 5414 14382 5466
rect 14382 5414 14394 5466
rect 14394 5414 14408 5466
rect 14432 5414 14446 5466
rect 14446 5414 14458 5466
rect 14458 5414 14488 5466
rect 14512 5414 14522 5466
rect 14522 5414 14568 5466
rect 14272 5412 14328 5414
rect 14352 5412 14408 5414
rect 14432 5412 14488 5414
rect 14512 5412 14568 5414
rect 13082 3984 13138 4040
rect 12053 2746 12109 2748
rect 12133 2746 12189 2748
rect 12213 2746 12269 2748
rect 12293 2746 12349 2748
rect 12053 2694 12099 2746
rect 12099 2694 12109 2746
rect 12133 2694 12163 2746
rect 12163 2694 12175 2746
rect 12175 2694 12189 2746
rect 12213 2694 12227 2746
rect 12227 2694 12239 2746
rect 12239 2694 12269 2746
rect 12293 2694 12303 2746
rect 12303 2694 12349 2746
rect 12053 2692 12109 2694
rect 12133 2692 12189 2694
rect 12213 2692 12269 2694
rect 12293 2692 12349 2694
rect 16492 4922 16548 4924
rect 16572 4922 16628 4924
rect 16652 4922 16708 4924
rect 16732 4922 16788 4924
rect 16492 4870 16538 4922
rect 16538 4870 16548 4922
rect 16572 4870 16602 4922
rect 16602 4870 16614 4922
rect 16614 4870 16628 4922
rect 16652 4870 16666 4922
rect 16666 4870 16678 4922
rect 16678 4870 16708 4922
rect 16732 4870 16742 4922
rect 16742 4870 16788 4922
rect 16492 4868 16548 4870
rect 16572 4868 16628 4870
rect 16652 4868 16708 4870
rect 16732 4868 16788 4870
rect 18711 6554 18767 6556
rect 18791 6554 18847 6556
rect 18871 6554 18927 6556
rect 18951 6554 19007 6556
rect 18711 6502 18757 6554
rect 18757 6502 18767 6554
rect 18791 6502 18821 6554
rect 18821 6502 18833 6554
rect 18833 6502 18847 6554
rect 18871 6502 18885 6554
rect 18885 6502 18897 6554
rect 18897 6502 18927 6554
rect 18951 6502 18961 6554
rect 18961 6502 19007 6554
rect 18711 6500 18767 6502
rect 18791 6500 18847 6502
rect 18871 6500 18927 6502
rect 18951 6500 19007 6502
rect 18711 5466 18767 5468
rect 18791 5466 18847 5468
rect 18871 5466 18927 5468
rect 18951 5466 19007 5468
rect 18711 5414 18757 5466
rect 18757 5414 18767 5466
rect 18791 5414 18821 5466
rect 18821 5414 18833 5466
rect 18833 5414 18847 5466
rect 18871 5414 18885 5466
rect 18885 5414 18897 5466
rect 18897 5414 18927 5466
rect 18951 5414 18961 5466
rect 18961 5414 19007 5466
rect 18711 5412 18767 5414
rect 18791 5412 18847 5414
rect 18871 5412 18927 5414
rect 18951 5412 19007 5414
rect 14272 4378 14328 4380
rect 14352 4378 14408 4380
rect 14432 4378 14488 4380
rect 14512 4378 14568 4380
rect 14272 4326 14318 4378
rect 14318 4326 14328 4378
rect 14352 4326 14382 4378
rect 14382 4326 14394 4378
rect 14394 4326 14408 4378
rect 14432 4326 14446 4378
rect 14446 4326 14458 4378
rect 14458 4326 14488 4378
rect 14512 4326 14522 4378
rect 14522 4326 14568 4378
rect 14272 4324 14328 4326
rect 14352 4324 14408 4326
rect 14432 4324 14488 4326
rect 14512 4324 14568 4326
rect 14272 3290 14328 3292
rect 14352 3290 14408 3292
rect 14432 3290 14488 3292
rect 14512 3290 14568 3292
rect 14272 3238 14318 3290
rect 14318 3238 14328 3290
rect 14352 3238 14382 3290
rect 14382 3238 14394 3290
rect 14394 3238 14408 3290
rect 14432 3238 14446 3290
rect 14446 3238 14458 3290
rect 14458 3238 14488 3290
rect 14512 3238 14522 3290
rect 14522 3238 14568 3290
rect 14272 3236 14328 3238
rect 14352 3236 14408 3238
rect 14432 3236 14488 3238
rect 14512 3236 14568 3238
rect 16492 3834 16548 3836
rect 16572 3834 16628 3836
rect 16652 3834 16708 3836
rect 16732 3834 16788 3836
rect 16492 3782 16538 3834
rect 16538 3782 16548 3834
rect 16572 3782 16602 3834
rect 16602 3782 16614 3834
rect 16614 3782 16628 3834
rect 16652 3782 16666 3834
rect 16666 3782 16678 3834
rect 16678 3782 16708 3834
rect 16732 3782 16742 3834
rect 16742 3782 16788 3834
rect 16492 3780 16548 3782
rect 16572 3780 16628 3782
rect 16652 3780 16708 3782
rect 16732 3780 16788 3782
rect 18711 4378 18767 4380
rect 18791 4378 18847 4380
rect 18871 4378 18927 4380
rect 18951 4378 19007 4380
rect 18711 4326 18757 4378
rect 18757 4326 18767 4378
rect 18791 4326 18821 4378
rect 18821 4326 18833 4378
rect 18833 4326 18847 4378
rect 18871 4326 18885 4378
rect 18885 4326 18897 4378
rect 18897 4326 18927 4378
rect 18951 4326 18961 4378
rect 18961 4326 19007 4378
rect 18711 4324 18767 4326
rect 18791 4324 18847 4326
rect 18871 4324 18927 4326
rect 18951 4324 19007 4326
rect 18711 3290 18767 3292
rect 18791 3290 18847 3292
rect 18871 3290 18927 3292
rect 18951 3290 19007 3292
rect 18711 3238 18757 3290
rect 18757 3238 18767 3290
rect 18791 3238 18821 3290
rect 18821 3238 18833 3290
rect 18833 3238 18847 3290
rect 18871 3238 18885 3290
rect 18885 3238 18897 3290
rect 18897 3238 18927 3290
rect 18951 3238 18961 3290
rect 18961 3238 19007 3290
rect 18711 3236 18767 3238
rect 18791 3236 18847 3238
rect 18871 3236 18927 3238
rect 18951 3236 19007 3238
rect 16492 2746 16548 2748
rect 16572 2746 16628 2748
rect 16652 2746 16708 2748
rect 16732 2746 16788 2748
rect 16492 2694 16538 2746
rect 16538 2694 16548 2746
rect 16572 2694 16602 2746
rect 16602 2694 16614 2746
rect 16614 2694 16628 2746
rect 16652 2694 16666 2746
rect 16666 2694 16678 2746
rect 16678 2694 16708 2746
rect 16732 2694 16742 2746
rect 16742 2694 16788 2746
rect 16492 2692 16548 2694
rect 16572 2692 16628 2694
rect 16652 2692 16708 2694
rect 16732 2692 16788 2694
rect 14272 2202 14328 2204
rect 14352 2202 14408 2204
rect 14432 2202 14488 2204
rect 14512 2202 14568 2204
rect 14272 2150 14318 2202
rect 14318 2150 14328 2202
rect 14352 2150 14382 2202
rect 14382 2150 14394 2202
rect 14394 2150 14408 2202
rect 14432 2150 14446 2202
rect 14446 2150 14458 2202
rect 14458 2150 14488 2202
rect 14512 2150 14522 2202
rect 14522 2150 14568 2202
rect 14272 2148 14328 2150
rect 14352 2148 14408 2150
rect 14432 2148 14488 2150
rect 14512 2148 14568 2150
rect 18711 2202 18767 2204
rect 18791 2202 18847 2204
rect 18871 2202 18927 2204
rect 18951 2202 19007 2204
rect 18711 2150 18757 2202
rect 18757 2150 18767 2202
rect 18791 2150 18821 2202
rect 18821 2150 18833 2202
rect 18833 2150 18847 2202
rect 18871 2150 18885 2202
rect 18885 2150 18897 2202
rect 18897 2150 18927 2202
rect 18951 2150 18961 2202
rect 18961 2150 19007 2202
rect 18711 2148 18767 2150
rect 18791 2148 18847 2150
rect 18871 2148 18927 2150
rect 18951 2148 19007 2150
<< metal3 >>
rect 5384 7648 5700 7649
rect 5384 7584 5390 7648
rect 5454 7584 5470 7648
rect 5534 7584 5550 7648
rect 5614 7584 5630 7648
rect 5694 7584 5700 7648
rect 5384 7583 5700 7584
rect 9823 7648 10139 7649
rect 9823 7584 9829 7648
rect 9893 7584 9909 7648
rect 9973 7584 9989 7648
rect 10053 7584 10069 7648
rect 10133 7584 10139 7648
rect 9823 7583 10139 7584
rect 14262 7648 14578 7649
rect 14262 7584 14268 7648
rect 14332 7584 14348 7648
rect 14412 7584 14428 7648
rect 14492 7584 14508 7648
rect 14572 7584 14578 7648
rect 14262 7583 14578 7584
rect 18701 7648 19017 7649
rect 18701 7584 18707 7648
rect 18771 7584 18787 7648
rect 18851 7584 18867 7648
rect 18931 7584 18947 7648
rect 19011 7584 19017 7648
rect 18701 7583 19017 7584
rect 3165 7104 3481 7105
rect 3165 7040 3171 7104
rect 3235 7040 3251 7104
rect 3315 7040 3331 7104
rect 3395 7040 3411 7104
rect 3475 7040 3481 7104
rect 3165 7039 3481 7040
rect 7604 7104 7920 7105
rect 7604 7040 7610 7104
rect 7674 7040 7690 7104
rect 7754 7040 7770 7104
rect 7834 7040 7850 7104
rect 7914 7040 7920 7104
rect 7604 7039 7920 7040
rect 12043 7104 12359 7105
rect 12043 7040 12049 7104
rect 12113 7040 12129 7104
rect 12193 7040 12209 7104
rect 12273 7040 12289 7104
rect 12353 7040 12359 7104
rect 12043 7039 12359 7040
rect 16482 7104 16798 7105
rect 16482 7040 16488 7104
rect 16552 7040 16568 7104
rect 16632 7040 16648 7104
rect 16712 7040 16728 7104
rect 16792 7040 16798 7104
rect 16482 7039 16798 7040
rect 5384 6560 5700 6561
rect 5384 6496 5390 6560
rect 5454 6496 5470 6560
rect 5534 6496 5550 6560
rect 5614 6496 5630 6560
rect 5694 6496 5700 6560
rect 5384 6495 5700 6496
rect 9823 6560 10139 6561
rect 9823 6496 9829 6560
rect 9893 6496 9909 6560
rect 9973 6496 9989 6560
rect 10053 6496 10069 6560
rect 10133 6496 10139 6560
rect 9823 6495 10139 6496
rect 14262 6560 14578 6561
rect 14262 6496 14268 6560
rect 14332 6496 14348 6560
rect 14412 6496 14428 6560
rect 14492 6496 14508 6560
rect 14572 6496 14578 6560
rect 14262 6495 14578 6496
rect 18701 6560 19017 6561
rect 18701 6496 18707 6560
rect 18771 6496 18787 6560
rect 18851 6496 18867 6560
rect 18931 6496 18947 6560
rect 19011 6496 19017 6560
rect 18701 6495 19017 6496
rect 3165 6016 3481 6017
rect 3165 5952 3171 6016
rect 3235 5952 3251 6016
rect 3315 5952 3331 6016
rect 3395 5952 3411 6016
rect 3475 5952 3481 6016
rect 3165 5951 3481 5952
rect 7604 6016 7920 6017
rect 7604 5952 7610 6016
rect 7674 5952 7690 6016
rect 7754 5952 7770 6016
rect 7834 5952 7850 6016
rect 7914 5952 7920 6016
rect 7604 5951 7920 5952
rect 12043 6016 12359 6017
rect 12043 5952 12049 6016
rect 12113 5952 12129 6016
rect 12193 5952 12209 6016
rect 12273 5952 12289 6016
rect 12353 5952 12359 6016
rect 12043 5951 12359 5952
rect 16482 6016 16798 6017
rect 16482 5952 16488 6016
rect 16552 5952 16568 6016
rect 16632 5952 16648 6016
rect 16712 5952 16728 6016
rect 16792 5952 16798 6016
rect 16482 5951 16798 5952
rect 5384 5472 5700 5473
rect 5384 5408 5390 5472
rect 5454 5408 5470 5472
rect 5534 5408 5550 5472
rect 5614 5408 5630 5472
rect 5694 5408 5700 5472
rect 5384 5407 5700 5408
rect 9823 5472 10139 5473
rect 9823 5408 9829 5472
rect 9893 5408 9909 5472
rect 9973 5408 9989 5472
rect 10053 5408 10069 5472
rect 10133 5408 10139 5472
rect 9823 5407 10139 5408
rect 14262 5472 14578 5473
rect 14262 5408 14268 5472
rect 14332 5408 14348 5472
rect 14412 5408 14428 5472
rect 14492 5408 14508 5472
rect 14572 5408 14578 5472
rect 14262 5407 14578 5408
rect 18701 5472 19017 5473
rect 18701 5408 18707 5472
rect 18771 5408 18787 5472
rect 18851 5408 18867 5472
rect 18931 5408 18947 5472
rect 19011 5408 19017 5472
rect 18701 5407 19017 5408
rect 3165 4928 3481 4929
rect 3165 4864 3171 4928
rect 3235 4864 3251 4928
rect 3315 4864 3331 4928
rect 3395 4864 3411 4928
rect 3475 4864 3481 4928
rect 3165 4863 3481 4864
rect 7604 4928 7920 4929
rect 7604 4864 7610 4928
rect 7674 4864 7690 4928
rect 7754 4864 7770 4928
rect 7834 4864 7850 4928
rect 7914 4864 7920 4928
rect 7604 4863 7920 4864
rect 12043 4928 12359 4929
rect 12043 4864 12049 4928
rect 12113 4864 12129 4928
rect 12193 4864 12209 4928
rect 12273 4864 12289 4928
rect 12353 4864 12359 4928
rect 12043 4863 12359 4864
rect 16482 4928 16798 4929
rect 16482 4864 16488 4928
rect 16552 4864 16568 4928
rect 16632 4864 16648 4928
rect 16712 4864 16728 4928
rect 16792 4864 16798 4928
rect 16482 4863 16798 4864
rect 5384 4384 5700 4385
rect 5384 4320 5390 4384
rect 5454 4320 5470 4384
rect 5534 4320 5550 4384
rect 5614 4320 5630 4384
rect 5694 4320 5700 4384
rect 5384 4319 5700 4320
rect 9823 4384 10139 4385
rect 9823 4320 9829 4384
rect 9893 4320 9909 4384
rect 9973 4320 9989 4384
rect 10053 4320 10069 4384
rect 10133 4320 10139 4384
rect 9823 4319 10139 4320
rect 14262 4384 14578 4385
rect 14262 4320 14268 4384
rect 14332 4320 14348 4384
rect 14412 4320 14428 4384
rect 14492 4320 14508 4384
rect 14572 4320 14578 4384
rect 14262 4319 14578 4320
rect 18701 4384 19017 4385
rect 18701 4320 18707 4384
rect 18771 4320 18787 4384
rect 18851 4320 18867 4384
rect 18931 4320 18947 4384
rect 19011 4320 19017 4384
rect 18701 4319 19017 4320
rect 11881 4042 11947 4045
rect 13077 4042 13143 4045
rect 11881 4040 13143 4042
rect 11881 3984 11886 4040
rect 11942 3984 13082 4040
rect 13138 3984 13143 4040
rect 11881 3982 13143 3984
rect 11881 3979 11947 3982
rect 13077 3979 13143 3982
rect 3165 3840 3481 3841
rect 3165 3776 3171 3840
rect 3235 3776 3251 3840
rect 3315 3776 3331 3840
rect 3395 3776 3411 3840
rect 3475 3776 3481 3840
rect 3165 3775 3481 3776
rect 7604 3840 7920 3841
rect 7604 3776 7610 3840
rect 7674 3776 7690 3840
rect 7754 3776 7770 3840
rect 7834 3776 7850 3840
rect 7914 3776 7920 3840
rect 7604 3775 7920 3776
rect 12043 3840 12359 3841
rect 12043 3776 12049 3840
rect 12113 3776 12129 3840
rect 12193 3776 12209 3840
rect 12273 3776 12289 3840
rect 12353 3776 12359 3840
rect 12043 3775 12359 3776
rect 16482 3840 16798 3841
rect 16482 3776 16488 3840
rect 16552 3776 16568 3840
rect 16632 3776 16648 3840
rect 16712 3776 16728 3840
rect 16792 3776 16798 3840
rect 16482 3775 16798 3776
rect 7373 3362 7439 3365
rect 8293 3362 8359 3365
rect 7373 3360 8359 3362
rect 7373 3304 7378 3360
rect 7434 3304 8298 3360
rect 8354 3304 8359 3360
rect 7373 3302 8359 3304
rect 7373 3299 7439 3302
rect 8293 3299 8359 3302
rect 5384 3296 5700 3297
rect 5384 3232 5390 3296
rect 5454 3232 5470 3296
rect 5534 3232 5550 3296
rect 5614 3232 5630 3296
rect 5694 3232 5700 3296
rect 5384 3231 5700 3232
rect 9823 3296 10139 3297
rect 9823 3232 9829 3296
rect 9893 3232 9909 3296
rect 9973 3232 9989 3296
rect 10053 3232 10069 3296
rect 10133 3232 10139 3296
rect 9823 3231 10139 3232
rect 14262 3296 14578 3297
rect 14262 3232 14268 3296
rect 14332 3232 14348 3296
rect 14412 3232 14428 3296
rect 14492 3232 14508 3296
rect 14572 3232 14578 3296
rect 14262 3231 14578 3232
rect 18701 3296 19017 3297
rect 18701 3232 18707 3296
rect 18771 3232 18787 3296
rect 18851 3232 18867 3296
rect 18931 3232 18947 3296
rect 19011 3232 19017 3296
rect 18701 3231 19017 3232
rect 7097 3090 7163 3093
rect 9029 3090 9095 3093
rect 7097 3088 9095 3090
rect 7097 3032 7102 3088
rect 7158 3032 9034 3088
rect 9090 3032 9095 3088
rect 7097 3030 9095 3032
rect 7097 3027 7163 3030
rect 9029 3027 9095 3030
rect 3165 2752 3481 2753
rect 3165 2688 3171 2752
rect 3235 2688 3251 2752
rect 3315 2688 3331 2752
rect 3395 2688 3411 2752
rect 3475 2688 3481 2752
rect 3165 2687 3481 2688
rect 7604 2752 7920 2753
rect 7604 2688 7610 2752
rect 7674 2688 7690 2752
rect 7754 2688 7770 2752
rect 7834 2688 7850 2752
rect 7914 2688 7920 2752
rect 7604 2687 7920 2688
rect 12043 2752 12359 2753
rect 12043 2688 12049 2752
rect 12113 2688 12129 2752
rect 12193 2688 12209 2752
rect 12273 2688 12289 2752
rect 12353 2688 12359 2752
rect 12043 2687 12359 2688
rect 16482 2752 16798 2753
rect 16482 2688 16488 2752
rect 16552 2688 16568 2752
rect 16632 2688 16648 2752
rect 16712 2688 16728 2752
rect 16792 2688 16798 2752
rect 16482 2687 16798 2688
rect 5384 2208 5700 2209
rect 5384 2144 5390 2208
rect 5454 2144 5470 2208
rect 5534 2144 5550 2208
rect 5614 2144 5630 2208
rect 5694 2144 5700 2208
rect 5384 2143 5700 2144
rect 9823 2208 10139 2209
rect 9823 2144 9829 2208
rect 9893 2144 9909 2208
rect 9973 2144 9989 2208
rect 10053 2144 10069 2208
rect 10133 2144 10139 2208
rect 9823 2143 10139 2144
rect 14262 2208 14578 2209
rect 14262 2144 14268 2208
rect 14332 2144 14348 2208
rect 14412 2144 14428 2208
rect 14492 2144 14508 2208
rect 14572 2144 14578 2208
rect 14262 2143 14578 2144
rect 18701 2208 19017 2209
rect 18701 2144 18707 2208
rect 18771 2144 18787 2208
rect 18851 2144 18867 2208
rect 18931 2144 18947 2208
rect 19011 2144 19017 2208
rect 18701 2143 19017 2144
<< via3 >>
rect 5390 7644 5454 7648
rect 5390 7588 5394 7644
rect 5394 7588 5450 7644
rect 5450 7588 5454 7644
rect 5390 7584 5454 7588
rect 5470 7644 5534 7648
rect 5470 7588 5474 7644
rect 5474 7588 5530 7644
rect 5530 7588 5534 7644
rect 5470 7584 5534 7588
rect 5550 7644 5614 7648
rect 5550 7588 5554 7644
rect 5554 7588 5610 7644
rect 5610 7588 5614 7644
rect 5550 7584 5614 7588
rect 5630 7644 5694 7648
rect 5630 7588 5634 7644
rect 5634 7588 5690 7644
rect 5690 7588 5694 7644
rect 5630 7584 5694 7588
rect 9829 7644 9893 7648
rect 9829 7588 9833 7644
rect 9833 7588 9889 7644
rect 9889 7588 9893 7644
rect 9829 7584 9893 7588
rect 9909 7644 9973 7648
rect 9909 7588 9913 7644
rect 9913 7588 9969 7644
rect 9969 7588 9973 7644
rect 9909 7584 9973 7588
rect 9989 7644 10053 7648
rect 9989 7588 9993 7644
rect 9993 7588 10049 7644
rect 10049 7588 10053 7644
rect 9989 7584 10053 7588
rect 10069 7644 10133 7648
rect 10069 7588 10073 7644
rect 10073 7588 10129 7644
rect 10129 7588 10133 7644
rect 10069 7584 10133 7588
rect 14268 7644 14332 7648
rect 14268 7588 14272 7644
rect 14272 7588 14328 7644
rect 14328 7588 14332 7644
rect 14268 7584 14332 7588
rect 14348 7644 14412 7648
rect 14348 7588 14352 7644
rect 14352 7588 14408 7644
rect 14408 7588 14412 7644
rect 14348 7584 14412 7588
rect 14428 7644 14492 7648
rect 14428 7588 14432 7644
rect 14432 7588 14488 7644
rect 14488 7588 14492 7644
rect 14428 7584 14492 7588
rect 14508 7644 14572 7648
rect 14508 7588 14512 7644
rect 14512 7588 14568 7644
rect 14568 7588 14572 7644
rect 14508 7584 14572 7588
rect 18707 7644 18771 7648
rect 18707 7588 18711 7644
rect 18711 7588 18767 7644
rect 18767 7588 18771 7644
rect 18707 7584 18771 7588
rect 18787 7644 18851 7648
rect 18787 7588 18791 7644
rect 18791 7588 18847 7644
rect 18847 7588 18851 7644
rect 18787 7584 18851 7588
rect 18867 7644 18931 7648
rect 18867 7588 18871 7644
rect 18871 7588 18927 7644
rect 18927 7588 18931 7644
rect 18867 7584 18931 7588
rect 18947 7644 19011 7648
rect 18947 7588 18951 7644
rect 18951 7588 19007 7644
rect 19007 7588 19011 7644
rect 18947 7584 19011 7588
rect 3171 7100 3235 7104
rect 3171 7044 3175 7100
rect 3175 7044 3231 7100
rect 3231 7044 3235 7100
rect 3171 7040 3235 7044
rect 3251 7100 3315 7104
rect 3251 7044 3255 7100
rect 3255 7044 3311 7100
rect 3311 7044 3315 7100
rect 3251 7040 3315 7044
rect 3331 7100 3395 7104
rect 3331 7044 3335 7100
rect 3335 7044 3391 7100
rect 3391 7044 3395 7100
rect 3331 7040 3395 7044
rect 3411 7100 3475 7104
rect 3411 7044 3415 7100
rect 3415 7044 3471 7100
rect 3471 7044 3475 7100
rect 3411 7040 3475 7044
rect 7610 7100 7674 7104
rect 7610 7044 7614 7100
rect 7614 7044 7670 7100
rect 7670 7044 7674 7100
rect 7610 7040 7674 7044
rect 7690 7100 7754 7104
rect 7690 7044 7694 7100
rect 7694 7044 7750 7100
rect 7750 7044 7754 7100
rect 7690 7040 7754 7044
rect 7770 7100 7834 7104
rect 7770 7044 7774 7100
rect 7774 7044 7830 7100
rect 7830 7044 7834 7100
rect 7770 7040 7834 7044
rect 7850 7100 7914 7104
rect 7850 7044 7854 7100
rect 7854 7044 7910 7100
rect 7910 7044 7914 7100
rect 7850 7040 7914 7044
rect 12049 7100 12113 7104
rect 12049 7044 12053 7100
rect 12053 7044 12109 7100
rect 12109 7044 12113 7100
rect 12049 7040 12113 7044
rect 12129 7100 12193 7104
rect 12129 7044 12133 7100
rect 12133 7044 12189 7100
rect 12189 7044 12193 7100
rect 12129 7040 12193 7044
rect 12209 7100 12273 7104
rect 12209 7044 12213 7100
rect 12213 7044 12269 7100
rect 12269 7044 12273 7100
rect 12209 7040 12273 7044
rect 12289 7100 12353 7104
rect 12289 7044 12293 7100
rect 12293 7044 12349 7100
rect 12349 7044 12353 7100
rect 12289 7040 12353 7044
rect 16488 7100 16552 7104
rect 16488 7044 16492 7100
rect 16492 7044 16548 7100
rect 16548 7044 16552 7100
rect 16488 7040 16552 7044
rect 16568 7100 16632 7104
rect 16568 7044 16572 7100
rect 16572 7044 16628 7100
rect 16628 7044 16632 7100
rect 16568 7040 16632 7044
rect 16648 7100 16712 7104
rect 16648 7044 16652 7100
rect 16652 7044 16708 7100
rect 16708 7044 16712 7100
rect 16648 7040 16712 7044
rect 16728 7100 16792 7104
rect 16728 7044 16732 7100
rect 16732 7044 16788 7100
rect 16788 7044 16792 7100
rect 16728 7040 16792 7044
rect 5390 6556 5454 6560
rect 5390 6500 5394 6556
rect 5394 6500 5450 6556
rect 5450 6500 5454 6556
rect 5390 6496 5454 6500
rect 5470 6556 5534 6560
rect 5470 6500 5474 6556
rect 5474 6500 5530 6556
rect 5530 6500 5534 6556
rect 5470 6496 5534 6500
rect 5550 6556 5614 6560
rect 5550 6500 5554 6556
rect 5554 6500 5610 6556
rect 5610 6500 5614 6556
rect 5550 6496 5614 6500
rect 5630 6556 5694 6560
rect 5630 6500 5634 6556
rect 5634 6500 5690 6556
rect 5690 6500 5694 6556
rect 5630 6496 5694 6500
rect 9829 6556 9893 6560
rect 9829 6500 9833 6556
rect 9833 6500 9889 6556
rect 9889 6500 9893 6556
rect 9829 6496 9893 6500
rect 9909 6556 9973 6560
rect 9909 6500 9913 6556
rect 9913 6500 9969 6556
rect 9969 6500 9973 6556
rect 9909 6496 9973 6500
rect 9989 6556 10053 6560
rect 9989 6500 9993 6556
rect 9993 6500 10049 6556
rect 10049 6500 10053 6556
rect 9989 6496 10053 6500
rect 10069 6556 10133 6560
rect 10069 6500 10073 6556
rect 10073 6500 10129 6556
rect 10129 6500 10133 6556
rect 10069 6496 10133 6500
rect 14268 6556 14332 6560
rect 14268 6500 14272 6556
rect 14272 6500 14328 6556
rect 14328 6500 14332 6556
rect 14268 6496 14332 6500
rect 14348 6556 14412 6560
rect 14348 6500 14352 6556
rect 14352 6500 14408 6556
rect 14408 6500 14412 6556
rect 14348 6496 14412 6500
rect 14428 6556 14492 6560
rect 14428 6500 14432 6556
rect 14432 6500 14488 6556
rect 14488 6500 14492 6556
rect 14428 6496 14492 6500
rect 14508 6556 14572 6560
rect 14508 6500 14512 6556
rect 14512 6500 14568 6556
rect 14568 6500 14572 6556
rect 14508 6496 14572 6500
rect 18707 6556 18771 6560
rect 18707 6500 18711 6556
rect 18711 6500 18767 6556
rect 18767 6500 18771 6556
rect 18707 6496 18771 6500
rect 18787 6556 18851 6560
rect 18787 6500 18791 6556
rect 18791 6500 18847 6556
rect 18847 6500 18851 6556
rect 18787 6496 18851 6500
rect 18867 6556 18931 6560
rect 18867 6500 18871 6556
rect 18871 6500 18927 6556
rect 18927 6500 18931 6556
rect 18867 6496 18931 6500
rect 18947 6556 19011 6560
rect 18947 6500 18951 6556
rect 18951 6500 19007 6556
rect 19007 6500 19011 6556
rect 18947 6496 19011 6500
rect 3171 6012 3235 6016
rect 3171 5956 3175 6012
rect 3175 5956 3231 6012
rect 3231 5956 3235 6012
rect 3171 5952 3235 5956
rect 3251 6012 3315 6016
rect 3251 5956 3255 6012
rect 3255 5956 3311 6012
rect 3311 5956 3315 6012
rect 3251 5952 3315 5956
rect 3331 6012 3395 6016
rect 3331 5956 3335 6012
rect 3335 5956 3391 6012
rect 3391 5956 3395 6012
rect 3331 5952 3395 5956
rect 3411 6012 3475 6016
rect 3411 5956 3415 6012
rect 3415 5956 3471 6012
rect 3471 5956 3475 6012
rect 3411 5952 3475 5956
rect 7610 6012 7674 6016
rect 7610 5956 7614 6012
rect 7614 5956 7670 6012
rect 7670 5956 7674 6012
rect 7610 5952 7674 5956
rect 7690 6012 7754 6016
rect 7690 5956 7694 6012
rect 7694 5956 7750 6012
rect 7750 5956 7754 6012
rect 7690 5952 7754 5956
rect 7770 6012 7834 6016
rect 7770 5956 7774 6012
rect 7774 5956 7830 6012
rect 7830 5956 7834 6012
rect 7770 5952 7834 5956
rect 7850 6012 7914 6016
rect 7850 5956 7854 6012
rect 7854 5956 7910 6012
rect 7910 5956 7914 6012
rect 7850 5952 7914 5956
rect 12049 6012 12113 6016
rect 12049 5956 12053 6012
rect 12053 5956 12109 6012
rect 12109 5956 12113 6012
rect 12049 5952 12113 5956
rect 12129 6012 12193 6016
rect 12129 5956 12133 6012
rect 12133 5956 12189 6012
rect 12189 5956 12193 6012
rect 12129 5952 12193 5956
rect 12209 6012 12273 6016
rect 12209 5956 12213 6012
rect 12213 5956 12269 6012
rect 12269 5956 12273 6012
rect 12209 5952 12273 5956
rect 12289 6012 12353 6016
rect 12289 5956 12293 6012
rect 12293 5956 12349 6012
rect 12349 5956 12353 6012
rect 12289 5952 12353 5956
rect 16488 6012 16552 6016
rect 16488 5956 16492 6012
rect 16492 5956 16548 6012
rect 16548 5956 16552 6012
rect 16488 5952 16552 5956
rect 16568 6012 16632 6016
rect 16568 5956 16572 6012
rect 16572 5956 16628 6012
rect 16628 5956 16632 6012
rect 16568 5952 16632 5956
rect 16648 6012 16712 6016
rect 16648 5956 16652 6012
rect 16652 5956 16708 6012
rect 16708 5956 16712 6012
rect 16648 5952 16712 5956
rect 16728 6012 16792 6016
rect 16728 5956 16732 6012
rect 16732 5956 16788 6012
rect 16788 5956 16792 6012
rect 16728 5952 16792 5956
rect 5390 5468 5454 5472
rect 5390 5412 5394 5468
rect 5394 5412 5450 5468
rect 5450 5412 5454 5468
rect 5390 5408 5454 5412
rect 5470 5468 5534 5472
rect 5470 5412 5474 5468
rect 5474 5412 5530 5468
rect 5530 5412 5534 5468
rect 5470 5408 5534 5412
rect 5550 5468 5614 5472
rect 5550 5412 5554 5468
rect 5554 5412 5610 5468
rect 5610 5412 5614 5468
rect 5550 5408 5614 5412
rect 5630 5468 5694 5472
rect 5630 5412 5634 5468
rect 5634 5412 5690 5468
rect 5690 5412 5694 5468
rect 5630 5408 5694 5412
rect 9829 5468 9893 5472
rect 9829 5412 9833 5468
rect 9833 5412 9889 5468
rect 9889 5412 9893 5468
rect 9829 5408 9893 5412
rect 9909 5468 9973 5472
rect 9909 5412 9913 5468
rect 9913 5412 9969 5468
rect 9969 5412 9973 5468
rect 9909 5408 9973 5412
rect 9989 5468 10053 5472
rect 9989 5412 9993 5468
rect 9993 5412 10049 5468
rect 10049 5412 10053 5468
rect 9989 5408 10053 5412
rect 10069 5468 10133 5472
rect 10069 5412 10073 5468
rect 10073 5412 10129 5468
rect 10129 5412 10133 5468
rect 10069 5408 10133 5412
rect 14268 5468 14332 5472
rect 14268 5412 14272 5468
rect 14272 5412 14328 5468
rect 14328 5412 14332 5468
rect 14268 5408 14332 5412
rect 14348 5468 14412 5472
rect 14348 5412 14352 5468
rect 14352 5412 14408 5468
rect 14408 5412 14412 5468
rect 14348 5408 14412 5412
rect 14428 5468 14492 5472
rect 14428 5412 14432 5468
rect 14432 5412 14488 5468
rect 14488 5412 14492 5468
rect 14428 5408 14492 5412
rect 14508 5468 14572 5472
rect 14508 5412 14512 5468
rect 14512 5412 14568 5468
rect 14568 5412 14572 5468
rect 14508 5408 14572 5412
rect 18707 5468 18771 5472
rect 18707 5412 18711 5468
rect 18711 5412 18767 5468
rect 18767 5412 18771 5468
rect 18707 5408 18771 5412
rect 18787 5468 18851 5472
rect 18787 5412 18791 5468
rect 18791 5412 18847 5468
rect 18847 5412 18851 5468
rect 18787 5408 18851 5412
rect 18867 5468 18931 5472
rect 18867 5412 18871 5468
rect 18871 5412 18927 5468
rect 18927 5412 18931 5468
rect 18867 5408 18931 5412
rect 18947 5468 19011 5472
rect 18947 5412 18951 5468
rect 18951 5412 19007 5468
rect 19007 5412 19011 5468
rect 18947 5408 19011 5412
rect 3171 4924 3235 4928
rect 3171 4868 3175 4924
rect 3175 4868 3231 4924
rect 3231 4868 3235 4924
rect 3171 4864 3235 4868
rect 3251 4924 3315 4928
rect 3251 4868 3255 4924
rect 3255 4868 3311 4924
rect 3311 4868 3315 4924
rect 3251 4864 3315 4868
rect 3331 4924 3395 4928
rect 3331 4868 3335 4924
rect 3335 4868 3391 4924
rect 3391 4868 3395 4924
rect 3331 4864 3395 4868
rect 3411 4924 3475 4928
rect 3411 4868 3415 4924
rect 3415 4868 3471 4924
rect 3471 4868 3475 4924
rect 3411 4864 3475 4868
rect 7610 4924 7674 4928
rect 7610 4868 7614 4924
rect 7614 4868 7670 4924
rect 7670 4868 7674 4924
rect 7610 4864 7674 4868
rect 7690 4924 7754 4928
rect 7690 4868 7694 4924
rect 7694 4868 7750 4924
rect 7750 4868 7754 4924
rect 7690 4864 7754 4868
rect 7770 4924 7834 4928
rect 7770 4868 7774 4924
rect 7774 4868 7830 4924
rect 7830 4868 7834 4924
rect 7770 4864 7834 4868
rect 7850 4924 7914 4928
rect 7850 4868 7854 4924
rect 7854 4868 7910 4924
rect 7910 4868 7914 4924
rect 7850 4864 7914 4868
rect 12049 4924 12113 4928
rect 12049 4868 12053 4924
rect 12053 4868 12109 4924
rect 12109 4868 12113 4924
rect 12049 4864 12113 4868
rect 12129 4924 12193 4928
rect 12129 4868 12133 4924
rect 12133 4868 12189 4924
rect 12189 4868 12193 4924
rect 12129 4864 12193 4868
rect 12209 4924 12273 4928
rect 12209 4868 12213 4924
rect 12213 4868 12269 4924
rect 12269 4868 12273 4924
rect 12209 4864 12273 4868
rect 12289 4924 12353 4928
rect 12289 4868 12293 4924
rect 12293 4868 12349 4924
rect 12349 4868 12353 4924
rect 12289 4864 12353 4868
rect 16488 4924 16552 4928
rect 16488 4868 16492 4924
rect 16492 4868 16548 4924
rect 16548 4868 16552 4924
rect 16488 4864 16552 4868
rect 16568 4924 16632 4928
rect 16568 4868 16572 4924
rect 16572 4868 16628 4924
rect 16628 4868 16632 4924
rect 16568 4864 16632 4868
rect 16648 4924 16712 4928
rect 16648 4868 16652 4924
rect 16652 4868 16708 4924
rect 16708 4868 16712 4924
rect 16648 4864 16712 4868
rect 16728 4924 16792 4928
rect 16728 4868 16732 4924
rect 16732 4868 16788 4924
rect 16788 4868 16792 4924
rect 16728 4864 16792 4868
rect 5390 4380 5454 4384
rect 5390 4324 5394 4380
rect 5394 4324 5450 4380
rect 5450 4324 5454 4380
rect 5390 4320 5454 4324
rect 5470 4380 5534 4384
rect 5470 4324 5474 4380
rect 5474 4324 5530 4380
rect 5530 4324 5534 4380
rect 5470 4320 5534 4324
rect 5550 4380 5614 4384
rect 5550 4324 5554 4380
rect 5554 4324 5610 4380
rect 5610 4324 5614 4380
rect 5550 4320 5614 4324
rect 5630 4380 5694 4384
rect 5630 4324 5634 4380
rect 5634 4324 5690 4380
rect 5690 4324 5694 4380
rect 5630 4320 5694 4324
rect 9829 4380 9893 4384
rect 9829 4324 9833 4380
rect 9833 4324 9889 4380
rect 9889 4324 9893 4380
rect 9829 4320 9893 4324
rect 9909 4380 9973 4384
rect 9909 4324 9913 4380
rect 9913 4324 9969 4380
rect 9969 4324 9973 4380
rect 9909 4320 9973 4324
rect 9989 4380 10053 4384
rect 9989 4324 9993 4380
rect 9993 4324 10049 4380
rect 10049 4324 10053 4380
rect 9989 4320 10053 4324
rect 10069 4380 10133 4384
rect 10069 4324 10073 4380
rect 10073 4324 10129 4380
rect 10129 4324 10133 4380
rect 10069 4320 10133 4324
rect 14268 4380 14332 4384
rect 14268 4324 14272 4380
rect 14272 4324 14328 4380
rect 14328 4324 14332 4380
rect 14268 4320 14332 4324
rect 14348 4380 14412 4384
rect 14348 4324 14352 4380
rect 14352 4324 14408 4380
rect 14408 4324 14412 4380
rect 14348 4320 14412 4324
rect 14428 4380 14492 4384
rect 14428 4324 14432 4380
rect 14432 4324 14488 4380
rect 14488 4324 14492 4380
rect 14428 4320 14492 4324
rect 14508 4380 14572 4384
rect 14508 4324 14512 4380
rect 14512 4324 14568 4380
rect 14568 4324 14572 4380
rect 14508 4320 14572 4324
rect 18707 4380 18771 4384
rect 18707 4324 18711 4380
rect 18711 4324 18767 4380
rect 18767 4324 18771 4380
rect 18707 4320 18771 4324
rect 18787 4380 18851 4384
rect 18787 4324 18791 4380
rect 18791 4324 18847 4380
rect 18847 4324 18851 4380
rect 18787 4320 18851 4324
rect 18867 4380 18931 4384
rect 18867 4324 18871 4380
rect 18871 4324 18927 4380
rect 18927 4324 18931 4380
rect 18867 4320 18931 4324
rect 18947 4380 19011 4384
rect 18947 4324 18951 4380
rect 18951 4324 19007 4380
rect 19007 4324 19011 4380
rect 18947 4320 19011 4324
rect 3171 3836 3235 3840
rect 3171 3780 3175 3836
rect 3175 3780 3231 3836
rect 3231 3780 3235 3836
rect 3171 3776 3235 3780
rect 3251 3836 3315 3840
rect 3251 3780 3255 3836
rect 3255 3780 3311 3836
rect 3311 3780 3315 3836
rect 3251 3776 3315 3780
rect 3331 3836 3395 3840
rect 3331 3780 3335 3836
rect 3335 3780 3391 3836
rect 3391 3780 3395 3836
rect 3331 3776 3395 3780
rect 3411 3836 3475 3840
rect 3411 3780 3415 3836
rect 3415 3780 3471 3836
rect 3471 3780 3475 3836
rect 3411 3776 3475 3780
rect 7610 3836 7674 3840
rect 7610 3780 7614 3836
rect 7614 3780 7670 3836
rect 7670 3780 7674 3836
rect 7610 3776 7674 3780
rect 7690 3836 7754 3840
rect 7690 3780 7694 3836
rect 7694 3780 7750 3836
rect 7750 3780 7754 3836
rect 7690 3776 7754 3780
rect 7770 3836 7834 3840
rect 7770 3780 7774 3836
rect 7774 3780 7830 3836
rect 7830 3780 7834 3836
rect 7770 3776 7834 3780
rect 7850 3836 7914 3840
rect 7850 3780 7854 3836
rect 7854 3780 7910 3836
rect 7910 3780 7914 3836
rect 7850 3776 7914 3780
rect 12049 3836 12113 3840
rect 12049 3780 12053 3836
rect 12053 3780 12109 3836
rect 12109 3780 12113 3836
rect 12049 3776 12113 3780
rect 12129 3836 12193 3840
rect 12129 3780 12133 3836
rect 12133 3780 12189 3836
rect 12189 3780 12193 3836
rect 12129 3776 12193 3780
rect 12209 3836 12273 3840
rect 12209 3780 12213 3836
rect 12213 3780 12269 3836
rect 12269 3780 12273 3836
rect 12209 3776 12273 3780
rect 12289 3836 12353 3840
rect 12289 3780 12293 3836
rect 12293 3780 12349 3836
rect 12349 3780 12353 3836
rect 12289 3776 12353 3780
rect 16488 3836 16552 3840
rect 16488 3780 16492 3836
rect 16492 3780 16548 3836
rect 16548 3780 16552 3836
rect 16488 3776 16552 3780
rect 16568 3836 16632 3840
rect 16568 3780 16572 3836
rect 16572 3780 16628 3836
rect 16628 3780 16632 3836
rect 16568 3776 16632 3780
rect 16648 3836 16712 3840
rect 16648 3780 16652 3836
rect 16652 3780 16708 3836
rect 16708 3780 16712 3836
rect 16648 3776 16712 3780
rect 16728 3836 16792 3840
rect 16728 3780 16732 3836
rect 16732 3780 16788 3836
rect 16788 3780 16792 3836
rect 16728 3776 16792 3780
rect 5390 3292 5454 3296
rect 5390 3236 5394 3292
rect 5394 3236 5450 3292
rect 5450 3236 5454 3292
rect 5390 3232 5454 3236
rect 5470 3292 5534 3296
rect 5470 3236 5474 3292
rect 5474 3236 5530 3292
rect 5530 3236 5534 3292
rect 5470 3232 5534 3236
rect 5550 3292 5614 3296
rect 5550 3236 5554 3292
rect 5554 3236 5610 3292
rect 5610 3236 5614 3292
rect 5550 3232 5614 3236
rect 5630 3292 5694 3296
rect 5630 3236 5634 3292
rect 5634 3236 5690 3292
rect 5690 3236 5694 3292
rect 5630 3232 5694 3236
rect 9829 3292 9893 3296
rect 9829 3236 9833 3292
rect 9833 3236 9889 3292
rect 9889 3236 9893 3292
rect 9829 3232 9893 3236
rect 9909 3292 9973 3296
rect 9909 3236 9913 3292
rect 9913 3236 9969 3292
rect 9969 3236 9973 3292
rect 9909 3232 9973 3236
rect 9989 3292 10053 3296
rect 9989 3236 9993 3292
rect 9993 3236 10049 3292
rect 10049 3236 10053 3292
rect 9989 3232 10053 3236
rect 10069 3292 10133 3296
rect 10069 3236 10073 3292
rect 10073 3236 10129 3292
rect 10129 3236 10133 3292
rect 10069 3232 10133 3236
rect 14268 3292 14332 3296
rect 14268 3236 14272 3292
rect 14272 3236 14328 3292
rect 14328 3236 14332 3292
rect 14268 3232 14332 3236
rect 14348 3292 14412 3296
rect 14348 3236 14352 3292
rect 14352 3236 14408 3292
rect 14408 3236 14412 3292
rect 14348 3232 14412 3236
rect 14428 3292 14492 3296
rect 14428 3236 14432 3292
rect 14432 3236 14488 3292
rect 14488 3236 14492 3292
rect 14428 3232 14492 3236
rect 14508 3292 14572 3296
rect 14508 3236 14512 3292
rect 14512 3236 14568 3292
rect 14568 3236 14572 3292
rect 14508 3232 14572 3236
rect 18707 3292 18771 3296
rect 18707 3236 18711 3292
rect 18711 3236 18767 3292
rect 18767 3236 18771 3292
rect 18707 3232 18771 3236
rect 18787 3292 18851 3296
rect 18787 3236 18791 3292
rect 18791 3236 18847 3292
rect 18847 3236 18851 3292
rect 18787 3232 18851 3236
rect 18867 3292 18931 3296
rect 18867 3236 18871 3292
rect 18871 3236 18927 3292
rect 18927 3236 18931 3292
rect 18867 3232 18931 3236
rect 18947 3292 19011 3296
rect 18947 3236 18951 3292
rect 18951 3236 19007 3292
rect 19007 3236 19011 3292
rect 18947 3232 19011 3236
rect 3171 2748 3235 2752
rect 3171 2692 3175 2748
rect 3175 2692 3231 2748
rect 3231 2692 3235 2748
rect 3171 2688 3235 2692
rect 3251 2748 3315 2752
rect 3251 2692 3255 2748
rect 3255 2692 3311 2748
rect 3311 2692 3315 2748
rect 3251 2688 3315 2692
rect 3331 2748 3395 2752
rect 3331 2692 3335 2748
rect 3335 2692 3391 2748
rect 3391 2692 3395 2748
rect 3331 2688 3395 2692
rect 3411 2748 3475 2752
rect 3411 2692 3415 2748
rect 3415 2692 3471 2748
rect 3471 2692 3475 2748
rect 3411 2688 3475 2692
rect 7610 2748 7674 2752
rect 7610 2692 7614 2748
rect 7614 2692 7670 2748
rect 7670 2692 7674 2748
rect 7610 2688 7674 2692
rect 7690 2748 7754 2752
rect 7690 2692 7694 2748
rect 7694 2692 7750 2748
rect 7750 2692 7754 2748
rect 7690 2688 7754 2692
rect 7770 2748 7834 2752
rect 7770 2692 7774 2748
rect 7774 2692 7830 2748
rect 7830 2692 7834 2748
rect 7770 2688 7834 2692
rect 7850 2748 7914 2752
rect 7850 2692 7854 2748
rect 7854 2692 7910 2748
rect 7910 2692 7914 2748
rect 7850 2688 7914 2692
rect 12049 2748 12113 2752
rect 12049 2692 12053 2748
rect 12053 2692 12109 2748
rect 12109 2692 12113 2748
rect 12049 2688 12113 2692
rect 12129 2748 12193 2752
rect 12129 2692 12133 2748
rect 12133 2692 12189 2748
rect 12189 2692 12193 2748
rect 12129 2688 12193 2692
rect 12209 2748 12273 2752
rect 12209 2692 12213 2748
rect 12213 2692 12269 2748
rect 12269 2692 12273 2748
rect 12209 2688 12273 2692
rect 12289 2748 12353 2752
rect 12289 2692 12293 2748
rect 12293 2692 12349 2748
rect 12349 2692 12353 2748
rect 12289 2688 12353 2692
rect 16488 2748 16552 2752
rect 16488 2692 16492 2748
rect 16492 2692 16548 2748
rect 16548 2692 16552 2748
rect 16488 2688 16552 2692
rect 16568 2748 16632 2752
rect 16568 2692 16572 2748
rect 16572 2692 16628 2748
rect 16628 2692 16632 2748
rect 16568 2688 16632 2692
rect 16648 2748 16712 2752
rect 16648 2692 16652 2748
rect 16652 2692 16708 2748
rect 16708 2692 16712 2748
rect 16648 2688 16712 2692
rect 16728 2748 16792 2752
rect 16728 2692 16732 2748
rect 16732 2692 16788 2748
rect 16788 2692 16792 2748
rect 16728 2688 16792 2692
rect 5390 2204 5454 2208
rect 5390 2148 5394 2204
rect 5394 2148 5450 2204
rect 5450 2148 5454 2204
rect 5390 2144 5454 2148
rect 5470 2204 5534 2208
rect 5470 2148 5474 2204
rect 5474 2148 5530 2204
rect 5530 2148 5534 2204
rect 5470 2144 5534 2148
rect 5550 2204 5614 2208
rect 5550 2148 5554 2204
rect 5554 2148 5610 2204
rect 5610 2148 5614 2204
rect 5550 2144 5614 2148
rect 5630 2204 5694 2208
rect 5630 2148 5634 2204
rect 5634 2148 5690 2204
rect 5690 2148 5694 2204
rect 5630 2144 5694 2148
rect 9829 2204 9893 2208
rect 9829 2148 9833 2204
rect 9833 2148 9889 2204
rect 9889 2148 9893 2204
rect 9829 2144 9893 2148
rect 9909 2204 9973 2208
rect 9909 2148 9913 2204
rect 9913 2148 9969 2204
rect 9969 2148 9973 2204
rect 9909 2144 9973 2148
rect 9989 2204 10053 2208
rect 9989 2148 9993 2204
rect 9993 2148 10049 2204
rect 10049 2148 10053 2204
rect 9989 2144 10053 2148
rect 10069 2204 10133 2208
rect 10069 2148 10073 2204
rect 10073 2148 10129 2204
rect 10129 2148 10133 2204
rect 10069 2144 10133 2148
rect 14268 2204 14332 2208
rect 14268 2148 14272 2204
rect 14272 2148 14328 2204
rect 14328 2148 14332 2204
rect 14268 2144 14332 2148
rect 14348 2204 14412 2208
rect 14348 2148 14352 2204
rect 14352 2148 14408 2204
rect 14408 2148 14412 2204
rect 14348 2144 14412 2148
rect 14428 2204 14492 2208
rect 14428 2148 14432 2204
rect 14432 2148 14488 2204
rect 14488 2148 14492 2204
rect 14428 2144 14492 2148
rect 14508 2204 14572 2208
rect 14508 2148 14512 2204
rect 14512 2148 14568 2204
rect 14568 2148 14572 2204
rect 14508 2144 14572 2148
rect 18707 2204 18771 2208
rect 18707 2148 18711 2204
rect 18711 2148 18767 2204
rect 18767 2148 18771 2204
rect 18707 2144 18771 2148
rect 18787 2204 18851 2208
rect 18787 2148 18791 2204
rect 18791 2148 18847 2204
rect 18847 2148 18851 2204
rect 18787 2144 18851 2148
rect 18867 2204 18931 2208
rect 18867 2148 18871 2204
rect 18871 2148 18927 2204
rect 18927 2148 18931 2204
rect 18867 2144 18931 2148
rect 18947 2204 19011 2208
rect 18947 2148 18951 2204
rect 18951 2148 19007 2204
rect 19007 2148 19011 2204
rect 18947 2144 19011 2148
<< metal4 >>
rect 3163 7104 3483 7664
rect 3163 7040 3171 7104
rect 3235 7040 3251 7104
rect 3315 7040 3331 7104
rect 3395 7040 3411 7104
rect 3475 7040 3483 7104
rect 3163 6016 3483 7040
rect 3163 5952 3171 6016
rect 3235 5952 3251 6016
rect 3315 5952 3331 6016
rect 3395 5952 3411 6016
rect 3475 5952 3483 6016
rect 3163 4928 3483 5952
rect 3163 4864 3171 4928
rect 3235 4864 3251 4928
rect 3315 4864 3331 4928
rect 3395 4864 3411 4928
rect 3475 4864 3483 4928
rect 3163 3840 3483 4864
rect 3163 3776 3171 3840
rect 3235 3776 3251 3840
rect 3315 3776 3331 3840
rect 3395 3776 3411 3840
rect 3475 3776 3483 3840
rect 3163 2752 3483 3776
rect 3163 2688 3171 2752
rect 3235 2688 3251 2752
rect 3315 2688 3331 2752
rect 3395 2688 3411 2752
rect 3475 2688 3483 2752
rect 3163 2128 3483 2688
rect 5382 7648 5702 7664
rect 5382 7584 5390 7648
rect 5454 7584 5470 7648
rect 5534 7584 5550 7648
rect 5614 7584 5630 7648
rect 5694 7584 5702 7648
rect 5382 6560 5702 7584
rect 5382 6496 5390 6560
rect 5454 6496 5470 6560
rect 5534 6496 5550 6560
rect 5614 6496 5630 6560
rect 5694 6496 5702 6560
rect 5382 5472 5702 6496
rect 5382 5408 5390 5472
rect 5454 5408 5470 5472
rect 5534 5408 5550 5472
rect 5614 5408 5630 5472
rect 5694 5408 5702 5472
rect 5382 4384 5702 5408
rect 5382 4320 5390 4384
rect 5454 4320 5470 4384
rect 5534 4320 5550 4384
rect 5614 4320 5630 4384
rect 5694 4320 5702 4384
rect 5382 3296 5702 4320
rect 5382 3232 5390 3296
rect 5454 3232 5470 3296
rect 5534 3232 5550 3296
rect 5614 3232 5630 3296
rect 5694 3232 5702 3296
rect 5382 2208 5702 3232
rect 5382 2144 5390 2208
rect 5454 2144 5470 2208
rect 5534 2144 5550 2208
rect 5614 2144 5630 2208
rect 5694 2144 5702 2208
rect 5382 2128 5702 2144
rect 7602 7104 7922 7664
rect 7602 7040 7610 7104
rect 7674 7040 7690 7104
rect 7754 7040 7770 7104
rect 7834 7040 7850 7104
rect 7914 7040 7922 7104
rect 7602 6016 7922 7040
rect 7602 5952 7610 6016
rect 7674 5952 7690 6016
rect 7754 5952 7770 6016
rect 7834 5952 7850 6016
rect 7914 5952 7922 6016
rect 7602 4928 7922 5952
rect 7602 4864 7610 4928
rect 7674 4864 7690 4928
rect 7754 4864 7770 4928
rect 7834 4864 7850 4928
rect 7914 4864 7922 4928
rect 7602 3840 7922 4864
rect 7602 3776 7610 3840
rect 7674 3776 7690 3840
rect 7754 3776 7770 3840
rect 7834 3776 7850 3840
rect 7914 3776 7922 3840
rect 7602 2752 7922 3776
rect 7602 2688 7610 2752
rect 7674 2688 7690 2752
rect 7754 2688 7770 2752
rect 7834 2688 7850 2752
rect 7914 2688 7922 2752
rect 7602 2128 7922 2688
rect 9821 7648 10141 7664
rect 9821 7584 9829 7648
rect 9893 7584 9909 7648
rect 9973 7584 9989 7648
rect 10053 7584 10069 7648
rect 10133 7584 10141 7648
rect 9821 6560 10141 7584
rect 9821 6496 9829 6560
rect 9893 6496 9909 6560
rect 9973 6496 9989 6560
rect 10053 6496 10069 6560
rect 10133 6496 10141 6560
rect 9821 5472 10141 6496
rect 9821 5408 9829 5472
rect 9893 5408 9909 5472
rect 9973 5408 9989 5472
rect 10053 5408 10069 5472
rect 10133 5408 10141 5472
rect 9821 4384 10141 5408
rect 9821 4320 9829 4384
rect 9893 4320 9909 4384
rect 9973 4320 9989 4384
rect 10053 4320 10069 4384
rect 10133 4320 10141 4384
rect 9821 3296 10141 4320
rect 9821 3232 9829 3296
rect 9893 3232 9909 3296
rect 9973 3232 9989 3296
rect 10053 3232 10069 3296
rect 10133 3232 10141 3296
rect 9821 2208 10141 3232
rect 9821 2144 9829 2208
rect 9893 2144 9909 2208
rect 9973 2144 9989 2208
rect 10053 2144 10069 2208
rect 10133 2144 10141 2208
rect 9821 2128 10141 2144
rect 12041 7104 12361 7664
rect 12041 7040 12049 7104
rect 12113 7040 12129 7104
rect 12193 7040 12209 7104
rect 12273 7040 12289 7104
rect 12353 7040 12361 7104
rect 12041 6016 12361 7040
rect 12041 5952 12049 6016
rect 12113 5952 12129 6016
rect 12193 5952 12209 6016
rect 12273 5952 12289 6016
rect 12353 5952 12361 6016
rect 12041 4928 12361 5952
rect 12041 4864 12049 4928
rect 12113 4864 12129 4928
rect 12193 4864 12209 4928
rect 12273 4864 12289 4928
rect 12353 4864 12361 4928
rect 12041 3840 12361 4864
rect 12041 3776 12049 3840
rect 12113 3776 12129 3840
rect 12193 3776 12209 3840
rect 12273 3776 12289 3840
rect 12353 3776 12361 3840
rect 12041 2752 12361 3776
rect 12041 2688 12049 2752
rect 12113 2688 12129 2752
rect 12193 2688 12209 2752
rect 12273 2688 12289 2752
rect 12353 2688 12361 2752
rect 12041 2128 12361 2688
rect 14260 7648 14580 7664
rect 14260 7584 14268 7648
rect 14332 7584 14348 7648
rect 14412 7584 14428 7648
rect 14492 7584 14508 7648
rect 14572 7584 14580 7648
rect 14260 6560 14580 7584
rect 14260 6496 14268 6560
rect 14332 6496 14348 6560
rect 14412 6496 14428 6560
rect 14492 6496 14508 6560
rect 14572 6496 14580 6560
rect 14260 5472 14580 6496
rect 14260 5408 14268 5472
rect 14332 5408 14348 5472
rect 14412 5408 14428 5472
rect 14492 5408 14508 5472
rect 14572 5408 14580 5472
rect 14260 4384 14580 5408
rect 14260 4320 14268 4384
rect 14332 4320 14348 4384
rect 14412 4320 14428 4384
rect 14492 4320 14508 4384
rect 14572 4320 14580 4384
rect 14260 3296 14580 4320
rect 14260 3232 14268 3296
rect 14332 3232 14348 3296
rect 14412 3232 14428 3296
rect 14492 3232 14508 3296
rect 14572 3232 14580 3296
rect 14260 2208 14580 3232
rect 14260 2144 14268 2208
rect 14332 2144 14348 2208
rect 14412 2144 14428 2208
rect 14492 2144 14508 2208
rect 14572 2144 14580 2208
rect 14260 2128 14580 2144
rect 16480 7104 16800 7664
rect 16480 7040 16488 7104
rect 16552 7040 16568 7104
rect 16632 7040 16648 7104
rect 16712 7040 16728 7104
rect 16792 7040 16800 7104
rect 16480 6016 16800 7040
rect 16480 5952 16488 6016
rect 16552 5952 16568 6016
rect 16632 5952 16648 6016
rect 16712 5952 16728 6016
rect 16792 5952 16800 6016
rect 16480 4928 16800 5952
rect 16480 4864 16488 4928
rect 16552 4864 16568 4928
rect 16632 4864 16648 4928
rect 16712 4864 16728 4928
rect 16792 4864 16800 4928
rect 16480 3840 16800 4864
rect 16480 3776 16488 3840
rect 16552 3776 16568 3840
rect 16632 3776 16648 3840
rect 16712 3776 16728 3840
rect 16792 3776 16800 3840
rect 16480 2752 16800 3776
rect 16480 2688 16488 2752
rect 16552 2688 16568 2752
rect 16632 2688 16648 2752
rect 16712 2688 16728 2752
rect 16792 2688 16800 2752
rect 16480 2128 16800 2688
rect 18699 7648 19019 7664
rect 18699 7584 18707 7648
rect 18771 7584 18787 7648
rect 18851 7584 18867 7648
rect 18931 7584 18947 7648
rect 19011 7584 19019 7648
rect 18699 6560 19019 7584
rect 18699 6496 18707 6560
rect 18771 6496 18787 6560
rect 18851 6496 18867 6560
rect 18931 6496 18947 6560
rect 19011 6496 19019 6560
rect 18699 5472 19019 6496
rect 18699 5408 18707 5472
rect 18771 5408 18787 5472
rect 18851 5408 18867 5472
rect 18931 5408 18947 5472
rect 19011 5408 19019 5472
rect 18699 4384 19019 5408
rect 18699 4320 18707 4384
rect 18771 4320 18787 4384
rect 18851 4320 18867 4384
rect 18931 4320 18947 4384
rect 19011 4320 19019 4384
rect 18699 3296 19019 4320
rect 18699 3232 18707 3296
rect 18771 3232 18787 3296
rect 18851 3232 18867 3296
rect 18931 3232 18947 3296
rect 19011 3232 19019 3296
rect 18699 2208 19019 3232
rect 18699 2144 18707 2208
rect 18771 2144 18787 2208
rect 18851 2144 18867 2208
rect 18931 2144 18947 2208
rect 19011 2144 19019 2208
rect 18699 2128 19019 2144
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 10120 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold1_A
timestamp 1667941163
transform -1 0 5060 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1667941163
transform -1 0 9660 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3 pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26 pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29 pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33 pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 4140 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1667941163
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57 pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1667941163
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1667941163
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1667941163
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_107
timestamp 1667941163
transform 1 0 10948 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1667941163
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_113
timestamp 1667941163
transform 1 0 11500 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117
timestamp 1667941163
transform 1 0 11868 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1667941163
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1667941163
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_163
timestamp 1667941163
transform 1 0 16100 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1667941163
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_169 pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 16652 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_177
timestamp 1667941163
transform 1 0 17388 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_182
timestamp 1667941163
transform 1 0 17848 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3 pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1380 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_29
timestamp 1667941163
transform 1 0 3772 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1667941163
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_57
timestamp 1667941163
transform 1 0 6348 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_65
timestamp 1667941163
transform 1 0 7084 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_86
timestamp 1667941163
transform 1 0 9016 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1667941163
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_113
timestamp 1667941163
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_135
timestamp 1667941163
transform 1 0 13524 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_143
timestamp 1667941163
transform 1 0 14260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_155
timestamp 1667941163
transform 1 0 15364 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1667941163
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1667941163
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_181
timestamp 1667941163
transform 1 0 17756 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_189
timestamp 1667941163
transform 1 0 18492 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_3
timestamp 1667941163
transform 1 0 1380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1667941163
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_29
timestamp 1667941163
transform 1 0 3772 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_57
timestamp 1667941163
transform 1 0 6348 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_81
timestamp 1667941163
transform 1 0 8556 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_85
timestamp 1667941163
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_91
timestamp 1667941163
transform 1 0 9476 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_100
timestamp 1667941163
transform 1 0 10304 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_106
timestamp 1667941163
transform 1 0 10856 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_110
timestamp 1667941163
transform 1 0 11224 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1667941163
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1667941163
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1667941163
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1667941163
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1667941163
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_189
timestamp 1667941163
transform 1 0 18492 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_3
timestamp 1667941163
transform 1 0 1380 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_11
timestamp 1667941163
transform 1 0 2116 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_15
timestamp 1667941163
transform 1 0 2484 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_39
timestamp 1667941163
transform 1 0 4692 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_46
timestamp 1667941163
transform 1 0 5336 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 1667941163
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_57
timestamp 1667941163
transform 1 0 6348 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_63
timestamp 1667941163
transform 1 0 6900 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_80
timestamp 1667941163
transform 1 0 8464 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_84
timestamp 1667941163
transform 1 0 8832 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1667941163
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1667941163
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_113
timestamp 1667941163
transform 1 0 11500 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_135
timestamp 1667941163
transform 1 0 13524 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_159
timestamp 1667941163
transform 1 0 15732 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1667941163
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1667941163
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_181
timestamp 1667941163
transform 1 0 17756 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_189
timestamp 1667941163
transform 1 0 18492 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_3
timestamp 1667941163
transform 1 0 1380 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_11
timestamp 1667941163
transform 1 0 2116 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_22
timestamp 1667941163
transform 1 0 3128 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp 1667941163
transform 1 0 3772 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_37
timestamp 1667941163
transform 1 0 4508 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_43
timestamp 1667941163
transform 1 0 5060 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_51
timestamp 1667941163
transform 1 0 5796 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_58
timestamp 1667941163
transform 1 0 6440 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_67
timestamp 1667941163
transform 1 0 7268 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp 1667941163
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_85
timestamp 1667941163
transform 1 0 8924 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_92
timestamp 1667941163
transform 1 0 9568 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_98
timestamp 1667941163
transform 1 0 10120 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_107
timestamp 1667941163
transform 1 0 10948 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_114
timestamp 1667941163
transform 1 0 11592 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_127
timestamp 1667941163
transform 1 0 12788 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_134
timestamp 1667941163
transform 1 0 13432 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1667941163
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_158
timestamp 1667941163
transform 1 0 15640 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_165
timestamp 1667941163
transform 1 0 16284 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_172
timestamp 1667941163
transform 1 0 16928 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_184
timestamp 1667941163
transform 1 0 18032 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1667941163
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_15
timestamp 1667941163
transform 1 0 2484 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_38
timestamp 1667941163
transform 1 0 4600 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_50
timestamp 1667941163
transform 1 0 5704 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_5_57
timestamp 1667941163
transform 1 0 6348 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_69
timestamp 1667941163
transform 1 0 7452 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_93
timestamp 1667941163
transform 1 0 9660 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_106
timestamp 1667941163
transform 1 0 10856 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_113
timestamp 1667941163
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_124
timestamp 1667941163
transform 1 0 12512 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1667941163
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1667941163
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1667941163
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1667941163
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1667941163
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_181
timestamp 1667941163
transform 1 0 17756 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_189
timestamp 1667941163
transform 1 0 18492 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1667941163
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1667941163
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1667941163
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1667941163
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1667941163
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_53
timestamp 1667941163
transform 1 0 5980 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_6_64
timestamp 1667941163
transform 1 0 6992 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_79
timestamp 1667941163
transform 1 0 8372 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1667941163
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1667941163
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1667941163
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_109
timestamp 1667941163
transform 1 0 11132 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_118
timestamp 1667941163
transform 1 0 11960 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_126
timestamp 1667941163
transform 1 0 12696 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_132
timestamp 1667941163
transform 1 0 13248 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1667941163
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1667941163
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1667941163
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1667941163
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_189
timestamp 1667941163
transform 1 0 18492 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1667941163
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1667941163
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1667941163
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1667941163
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1667941163
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1667941163
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1667941163
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_69
timestamp 1667941163
transform 1 0 7452 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_80
timestamp 1667941163
transform 1 0 8464 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_92
timestamp 1667941163
transform 1 0 9568 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_104
timestamp 1667941163
transform 1 0 10672 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1667941163
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1667941163
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1667941163
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1667941163
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1667941163
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1667941163
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1667941163
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_181
timestamp 1667941163
transform 1 0 17756 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_189
timestamp 1667941163
transform 1 0 18492 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1667941163
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1667941163
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1667941163
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1667941163
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1667941163
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1667941163
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1667941163
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1667941163
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1667941163
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1667941163
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1667941163
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1667941163
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1667941163
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1667941163
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1667941163
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1667941163
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1667941163
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1667941163
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1667941163
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_189
timestamp 1667941163
transform 1 0 18492 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1667941163
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_9
timestamp 1667941163
transform 1 0 1932 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_21
timestamp 1667941163
transform 1 0 3036 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_27
timestamp 1667941163
transform 1 0 3588 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_29
timestamp 1667941163
transform 1 0 3772 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_35
timestamp 1667941163
transform 1 0 4324 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_47
timestamp 1667941163
transform 1 0 5428 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_53
timestamp 1667941163
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1667941163
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_69
timestamp 1667941163
transform 1 0 7452 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_77
timestamp 1667941163
transform 1 0 8188 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_83
timestamp 1667941163
transform 1 0 8740 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_85
timestamp 1667941163
transform 1 0 8924 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_93
timestamp 1667941163
transform 1 0 9660 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_101
timestamp 1667941163
transform 1 0 10396 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_109
timestamp 1667941163
transform 1 0 11132 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_113
timestamp 1667941163
transform 1 0 11500 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1667941163
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_137
timestamp 1667941163
transform 1 0 13708 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_141
timestamp 1667941163
transform 1 0 14076 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1667941163
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1667941163
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1667941163
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_169
timestamp 1667941163
transform 1 0 16652 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_175
timestamp 1667941163
transform 1 0 17204 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_183
timestamp 1667941163
transform 1 0 17940 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_188
timestamp 1667941163
transform 1 0 18400 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1667941163
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1667941163
transform -1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1667941163
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1667941163
transform -1 0 18860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1667941163
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1667941163
transform -1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1667941163
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1667941163
transform -1 0 18860 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1667941163
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1667941163
transform -1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1667941163
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1667941163
transform -1 0 18860 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1667941163
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1667941163
transform -1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1667941163
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1667941163
transform -1 0 18860 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1667941163
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1667941163
transform -1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1667941163
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1667941163
transform -1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_20 pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_21
timestamp 1667941163
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_22
timestamp 1667941163
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_23
timestamp 1667941163
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_24
timestamp 1667941163
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_25
timestamp 1667941163
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_26
timestamp 1667941163
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_27
timestamp 1667941163
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28
timestamp 1667941163
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1667941163
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1667941163
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1667941163
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1667941163
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1667941163
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1667941163
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1667941163
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1667941163
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1667941163
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1667941163
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1667941163
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1667941163
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1667941163
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1667941163
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1667941163
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1667941163
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1667941163
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1667941163
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1667941163
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1667941163
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1667941163
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1667941163
transform 1 0 3680 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1667941163
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1667941163
transform 1 0 8832 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1667941163
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1667941163
transform 1 0 13984 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1667941163
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _25_ pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 10856 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _26_ pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 10488 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _27_ pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 11224 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _28_
timestamp 1667941163
transform -1 0 13708 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _29_
timestamp 1667941163
transform 1 0 15180 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _30_
timestamp 1667941163
transform 1 0 16652 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _31_
timestamp 1667941163
transform -1 0 12788 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _32_
timestamp 1667941163
transform 1 0 12788 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _33_
timestamp 1667941163
transform 1 0 16008 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _34_
timestamp 1667941163
transform 1 0 11684 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _35_
timestamp 1667941163
transform 1 0 11500 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _36_
timestamp 1667941163
transform 1 0 13156 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _37_
timestamp 1667941163
transform 1 0 7820 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _38_
timestamp 1667941163
transform -1 0 6440 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _39_
timestamp 1667941163
transform 1 0 6624 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _40_
timestamp 1667941163
transform -1 0 8372 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _41_
timestamp 1667941163
transform 1 0 8004 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _42_
timestamp 1667941163
transform -1 0 11592 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _43_
timestamp 1667941163
transform 1 0 6624 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _44_
timestamp 1667941163
transform 1 0 6808 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _45_
timestamp 1667941163
transform 1 0 6716 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _46_
timestamp 1667941163
transform -1 0 8464 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _47_
timestamp 1667941163
transform 1 0 9108 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _48_
timestamp 1667941163
transform 1 0 10028 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _49_ pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 13524 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _50_
timestamp 1667941163
transform 1 0 6716 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _51_
timestamp 1667941163
transform 1 0 1656 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _52_
timestamp 1667941163
transform 1 0 2760 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _53_
timestamp 1667941163
transform 1 0 2852 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _54_
timestamp 1667941163
transform 1 0 13892 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _55_
timestamp 1667941163
transform 1 0 4232 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _56_
timestamp 1667941163
transform -1 0 9016 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _57_
timestamp 1667941163
transform -1 0 10948 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _58_
timestamp 1667941163
transform -1 0 13800 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _59_
timestamp 1667941163
transform -1 0 16100 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  _60__15 pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 5336 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  _60_ pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 4140 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _61_
timestamp 1667941163
transform 1 0 1656 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _62_
timestamp 1667941163
transform -1 0 3772 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _63_
timestamp 1667941163
transform 1 0 7820 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _64_
timestamp 1667941163
transform -1 0 13800 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _65_
timestamp 1667941163
transform -1 0 13524 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 8924 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1667941163
transform -1 0 6348 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1667941163
transform 1 0 9384 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_4  fanout13 pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 4508 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout14 pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 9108 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform -1 0 3128 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  input1 pdk_1/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 10028 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1667941163
transform -1 0 2484 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output3
timestamp 1667941163
transform -1 0 1932 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output4
timestamp 1667941163
transform -1 0 4324 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output5
timestamp 1667941163
transform -1 0 5980 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp 1667941163
transform -1 0 8188 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp 1667941163
transform 1 0 12236 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp 1667941163
transform 1 0 14444 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 1667941163
transform 1 0 16836 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1667941163
transform 1 0 18032 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 1667941163
transform 1 0 17480 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1667941163
transform 1 0 13892 0 -1 3264
box -38 -48 406 592
<< labels >>
flabel metal2 s 7470 0 7526 800 0 FreeSans 224 90 0 0 clk
port 0 nsew signal input
flabel metal2 s 9954 9200 10010 10000 0 FreeSans 224 90 0 0 comp
port 1 nsew signal input
flabel metal2 s 1122 9200 1178 10000 0 FreeSans 224 90 0 0 dq[0]
port 2 nsew signal tristate
flabel metal2 s 3330 9200 3386 10000 0 FreeSans 224 90 0 0 dq[1]
port 3 nsew signal tristate
flabel metal2 s 5538 9200 5594 10000 0 FreeSans 224 90 0 0 dq[2]
port 4 nsew signal tristate
flabel metal2 s 7746 9200 7802 10000 0 FreeSans 224 90 0 0 dq[3]
port 5 nsew signal tristate
flabel metal2 s 12162 9200 12218 10000 0 FreeSans 224 90 0 0 dq[4]
port 6 nsew signal tristate
flabel metal2 s 14370 9200 14426 10000 0 FreeSans 224 90 0 0 dq[5]
port 7 nsew signal tristate
flabel metal2 s 16578 9200 16634 10000 0 FreeSans 224 90 0 0 dq[6]
port 8 nsew signal tristate
flabel metal2 s 18786 9200 18842 10000 0 FreeSans 224 90 0 0 dq[7]
port 9 nsew signal tristate
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 last_cycle
port 10 nsew signal tristate
flabel metal2 s 2502 0 2558 800 0 FreeSans 224 90 0 0 rst_n
port 11 nsew signal input
flabel metal2 s 12438 0 12494 800 0 FreeSans 224 90 0 0 valid
port 12 nsew signal tristate
flabel metal4 s 3163 2128 3483 7664 0 FreeSans 1920 90 0 0 vccd1
port 13 nsew power bidirectional
flabel metal4 s 7602 2128 7922 7664 0 FreeSans 1920 90 0 0 vccd1
port 13 nsew power bidirectional
flabel metal4 s 12041 2128 12361 7664 0 FreeSans 1920 90 0 0 vccd1
port 13 nsew power bidirectional
flabel metal4 s 16480 2128 16800 7664 0 FreeSans 1920 90 0 0 vccd1
port 13 nsew power bidirectional
flabel metal4 s 5382 2128 5702 7664 0 FreeSans 1920 90 0 0 vssd1
port 14 nsew ground bidirectional
flabel metal4 s 9821 2128 10141 7664 0 FreeSans 1920 90 0 0 vssd1
port 14 nsew ground bidirectional
flabel metal4 s 14260 2128 14580 7664 0 FreeSans 1920 90 0 0 vssd1
port 14 nsew ground bidirectional
flabel metal4 s 18699 2128 19019 7664 0 FreeSans 1920 90 0 0 vssd1
port 14 nsew ground bidirectional
rlabel metal1 9982 7072 9982 7072 0 vccd1
rlabel via1 10061 7616 10061 7616 0 vssd1
rlabel metal2 11178 3842 11178 3842 0 _00_
rlabel metal2 16882 3672 16882 3672 0 _01_
rlabel metal2 16054 4080 16054 4080 0 _02_
rlabel metal1 13202 4488 13202 4488 0 _03_
rlabel metal1 4922 4046 4922 4046 0 _04_
rlabel metal1 14122 4046 14122 4046 0 _05_
rlabel metal1 4600 2482 4600 2482 0 _06_
rlabel via1 8700 3094 8700 3094 0 _07_
rlabel metal2 10534 4794 10534 4794 0 _08_
rlabel metal2 10994 3978 10994 3978 0 _09_
rlabel metal2 15226 4794 15226 4794 0 _10_
rlabel metal1 16721 4590 16721 4590 0 _11_
rlabel metal1 12788 4794 12788 4794 0 _12_
rlabel metal1 16238 4624 16238 4624 0 _13_
rlabel metal1 11638 5338 11638 5338 0 _14_
rlabel metal1 13248 4590 13248 4590 0 _15_
rlabel metal1 6394 4624 6394 4624 0 _16_
rlabel metal2 6854 4284 6854 4284 0 _17_
rlabel metal1 8188 5882 8188 5882 0 _18_
rlabel metal1 11178 4590 11178 4590 0 _19_
rlabel metal2 6854 4794 6854 4794 0 _20_
rlabel metal1 7084 4794 7084 4794 0 _21_
rlabel metal2 8418 4386 8418 4386 0 _22_
rlabel metal2 10258 3978 10258 3978 0 _23_
rlabel metal1 9798 4590 9798 4590 0 clk
rlabel metal2 9430 3502 9430 3502 0 clknet_0_clk
rlabel metal1 2116 2482 2116 2482 0 clknet_1_0__leaf_clk
rlabel metal1 14904 2482 14904 2482 0 clknet_1_1__leaf_clk
rlabel metal1 10212 7446 10212 7446 0 comp
rlabel metal1 1426 7514 1426 7514 0 dq[0]
rlabel metal1 3726 7514 3726 7514 0 dq[1]
rlabel metal2 5750 8415 5750 8415 0 dq[2]
rlabel metal2 7958 8415 7958 8415 0 dq[3]
rlabel metal2 12374 8415 12374 8415 0 dq[4]
rlabel metal2 14674 8415 14674 8415 0 dq[5]
rlabel metal1 16836 7514 16836 7514 0 dq[6]
rlabel metal1 18354 7514 18354 7514 0 dq[7]
rlabel metal2 17434 1520 17434 1520 0 last_cycle
rlabel metal2 12466 4998 12466 4998 0 net1
rlabel metal1 18078 7344 18078 7344 0 net10
rlabel metal2 1978 2754 1978 2754 0 net11
rlabel metal2 13938 4046 13938 4046 0 net12
rlabel metal1 13708 4182 13708 4182 0 net13
rlabel metal2 9338 2519 9338 2519 0 net14
rlabel metal2 4554 3502 4554 3502 0 net15
rlabel metal2 2254 4284 2254 4284 0 net16
rlabel metal1 4692 4522 4692 4522 0 net2
rlabel metal1 1886 7344 1886 7344 0 net3
rlabel metal1 8004 4250 8004 4250 0 net4
rlabel metal1 6532 2618 6532 2618 0 net5
rlabel metal2 13110 3961 13110 3961 0 net6
rlabel metal1 7774 4454 7774 4454 0 net7
rlabel metal1 14168 7378 14168 7378 0 net8
rlabel metal2 16882 6052 16882 6052 0 net9
rlabel metal2 2714 3213 2714 3213 0 rst_n
rlabel metal1 7222 5100 7222 5100 0 sr\[1\]
rlabel metal1 8694 2618 8694 2618 0 sr\[2\]
rlabel metal1 9338 2482 9338 2482 0 sr\[3\]
rlabel metal1 12604 2482 12604 2482 0 sr\[4\]
rlabel metal1 13478 3400 13478 3400 0 sr\[5\]
rlabel metal1 13064 3094 13064 3094 0 sr\[6\]
rlabel metal2 15778 2618 15778 2618 0 sr\[7\]
rlabel metal2 12466 1792 12466 1792 0 valid
<< properties >>
string FIXED_BBOX 0 0 20000 10000
<< end >>
