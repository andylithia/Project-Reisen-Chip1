magic
tech sky130A
magscale 1 2
timestamp 1670863290
<< nwell >>
rect 1066 6789 18898 7355
rect 1066 5701 18898 6267
rect 1066 4613 18898 5179
rect 1066 3525 18898 4091
rect 1066 2437 18898 3003
<< pwell >>
rect 1133 7595 1167 7633
rect 1411 7604 1443 7626
rect 1869 7595 1903 7633
rect 1961 7595 1995 7633
rect 3065 7595 3099 7633
rect 3616 7605 3640 7627
rect 3803 7604 3835 7626
rect 4261 7595 4295 7633
rect 4353 7595 4387 7633
rect 5459 7604 5491 7626
rect 5917 7595 5951 7633
rect 6009 7595 6043 7633
rect 6377 7595 6411 7633
rect 7481 7595 7515 7633
rect 8125 7595 8159 7633
rect 8217 7595 8251 7633
rect 8768 7605 8792 7627
rect 8953 7595 8987 7633
rect 9597 7603 9631 7633
rect 1105 7433 1379 7595
rect 1565 7459 1931 7595
rect 1565 7413 1834 7459
rect 1933 7433 3035 7595
rect 3037 7433 3587 7595
rect 3683 7421 3769 7578
rect 3957 7459 4323 7595
rect 3957 7413 4226 7459
rect 4325 7433 5427 7595
rect 5613 7459 5979 7595
rect 5613 7413 5882 7459
rect 5981 7433 6255 7595
rect 6259 7421 6345 7578
rect 6349 7433 7451 7595
rect 7453 7433 7819 7595
rect 7821 7459 8187 7595
rect 7821 7413 8090 7459
rect 8189 7433 8739 7595
rect 8835 7421 8921 7578
rect 8925 7433 9475 7595
rect 9477 7413 9655 7603
rect 9689 7595 9723 7633
rect 10057 7595 10091 7633
rect 10425 7595 10459 7633
rect 11161 7595 11195 7633
rect 11529 7595 11563 7633
rect 12265 7595 12299 7633
rect 12633 7595 12667 7633
rect 13737 7595 13771 7633
rect 14105 7595 14139 7633
rect 14473 7595 14507 7633
rect 14841 7595 14875 7633
rect 15945 7595 15979 7633
rect 16496 7605 16520 7627
rect 16683 7604 16715 7626
rect 16865 7595 16899 7633
rect 17233 7595 17267 7633
rect 17968 7605 17992 7627
rect 18061 7595 18095 7633
rect 18431 7604 18463 7626
rect 18797 7595 18831 7633
rect 9661 7433 10027 7595
rect 10029 7459 10395 7595
rect 10397 7433 11131 7595
rect 11133 7433 11407 7595
rect 11411 7421 11497 7578
rect 11501 7433 12235 7595
rect 12237 7459 12603 7595
rect 12334 7413 12603 7459
rect 12605 7433 13707 7595
rect 13709 7433 13983 7595
rect 13987 7421 14073 7578
rect 14077 7433 14443 7595
rect 14445 7459 14811 7595
rect 14542 7413 14811 7459
rect 14813 7433 15915 7595
rect 15917 7433 16467 7595
rect 16563 7421 16649 7578
rect 16837 7459 17203 7595
rect 16934 7413 17203 7459
rect 17205 7433 17939 7595
rect 18033 7459 18399 7595
rect 18130 7413 18399 7459
rect 18585 7433 18859 7595
rect 1105 6549 1379 6711
rect 1381 6549 2483 6711
rect 2485 6549 3587 6711
rect 3683 6566 3769 6723
rect 3773 6549 4875 6711
rect 4877 6549 5979 6711
rect 5981 6549 7083 6711
rect 7085 6549 8187 6711
rect 8189 6549 8739 6711
rect 8835 6566 8921 6723
rect 8925 6549 10027 6711
rect 10029 6549 11131 6711
rect 11133 6549 12235 6711
rect 12237 6549 13339 6711
rect 13341 6549 13891 6711
rect 13987 6566 14073 6723
rect 14077 6549 15179 6711
rect 15181 6549 16283 6711
rect 16285 6549 17387 6711
rect 17389 6549 18491 6711
rect 18585 6549 18859 6711
rect 1133 6507 1167 6549
rect 1409 6507 1443 6549
rect 2513 6507 2547 6549
rect 3617 6539 3651 6545
rect 3616 6517 3651 6539
rect 3617 6507 3651 6517
rect 3801 6511 3835 6549
rect 4721 6507 4755 6545
rect 4905 6511 4939 6549
rect 5825 6507 5859 6545
rect 6009 6511 6043 6549
rect 6192 6517 6216 6539
rect 6377 6507 6411 6545
rect 7113 6511 7147 6549
rect 7481 6507 7515 6545
rect 8033 6511 8067 6545
rect 8217 6511 8251 6549
rect 8034 6507 8067 6511
rect 8493 6507 8527 6545
rect 8768 6517 8792 6539
rect 8953 6511 8987 6549
rect 9597 6507 9631 6545
rect 10057 6511 10091 6549
rect 10701 6507 10735 6545
rect 11161 6511 11195 6549
rect 11529 6507 11563 6545
rect 12265 6511 12299 6549
rect 12633 6507 12667 6545
rect 13369 6511 13403 6549
rect 13737 6507 13771 6545
rect 13920 6517 13944 6539
rect 14105 6511 14139 6549
rect 14841 6507 14875 6545
rect 15209 6511 15243 6549
rect 15945 6507 15979 6545
rect 16313 6511 16347 6549
rect 16496 6517 16520 6539
rect 16681 6507 16715 6545
rect 17417 6511 17451 6549
rect 17785 6507 17819 6545
rect 18520 6517 18544 6539
rect 18797 6507 18831 6549
rect 1105 6345 1379 6507
rect 1381 6345 2483 6507
rect 2485 6345 3587 6507
rect 3589 6345 4691 6507
rect 4693 6345 5795 6507
rect 5797 6345 6163 6507
rect 6259 6333 6345 6490
rect 6349 6345 7451 6507
rect 7453 6345 8003 6507
rect 8034 6371 8401 6507
rect 8215 6325 8401 6371
rect 8465 6345 9567 6507
rect 9569 6345 10671 6507
rect 10673 6345 11407 6507
rect 11411 6333 11497 6490
rect 11501 6345 12603 6507
rect 12605 6345 13707 6507
rect 13709 6345 14811 6507
rect 14813 6345 15915 6507
rect 15917 6345 16467 6507
rect 16563 6333 16649 6490
rect 16653 6345 17755 6507
rect 17757 6345 18491 6507
rect 18585 6345 18859 6507
rect 1105 5461 1379 5623
rect 1381 5461 2483 5623
rect 2485 5461 3587 5623
rect 3683 5478 3769 5635
rect 3773 5461 4875 5623
rect 4877 5461 5979 5623
rect 5981 5461 6715 5623
rect 6717 5461 6991 5617
rect 6993 5461 7543 5623
rect 8185 5597 8371 5643
rect 7591 5461 8371 5597
rect 8373 5461 8739 5623
rect 8835 5478 8921 5635
rect 8925 5461 10027 5623
rect 10029 5461 11131 5623
rect 11133 5461 11499 5623
rect 11711 5597 11897 5643
rect 11530 5461 11897 5597
rect 11961 5461 12695 5623
rect 12999 5597 13185 5643
rect 12818 5461 13185 5597
rect 13249 5461 13983 5623
rect 13987 5478 14073 5635
rect 14077 5461 15179 5623
rect 15181 5461 16283 5623
rect 16285 5461 17387 5623
rect 17389 5461 18491 5623
rect 18585 5461 18859 5623
rect 1133 5419 1167 5461
rect 1409 5419 1443 5461
rect 2513 5419 2547 5461
rect 2789 5419 2823 5457
rect 3616 5429 3640 5451
rect 3801 5423 3835 5461
rect 4629 5419 4663 5457
rect 4905 5423 4939 5461
rect 5733 5419 5767 5457
rect 6009 5423 6043 5461
rect 6377 5419 6411 5457
rect 6708 5419 6742 5457
rect 6929 5423 6963 5461
rect 7021 5423 7055 5461
rect 7481 5419 7515 5457
rect 7849 5419 7883 5457
rect 8254 5423 8288 5461
rect 8401 5423 8435 5461
rect 8768 5429 8792 5451
rect 8953 5423 8987 5461
rect 9689 5419 9723 5457
rect 10057 5423 10091 5461
rect 10738 5419 10772 5457
rect 10885 5419 10919 5457
rect 11161 5423 11195 5461
rect 11530 5457 11563 5461
rect 11529 5423 11563 5457
rect 11768 5419 11802 5457
rect 11989 5423 12023 5461
rect 12818 5457 12851 5461
rect 12541 5419 12575 5457
rect 12724 5429 12748 5451
rect 12817 5423 12851 5457
rect 13277 5423 13311 5461
rect 13590 5419 13624 5457
rect 13737 5419 13771 5457
rect 14105 5423 14139 5461
rect 14841 5419 14875 5457
rect 15209 5423 15243 5461
rect 15945 5419 15979 5457
rect 16313 5423 16347 5461
rect 16496 5429 16520 5451
rect 16681 5419 16715 5457
rect 17417 5423 17451 5461
rect 17785 5419 17819 5457
rect 18520 5429 18544 5451
rect 18797 5419 18831 5461
rect 1105 5257 1379 5419
rect 1381 5257 2483 5419
rect 2485 5257 2759 5419
rect 2761 5283 4599 5419
rect 3663 5239 3849 5283
rect 4415 5237 4599 5283
rect 4601 5257 5703 5419
rect 5705 5257 6255 5419
rect 6259 5245 6345 5402
rect 6349 5257 6623 5419
rect 6625 5283 7405 5419
rect 6625 5237 6811 5283
rect 7453 5257 7819 5419
rect 7821 5283 9659 5419
rect 8723 5239 8909 5283
rect 9475 5237 9659 5283
rect 9661 5257 10027 5419
rect 10075 5283 10855 5419
rect 10669 5237 10855 5283
rect 10857 5257 11407 5419
rect 11411 5245 11497 5402
rect 11685 5283 12465 5419
rect 11685 5237 11871 5283
rect 12513 5257 12879 5419
rect 12927 5283 13707 5419
rect 13521 5237 13707 5283
rect 13709 5257 14811 5419
rect 14813 5257 15915 5419
rect 15917 5257 16467 5419
rect 16563 5245 16649 5402
rect 16653 5257 17755 5419
rect 17757 5257 18491 5419
rect 18585 5257 18859 5419
rect 1105 4373 1379 4535
rect 1381 4373 2115 4535
rect 2117 4373 2391 4535
rect 2412 4509 2596 4555
rect 2412 4373 3105 4509
rect 3129 4373 3679 4535
rect 3683 4390 3769 4547
rect 3959 4373 4507 4509
rect 4509 4373 4875 4535
rect 1133 4331 1167 4373
rect 1409 4331 1443 4373
rect 2145 4363 2179 4373
rect 2144 4341 2179 4363
rect 2145 4335 2179 4341
rect 2237 4331 2271 4369
rect 2513 4331 2547 4369
rect 2881 4331 2915 4369
rect 3065 4335 3099 4373
rect 3157 4335 3191 4373
rect 3803 4342 3835 4364
rect 4445 4335 4479 4373
rect 4537 4335 4571 4373
rect 4721 4331 4755 4369
rect 4877 4365 5055 4555
rect 5061 4373 5795 4535
rect 6043 4509 6229 4555
rect 6043 4373 6410 4509
rect 6441 4373 6807 4535
rect 7019 4509 7205 4555
rect 6838 4373 7205 4509
rect 7269 4373 7819 4535
rect 7821 4509 8007 4555
rect 7821 4373 8601 4509
rect 8835 4390 8921 4547
rect 9319 4509 9505 4555
rect 9138 4373 9505 4509
rect 9569 4373 9935 4535
rect 4997 4335 5031 4365
rect 5089 4335 5123 4373
rect 6377 4369 6410 4373
rect 5273 4335 5307 4369
rect 5365 4331 5399 4369
rect 5827 4342 5859 4364
rect 6103 4340 6135 4362
rect 6377 4331 6411 4369
rect 6469 4335 6503 4373
rect 6838 4369 6871 4373
rect 6837 4331 6871 4369
rect 6929 4331 6963 4369
rect 7297 4335 7331 4373
rect 7904 4335 7938 4373
rect 9138 4369 9171 4373
rect 8346 4331 8380 4369
rect 8493 4331 8527 4369
rect 8679 4342 8711 4364
rect 8860 4341 8884 4363
rect 8953 4331 8987 4369
rect 9137 4335 9171 4369
rect 9597 4335 9631 4373
rect 9937 4365 10115 4555
rect 10121 4373 10487 4535
rect 10699 4509 10885 4555
rect 10518 4373 10885 4509
rect 10949 4373 11315 4535
rect 11317 4373 11591 4529
rect 11593 4373 11959 4535
rect 12601 4509 12787 4555
rect 12007 4373 12787 4509
rect 12789 4373 13155 4535
rect 13157 4373 13431 4529
rect 13433 4373 13983 4535
rect 13987 4390 14073 4547
rect 14077 4373 15179 4535
rect 15391 4509 15577 4555
rect 15210 4373 15577 4509
rect 15641 4373 16007 4535
rect 16009 4373 16283 4529
rect 16285 4373 16651 4535
rect 16653 4373 16927 4529
rect 16929 4373 18031 4535
rect 18033 4373 18583 4535
rect 18585 4373 18859 4535
rect 10057 4335 10091 4365
rect 10149 4335 10183 4373
rect 10518 4369 10551 4373
rect 10517 4335 10551 4369
rect 10793 4331 10827 4369
rect 10977 4335 11011 4373
rect 11345 4363 11379 4373
rect 11344 4341 11379 4363
rect 11345 4335 11379 4341
rect 11531 4340 11563 4362
rect 11621 4335 11655 4373
rect 12670 4335 12704 4373
rect 12817 4335 12851 4373
rect 13369 4335 13403 4373
rect 13461 4331 13495 4373
rect 13553 4331 13587 4369
rect 13921 4331 13955 4369
rect 14105 4335 14139 4373
rect 15210 4369 15243 4373
rect 15209 4335 15243 4369
rect 15669 4335 15703 4373
rect 15761 4331 15795 4369
rect 16221 4335 16255 4373
rect 16313 4335 16347 4373
rect 16496 4341 16520 4363
rect 16681 4331 16715 4369
rect 16865 4335 16899 4373
rect 16957 4335 16991 4373
rect 17785 4331 17819 4369
rect 18061 4335 18095 4373
rect 18520 4341 18544 4363
rect 18797 4331 18831 4373
rect 1105 4169 1379 4331
rect 1381 4169 2115 4331
rect 2209 4175 2483 4331
rect 2485 4169 2851 4331
rect 2853 4195 4691 4331
rect 3755 4151 3941 4195
rect 4507 4149 4691 4195
rect 4693 4169 5059 4331
rect 5337 4169 6071 4331
rect 6259 4157 6345 4314
rect 6349 4169 6623 4331
rect 6625 4175 6899 4331
rect 6901 4169 7635 4331
rect 7683 4195 8463 4331
rect 8277 4149 8463 4195
rect 8465 4169 8831 4331
rect 8925 4195 10746 4331
rect 10765 4169 11315 4331
rect 11411 4157 11497 4314
rect 11685 4195 13523 4331
rect 11685 4149 11869 4195
rect 12435 4151 12621 4195
rect 13525 4169 13891 4331
rect 13893 4195 15731 4331
rect 14795 4151 14981 4195
rect 15547 4149 15731 4195
rect 15733 4169 16467 4331
rect 16563 4157 16649 4314
rect 16653 4169 17755 4331
rect 17757 4169 18491 4331
rect 18585 4169 18859 4331
rect 1105 3285 1379 3447
rect 1381 3285 1655 3447
rect 2559 3421 2745 3465
rect 3311 3421 3495 3467
rect 1657 3285 3495 3421
rect 3683 3302 3769 3459
rect 3773 3285 4507 3447
rect 4526 3285 6347 3421
rect 6349 3285 6715 3447
rect 7619 3421 7805 3465
rect 8371 3421 8555 3467
rect 6717 3285 8555 3421
rect 8557 3285 8831 3447
rect 8835 3302 8921 3459
rect 9206 3421 9475 3467
rect 9109 3285 9475 3421
rect 9477 3285 10027 3447
rect 10029 3285 10303 3441
rect 10305 3285 10855 3447
rect 10949 3285 11223 3441
rect 11225 3285 11959 3447
rect 11961 3421 12145 3467
rect 12711 3421 12897 3465
rect 11961 3285 13799 3421
rect 13987 3302 14073 3459
rect 14077 3285 15179 3447
rect 15181 3285 16283 3447
rect 16285 3285 17387 3447
rect 17389 3285 18491 3447
rect 18585 3285 18859 3447
rect 1133 3243 1167 3285
rect 1409 3243 1443 3285
rect 1685 3247 1719 3285
rect 3527 3254 3559 3276
rect 3709 3243 3743 3281
rect 3801 3243 3835 3285
rect 4169 3243 4203 3281
rect 6103 3252 6135 3274
rect 6285 3247 6319 3285
rect 6377 3243 6411 3285
rect 6745 3247 6779 3285
rect 7112 3253 7136 3275
rect 8585 3247 8619 3285
rect 8953 3243 8987 3281
rect 9045 3243 9079 3281
rect 9137 3247 9171 3285
rect 9413 3243 9447 3281
rect 9505 3247 9539 3285
rect 10241 3247 10275 3285
rect 10333 3247 10367 3285
rect 10884 3253 10908 3275
rect 10977 3247 11011 3285
rect 11253 3247 11287 3285
rect 11531 3252 11563 3274
rect 13461 3243 13495 3281
rect 13553 3243 13587 3281
rect 13737 3247 13771 3285
rect 13831 3254 13863 3276
rect 13921 3243 13955 3281
rect 14105 3247 14139 3285
rect 14289 3243 14323 3281
rect 15209 3247 15243 3285
rect 15393 3243 15427 3281
rect 16313 3247 16347 3285
rect 16496 3253 16520 3275
rect 16681 3243 16715 3281
rect 17417 3247 17451 3285
rect 17785 3243 17819 3281
rect 18520 3253 18544 3275
rect 18797 3243 18831 3285
rect 1105 3081 1379 3243
rect 1381 3081 1931 3243
rect 1933 3107 3771 3243
rect 1933 3061 2117 3107
rect 2683 3063 2869 3107
rect 3773 3081 4139 3243
rect 4141 3107 5997 3243
rect 4413 3063 4597 3107
rect 5530 3083 5997 3107
rect 5813 3061 5997 3083
rect 6259 3069 6345 3226
rect 6349 3081 7083 3243
rect 7177 3107 9015 3243
rect 7177 3061 7361 3107
rect 7927 3063 8113 3107
rect 9017 3081 9383 3243
rect 9385 3107 11206 3243
rect 11411 3069 11497 3226
rect 11685 3107 13523 3243
rect 11685 3061 11869 3107
rect 12435 3063 12621 3107
rect 13525 3081 13891 3243
rect 13893 3107 14259 3243
rect 13990 3061 14259 3107
rect 14261 3081 15363 3243
rect 15365 3081 16467 3243
rect 16563 3069 16649 3226
rect 16653 3081 17755 3243
rect 17757 3081 18491 3243
rect 18585 3081 18859 3243
rect 1105 2197 1379 2359
rect 1381 2197 1655 2359
rect 2559 2333 2745 2377
rect 3311 2333 3495 2379
rect 1657 2197 3495 2333
rect 3683 2214 3769 2371
rect 3773 2197 4139 2359
rect 5135 2333 5321 2377
rect 5887 2333 6071 2379
rect 4233 2197 6071 2333
rect 6259 2214 6345 2371
rect 6349 2197 7451 2359
rect 7453 2197 8555 2359
rect 8557 2197 8831 2359
rect 8835 2214 8921 2371
rect 9109 2333 9293 2379
rect 9859 2333 10045 2377
rect 9109 2197 10947 2333
rect 10949 2197 11315 2359
rect 11411 2214 11497 2371
rect 11501 2197 11867 2359
rect 11961 2333 12145 2379
rect 12711 2333 12897 2377
rect 11961 2197 13799 2333
rect 13987 2214 14073 2371
rect 14261 2333 14445 2379
rect 15011 2333 15197 2377
rect 14261 2197 16099 2333
rect 16101 2197 16467 2359
rect 16563 2214 16649 2371
rect 16653 2197 17387 2359
rect 17578 2333 17847 2379
rect 17481 2197 17847 2333
rect 17849 2197 18583 2359
rect 18585 2197 18859 2359
rect 1133 2159 1167 2197
rect 1409 2159 1443 2197
rect 1685 2159 1719 2197
rect 3527 2166 3559 2188
rect 3801 2159 3835 2197
rect 4168 2165 4192 2187
rect 4261 2159 4295 2197
rect 6103 2166 6135 2188
rect 6377 2159 6411 2197
rect 7481 2159 7515 2197
rect 8585 2159 8619 2197
rect 8955 2166 8987 2188
rect 10885 2159 10919 2197
rect 10977 2159 11011 2197
rect 11344 2165 11368 2187
rect 11529 2159 11563 2197
rect 11896 2165 11920 2187
rect 13737 2159 13771 2197
rect 13831 2166 13863 2188
rect 14107 2166 14139 2188
rect 16037 2159 16071 2197
rect 16129 2159 16163 2197
rect 16496 2165 16520 2187
rect 16681 2159 16715 2197
rect 17416 2165 17440 2187
rect 17509 2159 17543 2197
rect 17877 2159 17911 2197
rect 18797 2159 18831 2197
<< scnmos >>
rect 1183 7459 1301 7569
rect 1644 7439 1674 7569
rect 1728 7439 1758 7569
rect 1823 7485 1853 7569
rect 2011 7459 2957 7569
rect 3115 7459 3509 7569
rect 4036 7439 4066 7569
rect 4120 7439 4150 7569
rect 4215 7485 4245 7569
rect 4403 7459 5349 7569
rect 5692 7439 5722 7569
rect 5776 7439 5806 7569
rect 5871 7485 5901 7569
rect 6059 7459 6177 7569
rect 6427 7459 7373 7569
rect 7531 7459 7741 7569
rect 7900 7439 7930 7569
rect 7984 7439 8014 7569
rect 8079 7485 8109 7569
rect 8267 7459 8661 7569
rect 9003 7459 9397 7569
rect 9739 7459 9949 7569
rect 10108 7485 10138 7569
rect 10203 7485 10233 7569
rect 10287 7485 10317 7569
rect 10475 7459 11053 7569
rect 11211 7459 11329 7569
rect 11579 7459 12157 7569
rect 12315 7485 12345 7569
rect 12410 7439 12440 7569
rect 12494 7439 12524 7569
rect 12683 7459 13629 7569
rect 13787 7459 13905 7569
rect 14155 7459 14365 7569
rect 14523 7485 14553 7569
rect 14618 7439 14648 7569
rect 14702 7439 14732 7569
rect 14891 7459 15837 7569
rect 15995 7459 16389 7569
rect 16915 7485 16945 7569
rect 17010 7439 17040 7569
rect 17094 7439 17124 7569
rect 17283 7459 17861 7569
rect 18111 7485 18141 7569
rect 18206 7439 18236 7569
rect 18290 7439 18320 7569
rect 18663 7459 18781 7569
rect 1183 6575 1301 6685
rect 1459 6575 2405 6685
rect 2563 6575 3509 6685
rect 3851 6575 4797 6685
rect 4955 6575 5901 6685
rect 6059 6575 7005 6685
rect 7163 6575 8109 6685
rect 8267 6575 8661 6685
rect 9003 6575 9949 6685
rect 10107 6575 11053 6685
rect 11211 6575 12157 6685
rect 12315 6575 13261 6685
rect 13419 6575 13813 6685
rect 14155 6575 15101 6685
rect 15259 6575 16205 6685
rect 16363 6575 17309 6685
rect 17467 6575 18413 6685
rect 18663 6575 18781 6685
rect 1183 6371 1301 6481
rect 1459 6371 2405 6481
rect 2563 6371 3509 6481
rect 3667 6371 4613 6481
rect 4771 6371 5717 6481
rect 5875 6371 6085 6481
rect 6427 6371 7373 6481
rect 7531 6371 7925 6481
rect 8112 6397 8142 6481
rect 8196 6397 8226 6481
rect 8293 6351 8323 6481
rect 8543 6371 9489 6481
rect 9647 6371 10593 6481
rect 10751 6371 11329 6481
rect 11579 6371 12525 6481
rect 12683 6371 13629 6481
rect 13787 6371 14733 6481
rect 14891 6371 15837 6481
rect 15995 6371 16389 6481
rect 16731 6371 17677 6481
rect 17835 6371 18413 6481
rect 18663 6371 18781 6481
rect 1183 5487 1301 5597
rect 1459 5487 2405 5597
rect 2563 5487 3509 5597
rect 3851 5487 4797 5597
rect 4955 5487 5901 5597
rect 6059 5487 6637 5597
rect 6795 5487 6825 5591
rect 6883 5487 6913 5591
rect 7071 5487 7465 5597
rect 7669 5487 7699 5571
rect 7837 5487 7867 5571
rect 7933 5487 7963 5571
rect 8058 5487 8088 5571
rect 8154 5487 8184 5571
rect 8263 5487 8293 5617
rect 8451 5487 8661 5597
rect 9003 5487 9949 5597
rect 10107 5487 11053 5597
rect 11211 5487 11421 5597
rect 11608 5487 11638 5571
rect 11692 5487 11722 5571
rect 11789 5487 11819 5617
rect 12039 5487 12617 5597
rect 12896 5487 12926 5571
rect 12980 5487 13010 5571
rect 13077 5487 13107 5617
rect 13327 5487 13905 5597
rect 14155 5487 15101 5597
rect 15259 5487 16205 5597
rect 16363 5487 17309 5597
rect 17467 5487 18413 5597
rect 18663 5487 18781 5597
rect 1183 5283 1301 5393
rect 1459 5283 2405 5393
rect 2563 5283 2681 5393
rect 2839 5309 2869 5393
rect 2923 5309 2953 5393
rect 3178 5309 3208 5393
rect 3273 5321 3303 5393
rect 3369 5321 3399 5393
rect 3535 5309 3565 5393
rect 3607 5309 3637 5393
rect 3739 5265 3769 5393
rect 3838 5321 3868 5393
rect 3947 5321 3977 5393
rect 4043 5309 4073 5393
rect 4192 5309 4222 5393
rect 4283 5309 4313 5393
rect 4491 5263 4521 5393
rect 4679 5283 5625 5393
rect 5783 5283 6177 5393
rect 6427 5283 6545 5393
rect 6703 5263 6733 5393
rect 6812 5309 6842 5393
rect 6908 5309 6938 5393
rect 7033 5309 7063 5393
rect 7129 5309 7159 5393
rect 7297 5309 7327 5393
rect 7531 5283 7741 5393
rect 7899 5309 7929 5393
rect 7983 5309 8013 5393
rect 8238 5309 8268 5393
rect 8333 5321 8363 5393
rect 8429 5321 8459 5393
rect 8595 5309 8625 5393
rect 8667 5309 8697 5393
rect 8799 5265 8829 5393
rect 8898 5321 8928 5393
rect 9007 5321 9037 5393
rect 9103 5309 9133 5393
rect 9252 5309 9282 5393
rect 9343 5309 9373 5393
rect 9551 5263 9581 5393
rect 9739 5283 9949 5393
rect 10153 5309 10183 5393
rect 10321 5309 10351 5393
rect 10417 5309 10447 5393
rect 10542 5309 10572 5393
rect 10638 5309 10668 5393
rect 10747 5263 10777 5393
rect 10935 5283 11329 5393
rect 11763 5263 11793 5393
rect 11872 5309 11902 5393
rect 11968 5309 11998 5393
rect 12093 5309 12123 5393
rect 12189 5309 12219 5393
rect 12357 5309 12387 5393
rect 12591 5283 12801 5393
rect 13005 5309 13035 5393
rect 13173 5309 13203 5393
rect 13269 5309 13299 5393
rect 13394 5309 13424 5393
rect 13490 5309 13520 5393
rect 13599 5263 13629 5393
rect 13787 5283 14733 5393
rect 14891 5283 15837 5393
rect 15995 5283 16389 5393
rect 16731 5283 17677 5393
rect 17835 5283 18413 5393
rect 18663 5283 18781 5393
rect 1183 4399 1301 4509
rect 1459 4399 2037 4509
rect 2195 4399 2313 4509
rect 2490 4399 2520 4529
rect 2585 4399 2685 4483
rect 2843 4399 2943 4483
rect 2997 4399 3027 4483
rect 3207 4399 3601 4509
rect 4043 4399 4073 4483
rect 4129 4399 4159 4483
rect 4215 4399 4245 4483
rect 4301 4399 4331 4483
rect 4398 4399 4428 4483
rect 4587 4399 4797 4509
rect 5139 4399 5717 4509
rect 6121 4399 6151 4529
rect 6218 4399 6248 4483
rect 6302 4399 6332 4483
rect 6519 4399 6729 4509
rect 6916 4399 6946 4483
rect 7000 4399 7030 4483
rect 7097 4399 7127 4529
rect 7347 4399 7741 4509
rect 7899 4399 7929 4529
rect 8008 4399 8038 4483
rect 8104 4399 8134 4483
rect 8229 4399 8259 4483
rect 8325 4399 8355 4483
rect 8493 4399 8523 4483
rect 9216 4399 9246 4483
rect 9300 4399 9330 4483
rect 9397 4399 9427 4529
rect 9647 4399 9857 4509
rect 10199 4399 10409 4509
rect 10596 4399 10626 4483
rect 10680 4399 10710 4483
rect 10777 4399 10807 4529
rect 11027 4399 11237 4509
rect 11395 4399 11425 4503
rect 11483 4399 11513 4503
rect 11671 4399 11881 4509
rect 12085 4399 12115 4483
rect 12253 4399 12283 4483
rect 12349 4399 12379 4483
rect 12474 4399 12504 4483
rect 12570 4399 12600 4483
rect 12679 4399 12709 4529
rect 12867 4399 13077 4509
rect 13235 4399 13265 4503
rect 13323 4399 13353 4503
rect 13511 4399 13905 4509
rect 14155 4399 15101 4509
rect 15288 4399 15318 4483
rect 15372 4399 15402 4483
rect 15469 4399 15499 4529
rect 15719 4399 15929 4509
rect 16087 4399 16117 4503
rect 16175 4399 16205 4503
rect 16363 4399 16573 4509
rect 16731 4399 16761 4503
rect 16819 4399 16849 4503
rect 17007 4399 17953 4509
rect 18111 4399 18505 4509
rect 18663 4399 18781 4509
rect 1183 4195 1301 4305
rect 1459 4195 2037 4305
rect 2287 4201 2317 4305
rect 2375 4201 2405 4305
rect 2563 4195 2773 4305
rect 2931 4221 2961 4305
rect 3015 4221 3045 4305
rect 3270 4221 3300 4305
rect 3365 4233 3395 4305
rect 3461 4233 3491 4305
rect 3627 4221 3657 4305
rect 3699 4221 3729 4305
rect 3831 4177 3861 4305
rect 3930 4233 3960 4305
rect 4039 4233 4069 4305
rect 4135 4221 4165 4305
rect 4284 4221 4314 4305
rect 4375 4221 4405 4305
rect 4583 4175 4613 4305
rect 4771 4195 4981 4305
rect 5415 4195 5993 4305
rect 6427 4195 6545 4305
rect 6703 4201 6733 4305
rect 6791 4201 6821 4305
rect 6979 4195 7557 4305
rect 7761 4221 7791 4305
rect 7929 4221 7959 4305
rect 8025 4221 8055 4305
rect 8150 4221 8180 4305
rect 8246 4221 8276 4305
rect 8355 4175 8385 4305
rect 8543 4195 8753 4305
rect 9004 4221 9034 4305
rect 9090 4221 9120 4305
rect 9176 4221 9206 4305
rect 9262 4221 9292 4305
rect 9348 4221 9378 4305
rect 9434 4221 9464 4305
rect 9520 4221 9550 4305
rect 9606 4221 9636 4305
rect 9692 4221 9722 4305
rect 9778 4221 9808 4305
rect 9864 4221 9894 4305
rect 9950 4221 9980 4305
rect 10035 4221 10065 4305
rect 10121 4221 10151 4305
rect 10207 4221 10237 4305
rect 10293 4221 10323 4305
rect 10379 4221 10409 4305
rect 10465 4221 10495 4305
rect 10551 4221 10581 4305
rect 10637 4221 10667 4305
rect 10843 4195 11237 4305
rect 11763 4175 11793 4305
rect 11971 4221 12001 4305
rect 12062 4221 12092 4305
rect 12211 4221 12241 4305
rect 12307 4233 12337 4305
rect 12416 4233 12446 4305
rect 12515 4177 12545 4305
rect 12647 4221 12677 4305
rect 12719 4221 12749 4305
rect 12885 4233 12915 4305
rect 12981 4233 13011 4305
rect 13076 4221 13106 4305
rect 13331 4221 13361 4305
rect 13415 4221 13445 4305
rect 13603 4195 13813 4305
rect 13971 4221 14001 4305
rect 14055 4221 14085 4305
rect 14310 4221 14340 4305
rect 14405 4233 14435 4305
rect 14501 4233 14531 4305
rect 14667 4221 14697 4305
rect 14739 4221 14769 4305
rect 14871 4177 14901 4305
rect 14970 4233 15000 4305
rect 15079 4233 15109 4305
rect 15175 4221 15205 4305
rect 15324 4221 15354 4305
rect 15415 4221 15445 4305
rect 15623 4175 15653 4305
rect 15811 4195 16389 4305
rect 16731 4195 17677 4305
rect 17835 4195 18413 4305
rect 18663 4195 18781 4305
rect 1183 3311 1301 3421
rect 1459 3311 1577 3421
rect 1735 3311 1765 3395
rect 1819 3311 1849 3395
rect 2074 3311 2104 3395
rect 2169 3311 2199 3383
rect 2265 3311 2295 3383
rect 2431 3311 2461 3395
rect 2503 3311 2533 3395
rect 2635 3311 2665 3439
rect 2734 3311 2764 3383
rect 2843 3311 2873 3383
rect 2939 3311 2969 3395
rect 3088 3311 3118 3395
rect 3179 3311 3209 3395
rect 3387 3311 3417 3441
rect 3851 3311 4429 3421
rect 4605 3311 4635 3395
rect 4691 3311 4721 3395
rect 4777 3311 4807 3395
rect 4863 3311 4893 3395
rect 4949 3311 4979 3395
rect 5035 3311 5065 3395
rect 5121 3311 5151 3395
rect 5207 3311 5237 3395
rect 5292 3311 5322 3395
rect 5378 3311 5408 3395
rect 5464 3311 5494 3395
rect 5550 3311 5580 3395
rect 5636 3311 5666 3395
rect 5722 3311 5752 3395
rect 5808 3311 5838 3395
rect 5894 3311 5924 3395
rect 5980 3311 6010 3395
rect 6066 3311 6096 3395
rect 6152 3311 6182 3395
rect 6238 3311 6268 3395
rect 6427 3311 6637 3421
rect 6795 3311 6825 3395
rect 6879 3311 6909 3395
rect 7134 3311 7164 3395
rect 7229 3311 7259 3383
rect 7325 3311 7355 3383
rect 7491 3311 7521 3395
rect 7563 3311 7593 3395
rect 7695 3311 7725 3439
rect 7794 3311 7824 3383
rect 7903 3311 7933 3383
rect 7999 3311 8029 3395
rect 8148 3311 8178 3395
rect 8239 3311 8269 3395
rect 8447 3311 8477 3441
rect 8635 3311 8753 3421
rect 9187 3311 9217 3395
rect 9282 3311 9312 3441
rect 9366 3311 9396 3441
rect 9555 3311 9949 3421
rect 10107 3311 10137 3415
rect 10195 3311 10225 3415
rect 10383 3311 10777 3421
rect 11027 3311 11057 3415
rect 11115 3311 11145 3415
rect 11303 3311 11881 3421
rect 12039 3311 12069 3441
rect 12247 3311 12277 3395
rect 12338 3311 12368 3395
rect 12487 3311 12517 3395
rect 12583 3311 12613 3383
rect 12692 3311 12722 3383
rect 12791 3311 12821 3439
rect 12923 3311 12953 3395
rect 12995 3311 13025 3395
rect 13161 3311 13191 3383
rect 13257 3311 13287 3383
rect 13352 3311 13382 3395
rect 13607 3311 13637 3395
rect 13691 3311 13721 3395
rect 14155 3311 15101 3421
rect 15259 3311 16205 3421
rect 16363 3311 17309 3421
rect 17467 3311 18413 3421
rect 18663 3311 18781 3421
rect 1183 3107 1301 3217
rect 1459 3107 1853 3217
rect 2011 3087 2041 3217
rect 2219 3133 2249 3217
rect 2310 3133 2340 3217
rect 2459 3133 2489 3217
rect 2555 3145 2585 3217
rect 2664 3145 2694 3217
rect 2763 3089 2793 3217
rect 2895 3133 2925 3217
rect 2967 3133 2997 3217
rect 3133 3145 3163 3217
rect 3229 3145 3259 3217
rect 3324 3133 3354 3217
rect 3579 3133 3609 3217
rect 3663 3133 3693 3217
rect 3851 3107 4061 3217
rect 4219 3133 4249 3217
rect 4303 3133 4333 3217
rect 4491 3089 4521 3217
rect 4586 3145 4616 3217
rect 4696 3145 4726 3217
rect 4792 3133 4822 3217
rect 4906 3133 4936 3217
rect 4978 3133 5008 3217
rect 5166 3133 5196 3217
rect 5238 3133 5268 3217
rect 5334 3133 5364 3217
rect 5406 3133 5436 3217
rect 5482 3133 5512 3217
rect 5606 3109 5636 3217
rect 5794 3133 5824 3217
rect 5889 3087 5919 3217
rect 6427 3107 7005 3217
rect 7255 3087 7285 3217
rect 7463 3133 7493 3217
rect 7554 3133 7584 3217
rect 7703 3133 7733 3217
rect 7799 3145 7829 3217
rect 7908 3145 7938 3217
rect 8007 3089 8037 3217
rect 8139 3133 8169 3217
rect 8211 3133 8241 3217
rect 8377 3145 8407 3217
rect 8473 3145 8503 3217
rect 8568 3133 8598 3217
rect 8823 3133 8853 3217
rect 8907 3133 8937 3217
rect 9095 3107 9305 3217
rect 9464 3133 9494 3217
rect 9550 3133 9580 3217
rect 9636 3133 9666 3217
rect 9722 3133 9752 3217
rect 9808 3133 9838 3217
rect 9894 3133 9924 3217
rect 9980 3133 10010 3217
rect 10066 3133 10096 3217
rect 10152 3133 10182 3217
rect 10238 3133 10268 3217
rect 10324 3133 10354 3217
rect 10410 3133 10440 3217
rect 10495 3133 10525 3217
rect 10581 3133 10611 3217
rect 10667 3133 10697 3217
rect 10753 3133 10783 3217
rect 10839 3133 10869 3217
rect 10925 3133 10955 3217
rect 11011 3133 11041 3217
rect 11097 3133 11127 3217
rect 11763 3087 11793 3217
rect 11971 3133 12001 3217
rect 12062 3133 12092 3217
rect 12211 3133 12241 3217
rect 12307 3145 12337 3217
rect 12416 3145 12446 3217
rect 12515 3089 12545 3217
rect 12647 3133 12677 3217
rect 12719 3133 12749 3217
rect 12885 3145 12915 3217
rect 12981 3145 13011 3217
rect 13076 3133 13106 3217
rect 13331 3133 13361 3217
rect 13415 3133 13445 3217
rect 13603 3107 13813 3217
rect 13971 3133 14001 3217
rect 14066 3087 14096 3217
rect 14150 3087 14180 3217
rect 14339 3107 15285 3217
rect 15443 3107 16389 3217
rect 16731 3107 17677 3217
rect 17835 3107 18413 3217
rect 18663 3107 18781 3217
rect 1183 2223 1301 2333
rect 1459 2223 1577 2333
rect 1735 2223 1765 2307
rect 1819 2223 1849 2307
rect 2074 2223 2104 2307
rect 2169 2223 2199 2295
rect 2265 2223 2295 2295
rect 2431 2223 2461 2307
rect 2503 2223 2533 2307
rect 2635 2223 2665 2351
rect 2734 2223 2764 2295
rect 2843 2223 2873 2295
rect 2939 2223 2969 2307
rect 3088 2223 3118 2307
rect 3179 2223 3209 2307
rect 3387 2223 3417 2353
rect 3851 2223 4061 2333
rect 4311 2223 4341 2307
rect 4395 2223 4425 2307
rect 4650 2223 4680 2307
rect 4745 2223 4775 2295
rect 4841 2223 4871 2295
rect 5007 2223 5037 2307
rect 5079 2223 5109 2307
rect 5211 2223 5241 2351
rect 5310 2223 5340 2295
rect 5419 2223 5449 2295
rect 5515 2223 5545 2307
rect 5664 2223 5694 2307
rect 5755 2223 5785 2307
rect 5963 2223 5993 2353
rect 6427 2223 7373 2333
rect 7531 2223 8477 2333
rect 8635 2223 8753 2333
rect 9187 2223 9217 2353
rect 9395 2223 9425 2307
rect 9486 2223 9516 2307
rect 9635 2223 9665 2307
rect 9731 2223 9761 2295
rect 9840 2223 9870 2295
rect 9939 2223 9969 2351
rect 10071 2223 10101 2307
rect 10143 2223 10173 2307
rect 10309 2223 10339 2295
rect 10405 2223 10435 2295
rect 10500 2223 10530 2307
rect 10755 2223 10785 2307
rect 10839 2223 10869 2307
rect 11027 2223 11237 2333
rect 11579 2223 11789 2333
rect 12039 2223 12069 2353
rect 12247 2223 12277 2307
rect 12338 2223 12368 2307
rect 12487 2223 12517 2307
rect 12583 2223 12613 2295
rect 12692 2223 12722 2295
rect 12791 2223 12821 2351
rect 12923 2223 12953 2307
rect 12995 2223 13025 2307
rect 13161 2223 13191 2295
rect 13257 2223 13287 2295
rect 13352 2223 13382 2307
rect 13607 2223 13637 2307
rect 13691 2223 13721 2307
rect 14339 2223 14369 2353
rect 14547 2223 14577 2307
rect 14638 2223 14668 2307
rect 14787 2223 14817 2307
rect 14883 2223 14913 2295
rect 14992 2223 15022 2295
rect 15091 2223 15121 2351
rect 15223 2223 15253 2307
rect 15295 2223 15325 2307
rect 15461 2223 15491 2295
rect 15557 2223 15587 2295
rect 15652 2223 15682 2307
rect 15907 2223 15937 2307
rect 15991 2223 16021 2307
rect 16179 2223 16389 2333
rect 16731 2223 17309 2333
rect 17559 2223 17589 2307
rect 17654 2223 17684 2353
rect 17738 2223 17768 2353
rect 17927 2223 18505 2333
rect 18663 2223 18781 2333
<< scpmoshvt >>
rect 1183 7119 1301 7293
rect 1644 7119 1674 7319
rect 1728 7119 1758 7319
rect 1823 7127 1853 7255
rect 2011 7119 2957 7293
rect 3115 7119 3509 7293
rect 4036 7119 4066 7319
rect 4120 7119 4150 7319
rect 4215 7127 4245 7255
rect 4403 7119 5349 7293
rect 5692 7119 5722 7319
rect 5776 7119 5806 7319
rect 5871 7127 5901 7255
rect 6059 7119 6177 7293
rect 6427 7119 7373 7293
rect 7531 7119 7741 7293
rect 7900 7119 7930 7319
rect 7984 7119 8014 7319
rect 8079 7127 8109 7255
rect 8267 7119 8661 7293
rect 9003 7119 9397 7293
rect 9739 7119 9949 7293
rect 10108 7119 10138 7319
rect 10203 7119 10233 7319
rect 10287 7119 10317 7319
rect 10475 7119 11053 7293
rect 11211 7119 11329 7293
rect 11579 7119 12157 7293
rect 12315 7127 12345 7255
rect 12410 7119 12440 7319
rect 12494 7119 12524 7319
rect 12683 7119 13629 7293
rect 13787 7119 13905 7293
rect 14155 7119 14365 7293
rect 14523 7127 14553 7255
rect 14618 7119 14648 7319
rect 14702 7119 14732 7319
rect 14891 7119 15837 7293
rect 15995 7119 16389 7293
rect 16915 7127 16945 7255
rect 17010 7119 17040 7319
rect 17094 7119 17124 7319
rect 17283 7119 17861 7293
rect 18111 7127 18141 7255
rect 18206 7119 18236 7319
rect 18290 7119 18320 7319
rect 18663 7119 18781 7293
rect 1183 6851 1301 7025
rect 1459 6851 2405 7025
rect 2563 6851 3509 7025
rect 3851 6851 4797 7025
rect 4955 6851 5901 7025
rect 6059 6851 7005 7025
rect 7163 6851 8109 7025
rect 8267 6851 8661 7025
rect 9003 6851 9949 7025
rect 10107 6851 11053 7025
rect 11211 6851 12157 7025
rect 12315 6851 13261 7025
rect 13419 6851 13813 7025
rect 14155 6851 15101 7025
rect 15259 6851 16205 7025
rect 16363 6851 17309 7025
rect 17467 6851 18413 7025
rect 18663 6851 18781 7025
rect 1183 6031 1301 6205
rect 1459 6031 2405 6205
rect 2563 6031 3509 6205
rect 3667 6031 4613 6205
rect 4771 6031 5717 6205
rect 5875 6031 6085 6205
rect 6427 6031 7373 6205
rect 7531 6031 7925 6205
rect 8124 6147 8154 6231
rect 8196 6147 8226 6231
rect 8293 6031 8323 6231
rect 8543 6031 9489 6205
rect 9647 6031 10593 6205
rect 10751 6031 11329 6205
rect 11579 6031 12525 6205
rect 12683 6031 13629 6205
rect 13787 6031 14733 6205
rect 14891 6031 15837 6205
rect 15995 6031 16389 6205
rect 16731 6031 17677 6205
rect 17835 6031 18413 6205
rect 18663 6031 18781 6205
rect 1183 5763 1301 5937
rect 1459 5763 2405 5937
rect 2563 5763 3509 5937
rect 3851 5763 4797 5937
rect 4955 5763 5901 5937
rect 6059 5763 6637 5937
rect 6795 5779 6825 5937
rect 6883 5779 6913 5937
rect 7071 5763 7465 5937
rect 7669 5814 7699 5898
rect 7765 5814 7795 5898
rect 7837 5814 7867 5898
rect 8051 5814 8081 5898
rect 8154 5814 8184 5898
rect 8263 5737 8293 5937
rect 8451 5763 8661 5937
rect 9003 5763 9949 5937
rect 10107 5763 11053 5937
rect 11211 5763 11421 5937
rect 11620 5737 11650 5821
rect 11692 5737 11722 5821
rect 11789 5737 11819 5937
rect 12039 5763 12617 5937
rect 12908 5737 12938 5821
rect 12980 5737 13010 5821
rect 13077 5737 13107 5937
rect 13327 5763 13905 5937
rect 14155 5763 15101 5937
rect 15259 5763 16205 5937
rect 16363 5763 17309 5937
rect 17467 5763 18413 5937
rect 18663 5763 18781 5937
rect 1183 4943 1301 5117
rect 1459 4943 2405 5117
rect 2563 4943 2681 5117
rect 2839 4949 2869 5077
rect 2923 4949 2953 5077
rect 3190 4943 3220 5027
rect 3282 4943 3312 5027
rect 3381 4943 3411 5027
rect 3521 4943 3551 5027
rect 3618 4943 3648 5027
rect 3815 4943 3845 5111
rect 3914 4943 3944 5027
rect 4000 4943 4030 5027
rect 4084 4943 4114 5027
rect 4192 4943 4222 5027
rect 4276 4943 4306 5027
rect 4491 4943 4521 5143
rect 4679 4943 5625 5117
rect 5783 4943 6177 5117
rect 6427 4943 6545 5117
rect 6703 4943 6733 5143
rect 6812 4982 6842 5066
rect 6915 4982 6945 5066
rect 7129 4982 7159 5066
rect 7201 4982 7231 5066
rect 7297 4982 7327 5066
rect 7531 4943 7741 5117
rect 7899 4949 7929 5077
rect 7983 4949 8013 5077
rect 8250 4943 8280 5027
rect 8342 4943 8372 5027
rect 8441 4943 8471 5027
rect 8581 4943 8611 5027
rect 8678 4943 8708 5027
rect 8875 4943 8905 5111
rect 8974 4943 9004 5027
rect 9060 4943 9090 5027
rect 9144 4943 9174 5027
rect 9252 4943 9282 5027
rect 9336 4943 9366 5027
rect 9551 4943 9581 5143
rect 9739 4943 9949 5117
rect 10153 4982 10183 5066
rect 10249 4982 10279 5066
rect 10321 4982 10351 5066
rect 10535 4982 10565 5066
rect 10638 4982 10668 5066
rect 10747 4943 10777 5143
rect 10935 4943 11329 5117
rect 11763 4943 11793 5143
rect 11872 4982 11902 5066
rect 11975 4982 12005 5066
rect 12189 4982 12219 5066
rect 12261 4982 12291 5066
rect 12357 4982 12387 5066
rect 12591 4943 12801 5117
rect 13005 4982 13035 5066
rect 13101 4982 13131 5066
rect 13173 4982 13203 5066
rect 13387 4982 13417 5066
rect 13490 4982 13520 5066
rect 13599 4943 13629 5143
rect 13787 4943 14733 5117
rect 14891 4943 15837 5117
rect 15995 4943 16389 5117
rect 16731 4943 17677 5117
rect 17835 4943 18413 5117
rect 18663 4943 18781 5117
rect 1183 4675 1301 4849
rect 1459 4675 2037 4849
rect 2195 4675 2313 4849
rect 2490 4649 2520 4849
rect 2585 4765 2685 4849
rect 2843 4765 2943 4849
rect 2997 4765 3027 4849
rect 3207 4675 3601 4849
rect 4044 4649 4074 4849
rect 4130 4649 4160 4849
rect 4216 4649 4246 4849
rect 4302 4649 4332 4849
rect 4398 4649 4428 4849
rect 4587 4675 4797 4849
rect 5139 4675 5717 4849
rect 6121 4649 6151 4849
rect 6218 4649 6248 4733
rect 6290 4649 6320 4733
rect 6519 4675 6729 4849
rect 6928 4649 6958 4733
rect 7000 4649 7030 4733
rect 7097 4649 7127 4849
rect 7347 4675 7741 4849
rect 7899 4649 7929 4849
rect 8008 4726 8038 4810
rect 8111 4726 8141 4810
rect 8325 4726 8355 4810
rect 8397 4726 8427 4810
rect 8493 4726 8523 4810
rect 9228 4649 9258 4733
rect 9300 4649 9330 4733
rect 9397 4649 9427 4849
rect 9647 4675 9857 4849
rect 10199 4675 10409 4849
rect 10608 4649 10638 4733
rect 10680 4649 10710 4733
rect 10777 4649 10807 4849
rect 11027 4675 11237 4849
rect 11395 4691 11425 4849
rect 11483 4691 11513 4849
rect 11671 4675 11881 4849
rect 12085 4726 12115 4810
rect 12181 4726 12211 4810
rect 12253 4726 12283 4810
rect 12467 4726 12497 4810
rect 12570 4726 12600 4810
rect 12679 4649 12709 4849
rect 12867 4675 13077 4849
rect 13235 4691 13265 4849
rect 13323 4691 13353 4849
rect 13511 4675 13905 4849
rect 14155 4675 15101 4849
rect 15300 4649 15330 4733
rect 15372 4649 15402 4733
rect 15469 4649 15499 4849
rect 15719 4675 15929 4849
rect 16087 4691 16117 4849
rect 16175 4691 16205 4849
rect 16363 4675 16573 4849
rect 16731 4691 16761 4849
rect 16819 4691 16849 4849
rect 17007 4675 17953 4849
rect 18111 4675 18505 4849
rect 18663 4675 18781 4849
rect 1183 3855 1301 4029
rect 1459 3855 2037 4029
rect 2287 3855 2317 4013
rect 2375 3855 2405 4013
rect 2563 3855 2773 4029
rect 2931 3861 2961 3989
rect 3015 3861 3045 3989
rect 3282 3855 3312 3939
rect 3374 3855 3404 3939
rect 3473 3855 3503 3939
rect 3613 3855 3643 3939
rect 3710 3855 3740 3939
rect 3907 3855 3937 4023
rect 4006 3855 4036 3939
rect 4092 3855 4122 3939
rect 4176 3855 4206 3939
rect 4284 3855 4314 3939
rect 4368 3855 4398 3939
rect 4583 3855 4613 4055
rect 4771 3855 4981 4029
rect 5415 3855 5993 4029
rect 6427 3855 6545 4029
rect 6703 3855 6733 4013
rect 6791 3855 6821 4013
rect 6979 3855 7557 4029
rect 7761 3894 7791 3978
rect 7857 3894 7887 3978
rect 7929 3894 7959 3978
rect 8143 3894 8173 3978
rect 8246 3894 8276 3978
rect 8355 3855 8385 4055
rect 8543 3855 8753 4029
rect 9004 3855 9034 4055
rect 9090 3855 9120 4055
rect 9176 3855 9206 4055
rect 9262 3855 9292 4055
rect 9348 3855 9378 4055
rect 9434 3855 9464 4055
rect 9520 3855 9550 4055
rect 9606 3855 9636 4055
rect 9692 3855 9722 4055
rect 9778 3855 9808 4055
rect 9864 3855 9894 4055
rect 9950 3855 9980 4055
rect 10035 3855 10065 4055
rect 10121 3855 10151 4055
rect 10207 3855 10237 4055
rect 10293 3855 10323 4055
rect 10379 3855 10409 4055
rect 10465 3855 10495 4055
rect 10551 3855 10581 4055
rect 10637 3855 10667 4055
rect 10843 3855 11237 4029
rect 11763 3855 11793 4055
rect 11978 3855 12008 3939
rect 12062 3855 12092 3939
rect 12170 3855 12200 3939
rect 12254 3855 12284 3939
rect 12340 3855 12370 3939
rect 12439 3855 12469 4023
rect 12636 3855 12666 3939
rect 12733 3855 12763 3939
rect 12873 3855 12903 3939
rect 12972 3855 13002 3939
rect 13064 3855 13094 3939
rect 13331 3861 13361 3989
rect 13415 3861 13445 3989
rect 13603 3855 13813 4029
rect 13971 3861 14001 3989
rect 14055 3861 14085 3989
rect 14322 3855 14352 3939
rect 14414 3855 14444 3939
rect 14513 3855 14543 3939
rect 14653 3855 14683 3939
rect 14750 3855 14780 3939
rect 14947 3855 14977 4023
rect 15046 3855 15076 3939
rect 15132 3855 15162 3939
rect 15216 3855 15246 3939
rect 15324 3855 15354 3939
rect 15408 3855 15438 3939
rect 15623 3855 15653 4055
rect 15811 3855 16389 4029
rect 16731 3855 17677 4029
rect 17835 3855 18413 4029
rect 18663 3855 18781 4029
rect 1183 3587 1301 3761
rect 1459 3587 1577 3761
rect 1735 3627 1765 3755
rect 1819 3627 1849 3755
rect 2086 3677 2116 3761
rect 2178 3677 2208 3761
rect 2277 3677 2307 3761
rect 2417 3677 2447 3761
rect 2514 3677 2544 3761
rect 2711 3593 2741 3761
rect 2810 3677 2840 3761
rect 2896 3677 2926 3761
rect 2980 3677 3010 3761
rect 3088 3677 3118 3761
rect 3172 3677 3202 3761
rect 3387 3561 3417 3761
rect 3851 3587 4429 3761
rect 4605 3561 4635 3761
rect 4691 3561 4721 3761
rect 4777 3561 4807 3761
rect 4863 3561 4893 3761
rect 4949 3561 4979 3761
rect 5035 3561 5065 3761
rect 5121 3561 5151 3761
rect 5207 3561 5237 3761
rect 5292 3561 5322 3761
rect 5378 3561 5408 3761
rect 5464 3561 5494 3761
rect 5550 3561 5580 3761
rect 5636 3561 5666 3761
rect 5722 3561 5752 3761
rect 5808 3561 5838 3761
rect 5894 3561 5924 3761
rect 5980 3561 6010 3761
rect 6066 3561 6096 3761
rect 6152 3561 6182 3761
rect 6238 3561 6268 3761
rect 6427 3587 6637 3761
rect 6795 3627 6825 3755
rect 6879 3627 6909 3755
rect 7146 3677 7176 3761
rect 7238 3677 7268 3761
rect 7337 3677 7367 3761
rect 7477 3677 7507 3761
rect 7574 3677 7604 3761
rect 7771 3593 7801 3761
rect 7870 3677 7900 3761
rect 7956 3677 7986 3761
rect 8040 3677 8070 3761
rect 8148 3677 8178 3761
rect 8232 3677 8262 3761
rect 8447 3561 8477 3761
rect 8635 3587 8753 3761
rect 9187 3625 9217 3753
rect 9282 3561 9312 3761
rect 9366 3561 9396 3761
rect 9555 3587 9949 3761
rect 10107 3603 10137 3761
rect 10195 3603 10225 3761
rect 10383 3587 10777 3761
rect 11027 3603 11057 3761
rect 11115 3603 11145 3761
rect 11303 3587 11881 3761
rect 12039 3561 12069 3761
rect 12254 3677 12284 3761
rect 12338 3677 12368 3761
rect 12446 3677 12476 3761
rect 12530 3677 12560 3761
rect 12616 3677 12646 3761
rect 12715 3593 12745 3761
rect 12912 3677 12942 3761
rect 13009 3677 13039 3761
rect 13149 3677 13179 3761
rect 13248 3677 13278 3761
rect 13340 3677 13370 3761
rect 13607 3627 13637 3755
rect 13691 3627 13721 3755
rect 14155 3587 15101 3761
rect 15259 3587 16205 3761
rect 16363 3587 17309 3761
rect 17467 3587 18413 3761
rect 18663 3587 18781 3761
rect 1183 2767 1301 2941
rect 1459 2767 1853 2941
rect 2011 2767 2041 2967
rect 2226 2767 2256 2851
rect 2310 2767 2340 2851
rect 2418 2767 2448 2851
rect 2502 2767 2532 2851
rect 2588 2767 2618 2851
rect 2687 2767 2717 2935
rect 2884 2767 2914 2851
rect 2981 2767 3011 2851
rect 3121 2767 3151 2851
rect 3220 2767 3250 2851
rect 3312 2767 3342 2851
rect 3579 2773 3609 2901
rect 3663 2773 3693 2901
rect 3851 2767 4061 2941
rect 4219 2773 4249 2901
rect 4303 2773 4333 2901
rect 4491 2767 4521 2935
rect 4588 2767 4618 2851
rect 4672 2767 4702 2851
rect 4792 2767 4822 2851
rect 4898 2767 4928 2851
rect 4982 2767 5012 2851
rect 5066 2767 5096 2851
rect 5142 2767 5172 2851
rect 5250 2767 5280 2851
rect 5322 2767 5352 2851
rect 5510 2767 5540 2851
rect 5606 2767 5636 2935
rect 5794 2767 5824 2895
rect 5889 2767 5919 2967
rect 6427 2767 7005 2941
rect 7255 2767 7285 2967
rect 7470 2767 7500 2851
rect 7554 2767 7584 2851
rect 7662 2767 7692 2851
rect 7746 2767 7776 2851
rect 7832 2767 7862 2851
rect 7931 2767 7961 2935
rect 8128 2767 8158 2851
rect 8225 2767 8255 2851
rect 8365 2767 8395 2851
rect 8464 2767 8494 2851
rect 8556 2767 8586 2851
rect 8823 2773 8853 2901
rect 8907 2773 8937 2901
rect 9095 2767 9305 2941
rect 9464 2767 9494 2967
rect 9550 2767 9580 2967
rect 9636 2767 9666 2967
rect 9722 2767 9752 2967
rect 9808 2767 9838 2967
rect 9894 2767 9924 2967
rect 9980 2767 10010 2967
rect 10066 2767 10096 2967
rect 10152 2767 10182 2967
rect 10238 2767 10268 2967
rect 10324 2767 10354 2967
rect 10410 2767 10440 2967
rect 10495 2767 10525 2967
rect 10581 2767 10611 2967
rect 10667 2767 10697 2967
rect 10753 2767 10783 2967
rect 10839 2767 10869 2967
rect 10925 2767 10955 2967
rect 11011 2767 11041 2967
rect 11097 2767 11127 2967
rect 11763 2767 11793 2967
rect 11978 2767 12008 2851
rect 12062 2767 12092 2851
rect 12170 2767 12200 2851
rect 12254 2767 12284 2851
rect 12340 2767 12370 2851
rect 12439 2767 12469 2935
rect 12636 2767 12666 2851
rect 12733 2767 12763 2851
rect 12873 2767 12903 2851
rect 12972 2767 13002 2851
rect 13064 2767 13094 2851
rect 13331 2773 13361 2901
rect 13415 2773 13445 2901
rect 13603 2767 13813 2941
rect 13971 2775 14001 2903
rect 14066 2767 14096 2967
rect 14150 2767 14180 2967
rect 14339 2767 15285 2941
rect 15443 2767 16389 2941
rect 16731 2767 17677 2941
rect 17835 2767 18413 2941
rect 18663 2767 18781 2941
rect 1183 2499 1301 2673
rect 1459 2499 1577 2673
rect 1735 2539 1765 2667
rect 1819 2539 1849 2667
rect 2086 2589 2116 2673
rect 2178 2589 2208 2673
rect 2277 2589 2307 2673
rect 2417 2589 2447 2673
rect 2514 2589 2544 2673
rect 2711 2505 2741 2673
rect 2810 2589 2840 2673
rect 2896 2589 2926 2673
rect 2980 2589 3010 2673
rect 3088 2589 3118 2673
rect 3172 2589 3202 2673
rect 3387 2473 3417 2673
rect 3851 2499 4061 2673
rect 4311 2539 4341 2667
rect 4395 2539 4425 2667
rect 4662 2589 4692 2673
rect 4754 2589 4784 2673
rect 4853 2589 4883 2673
rect 4993 2589 5023 2673
rect 5090 2589 5120 2673
rect 5287 2505 5317 2673
rect 5386 2589 5416 2673
rect 5472 2589 5502 2673
rect 5556 2589 5586 2673
rect 5664 2589 5694 2673
rect 5748 2589 5778 2673
rect 5963 2473 5993 2673
rect 6427 2499 7373 2673
rect 7531 2499 8477 2673
rect 8635 2499 8753 2673
rect 9187 2473 9217 2673
rect 9402 2589 9432 2673
rect 9486 2589 9516 2673
rect 9594 2589 9624 2673
rect 9678 2589 9708 2673
rect 9764 2589 9794 2673
rect 9863 2505 9893 2673
rect 10060 2589 10090 2673
rect 10157 2589 10187 2673
rect 10297 2589 10327 2673
rect 10396 2589 10426 2673
rect 10488 2589 10518 2673
rect 10755 2539 10785 2667
rect 10839 2539 10869 2667
rect 11027 2499 11237 2673
rect 11579 2499 11789 2673
rect 12039 2473 12069 2673
rect 12254 2589 12284 2673
rect 12338 2589 12368 2673
rect 12446 2589 12476 2673
rect 12530 2589 12560 2673
rect 12616 2589 12646 2673
rect 12715 2505 12745 2673
rect 12912 2589 12942 2673
rect 13009 2589 13039 2673
rect 13149 2589 13179 2673
rect 13248 2589 13278 2673
rect 13340 2589 13370 2673
rect 13607 2539 13637 2667
rect 13691 2539 13721 2667
rect 14339 2473 14369 2673
rect 14554 2589 14584 2673
rect 14638 2589 14668 2673
rect 14746 2589 14776 2673
rect 14830 2589 14860 2673
rect 14916 2589 14946 2673
rect 15015 2505 15045 2673
rect 15212 2589 15242 2673
rect 15309 2589 15339 2673
rect 15449 2589 15479 2673
rect 15548 2589 15578 2673
rect 15640 2589 15670 2673
rect 15907 2539 15937 2667
rect 15991 2539 16021 2667
rect 16179 2499 16389 2673
rect 16731 2499 17309 2673
rect 17559 2537 17589 2665
rect 17654 2473 17684 2673
rect 17738 2473 17768 2673
rect 17927 2499 18505 2673
rect 18663 2499 18781 2673
<< ndiff >>
rect 1131 7536 1183 7569
rect 1131 7502 1139 7536
rect 1173 7502 1183 7536
rect 1131 7459 1183 7502
rect 1301 7536 1353 7569
rect 1301 7502 1311 7536
rect 1345 7502 1353 7536
rect 1301 7459 1353 7502
rect 1591 7553 1644 7569
rect 1591 7519 1600 7553
rect 1634 7519 1644 7553
rect 1591 7485 1644 7519
rect 1591 7451 1600 7485
rect 1634 7451 1644 7485
rect 1591 7439 1644 7451
rect 1674 7527 1728 7569
rect 1674 7493 1684 7527
rect 1718 7493 1728 7527
rect 1674 7439 1728 7493
rect 1758 7557 1823 7569
rect 1758 7523 1770 7557
rect 1804 7523 1823 7557
rect 1758 7485 1823 7523
rect 1853 7544 1905 7569
rect 1853 7510 1863 7544
rect 1897 7510 1905 7544
rect 1853 7485 1905 7510
rect 1959 7538 2011 7569
rect 1959 7504 1967 7538
rect 2001 7504 2011 7538
rect 1758 7439 1808 7485
rect 1959 7459 2011 7504
rect 2957 7538 3009 7569
rect 2957 7504 2967 7538
rect 3001 7504 3009 7538
rect 2957 7459 3009 7504
rect 3063 7538 3115 7569
rect 3063 7504 3071 7538
rect 3105 7504 3115 7538
rect 3063 7459 3115 7504
rect 3509 7538 3561 7569
rect 3983 7553 4036 7569
rect 3509 7504 3519 7538
rect 3553 7504 3561 7538
rect 3509 7459 3561 7504
rect 3983 7519 3992 7553
rect 4026 7519 4036 7553
rect 3983 7485 4036 7519
rect 3983 7451 3992 7485
rect 4026 7451 4036 7485
rect 3983 7439 4036 7451
rect 4066 7527 4120 7569
rect 4066 7493 4076 7527
rect 4110 7493 4120 7527
rect 4066 7439 4120 7493
rect 4150 7557 4215 7569
rect 4150 7523 4162 7557
rect 4196 7523 4215 7557
rect 4150 7485 4215 7523
rect 4245 7544 4297 7569
rect 4245 7510 4255 7544
rect 4289 7510 4297 7544
rect 4245 7485 4297 7510
rect 4351 7538 4403 7569
rect 4351 7504 4359 7538
rect 4393 7504 4403 7538
rect 4150 7439 4200 7485
rect 4351 7459 4403 7504
rect 5349 7538 5401 7569
rect 5349 7504 5359 7538
rect 5393 7504 5401 7538
rect 5349 7459 5401 7504
rect 5639 7553 5692 7569
rect 5639 7519 5648 7553
rect 5682 7519 5692 7553
rect 5639 7485 5692 7519
rect 5639 7451 5648 7485
rect 5682 7451 5692 7485
rect 5639 7439 5692 7451
rect 5722 7527 5776 7569
rect 5722 7493 5732 7527
rect 5766 7493 5776 7527
rect 5722 7439 5776 7493
rect 5806 7557 5871 7569
rect 5806 7523 5818 7557
rect 5852 7523 5871 7557
rect 5806 7485 5871 7523
rect 5901 7544 5953 7569
rect 5901 7510 5911 7544
rect 5945 7510 5953 7544
rect 5901 7485 5953 7510
rect 6007 7536 6059 7569
rect 6007 7502 6015 7536
rect 6049 7502 6059 7536
rect 5806 7439 5856 7485
rect 6007 7459 6059 7502
rect 6177 7536 6229 7569
rect 6177 7502 6187 7536
rect 6221 7502 6229 7536
rect 6177 7459 6229 7502
rect 6375 7538 6427 7569
rect 6375 7504 6383 7538
rect 6417 7504 6427 7538
rect 6375 7459 6427 7504
rect 7373 7538 7425 7569
rect 7373 7504 7383 7538
rect 7417 7504 7425 7538
rect 7373 7459 7425 7504
rect 7479 7531 7531 7569
rect 7479 7497 7487 7531
rect 7521 7497 7531 7531
rect 7479 7459 7531 7497
rect 7741 7531 7793 7569
rect 7741 7497 7751 7531
rect 7785 7497 7793 7531
rect 7741 7459 7793 7497
rect 7847 7553 7900 7569
rect 7847 7519 7856 7553
rect 7890 7519 7900 7553
rect 7847 7485 7900 7519
rect 7847 7451 7856 7485
rect 7890 7451 7900 7485
rect 7847 7439 7900 7451
rect 7930 7527 7984 7569
rect 7930 7493 7940 7527
rect 7974 7493 7984 7527
rect 7930 7439 7984 7493
rect 8014 7557 8079 7569
rect 8014 7523 8026 7557
rect 8060 7523 8079 7557
rect 8014 7485 8079 7523
rect 8109 7544 8161 7569
rect 8109 7510 8119 7544
rect 8153 7510 8161 7544
rect 8109 7485 8161 7510
rect 8215 7538 8267 7569
rect 8215 7504 8223 7538
rect 8257 7504 8267 7538
rect 8014 7439 8064 7485
rect 8215 7459 8267 7504
rect 8661 7538 8713 7569
rect 8661 7504 8671 7538
rect 8705 7504 8713 7538
rect 8661 7459 8713 7504
rect 8951 7538 9003 7569
rect 8951 7504 8959 7538
rect 8993 7504 9003 7538
rect 8951 7459 9003 7504
rect 9397 7538 9449 7569
rect 9397 7504 9407 7538
rect 9441 7504 9449 7538
rect 9397 7459 9449 7504
rect 9687 7531 9739 7569
rect 9687 7497 9695 7531
rect 9729 7497 9739 7531
rect 9687 7459 9739 7497
rect 9949 7531 10001 7569
rect 9949 7497 9959 7531
rect 9993 7497 10001 7531
rect 9949 7459 10001 7497
rect 10055 7549 10108 7569
rect 10055 7515 10063 7549
rect 10097 7515 10108 7549
rect 10055 7485 10108 7515
rect 10138 7553 10203 7569
rect 10138 7519 10149 7553
rect 10183 7519 10203 7553
rect 10138 7485 10203 7519
rect 10233 7549 10287 7569
rect 10233 7515 10243 7549
rect 10277 7515 10287 7549
rect 10233 7485 10287 7515
rect 10317 7553 10369 7569
rect 10317 7519 10327 7553
rect 10361 7519 10369 7553
rect 10317 7485 10369 7519
rect 10423 7538 10475 7569
rect 10423 7504 10431 7538
rect 10465 7504 10475 7538
rect 10423 7459 10475 7504
rect 11053 7538 11105 7569
rect 11053 7504 11063 7538
rect 11097 7504 11105 7538
rect 11053 7459 11105 7504
rect 11159 7536 11211 7569
rect 11159 7502 11167 7536
rect 11201 7502 11211 7536
rect 11159 7459 11211 7502
rect 11329 7536 11381 7569
rect 11329 7502 11339 7536
rect 11373 7502 11381 7536
rect 11329 7459 11381 7502
rect 11527 7538 11579 7569
rect 11527 7504 11535 7538
rect 11569 7504 11579 7538
rect 11527 7459 11579 7504
rect 12157 7538 12209 7569
rect 12157 7504 12167 7538
rect 12201 7504 12209 7538
rect 12157 7459 12209 7504
rect 12263 7544 12315 7569
rect 12263 7510 12271 7544
rect 12305 7510 12315 7544
rect 12263 7485 12315 7510
rect 12345 7557 12410 7569
rect 12345 7523 12364 7557
rect 12398 7523 12410 7557
rect 12345 7485 12410 7523
rect 12360 7439 12410 7485
rect 12440 7527 12494 7569
rect 12440 7493 12450 7527
rect 12484 7493 12494 7527
rect 12440 7439 12494 7493
rect 12524 7553 12577 7569
rect 12524 7519 12534 7553
rect 12568 7519 12577 7553
rect 12524 7485 12577 7519
rect 12524 7451 12534 7485
rect 12568 7451 12577 7485
rect 12631 7538 12683 7569
rect 12631 7504 12639 7538
rect 12673 7504 12683 7538
rect 12631 7459 12683 7504
rect 13629 7538 13681 7569
rect 13629 7504 13639 7538
rect 13673 7504 13681 7538
rect 13629 7459 13681 7504
rect 13735 7536 13787 7569
rect 13735 7502 13743 7536
rect 13777 7502 13787 7536
rect 13735 7459 13787 7502
rect 13905 7536 13957 7569
rect 13905 7502 13915 7536
rect 13949 7502 13957 7536
rect 13905 7459 13957 7502
rect 12524 7439 12577 7451
rect 14103 7531 14155 7569
rect 14103 7497 14111 7531
rect 14145 7497 14155 7531
rect 14103 7459 14155 7497
rect 14365 7531 14417 7569
rect 14365 7497 14375 7531
rect 14409 7497 14417 7531
rect 14365 7459 14417 7497
rect 14471 7544 14523 7569
rect 14471 7510 14479 7544
rect 14513 7510 14523 7544
rect 14471 7485 14523 7510
rect 14553 7557 14618 7569
rect 14553 7523 14572 7557
rect 14606 7523 14618 7557
rect 14553 7485 14618 7523
rect 14568 7439 14618 7485
rect 14648 7527 14702 7569
rect 14648 7493 14658 7527
rect 14692 7493 14702 7527
rect 14648 7439 14702 7493
rect 14732 7553 14785 7569
rect 14732 7519 14742 7553
rect 14776 7519 14785 7553
rect 14732 7485 14785 7519
rect 14732 7451 14742 7485
rect 14776 7451 14785 7485
rect 14839 7538 14891 7569
rect 14839 7504 14847 7538
rect 14881 7504 14891 7538
rect 14839 7459 14891 7504
rect 15837 7538 15889 7569
rect 15837 7504 15847 7538
rect 15881 7504 15889 7538
rect 15837 7459 15889 7504
rect 15943 7538 15995 7569
rect 15943 7504 15951 7538
rect 15985 7504 15995 7538
rect 15943 7459 15995 7504
rect 16389 7538 16441 7569
rect 16389 7504 16399 7538
rect 16433 7504 16441 7538
rect 16389 7459 16441 7504
rect 16863 7544 16915 7569
rect 16863 7510 16871 7544
rect 16905 7510 16915 7544
rect 16863 7485 16915 7510
rect 16945 7557 17010 7569
rect 16945 7523 16964 7557
rect 16998 7523 17010 7557
rect 16945 7485 17010 7523
rect 14732 7439 14785 7451
rect 16960 7439 17010 7485
rect 17040 7527 17094 7569
rect 17040 7493 17050 7527
rect 17084 7493 17094 7527
rect 17040 7439 17094 7493
rect 17124 7553 17177 7569
rect 17124 7519 17134 7553
rect 17168 7519 17177 7553
rect 17124 7485 17177 7519
rect 17124 7451 17134 7485
rect 17168 7451 17177 7485
rect 17231 7538 17283 7569
rect 17231 7504 17239 7538
rect 17273 7504 17283 7538
rect 17231 7459 17283 7504
rect 17861 7538 17913 7569
rect 17861 7504 17871 7538
rect 17905 7504 17913 7538
rect 17861 7459 17913 7504
rect 18059 7544 18111 7569
rect 18059 7510 18067 7544
rect 18101 7510 18111 7544
rect 18059 7485 18111 7510
rect 18141 7557 18206 7569
rect 18141 7523 18160 7557
rect 18194 7523 18206 7557
rect 18141 7485 18206 7523
rect 17124 7439 17177 7451
rect 18156 7439 18206 7485
rect 18236 7527 18290 7569
rect 18236 7493 18246 7527
rect 18280 7493 18290 7527
rect 18236 7439 18290 7493
rect 18320 7553 18373 7569
rect 18320 7519 18330 7553
rect 18364 7519 18373 7553
rect 18320 7485 18373 7519
rect 18320 7451 18330 7485
rect 18364 7451 18373 7485
rect 18611 7536 18663 7569
rect 18611 7502 18619 7536
rect 18653 7502 18663 7536
rect 18611 7459 18663 7502
rect 18781 7536 18833 7569
rect 18781 7502 18791 7536
rect 18825 7502 18833 7536
rect 18781 7459 18833 7502
rect 18320 7439 18373 7451
rect 1131 6642 1183 6685
rect 1131 6608 1139 6642
rect 1173 6608 1183 6642
rect 1131 6575 1183 6608
rect 1301 6642 1353 6685
rect 1301 6608 1311 6642
rect 1345 6608 1353 6642
rect 1301 6575 1353 6608
rect 1407 6640 1459 6685
rect 1407 6606 1415 6640
rect 1449 6606 1459 6640
rect 1407 6575 1459 6606
rect 2405 6640 2457 6685
rect 2405 6606 2415 6640
rect 2449 6606 2457 6640
rect 2405 6575 2457 6606
rect 2511 6640 2563 6685
rect 2511 6606 2519 6640
rect 2553 6606 2563 6640
rect 2511 6575 2563 6606
rect 3509 6640 3561 6685
rect 3509 6606 3519 6640
rect 3553 6606 3561 6640
rect 3509 6575 3561 6606
rect 3799 6640 3851 6685
rect 3799 6606 3807 6640
rect 3841 6606 3851 6640
rect 3799 6575 3851 6606
rect 4797 6640 4849 6685
rect 4797 6606 4807 6640
rect 4841 6606 4849 6640
rect 4797 6575 4849 6606
rect 4903 6640 4955 6685
rect 4903 6606 4911 6640
rect 4945 6606 4955 6640
rect 4903 6575 4955 6606
rect 5901 6640 5953 6685
rect 5901 6606 5911 6640
rect 5945 6606 5953 6640
rect 5901 6575 5953 6606
rect 6007 6640 6059 6685
rect 6007 6606 6015 6640
rect 6049 6606 6059 6640
rect 6007 6575 6059 6606
rect 7005 6640 7057 6685
rect 7005 6606 7015 6640
rect 7049 6606 7057 6640
rect 7005 6575 7057 6606
rect 7111 6640 7163 6685
rect 7111 6606 7119 6640
rect 7153 6606 7163 6640
rect 7111 6575 7163 6606
rect 8109 6640 8161 6685
rect 8109 6606 8119 6640
rect 8153 6606 8161 6640
rect 8109 6575 8161 6606
rect 8215 6640 8267 6685
rect 8215 6606 8223 6640
rect 8257 6606 8267 6640
rect 8215 6575 8267 6606
rect 8661 6640 8713 6685
rect 8661 6606 8671 6640
rect 8705 6606 8713 6640
rect 8661 6575 8713 6606
rect 8951 6640 9003 6685
rect 8951 6606 8959 6640
rect 8993 6606 9003 6640
rect 8951 6575 9003 6606
rect 9949 6640 10001 6685
rect 9949 6606 9959 6640
rect 9993 6606 10001 6640
rect 9949 6575 10001 6606
rect 10055 6640 10107 6685
rect 10055 6606 10063 6640
rect 10097 6606 10107 6640
rect 10055 6575 10107 6606
rect 11053 6640 11105 6685
rect 11053 6606 11063 6640
rect 11097 6606 11105 6640
rect 11053 6575 11105 6606
rect 11159 6640 11211 6685
rect 11159 6606 11167 6640
rect 11201 6606 11211 6640
rect 11159 6575 11211 6606
rect 12157 6640 12209 6685
rect 12157 6606 12167 6640
rect 12201 6606 12209 6640
rect 12157 6575 12209 6606
rect 12263 6640 12315 6685
rect 12263 6606 12271 6640
rect 12305 6606 12315 6640
rect 12263 6575 12315 6606
rect 13261 6640 13313 6685
rect 13261 6606 13271 6640
rect 13305 6606 13313 6640
rect 13261 6575 13313 6606
rect 13367 6640 13419 6685
rect 13367 6606 13375 6640
rect 13409 6606 13419 6640
rect 13367 6575 13419 6606
rect 13813 6640 13865 6685
rect 13813 6606 13823 6640
rect 13857 6606 13865 6640
rect 13813 6575 13865 6606
rect 14103 6640 14155 6685
rect 14103 6606 14111 6640
rect 14145 6606 14155 6640
rect 14103 6575 14155 6606
rect 15101 6640 15153 6685
rect 15101 6606 15111 6640
rect 15145 6606 15153 6640
rect 15101 6575 15153 6606
rect 15207 6640 15259 6685
rect 15207 6606 15215 6640
rect 15249 6606 15259 6640
rect 15207 6575 15259 6606
rect 16205 6640 16257 6685
rect 16205 6606 16215 6640
rect 16249 6606 16257 6640
rect 16205 6575 16257 6606
rect 16311 6640 16363 6685
rect 16311 6606 16319 6640
rect 16353 6606 16363 6640
rect 16311 6575 16363 6606
rect 17309 6640 17361 6685
rect 17309 6606 17319 6640
rect 17353 6606 17361 6640
rect 17309 6575 17361 6606
rect 17415 6640 17467 6685
rect 17415 6606 17423 6640
rect 17457 6606 17467 6640
rect 17415 6575 17467 6606
rect 18413 6640 18465 6685
rect 18413 6606 18423 6640
rect 18457 6606 18465 6640
rect 18413 6575 18465 6606
rect 18611 6642 18663 6685
rect 18611 6608 18619 6642
rect 18653 6608 18663 6642
rect 18611 6575 18663 6608
rect 18781 6642 18833 6685
rect 18781 6608 18791 6642
rect 18825 6608 18833 6642
rect 18781 6575 18833 6608
rect 1131 6448 1183 6481
rect 1131 6414 1139 6448
rect 1173 6414 1183 6448
rect 1131 6371 1183 6414
rect 1301 6448 1353 6481
rect 1301 6414 1311 6448
rect 1345 6414 1353 6448
rect 1301 6371 1353 6414
rect 1407 6450 1459 6481
rect 1407 6416 1415 6450
rect 1449 6416 1459 6450
rect 1407 6371 1459 6416
rect 2405 6450 2457 6481
rect 2405 6416 2415 6450
rect 2449 6416 2457 6450
rect 2405 6371 2457 6416
rect 2511 6450 2563 6481
rect 2511 6416 2519 6450
rect 2553 6416 2563 6450
rect 2511 6371 2563 6416
rect 3509 6450 3561 6481
rect 3509 6416 3519 6450
rect 3553 6416 3561 6450
rect 3509 6371 3561 6416
rect 3615 6450 3667 6481
rect 3615 6416 3623 6450
rect 3657 6416 3667 6450
rect 3615 6371 3667 6416
rect 4613 6450 4665 6481
rect 4613 6416 4623 6450
rect 4657 6416 4665 6450
rect 4613 6371 4665 6416
rect 4719 6450 4771 6481
rect 4719 6416 4727 6450
rect 4761 6416 4771 6450
rect 4719 6371 4771 6416
rect 5717 6450 5769 6481
rect 5717 6416 5727 6450
rect 5761 6416 5769 6450
rect 5717 6371 5769 6416
rect 5823 6443 5875 6481
rect 5823 6409 5831 6443
rect 5865 6409 5875 6443
rect 5823 6371 5875 6409
rect 6085 6443 6137 6481
rect 6085 6409 6095 6443
rect 6129 6409 6137 6443
rect 6085 6371 6137 6409
rect 6375 6450 6427 6481
rect 6375 6416 6383 6450
rect 6417 6416 6427 6450
rect 6375 6371 6427 6416
rect 7373 6450 7425 6481
rect 7373 6416 7383 6450
rect 7417 6416 7425 6450
rect 7373 6371 7425 6416
rect 7479 6450 7531 6481
rect 7479 6416 7487 6450
rect 7521 6416 7531 6450
rect 7479 6371 7531 6416
rect 7925 6450 7977 6481
rect 7925 6416 7935 6450
rect 7969 6416 7977 6450
rect 7925 6371 7977 6416
rect 8060 6459 8112 6481
rect 8060 6425 8068 6459
rect 8102 6425 8112 6459
rect 8060 6397 8112 6425
rect 8142 6459 8196 6481
rect 8142 6425 8152 6459
rect 8186 6425 8196 6459
rect 8142 6397 8196 6425
rect 8226 6459 8293 6481
rect 8226 6425 8248 6459
rect 8282 6425 8293 6459
rect 8226 6397 8293 6425
rect 8241 6351 8293 6397
rect 8323 6467 8375 6481
rect 8323 6433 8333 6467
rect 8367 6433 8375 6467
rect 8323 6399 8375 6433
rect 8323 6365 8333 6399
rect 8367 6365 8375 6399
rect 8491 6450 8543 6481
rect 8491 6416 8499 6450
rect 8533 6416 8543 6450
rect 8491 6371 8543 6416
rect 9489 6450 9541 6481
rect 9489 6416 9499 6450
rect 9533 6416 9541 6450
rect 9489 6371 9541 6416
rect 9595 6450 9647 6481
rect 9595 6416 9603 6450
rect 9637 6416 9647 6450
rect 9595 6371 9647 6416
rect 10593 6450 10645 6481
rect 10593 6416 10603 6450
rect 10637 6416 10645 6450
rect 10593 6371 10645 6416
rect 10699 6450 10751 6481
rect 10699 6416 10707 6450
rect 10741 6416 10751 6450
rect 10699 6371 10751 6416
rect 11329 6450 11381 6481
rect 11329 6416 11339 6450
rect 11373 6416 11381 6450
rect 11329 6371 11381 6416
rect 8323 6351 8375 6365
rect 11527 6450 11579 6481
rect 11527 6416 11535 6450
rect 11569 6416 11579 6450
rect 11527 6371 11579 6416
rect 12525 6450 12577 6481
rect 12525 6416 12535 6450
rect 12569 6416 12577 6450
rect 12525 6371 12577 6416
rect 12631 6450 12683 6481
rect 12631 6416 12639 6450
rect 12673 6416 12683 6450
rect 12631 6371 12683 6416
rect 13629 6450 13681 6481
rect 13629 6416 13639 6450
rect 13673 6416 13681 6450
rect 13629 6371 13681 6416
rect 13735 6450 13787 6481
rect 13735 6416 13743 6450
rect 13777 6416 13787 6450
rect 13735 6371 13787 6416
rect 14733 6450 14785 6481
rect 14733 6416 14743 6450
rect 14777 6416 14785 6450
rect 14733 6371 14785 6416
rect 14839 6450 14891 6481
rect 14839 6416 14847 6450
rect 14881 6416 14891 6450
rect 14839 6371 14891 6416
rect 15837 6450 15889 6481
rect 15837 6416 15847 6450
rect 15881 6416 15889 6450
rect 15837 6371 15889 6416
rect 15943 6450 15995 6481
rect 15943 6416 15951 6450
rect 15985 6416 15995 6450
rect 15943 6371 15995 6416
rect 16389 6450 16441 6481
rect 16389 6416 16399 6450
rect 16433 6416 16441 6450
rect 16389 6371 16441 6416
rect 16679 6450 16731 6481
rect 16679 6416 16687 6450
rect 16721 6416 16731 6450
rect 16679 6371 16731 6416
rect 17677 6450 17729 6481
rect 17677 6416 17687 6450
rect 17721 6416 17729 6450
rect 17677 6371 17729 6416
rect 17783 6450 17835 6481
rect 17783 6416 17791 6450
rect 17825 6416 17835 6450
rect 17783 6371 17835 6416
rect 18413 6450 18465 6481
rect 18413 6416 18423 6450
rect 18457 6416 18465 6450
rect 18413 6371 18465 6416
rect 18611 6448 18663 6481
rect 18611 6414 18619 6448
rect 18653 6414 18663 6448
rect 18611 6371 18663 6414
rect 18781 6448 18833 6481
rect 18781 6414 18791 6448
rect 18825 6414 18833 6448
rect 18781 6371 18833 6414
rect 1131 5554 1183 5597
rect 1131 5520 1139 5554
rect 1173 5520 1183 5554
rect 1131 5487 1183 5520
rect 1301 5554 1353 5597
rect 1301 5520 1311 5554
rect 1345 5520 1353 5554
rect 1301 5487 1353 5520
rect 1407 5552 1459 5597
rect 1407 5518 1415 5552
rect 1449 5518 1459 5552
rect 1407 5487 1459 5518
rect 2405 5552 2457 5597
rect 2405 5518 2415 5552
rect 2449 5518 2457 5552
rect 2405 5487 2457 5518
rect 2511 5552 2563 5597
rect 2511 5518 2519 5552
rect 2553 5518 2563 5552
rect 2511 5487 2563 5518
rect 3509 5552 3561 5597
rect 3509 5518 3519 5552
rect 3553 5518 3561 5552
rect 3509 5487 3561 5518
rect 3799 5552 3851 5597
rect 3799 5518 3807 5552
rect 3841 5518 3851 5552
rect 3799 5487 3851 5518
rect 4797 5552 4849 5597
rect 4797 5518 4807 5552
rect 4841 5518 4849 5552
rect 4797 5487 4849 5518
rect 4903 5552 4955 5597
rect 4903 5518 4911 5552
rect 4945 5518 4955 5552
rect 4903 5487 4955 5518
rect 5901 5552 5953 5597
rect 5901 5518 5911 5552
rect 5945 5518 5953 5552
rect 5901 5487 5953 5518
rect 6007 5552 6059 5597
rect 6007 5518 6015 5552
rect 6049 5518 6059 5552
rect 6007 5487 6059 5518
rect 6637 5552 6689 5597
rect 6637 5518 6647 5552
rect 6681 5518 6689 5552
rect 6637 5487 6689 5518
rect 6743 5563 6795 5591
rect 6743 5529 6751 5563
rect 6785 5529 6795 5563
rect 6743 5487 6795 5529
rect 6825 5533 6883 5591
rect 6825 5499 6837 5533
rect 6871 5499 6883 5533
rect 6825 5487 6883 5499
rect 6913 5546 6965 5591
rect 6913 5512 6923 5546
rect 6957 5512 6965 5546
rect 6913 5487 6965 5512
rect 7019 5552 7071 5597
rect 7019 5518 7027 5552
rect 7061 5518 7071 5552
rect 7019 5487 7071 5518
rect 7465 5552 7517 5597
rect 8211 5571 8263 5617
rect 7465 5518 7475 5552
rect 7509 5518 7517 5552
rect 7465 5487 7517 5518
rect 7617 5548 7669 5571
rect 7617 5514 7625 5548
rect 7659 5514 7669 5548
rect 7617 5487 7669 5514
rect 7699 5548 7837 5571
rect 7699 5514 7709 5548
rect 7743 5514 7777 5548
rect 7811 5514 7837 5548
rect 7699 5487 7837 5514
rect 7867 5487 7933 5571
rect 7963 5548 8058 5571
rect 7963 5514 8012 5548
rect 8046 5514 8058 5548
rect 7963 5487 8058 5514
rect 8088 5487 8154 5571
rect 8184 5533 8263 5571
rect 8184 5499 8219 5533
rect 8253 5499 8263 5533
rect 8184 5487 8263 5499
rect 8293 5552 8345 5617
rect 8293 5518 8303 5552
rect 8337 5518 8345 5552
rect 8293 5487 8345 5518
rect 8399 5559 8451 5597
rect 8399 5525 8407 5559
rect 8441 5525 8451 5559
rect 8399 5487 8451 5525
rect 8661 5559 8713 5597
rect 8661 5525 8671 5559
rect 8705 5525 8713 5559
rect 8661 5487 8713 5525
rect 8951 5552 9003 5597
rect 8951 5518 8959 5552
rect 8993 5518 9003 5552
rect 8951 5487 9003 5518
rect 9949 5552 10001 5597
rect 9949 5518 9959 5552
rect 9993 5518 10001 5552
rect 9949 5487 10001 5518
rect 10055 5552 10107 5597
rect 10055 5518 10063 5552
rect 10097 5518 10107 5552
rect 10055 5487 10107 5518
rect 11053 5552 11105 5597
rect 11053 5518 11063 5552
rect 11097 5518 11105 5552
rect 11053 5487 11105 5518
rect 11159 5559 11211 5597
rect 11159 5525 11167 5559
rect 11201 5525 11211 5559
rect 11159 5487 11211 5525
rect 11421 5559 11473 5597
rect 11737 5571 11789 5617
rect 11421 5525 11431 5559
rect 11465 5525 11473 5559
rect 11421 5487 11473 5525
rect 11556 5543 11608 5571
rect 11556 5509 11564 5543
rect 11598 5509 11608 5543
rect 11556 5487 11608 5509
rect 11638 5543 11692 5571
rect 11638 5509 11648 5543
rect 11682 5509 11692 5543
rect 11638 5487 11692 5509
rect 11722 5543 11789 5571
rect 11722 5509 11744 5543
rect 11778 5509 11789 5543
rect 11722 5487 11789 5509
rect 11819 5603 11871 5617
rect 11819 5569 11829 5603
rect 11863 5569 11871 5603
rect 11819 5535 11871 5569
rect 11819 5501 11829 5535
rect 11863 5501 11871 5535
rect 11819 5487 11871 5501
rect 11987 5552 12039 5597
rect 11987 5518 11995 5552
rect 12029 5518 12039 5552
rect 11987 5487 12039 5518
rect 12617 5552 12669 5597
rect 13025 5571 13077 5617
rect 12617 5518 12627 5552
rect 12661 5518 12669 5552
rect 12617 5487 12669 5518
rect 12844 5543 12896 5571
rect 12844 5509 12852 5543
rect 12886 5509 12896 5543
rect 12844 5487 12896 5509
rect 12926 5543 12980 5571
rect 12926 5509 12936 5543
rect 12970 5509 12980 5543
rect 12926 5487 12980 5509
rect 13010 5543 13077 5571
rect 13010 5509 13032 5543
rect 13066 5509 13077 5543
rect 13010 5487 13077 5509
rect 13107 5603 13159 5617
rect 13107 5569 13117 5603
rect 13151 5569 13159 5603
rect 13107 5535 13159 5569
rect 13107 5501 13117 5535
rect 13151 5501 13159 5535
rect 13107 5487 13159 5501
rect 13275 5552 13327 5597
rect 13275 5518 13283 5552
rect 13317 5518 13327 5552
rect 13275 5487 13327 5518
rect 13905 5552 13957 5597
rect 13905 5518 13915 5552
rect 13949 5518 13957 5552
rect 13905 5487 13957 5518
rect 14103 5552 14155 5597
rect 14103 5518 14111 5552
rect 14145 5518 14155 5552
rect 14103 5487 14155 5518
rect 15101 5552 15153 5597
rect 15101 5518 15111 5552
rect 15145 5518 15153 5552
rect 15101 5487 15153 5518
rect 15207 5552 15259 5597
rect 15207 5518 15215 5552
rect 15249 5518 15259 5552
rect 15207 5487 15259 5518
rect 16205 5552 16257 5597
rect 16205 5518 16215 5552
rect 16249 5518 16257 5552
rect 16205 5487 16257 5518
rect 16311 5552 16363 5597
rect 16311 5518 16319 5552
rect 16353 5518 16363 5552
rect 16311 5487 16363 5518
rect 17309 5552 17361 5597
rect 17309 5518 17319 5552
rect 17353 5518 17361 5552
rect 17309 5487 17361 5518
rect 17415 5552 17467 5597
rect 17415 5518 17423 5552
rect 17457 5518 17467 5552
rect 17415 5487 17467 5518
rect 18413 5552 18465 5597
rect 18413 5518 18423 5552
rect 18457 5518 18465 5552
rect 18413 5487 18465 5518
rect 18611 5554 18663 5597
rect 18611 5520 18619 5554
rect 18653 5520 18663 5554
rect 18611 5487 18663 5520
rect 18781 5554 18833 5597
rect 18781 5520 18791 5554
rect 18825 5520 18833 5554
rect 18781 5487 18833 5520
rect 1131 5360 1183 5393
rect 1131 5326 1139 5360
rect 1173 5326 1183 5360
rect 1131 5283 1183 5326
rect 1301 5360 1353 5393
rect 1301 5326 1311 5360
rect 1345 5326 1353 5360
rect 1301 5283 1353 5326
rect 1407 5362 1459 5393
rect 1407 5328 1415 5362
rect 1449 5328 1459 5362
rect 1407 5283 1459 5328
rect 2405 5362 2457 5393
rect 2405 5328 2415 5362
rect 2449 5328 2457 5362
rect 2405 5283 2457 5328
rect 2511 5360 2563 5393
rect 2511 5326 2519 5360
rect 2553 5326 2563 5360
rect 2511 5283 2563 5326
rect 2681 5360 2733 5393
rect 2681 5326 2691 5360
rect 2725 5326 2733 5360
rect 2681 5283 2733 5326
rect 2787 5355 2839 5393
rect 2787 5321 2795 5355
rect 2829 5321 2839 5355
rect 2787 5309 2839 5321
rect 2869 5381 2923 5393
rect 2869 5347 2879 5381
rect 2913 5347 2923 5381
rect 2869 5309 2923 5347
rect 2953 5355 3005 5393
rect 2953 5321 2963 5355
rect 2997 5321 3005 5355
rect 2953 5309 3005 5321
rect 3073 5385 3178 5393
rect 3073 5351 3085 5385
rect 3119 5351 3178 5385
rect 3073 5309 3178 5351
rect 3208 5379 3273 5393
rect 3208 5345 3218 5379
rect 3252 5345 3273 5379
rect 3208 5321 3273 5345
rect 3303 5379 3369 5393
rect 3303 5345 3325 5379
rect 3359 5345 3369 5379
rect 3303 5321 3369 5345
rect 3399 5321 3535 5393
rect 3208 5309 3258 5321
rect 3417 5309 3535 5321
rect 3565 5309 3607 5393
rect 3637 5381 3739 5393
rect 3637 5347 3671 5381
rect 3705 5347 3739 5381
rect 3637 5309 3739 5347
rect 3689 5265 3739 5309
rect 3769 5385 3838 5393
rect 3769 5351 3783 5385
rect 3817 5351 3838 5385
rect 3769 5321 3838 5351
rect 3868 5381 3947 5393
rect 3868 5347 3893 5381
rect 3927 5347 3947 5381
rect 3868 5321 3947 5347
rect 3977 5321 4043 5393
rect 3769 5265 3823 5321
rect 3993 5309 4043 5321
rect 4073 5385 4192 5393
rect 4073 5351 4105 5385
rect 4139 5351 4192 5385
rect 4073 5309 4192 5351
rect 4222 5309 4283 5393
rect 4313 5365 4365 5393
rect 4313 5331 4323 5365
rect 4357 5331 4365 5365
rect 4313 5309 4365 5331
rect 4419 5381 4491 5393
rect 4419 5347 4447 5381
rect 4481 5347 4491 5381
rect 4419 5309 4491 5347
rect 4441 5263 4491 5309
rect 4521 5331 4573 5393
rect 4521 5297 4531 5331
rect 4565 5297 4573 5331
rect 4521 5263 4573 5297
rect 4627 5362 4679 5393
rect 4627 5328 4635 5362
rect 4669 5328 4679 5362
rect 4627 5283 4679 5328
rect 5625 5362 5677 5393
rect 5625 5328 5635 5362
rect 5669 5328 5677 5362
rect 5625 5283 5677 5328
rect 5731 5362 5783 5393
rect 5731 5328 5739 5362
rect 5773 5328 5783 5362
rect 5731 5283 5783 5328
rect 6177 5362 6229 5393
rect 6177 5328 6187 5362
rect 6221 5328 6229 5362
rect 6177 5283 6229 5328
rect 6375 5360 6427 5393
rect 6375 5326 6383 5360
rect 6417 5326 6427 5360
rect 6375 5283 6427 5326
rect 6545 5360 6597 5393
rect 6545 5326 6555 5360
rect 6589 5326 6597 5360
rect 6545 5283 6597 5326
rect 6651 5362 6703 5393
rect 6651 5328 6659 5362
rect 6693 5328 6703 5362
rect 6651 5263 6703 5328
rect 6733 5381 6812 5393
rect 6733 5347 6743 5381
rect 6777 5347 6812 5381
rect 6733 5309 6812 5347
rect 6842 5309 6908 5393
rect 6938 5366 7033 5393
rect 6938 5332 6950 5366
rect 6984 5332 7033 5366
rect 6938 5309 7033 5332
rect 7063 5309 7129 5393
rect 7159 5366 7297 5393
rect 7159 5332 7185 5366
rect 7219 5332 7253 5366
rect 7287 5332 7297 5366
rect 7159 5309 7297 5332
rect 7327 5366 7379 5393
rect 7327 5332 7337 5366
rect 7371 5332 7379 5366
rect 7327 5309 7379 5332
rect 7479 5355 7531 5393
rect 7479 5321 7487 5355
rect 7521 5321 7531 5355
rect 6733 5263 6785 5309
rect 7479 5283 7531 5321
rect 7741 5355 7793 5393
rect 7741 5321 7751 5355
rect 7785 5321 7793 5355
rect 7741 5283 7793 5321
rect 7847 5355 7899 5393
rect 7847 5321 7855 5355
rect 7889 5321 7899 5355
rect 7847 5309 7899 5321
rect 7929 5381 7983 5393
rect 7929 5347 7939 5381
rect 7973 5347 7983 5381
rect 7929 5309 7983 5347
rect 8013 5355 8065 5393
rect 8013 5321 8023 5355
rect 8057 5321 8065 5355
rect 8013 5309 8065 5321
rect 8133 5385 8238 5393
rect 8133 5351 8145 5385
rect 8179 5351 8238 5385
rect 8133 5309 8238 5351
rect 8268 5379 8333 5393
rect 8268 5345 8278 5379
rect 8312 5345 8333 5379
rect 8268 5321 8333 5345
rect 8363 5379 8429 5393
rect 8363 5345 8385 5379
rect 8419 5345 8429 5379
rect 8363 5321 8429 5345
rect 8459 5321 8595 5393
rect 8268 5309 8318 5321
rect 8477 5309 8595 5321
rect 8625 5309 8667 5393
rect 8697 5381 8799 5393
rect 8697 5347 8731 5381
rect 8765 5347 8799 5381
rect 8697 5309 8799 5347
rect 8749 5265 8799 5309
rect 8829 5385 8898 5393
rect 8829 5351 8843 5385
rect 8877 5351 8898 5385
rect 8829 5321 8898 5351
rect 8928 5381 9007 5393
rect 8928 5347 8953 5381
rect 8987 5347 9007 5381
rect 8928 5321 9007 5347
rect 9037 5321 9103 5393
rect 8829 5265 8883 5321
rect 9053 5309 9103 5321
rect 9133 5385 9252 5393
rect 9133 5351 9165 5385
rect 9199 5351 9252 5385
rect 9133 5309 9252 5351
rect 9282 5309 9343 5393
rect 9373 5365 9425 5393
rect 9373 5331 9383 5365
rect 9417 5331 9425 5365
rect 9373 5309 9425 5331
rect 9479 5381 9551 5393
rect 9479 5347 9507 5381
rect 9541 5347 9551 5381
rect 9479 5309 9551 5347
rect 9501 5263 9551 5309
rect 9581 5331 9633 5393
rect 9581 5297 9591 5331
rect 9625 5297 9633 5331
rect 9581 5263 9633 5297
rect 9687 5355 9739 5393
rect 9687 5321 9695 5355
rect 9729 5321 9739 5355
rect 9687 5283 9739 5321
rect 9949 5355 10001 5393
rect 9949 5321 9959 5355
rect 9993 5321 10001 5355
rect 9949 5283 10001 5321
rect 10101 5366 10153 5393
rect 10101 5332 10109 5366
rect 10143 5332 10153 5366
rect 10101 5309 10153 5332
rect 10183 5366 10321 5393
rect 10183 5332 10193 5366
rect 10227 5332 10261 5366
rect 10295 5332 10321 5366
rect 10183 5309 10321 5332
rect 10351 5309 10417 5393
rect 10447 5366 10542 5393
rect 10447 5332 10496 5366
rect 10530 5332 10542 5366
rect 10447 5309 10542 5332
rect 10572 5309 10638 5393
rect 10668 5381 10747 5393
rect 10668 5347 10703 5381
rect 10737 5347 10747 5381
rect 10668 5309 10747 5347
rect 10695 5263 10747 5309
rect 10777 5362 10829 5393
rect 10777 5328 10787 5362
rect 10821 5328 10829 5362
rect 10777 5263 10829 5328
rect 10883 5362 10935 5393
rect 10883 5328 10891 5362
rect 10925 5328 10935 5362
rect 10883 5283 10935 5328
rect 11329 5362 11381 5393
rect 11329 5328 11339 5362
rect 11373 5328 11381 5362
rect 11329 5283 11381 5328
rect 11711 5362 11763 5393
rect 11711 5328 11719 5362
rect 11753 5328 11763 5362
rect 11711 5263 11763 5328
rect 11793 5381 11872 5393
rect 11793 5347 11803 5381
rect 11837 5347 11872 5381
rect 11793 5309 11872 5347
rect 11902 5309 11968 5393
rect 11998 5366 12093 5393
rect 11998 5332 12010 5366
rect 12044 5332 12093 5366
rect 11998 5309 12093 5332
rect 12123 5309 12189 5393
rect 12219 5366 12357 5393
rect 12219 5332 12245 5366
rect 12279 5332 12313 5366
rect 12347 5332 12357 5366
rect 12219 5309 12357 5332
rect 12387 5366 12439 5393
rect 12387 5332 12397 5366
rect 12431 5332 12439 5366
rect 12387 5309 12439 5332
rect 12539 5355 12591 5393
rect 12539 5321 12547 5355
rect 12581 5321 12591 5355
rect 11793 5263 11845 5309
rect 12539 5283 12591 5321
rect 12801 5355 12853 5393
rect 12801 5321 12811 5355
rect 12845 5321 12853 5355
rect 12801 5283 12853 5321
rect 12953 5366 13005 5393
rect 12953 5332 12961 5366
rect 12995 5332 13005 5366
rect 12953 5309 13005 5332
rect 13035 5366 13173 5393
rect 13035 5332 13045 5366
rect 13079 5332 13113 5366
rect 13147 5332 13173 5366
rect 13035 5309 13173 5332
rect 13203 5309 13269 5393
rect 13299 5366 13394 5393
rect 13299 5332 13348 5366
rect 13382 5332 13394 5366
rect 13299 5309 13394 5332
rect 13424 5309 13490 5393
rect 13520 5381 13599 5393
rect 13520 5347 13555 5381
rect 13589 5347 13599 5381
rect 13520 5309 13599 5347
rect 13547 5263 13599 5309
rect 13629 5362 13681 5393
rect 13629 5328 13639 5362
rect 13673 5328 13681 5362
rect 13629 5263 13681 5328
rect 13735 5362 13787 5393
rect 13735 5328 13743 5362
rect 13777 5328 13787 5362
rect 13735 5283 13787 5328
rect 14733 5362 14785 5393
rect 14733 5328 14743 5362
rect 14777 5328 14785 5362
rect 14733 5283 14785 5328
rect 14839 5362 14891 5393
rect 14839 5328 14847 5362
rect 14881 5328 14891 5362
rect 14839 5283 14891 5328
rect 15837 5362 15889 5393
rect 15837 5328 15847 5362
rect 15881 5328 15889 5362
rect 15837 5283 15889 5328
rect 15943 5362 15995 5393
rect 15943 5328 15951 5362
rect 15985 5328 15995 5362
rect 15943 5283 15995 5328
rect 16389 5362 16441 5393
rect 16389 5328 16399 5362
rect 16433 5328 16441 5362
rect 16389 5283 16441 5328
rect 16679 5362 16731 5393
rect 16679 5328 16687 5362
rect 16721 5328 16731 5362
rect 16679 5283 16731 5328
rect 17677 5362 17729 5393
rect 17677 5328 17687 5362
rect 17721 5328 17729 5362
rect 17677 5283 17729 5328
rect 17783 5362 17835 5393
rect 17783 5328 17791 5362
rect 17825 5328 17835 5362
rect 17783 5283 17835 5328
rect 18413 5362 18465 5393
rect 18413 5328 18423 5362
rect 18457 5328 18465 5362
rect 18413 5283 18465 5328
rect 18611 5360 18663 5393
rect 18611 5326 18619 5360
rect 18653 5326 18663 5360
rect 18611 5283 18663 5326
rect 18781 5360 18833 5393
rect 18781 5326 18791 5360
rect 18825 5326 18833 5360
rect 18781 5283 18833 5326
rect 1131 4466 1183 4509
rect 1131 4432 1139 4466
rect 1173 4432 1183 4466
rect 1131 4399 1183 4432
rect 1301 4466 1353 4509
rect 1301 4432 1311 4466
rect 1345 4432 1353 4466
rect 1301 4399 1353 4432
rect 1407 4464 1459 4509
rect 1407 4430 1415 4464
rect 1449 4430 1459 4464
rect 1407 4399 1459 4430
rect 2037 4464 2089 4509
rect 2037 4430 2047 4464
rect 2081 4430 2089 4464
rect 2037 4399 2089 4430
rect 2143 4466 2195 4509
rect 2143 4432 2151 4466
rect 2185 4432 2195 4466
rect 2143 4399 2195 4432
rect 2313 4466 2365 4509
rect 2313 4432 2323 4466
rect 2357 4432 2365 4466
rect 2313 4399 2365 4432
rect 2438 4471 2490 4529
rect 2438 4437 2446 4471
rect 2480 4437 2490 4471
rect 2438 4399 2490 4437
rect 2520 4483 2570 4529
rect 2520 4445 2585 4483
rect 2520 4411 2536 4445
rect 2570 4411 2585 4445
rect 2520 4399 2585 4411
rect 2685 4471 2737 4483
rect 2685 4437 2695 4471
rect 2729 4437 2737 4471
rect 2685 4399 2737 4437
rect 2791 4471 2843 4483
rect 2791 4437 2799 4471
rect 2833 4437 2843 4471
rect 2791 4399 2843 4437
rect 2943 4445 2997 4483
rect 2943 4411 2953 4445
rect 2987 4411 2997 4445
rect 2943 4399 2997 4411
rect 3027 4471 3079 4483
rect 3027 4437 3037 4471
rect 3071 4437 3079 4471
rect 3027 4399 3079 4437
rect 3155 4464 3207 4509
rect 3155 4430 3163 4464
rect 3197 4430 3207 4464
rect 3155 4399 3207 4430
rect 3601 4464 3653 4509
rect 3601 4430 3611 4464
rect 3645 4430 3653 4464
rect 3601 4399 3653 4430
rect 3985 4449 4043 4483
rect 3985 4415 3998 4449
rect 4032 4415 4043 4449
rect 3985 4399 4043 4415
rect 4073 4471 4129 4483
rect 4073 4437 4084 4471
rect 4118 4437 4129 4471
rect 4073 4399 4129 4437
rect 4159 4449 4215 4483
rect 4159 4415 4170 4449
rect 4204 4415 4215 4449
rect 4159 4399 4215 4415
rect 4245 4471 4301 4483
rect 4245 4437 4256 4471
rect 4290 4437 4301 4471
rect 4245 4399 4301 4437
rect 4331 4449 4398 4483
rect 4331 4415 4353 4449
rect 4387 4415 4398 4449
rect 4331 4399 4398 4415
rect 4428 4453 4481 4483
rect 4428 4419 4439 4453
rect 4473 4419 4481 4453
rect 4428 4399 4481 4419
rect 4535 4471 4587 4509
rect 4535 4437 4543 4471
rect 4577 4437 4587 4471
rect 4535 4399 4587 4437
rect 4797 4471 4849 4509
rect 4797 4437 4807 4471
rect 4841 4437 4849 4471
rect 4797 4399 4849 4437
rect 6069 4515 6121 4529
rect 5087 4464 5139 4509
rect 5087 4430 5095 4464
rect 5129 4430 5139 4464
rect 5087 4399 5139 4430
rect 5717 4464 5769 4509
rect 5717 4430 5727 4464
rect 5761 4430 5769 4464
rect 5717 4399 5769 4430
rect 6069 4481 6077 4515
rect 6111 4481 6121 4515
rect 6069 4447 6121 4481
rect 6069 4413 6077 4447
rect 6111 4413 6121 4447
rect 6069 4399 6121 4413
rect 6151 4483 6203 4529
rect 6151 4455 6218 4483
rect 6151 4421 6162 4455
rect 6196 4421 6218 4455
rect 6151 4399 6218 4421
rect 6248 4455 6302 4483
rect 6248 4421 6258 4455
rect 6292 4421 6302 4455
rect 6248 4399 6302 4421
rect 6332 4455 6384 4483
rect 6332 4421 6342 4455
rect 6376 4421 6384 4455
rect 6332 4399 6384 4421
rect 6467 4471 6519 4509
rect 6467 4437 6475 4471
rect 6509 4437 6519 4471
rect 6467 4399 6519 4437
rect 6729 4471 6781 4509
rect 7045 4483 7097 4529
rect 6729 4437 6739 4471
rect 6773 4437 6781 4471
rect 6729 4399 6781 4437
rect 6864 4455 6916 4483
rect 6864 4421 6872 4455
rect 6906 4421 6916 4455
rect 6864 4399 6916 4421
rect 6946 4455 7000 4483
rect 6946 4421 6956 4455
rect 6990 4421 7000 4455
rect 6946 4399 7000 4421
rect 7030 4455 7097 4483
rect 7030 4421 7052 4455
rect 7086 4421 7097 4455
rect 7030 4399 7097 4421
rect 7127 4515 7179 4529
rect 7127 4481 7137 4515
rect 7171 4481 7179 4515
rect 7127 4447 7179 4481
rect 7127 4413 7137 4447
rect 7171 4413 7179 4447
rect 7127 4399 7179 4413
rect 7295 4464 7347 4509
rect 7295 4430 7303 4464
rect 7337 4430 7347 4464
rect 7295 4399 7347 4430
rect 7741 4464 7793 4509
rect 7741 4430 7751 4464
rect 7785 4430 7793 4464
rect 7741 4399 7793 4430
rect 7847 4464 7899 4529
rect 7847 4430 7855 4464
rect 7889 4430 7899 4464
rect 7847 4399 7899 4430
rect 7929 4483 7981 4529
rect 7929 4445 8008 4483
rect 7929 4411 7939 4445
rect 7973 4411 8008 4445
rect 7929 4399 8008 4411
rect 8038 4399 8104 4483
rect 8134 4460 8229 4483
rect 8134 4426 8146 4460
rect 8180 4426 8229 4460
rect 8134 4399 8229 4426
rect 8259 4399 8325 4483
rect 8355 4460 8493 4483
rect 8355 4426 8381 4460
rect 8415 4426 8449 4460
rect 8483 4426 8493 4460
rect 8355 4399 8493 4426
rect 8523 4460 8575 4483
rect 8523 4426 8533 4460
rect 8567 4426 8575 4460
rect 8523 4399 8575 4426
rect 9345 4483 9397 4529
rect 9164 4455 9216 4483
rect 9164 4421 9172 4455
rect 9206 4421 9216 4455
rect 9164 4399 9216 4421
rect 9246 4455 9300 4483
rect 9246 4421 9256 4455
rect 9290 4421 9300 4455
rect 9246 4399 9300 4421
rect 9330 4455 9397 4483
rect 9330 4421 9352 4455
rect 9386 4421 9397 4455
rect 9330 4399 9397 4421
rect 9427 4515 9479 4529
rect 9427 4481 9437 4515
rect 9471 4481 9479 4515
rect 9427 4447 9479 4481
rect 9427 4413 9437 4447
rect 9471 4413 9479 4447
rect 9427 4399 9479 4413
rect 9595 4471 9647 4509
rect 9595 4437 9603 4471
rect 9637 4437 9647 4471
rect 9595 4399 9647 4437
rect 9857 4471 9909 4509
rect 9857 4437 9867 4471
rect 9901 4437 9909 4471
rect 9857 4399 9909 4437
rect 10147 4471 10199 4509
rect 10147 4437 10155 4471
rect 10189 4437 10199 4471
rect 10147 4399 10199 4437
rect 10409 4471 10461 4509
rect 10725 4483 10777 4529
rect 10409 4437 10419 4471
rect 10453 4437 10461 4471
rect 10409 4399 10461 4437
rect 10544 4455 10596 4483
rect 10544 4421 10552 4455
rect 10586 4421 10596 4455
rect 10544 4399 10596 4421
rect 10626 4455 10680 4483
rect 10626 4421 10636 4455
rect 10670 4421 10680 4455
rect 10626 4399 10680 4421
rect 10710 4455 10777 4483
rect 10710 4421 10732 4455
rect 10766 4421 10777 4455
rect 10710 4399 10777 4421
rect 10807 4515 10859 4529
rect 10807 4481 10817 4515
rect 10851 4481 10859 4515
rect 10807 4447 10859 4481
rect 10807 4413 10817 4447
rect 10851 4413 10859 4447
rect 10807 4399 10859 4413
rect 10975 4471 11027 4509
rect 10975 4437 10983 4471
rect 11017 4437 11027 4471
rect 10975 4399 11027 4437
rect 11237 4471 11289 4509
rect 11237 4437 11247 4471
rect 11281 4437 11289 4471
rect 11237 4399 11289 4437
rect 11343 4458 11395 4503
rect 11343 4424 11351 4458
rect 11385 4424 11395 4458
rect 11343 4399 11395 4424
rect 11425 4445 11483 4503
rect 11425 4411 11437 4445
rect 11471 4411 11483 4445
rect 11425 4399 11483 4411
rect 11513 4475 11565 4503
rect 11513 4441 11523 4475
rect 11557 4441 11565 4475
rect 11513 4399 11565 4441
rect 11619 4471 11671 4509
rect 11619 4437 11627 4471
rect 11661 4437 11671 4471
rect 11619 4399 11671 4437
rect 11881 4471 11933 4509
rect 12627 4483 12679 4529
rect 11881 4437 11891 4471
rect 11925 4437 11933 4471
rect 11881 4399 11933 4437
rect 12033 4460 12085 4483
rect 12033 4426 12041 4460
rect 12075 4426 12085 4460
rect 12033 4399 12085 4426
rect 12115 4460 12253 4483
rect 12115 4426 12125 4460
rect 12159 4426 12193 4460
rect 12227 4426 12253 4460
rect 12115 4399 12253 4426
rect 12283 4399 12349 4483
rect 12379 4460 12474 4483
rect 12379 4426 12428 4460
rect 12462 4426 12474 4460
rect 12379 4399 12474 4426
rect 12504 4399 12570 4483
rect 12600 4445 12679 4483
rect 12600 4411 12635 4445
rect 12669 4411 12679 4445
rect 12600 4399 12679 4411
rect 12709 4464 12761 4529
rect 12709 4430 12719 4464
rect 12753 4430 12761 4464
rect 12709 4399 12761 4430
rect 12815 4471 12867 4509
rect 12815 4437 12823 4471
rect 12857 4437 12867 4471
rect 12815 4399 12867 4437
rect 13077 4471 13129 4509
rect 13077 4437 13087 4471
rect 13121 4437 13129 4471
rect 13077 4399 13129 4437
rect 13183 4475 13235 4503
rect 13183 4441 13191 4475
rect 13225 4441 13235 4475
rect 13183 4399 13235 4441
rect 13265 4445 13323 4503
rect 13265 4411 13277 4445
rect 13311 4411 13323 4445
rect 13265 4399 13323 4411
rect 13353 4458 13405 4503
rect 13353 4424 13363 4458
rect 13397 4424 13405 4458
rect 13353 4399 13405 4424
rect 13459 4464 13511 4509
rect 13459 4430 13467 4464
rect 13501 4430 13511 4464
rect 13459 4399 13511 4430
rect 13905 4464 13957 4509
rect 13905 4430 13915 4464
rect 13949 4430 13957 4464
rect 13905 4399 13957 4430
rect 14103 4464 14155 4509
rect 14103 4430 14111 4464
rect 14145 4430 14155 4464
rect 14103 4399 14155 4430
rect 15101 4464 15153 4509
rect 15417 4483 15469 4529
rect 15101 4430 15111 4464
rect 15145 4430 15153 4464
rect 15101 4399 15153 4430
rect 15236 4455 15288 4483
rect 15236 4421 15244 4455
rect 15278 4421 15288 4455
rect 15236 4399 15288 4421
rect 15318 4455 15372 4483
rect 15318 4421 15328 4455
rect 15362 4421 15372 4455
rect 15318 4399 15372 4421
rect 15402 4455 15469 4483
rect 15402 4421 15424 4455
rect 15458 4421 15469 4455
rect 15402 4399 15469 4421
rect 15499 4515 15551 4529
rect 15499 4481 15509 4515
rect 15543 4481 15551 4515
rect 15499 4447 15551 4481
rect 15499 4413 15509 4447
rect 15543 4413 15551 4447
rect 15499 4399 15551 4413
rect 15667 4471 15719 4509
rect 15667 4437 15675 4471
rect 15709 4437 15719 4471
rect 15667 4399 15719 4437
rect 15929 4471 15981 4509
rect 15929 4437 15939 4471
rect 15973 4437 15981 4471
rect 15929 4399 15981 4437
rect 16035 4475 16087 4503
rect 16035 4441 16043 4475
rect 16077 4441 16087 4475
rect 16035 4399 16087 4441
rect 16117 4445 16175 4503
rect 16117 4411 16129 4445
rect 16163 4411 16175 4445
rect 16117 4399 16175 4411
rect 16205 4458 16257 4503
rect 16205 4424 16215 4458
rect 16249 4424 16257 4458
rect 16205 4399 16257 4424
rect 16311 4471 16363 4509
rect 16311 4437 16319 4471
rect 16353 4437 16363 4471
rect 16311 4399 16363 4437
rect 16573 4471 16625 4509
rect 16573 4437 16583 4471
rect 16617 4437 16625 4471
rect 16573 4399 16625 4437
rect 16679 4475 16731 4503
rect 16679 4441 16687 4475
rect 16721 4441 16731 4475
rect 16679 4399 16731 4441
rect 16761 4445 16819 4503
rect 16761 4411 16773 4445
rect 16807 4411 16819 4445
rect 16761 4399 16819 4411
rect 16849 4458 16901 4503
rect 16849 4424 16859 4458
rect 16893 4424 16901 4458
rect 16849 4399 16901 4424
rect 16955 4464 17007 4509
rect 16955 4430 16963 4464
rect 16997 4430 17007 4464
rect 16955 4399 17007 4430
rect 17953 4464 18005 4509
rect 17953 4430 17963 4464
rect 17997 4430 18005 4464
rect 17953 4399 18005 4430
rect 18059 4464 18111 4509
rect 18059 4430 18067 4464
rect 18101 4430 18111 4464
rect 18059 4399 18111 4430
rect 18505 4464 18557 4509
rect 18505 4430 18515 4464
rect 18549 4430 18557 4464
rect 18505 4399 18557 4430
rect 18611 4466 18663 4509
rect 18611 4432 18619 4466
rect 18653 4432 18663 4466
rect 18611 4399 18663 4432
rect 18781 4466 18833 4509
rect 18781 4432 18791 4466
rect 18825 4432 18833 4466
rect 18781 4399 18833 4432
rect 1131 4272 1183 4305
rect 1131 4238 1139 4272
rect 1173 4238 1183 4272
rect 1131 4195 1183 4238
rect 1301 4272 1353 4305
rect 1301 4238 1311 4272
rect 1345 4238 1353 4272
rect 1301 4195 1353 4238
rect 1407 4274 1459 4305
rect 1407 4240 1415 4274
rect 1449 4240 1459 4274
rect 1407 4195 1459 4240
rect 2037 4274 2089 4305
rect 2037 4240 2047 4274
rect 2081 4240 2089 4274
rect 2037 4195 2089 4240
rect 2235 4280 2287 4305
rect 2235 4246 2243 4280
rect 2277 4246 2287 4280
rect 2235 4201 2287 4246
rect 2317 4293 2375 4305
rect 2317 4259 2329 4293
rect 2363 4259 2375 4293
rect 2317 4201 2375 4259
rect 2405 4263 2457 4305
rect 2405 4229 2415 4263
rect 2449 4229 2457 4263
rect 2405 4201 2457 4229
rect 2511 4267 2563 4305
rect 2511 4233 2519 4267
rect 2553 4233 2563 4267
rect 2511 4195 2563 4233
rect 2773 4267 2825 4305
rect 2773 4233 2783 4267
rect 2817 4233 2825 4267
rect 2773 4195 2825 4233
rect 2879 4267 2931 4305
rect 2879 4233 2887 4267
rect 2921 4233 2931 4267
rect 2879 4221 2931 4233
rect 2961 4293 3015 4305
rect 2961 4259 2971 4293
rect 3005 4259 3015 4293
rect 2961 4221 3015 4259
rect 3045 4267 3097 4305
rect 3045 4233 3055 4267
rect 3089 4233 3097 4267
rect 3045 4221 3097 4233
rect 3165 4297 3270 4305
rect 3165 4263 3177 4297
rect 3211 4263 3270 4297
rect 3165 4221 3270 4263
rect 3300 4291 3365 4305
rect 3300 4257 3310 4291
rect 3344 4257 3365 4291
rect 3300 4233 3365 4257
rect 3395 4291 3461 4305
rect 3395 4257 3417 4291
rect 3451 4257 3461 4291
rect 3395 4233 3461 4257
rect 3491 4233 3627 4305
rect 3300 4221 3350 4233
rect 3509 4221 3627 4233
rect 3657 4221 3699 4305
rect 3729 4293 3831 4305
rect 3729 4259 3763 4293
rect 3797 4259 3831 4293
rect 3729 4221 3831 4259
rect 3781 4177 3831 4221
rect 3861 4297 3930 4305
rect 3861 4263 3875 4297
rect 3909 4263 3930 4297
rect 3861 4233 3930 4263
rect 3960 4293 4039 4305
rect 3960 4259 3985 4293
rect 4019 4259 4039 4293
rect 3960 4233 4039 4259
rect 4069 4233 4135 4305
rect 3861 4177 3915 4233
rect 4085 4221 4135 4233
rect 4165 4297 4284 4305
rect 4165 4263 4197 4297
rect 4231 4263 4284 4297
rect 4165 4221 4284 4263
rect 4314 4221 4375 4305
rect 4405 4277 4457 4305
rect 4405 4243 4415 4277
rect 4449 4243 4457 4277
rect 4405 4221 4457 4243
rect 4511 4293 4583 4305
rect 4511 4259 4539 4293
rect 4573 4259 4583 4293
rect 4511 4221 4583 4259
rect 4533 4175 4583 4221
rect 4613 4243 4665 4305
rect 4613 4209 4623 4243
rect 4657 4209 4665 4243
rect 4613 4175 4665 4209
rect 4719 4267 4771 4305
rect 4719 4233 4727 4267
rect 4761 4233 4771 4267
rect 4719 4195 4771 4233
rect 4981 4267 5033 4305
rect 4981 4233 4991 4267
rect 5025 4233 5033 4267
rect 4981 4195 5033 4233
rect 5363 4274 5415 4305
rect 5363 4240 5371 4274
rect 5405 4240 5415 4274
rect 5363 4195 5415 4240
rect 5993 4274 6045 4305
rect 5993 4240 6003 4274
rect 6037 4240 6045 4274
rect 5993 4195 6045 4240
rect 6375 4272 6427 4305
rect 6375 4238 6383 4272
rect 6417 4238 6427 4272
rect 6375 4195 6427 4238
rect 6545 4272 6597 4305
rect 6545 4238 6555 4272
rect 6589 4238 6597 4272
rect 6545 4195 6597 4238
rect 6651 4263 6703 4305
rect 6651 4229 6659 4263
rect 6693 4229 6703 4263
rect 6651 4201 6703 4229
rect 6733 4293 6791 4305
rect 6733 4259 6745 4293
rect 6779 4259 6791 4293
rect 6733 4201 6791 4259
rect 6821 4280 6873 4305
rect 6821 4246 6831 4280
rect 6865 4246 6873 4280
rect 6821 4201 6873 4246
rect 6927 4274 6979 4305
rect 6927 4240 6935 4274
rect 6969 4240 6979 4274
rect 6927 4195 6979 4240
rect 7557 4274 7609 4305
rect 7557 4240 7567 4274
rect 7601 4240 7609 4274
rect 7557 4195 7609 4240
rect 7709 4278 7761 4305
rect 7709 4244 7717 4278
rect 7751 4244 7761 4278
rect 7709 4221 7761 4244
rect 7791 4278 7929 4305
rect 7791 4244 7801 4278
rect 7835 4244 7869 4278
rect 7903 4244 7929 4278
rect 7791 4221 7929 4244
rect 7959 4221 8025 4305
rect 8055 4278 8150 4305
rect 8055 4244 8104 4278
rect 8138 4244 8150 4278
rect 8055 4221 8150 4244
rect 8180 4221 8246 4305
rect 8276 4293 8355 4305
rect 8276 4259 8311 4293
rect 8345 4259 8355 4293
rect 8276 4221 8355 4259
rect 8303 4175 8355 4221
rect 8385 4274 8437 4305
rect 8385 4240 8395 4274
rect 8429 4240 8437 4274
rect 8385 4175 8437 4240
rect 8491 4267 8543 4305
rect 8491 4233 8499 4267
rect 8533 4233 8543 4267
rect 8491 4195 8543 4233
rect 8753 4267 8805 4305
rect 8753 4233 8763 4267
rect 8797 4233 8805 4267
rect 8753 4195 8805 4233
rect 8951 4293 9004 4305
rect 8951 4259 8959 4293
rect 8993 4259 9004 4293
rect 8951 4221 9004 4259
rect 9034 4280 9090 4305
rect 9034 4246 9045 4280
rect 9079 4246 9090 4280
rect 9034 4221 9090 4246
rect 9120 4280 9176 4305
rect 9120 4246 9131 4280
rect 9165 4246 9176 4280
rect 9120 4221 9176 4246
rect 9206 4280 9262 4305
rect 9206 4246 9217 4280
rect 9251 4246 9262 4280
rect 9206 4221 9262 4246
rect 9292 4280 9348 4305
rect 9292 4246 9303 4280
rect 9337 4246 9348 4280
rect 9292 4221 9348 4246
rect 9378 4280 9434 4305
rect 9378 4246 9389 4280
rect 9423 4246 9434 4280
rect 9378 4221 9434 4246
rect 9464 4289 9520 4305
rect 9464 4255 9475 4289
rect 9509 4255 9520 4289
rect 9464 4221 9520 4255
rect 9550 4280 9606 4305
rect 9550 4246 9561 4280
rect 9595 4246 9606 4280
rect 9550 4221 9606 4246
rect 9636 4289 9692 4305
rect 9636 4255 9647 4289
rect 9681 4255 9692 4289
rect 9636 4221 9692 4255
rect 9722 4280 9778 4305
rect 9722 4246 9733 4280
rect 9767 4246 9778 4280
rect 9722 4221 9778 4246
rect 9808 4289 9864 4305
rect 9808 4255 9819 4289
rect 9853 4255 9864 4289
rect 9808 4221 9864 4255
rect 9894 4280 9950 4305
rect 9894 4246 9905 4280
rect 9939 4246 9950 4280
rect 9894 4221 9950 4246
rect 9980 4289 10035 4305
rect 9980 4255 9991 4289
rect 10025 4255 10035 4289
rect 9980 4221 10035 4255
rect 10065 4280 10121 4305
rect 10065 4246 10076 4280
rect 10110 4246 10121 4280
rect 10065 4221 10121 4246
rect 10151 4289 10207 4305
rect 10151 4255 10162 4289
rect 10196 4255 10207 4289
rect 10151 4221 10207 4255
rect 10237 4280 10293 4305
rect 10237 4246 10248 4280
rect 10282 4246 10293 4280
rect 10237 4221 10293 4246
rect 10323 4289 10379 4305
rect 10323 4255 10334 4289
rect 10368 4255 10379 4289
rect 10323 4221 10379 4255
rect 10409 4280 10465 4305
rect 10409 4246 10420 4280
rect 10454 4246 10465 4280
rect 10409 4221 10465 4246
rect 10495 4289 10551 4305
rect 10495 4255 10506 4289
rect 10540 4255 10551 4289
rect 10495 4221 10551 4255
rect 10581 4280 10637 4305
rect 10581 4246 10592 4280
rect 10626 4246 10637 4280
rect 10581 4221 10637 4246
rect 10667 4289 10720 4305
rect 10667 4255 10678 4289
rect 10712 4255 10720 4289
rect 10667 4221 10720 4255
rect 10791 4274 10843 4305
rect 10791 4240 10799 4274
rect 10833 4240 10843 4274
rect 10791 4195 10843 4240
rect 11237 4274 11289 4305
rect 11237 4240 11247 4274
rect 11281 4240 11289 4274
rect 11237 4195 11289 4240
rect 11711 4243 11763 4305
rect 11711 4209 11719 4243
rect 11753 4209 11763 4243
rect 11711 4175 11763 4209
rect 11793 4293 11865 4305
rect 11793 4259 11803 4293
rect 11837 4259 11865 4293
rect 11793 4221 11865 4259
rect 11919 4277 11971 4305
rect 11919 4243 11927 4277
rect 11961 4243 11971 4277
rect 11919 4221 11971 4243
rect 12001 4221 12062 4305
rect 12092 4297 12211 4305
rect 12092 4263 12145 4297
rect 12179 4263 12211 4297
rect 12092 4221 12211 4263
rect 12241 4233 12307 4305
rect 12337 4293 12416 4305
rect 12337 4259 12357 4293
rect 12391 4259 12416 4293
rect 12337 4233 12416 4259
rect 12446 4297 12515 4305
rect 12446 4263 12467 4297
rect 12501 4263 12515 4297
rect 12446 4233 12515 4263
rect 12241 4221 12291 4233
rect 11793 4175 11843 4221
rect 12461 4177 12515 4233
rect 12545 4293 12647 4305
rect 12545 4259 12579 4293
rect 12613 4259 12647 4293
rect 12545 4221 12647 4259
rect 12677 4221 12719 4305
rect 12749 4233 12885 4305
rect 12915 4291 12981 4305
rect 12915 4257 12925 4291
rect 12959 4257 12981 4291
rect 12915 4233 12981 4257
rect 13011 4291 13076 4305
rect 13011 4257 13032 4291
rect 13066 4257 13076 4291
rect 13011 4233 13076 4257
rect 12749 4221 12867 4233
rect 12545 4177 12595 4221
rect 13026 4221 13076 4233
rect 13106 4297 13211 4305
rect 13106 4263 13165 4297
rect 13199 4263 13211 4297
rect 13106 4221 13211 4263
rect 13279 4267 13331 4305
rect 13279 4233 13287 4267
rect 13321 4233 13331 4267
rect 13279 4221 13331 4233
rect 13361 4293 13415 4305
rect 13361 4259 13371 4293
rect 13405 4259 13415 4293
rect 13361 4221 13415 4259
rect 13445 4267 13497 4305
rect 13445 4233 13455 4267
rect 13489 4233 13497 4267
rect 13445 4221 13497 4233
rect 13551 4267 13603 4305
rect 13551 4233 13559 4267
rect 13593 4233 13603 4267
rect 13551 4195 13603 4233
rect 13813 4267 13865 4305
rect 13813 4233 13823 4267
rect 13857 4233 13865 4267
rect 13813 4195 13865 4233
rect 13919 4267 13971 4305
rect 13919 4233 13927 4267
rect 13961 4233 13971 4267
rect 13919 4221 13971 4233
rect 14001 4293 14055 4305
rect 14001 4259 14011 4293
rect 14045 4259 14055 4293
rect 14001 4221 14055 4259
rect 14085 4267 14137 4305
rect 14085 4233 14095 4267
rect 14129 4233 14137 4267
rect 14085 4221 14137 4233
rect 14205 4297 14310 4305
rect 14205 4263 14217 4297
rect 14251 4263 14310 4297
rect 14205 4221 14310 4263
rect 14340 4291 14405 4305
rect 14340 4257 14350 4291
rect 14384 4257 14405 4291
rect 14340 4233 14405 4257
rect 14435 4291 14501 4305
rect 14435 4257 14457 4291
rect 14491 4257 14501 4291
rect 14435 4233 14501 4257
rect 14531 4233 14667 4305
rect 14340 4221 14390 4233
rect 14549 4221 14667 4233
rect 14697 4221 14739 4305
rect 14769 4293 14871 4305
rect 14769 4259 14803 4293
rect 14837 4259 14871 4293
rect 14769 4221 14871 4259
rect 14821 4177 14871 4221
rect 14901 4297 14970 4305
rect 14901 4263 14915 4297
rect 14949 4263 14970 4297
rect 14901 4233 14970 4263
rect 15000 4293 15079 4305
rect 15000 4259 15025 4293
rect 15059 4259 15079 4293
rect 15000 4233 15079 4259
rect 15109 4233 15175 4305
rect 14901 4177 14955 4233
rect 15125 4221 15175 4233
rect 15205 4297 15324 4305
rect 15205 4263 15237 4297
rect 15271 4263 15324 4297
rect 15205 4221 15324 4263
rect 15354 4221 15415 4305
rect 15445 4277 15497 4305
rect 15445 4243 15455 4277
rect 15489 4243 15497 4277
rect 15445 4221 15497 4243
rect 15551 4293 15623 4305
rect 15551 4259 15579 4293
rect 15613 4259 15623 4293
rect 15551 4221 15623 4259
rect 15573 4175 15623 4221
rect 15653 4243 15705 4305
rect 15653 4209 15663 4243
rect 15697 4209 15705 4243
rect 15653 4175 15705 4209
rect 15759 4274 15811 4305
rect 15759 4240 15767 4274
rect 15801 4240 15811 4274
rect 15759 4195 15811 4240
rect 16389 4274 16441 4305
rect 16389 4240 16399 4274
rect 16433 4240 16441 4274
rect 16389 4195 16441 4240
rect 16679 4274 16731 4305
rect 16679 4240 16687 4274
rect 16721 4240 16731 4274
rect 16679 4195 16731 4240
rect 17677 4274 17729 4305
rect 17677 4240 17687 4274
rect 17721 4240 17729 4274
rect 17677 4195 17729 4240
rect 17783 4274 17835 4305
rect 17783 4240 17791 4274
rect 17825 4240 17835 4274
rect 17783 4195 17835 4240
rect 18413 4274 18465 4305
rect 18413 4240 18423 4274
rect 18457 4240 18465 4274
rect 18413 4195 18465 4240
rect 18611 4272 18663 4305
rect 18611 4238 18619 4272
rect 18653 4238 18663 4272
rect 18611 4195 18663 4238
rect 18781 4272 18833 4305
rect 18781 4238 18791 4272
rect 18825 4238 18833 4272
rect 18781 4195 18833 4238
rect 1131 3378 1183 3421
rect 1131 3344 1139 3378
rect 1173 3344 1183 3378
rect 1131 3311 1183 3344
rect 1301 3378 1353 3421
rect 1301 3344 1311 3378
rect 1345 3344 1353 3378
rect 1301 3311 1353 3344
rect 1407 3378 1459 3421
rect 1407 3344 1415 3378
rect 1449 3344 1459 3378
rect 1407 3311 1459 3344
rect 1577 3378 1629 3421
rect 1577 3344 1587 3378
rect 1621 3344 1629 3378
rect 1577 3311 1629 3344
rect 1683 3383 1735 3395
rect 1683 3349 1691 3383
rect 1725 3349 1735 3383
rect 1683 3311 1735 3349
rect 1765 3357 1819 3395
rect 1765 3323 1775 3357
rect 1809 3323 1819 3357
rect 1765 3311 1819 3323
rect 1849 3383 1901 3395
rect 1849 3349 1859 3383
rect 1893 3349 1901 3383
rect 1849 3311 1901 3349
rect 1969 3353 2074 3395
rect 1969 3319 1981 3353
rect 2015 3319 2074 3353
rect 1969 3311 2074 3319
rect 2104 3383 2154 3395
rect 2585 3395 2635 3439
rect 2313 3383 2431 3395
rect 2104 3359 2169 3383
rect 2104 3325 2114 3359
rect 2148 3325 2169 3359
rect 2104 3311 2169 3325
rect 2199 3359 2265 3383
rect 2199 3325 2221 3359
rect 2255 3325 2265 3359
rect 2199 3311 2265 3325
rect 2295 3311 2431 3383
rect 2461 3311 2503 3395
rect 2533 3357 2635 3395
rect 2533 3323 2567 3357
rect 2601 3323 2635 3357
rect 2533 3311 2635 3323
rect 2665 3383 2719 3439
rect 3337 3395 3387 3441
rect 2889 3383 2939 3395
rect 2665 3353 2734 3383
rect 2665 3319 2679 3353
rect 2713 3319 2734 3353
rect 2665 3311 2734 3319
rect 2764 3357 2843 3383
rect 2764 3323 2789 3357
rect 2823 3323 2843 3357
rect 2764 3311 2843 3323
rect 2873 3311 2939 3383
rect 2969 3353 3088 3395
rect 2969 3319 3001 3353
rect 3035 3319 3088 3353
rect 2969 3311 3088 3319
rect 3118 3311 3179 3395
rect 3209 3373 3261 3395
rect 3209 3339 3219 3373
rect 3253 3339 3261 3373
rect 3209 3311 3261 3339
rect 3315 3357 3387 3395
rect 3315 3323 3343 3357
rect 3377 3323 3387 3357
rect 3315 3311 3387 3323
rect 3417 3407 3469 3441
rect 3417 3373 3427 3407
rect 3461 3373 3469 3407
rect 3417 3311 3469 3373
rect 3799 3376 3851 3421
rect 3799 3342 3807 3376
rect 3841 3342 3851 3376
rect 3799 3311 3851 3342
rect 4429 3376 4481 3421
rect 4429 3342 4439 3376
rect 4473 3342 4481 3376
rect 4429 3311 4481 3342
rect 4552 3361 4605 3395
rect 4552 3327 4560 3361
rect 4594 3327 4605 3361
rect 4552 3311 4605 3327
rect 4635 3370 4691 3395
rect 4635 3336 4646 3370
rect 4680 3336 4691 3370
rect 4635 3311 4691 3336
rect 4721 3361 4777 3395
rect 4721 3327 4732 3361
rect 4766 3327 4777 3361
rect 4721 3311 4777 3327
rect 4807 3370 4863 3395
rect 4807 3336 4818 3370
rect 4852 3336 4863 3370
rect 4807 3311 4863 3336
rect 4893 3361 4949 3395
rect 4893 3327 4904 3361
rect 4938 3327 4949 3361
rect 4893 3311 4949 3327
rect 4979 3370 5035 3395
rect 4979 3336 4990 3370
rect 5024 3336 5035 3370
rect 4979 3311 5035 3336
rect 5065 3361 5121 3395
rect 5065 3327 5076 3361
rect 5110 3327 5121 3361
rect 5065 3311 5121 3327
rect 5151 3370 5207 3395
rect 5151 3336 5162 3370
rect 5196 3336 5207 3370
rect 5151 3311 5207 3336
rect 5237 3361 5292 3395
rect 5237 3327 5247 3361
rect 5281 3327 5292 3361
rect 5237 3311 5292 3327
rect 5322 3370 5378 3395
rect 5322 3336 5333 3370
rect 5367 3336 5378 3370
rect 5322 3311 5378 3336
rect 5408 3361 5464 3395
rect 5408 3327 5419 3361
rect 5453 3327 5464 3361
rect 5408 3311 5464 3327
rect 5494 3370 5550 3395
rect 5494 3336 5505 3370
rect 5539 3336 5550 3370
rect 5494 3311 5550 3336
rect 5580 3361 5636 3395
rect 5580 3327 5591 3361
rect 5625 3327 5636 3361
rect 5580 3311 5636 3327
rect 5666 3370 5722 3395
rect 5666 3336 5677 3370
rect 5711 3336 5722 3370
rect 5666 3311 5722 3336
rect 5752 3361 5808 3395
rect 5752 3327 5763 3361
rect 5797 3327 5808 3361
rect 5752 3311 5808 3327
rect 5838 3370 5894 3395
rect 5838 3336 5849 3370
rect 5883 3336 5894 3370
rect 5838 3311 5894 3336
rect 5924 3370 5980 3395
rect 5924 3336 5935 3370
rect 5969 3336 5980 3370
rect 5924 3311 5980 3336
rect 6010 3370 6066 3395
rect 6010 3336 6021 3370
rect 6055 3336 6066 3370
rect 6010 3311 6066 3336
rect 6096 3370 6152 3395
rect 6096 3336 6107 3370
rect 6141 3336 6152 3370
rect 6096 3311 6152 3336
rect 6182 3370 6238 3395
rect 6182 3336 6193 3370
rect 6227 3336 6238 3370
rect 6182 3311 6238 3336
rect 6268 3357 6321 3395
rect 6268 3323 6279 3357
rect 6313 3323 6321 3357
rect 6268 3311 6321 3323
rect 6375 3383 6427 3421
rect 6375 3349 6383 3383
rect 6417 3349 6427 3383
rect 6375 3311 6427 3349
rect 6637 3383 6689 3421
rect 6637 3349 6647 3383
rect 6681 3349 6689 3383
rect 6637 3311 6689 3349
rect 6743 3383 6795 3395
rect 6743 3349 6751 3383
rect 6785 3349 6795 3383
rect 6743 3311 6795 3349
rect 6825 3357 6879 3395
rect 6825 3323 6835 3357
rect 6869 3323 6879 3357
rect 6825 3311 6879 3323
rect 6909 3383 6961 3395
rect 6909 3349 6919 3383
rect 6953 3349 6961 3383
rect 6909 3311 6961 3349
rect 7029 3353 7134 3395
rect 7029 3319 7041 3353
rect 7075 3319 7134 3353
rect 7029 3311 7134 3319
rect 7164 3383 7214 3395
rect 7645 3395 7695 3439
rect 7373 3383 7491 3395
rect 7164 3359 7229 3383
rect 7164 3325 7174 3359
rect 7208 3325 7229 3359
rect 7164 3311 7229 3325
rect 7259 3359 7325 3383
rect 7259 3325 7281 3359
rect 7315 3325 7325 3359
rect 7259 3311 7325 3325
rect 7355 3311 7491 3383
rect 7521 3311 7563 3395
rect 7593 3357 7695 3395
rect 7593 3323 7627 3357
rect 7661 3323 7695 3357
rect 7593 3311 7695 3323
rect 7725 3383 7779 3439
rect 8397 3395 8447 3441
rect 7949 3383 7999 3395
rect 7725 3353 7794 3383
rect 7725 3319 7739 3353
rect 7773 3319 7794 3353
rect 7725 3311 7794 3319
rect 7824 3357 7903 3383
rect 7824 3323 7849 3357
rect 7883 3323 7903 3357
rect 7824 3311 7903 3323
rect 7933 3311 7999 3383
rect 8029 3353 8148 3395
rect 8029 3319 8061 3353
rect 8095 3319 8148 3353
rect 8029 3311 8148 3319
rect 8178 3311 8239 3395
rect 8269 3373 8321 3395
rect 8269 3339 8279 3373
rect 8313 3339 8321 3373
rect 8269 3311 8321 3339
rect 8375 3357 8447 3395
rect 8375 3323 8403 3357
rect 8437 3323 8447 3357
rect 8375 3311 8447 3323
rect 8477 3407 8529 3441
rect 8477 3373 8487 3407
rect 8521 3373 8529 3407
rect 8477 3311 8529 3373
rect 8583 3378 8635 3421
rect 8583 3344 8591 3378
rect 8625 3344 8635 3378
rect 8583 3311 8635 3344
rect 8753 3378 8805 3421
rect 8753 3344 8763 3378
rect 8797 3344 8805 3378
rect 8753 3311 8805 3344
rect 9232 3395 9282 3441
rect 9135 3370 9187 3395
rect 9135 3336 9143 3370
rect 9177 3336 9187 3370
rect 9135 3311 9187 3336
rect 9217 3357 9282 3395
rect 9217 3323 9236 3357
rect 9270 3323 9282 3357
rect 9217 3311 9282 3323
rect 9312 3387 9366 3441
rect 9312 3353 9322 3387
rect 9356 3353 9366 3387
rect 9312 3311 9366 3353
rect 9396 3429 9449 3441
rect 9396 3395 9406 3429
rect 9440 3395 9449 3429
rect 9396 3361 9449 3395
rect 9396 3327 9406 3361
rect 9440 3327 9449 3361
rect 9396 3311 9449 3327
rect 9503 3376 9555 3421
rect 9503 3342 9511 3376
rect 9545 3342 9555 3376
rect 9503 3311 9555 3342
rect 9949 3376 10001 3421
rect 9949 3342 9959 3376
rect 9993 3342 10001 3376
rect 9949 3311 10001 3342
rect 10055 3387 10107 3415
rect 10055 3353 10063 3387
rect 10097 3353 10107 3387
rect 10055 3311 10107 3353
rect 10137 3357 10195 3415
rect 10137 3323 10149 3357
rect 10183 3323 10195 3357
rect 10137 3311 10195 3323
rect 10225 3370 10277 3415
rect 10225 3336 10235 3370
rect 10269 3336 10277 3370
rect 10225 3311 10277 3336
rect 10331 3376 10383 3421
rect 10331 3342 10339 3376
rect 10373 3342 10383 3376
rect 10331 3311 10383 3342
rect 10777 3376 10829 3421
rect 10777 3342 10787 3376
rect 10821 3342 10829 3376
rect 10777 3311 10829 3342
rect 10975 3370 11027 3415
rect 10975 3336 10983 3370
rect 11017 3336 11027 3370
rect 10975 3311 11027 3336
rect 11057 3357 11115 3415
rect 11057 3323 11069 3357
rect 11103 3323 11115 3357
rect 11057 3311 11115 3323
rect 11145 3387 11197 3415
rect 11145 3353 11155 3387
rect 11189 3353 11197 3387
rect 11145 3311 11197 3353
rect 11251 3376 11303 3421
rect 11251 3342 11259 3376
rect 11293 3342 11303 3376
rect 11251 3311 11303 3342
rect 11881 3376 11933 3421
rect 11881 3342 11891 3376
rect 11925 3342 11933 3376
rect 11881 3311 11933 3342
rect 11987 3407 12039 3441
rect 11987 3373 11995 3407
rect 12029 3373 12039 3407
rect 11987 3311 12039 3373
rect 12069 3395 12119 3441
rect 12069 3357 12141 3395
rect 12069 3323 12079 3357
rect 12113 3323 12141 3357
rect 12069 3311 12141 3323
rect 12195 3373 12247 3395
rect 12195 3339 12203 3373
rect 12237 3339 12247 3373
rect 12195 3311 12247 3339
rect 12277 3311 12338 3395
rect 12368 3353 12487 3395
rect 12368 3319 12421 3353
rect 12455 3319 12487 3353
rect 12368 3311 12487 3319
rect 12517 3383 12567 3395
rect 12737 3383 12791 3439
rect 12517 3311 12583 3383
rect 12613 3357 12692 3383
rect 12613 3323 12633 3357
rect 12667 3323 12692 3357
rect 12613 3311 12692 3323
rect 12722 3353 12791 3383
rect 12722 3319 12743 3353
rect 12777 3319 12791 3353
rect 12722 3311 12791 3319
rect 12821 3395 12871 3439
rect 12821 3357 12923 3395
rect 12821 3323 12855 3357
rect 12889 3323 12923 3357
rect 12821 3311 12923 3323
rect 12953 3311 12995 3395
rect 13025 3383 13143 3395
rect 13302 3383 13352 3395
rect 13025 3311 13161 3383
rect 13191 3359 13257 3383
rect 13191 3325 13201 3359
rect 13235 3325 13257 3359
rect 13191 3311 13257 3325
rect 13287 3359 13352 3383
rect 13287 3325 13308 3359
rect 13342 3325 13352 3359
rect 13287 3311 13352 3325
rect 13382 3353 13487 3395
rect 13382 3319 13441 3353
rect 13475 3319 13487 3353
rect 13382 3311 13487 3319
rect 13555 3383 13607 3395
rect 13555 3349 13563 3383
rect 13597 3349 13607 3383
rect 13555 3311 13607 3349
rect 13637 3357 13691 3395
rect 13637 3323 13647 3357
rect 13681 3323 13691 3357
rect 13637 3311 13691 3323
rect 13721 3383 13773 3395
rect 13721 3349 13731 3383
rect 13765 3349 13773 3383
rect 13721 3311 13773 3349
rect 14103 3376 14155 3421
rect 14103 3342 14111 3376
rect 14145 3342 14155 3376
rect 14103 3311 14155 3342
rect 15101 3376 15153 3421
rect 15101 3342 15111 3376
rect 15145 3342 15153 3376
rect 15101 3311 15153 3342
rect 15207 3376 15259 3421
rect 15207 3342 15215 3376
rect 15249 3342 15259 3376
rect 15207 3311 15259 3342
rect 16205 3376 16257 3421
rect 16205 3342 16215 3376
rect 16249 3342 16257 3376
rect 16205 3311 16257 3342
rect 16311 3376 16363 3421
rect 16311 3342 16319 3376
rect 16353 3342 16363 3376
rect 16311 3311 16363 3342
rect 17309 3376 17361 3421
rect 17309 3342 17319 3376
rect 17353 3342 17361 3376
rect 17309 3311 17361 3342
rect 17415 3376 17467 3421
rect 17415 3342 17423 3376
rect 17457 3342 17467 3376
rect 17415 3311 17467 3342
rect 18413 3376 18465 3421
rect 18413 3342 18423 3376
rect 18457 3342 18465 3376
rect 18413 3311 18465 3342
rect 18611 3378 18663 3421
rect 18611 3344 18619 3378
rect 18653 3344 18663 3378
rect 18611 3311 18663 3344
rect 18781 3378 18833 3421
rect 18781 3344 18791 3378
rect 18825 3344 18833 3378
rect 18781 3311 18833 3344
rect 1131 3184 1183 3217
rect 1131 3150 1139 3184
rect 1173 3150 1183 3184
rect 1131 3107 1183 3150
rect 1301 3184 1353 3217
rect 1301 3150 1311 3184
rect 1345 3150 1353 3184
rect 1301 3107 1353 3150
rect 1407 3186 1459 3217
rect 1407 3152 1415 3186
rect 1449 3152 1459 3186
rect 1407 3107 1459 3152
rect 1853 3186 1905 3217
rect 1853 3152 1863 3186
rect 1897 3152 1905 3186
rect 1853 3107 1905 3152
rect 1959 3155 2011 3217
rect 1959 3121 1967 3155
rect 2001 3121 2011 3155
rect 1959 3087 2011 3121
rect 2041 3205 2113 3217
rect 2041 3171 2051 3205
rect 2085 3171 2113 3205
rect 2041 3133 2113 3171
rect 2167 3189 2219 3217
rect 2167 3155 2175 3189
rect 2209 3155 2219 3189
rect 2167 3133 2219 3155
rect 2249 3133 2310 3217
rect 2340 3209 2459 3217
rect 2340 3175 2393 3209
rect 2427 3175 2459 3209
rect 2340 3133 2459 3175
rect 2489 3145 2555 3217
rect 2585 3205 2664 3217
rect 2585 3171 2605 3205
rect 2639 3171 2664 3205
rect 2585 3145 2664 3171
rect 2694 3209 2763 3217
rect 2694 3175 2715 3209
rect 2749 3175 2763 3209
rect 2694 3145 2763 3175
rect 2489 3133 2539 3145
rect 2041 3087 2091 3133
rect 2709 3089 2763 3145
rect 2793 3205 2895 3217
rect 2793 3171 2827 3205
rect 2861 3171 2895 3205
rect 2793 3133 2895 3171
rect 2925 3133 2967 3217
rect 2997 3145 3133 3217
rect 3163 3203 3229 3217
rect 3163 3169 3173 3203
rect 3207 3169 3229 3203
rect 3163 3145 3229 3169
rect 3259 3203 3324 3217
rect 3259 3169 3280 3203
rect 3314 3169 3324 3203
rect 3259 3145 3324 3169
rect 2997 3133 3115 3145
rect 2793 3089 2843 3133
rect 3274 3133 3324 3145
rect 3354 3209 3459 3217
rect 3354 3175 3413 3209
rect 3447 3175 3459 3209
rect 3354 3133 3459 3175
rect 3527 3179 3579 3217
rect 3527 3145 3535 3179
rect 3569 3145 3579 3179
rect 3527 3133 3579 3145
rect 3609 3205 3663 3217
rect 3609 3171 3619 3205
rect 3653 3171 3663 3205
rect 3609 3133 3663 3171
rect 3693 3179 3745 3217
rect 3693 3145 3703 3179
rect 3737 3145 3745 3179
rect 3693 3133 3745 3145
rect 3799 3179 3851 3217
rect 3799 3145 3807 3179
rect 3841 3145 3851 3179
rect 3799 3107 3851 3145
rect 4061 3179 4113 3217
rect 4061 3145 4071 3179
rect 4105 3145 4113 3179
rect 4061 3107 4113 3145
rect 4167 3179 4219 3217
rect 4167 3145 4175 3179
rect 4209 3145 4219 3179
rect 4167 3133 4219 3145
rect 4249 3205 4303 3217
rect 4249 3171 4259 3205
rect 4293 3171 4303 3205
rect 4249 3133 4303 3171
rect 4333 3179 4385 3217
rect 4333 3145 4343 3179
rect 4377 3145 4385 3179
rect 4333 3133 4385 3145
rect 4439 3205 4491 3217
rect 4439 3171 4447 3205
rect 4481 3171 4491 3205
rect 4439 3089 4491 3171
rect 4521 3187 4586 3217
rect 4521 3153 4531 3187
rect 4565 3153 4586 3187
rect 4521 3145 4586 3153
rect 4616 3205 4696 3217
rect 4616 3171 4641 3205
rect 4675 3171 4696 3205
rect 4616 3145 4696 3171
rect 4726 3145 4792 3217
rect 4521 3089 4571 3145
rect 4741 3133 4792 3145
rect 4822 3209 4906 3217
rect 4822 3175 4862 3209
rect 4896 3175 4906 3209
rect 4822 3133 4906 3175
rect 4936 3133 4978 3217
rect 5008 3189 5060 3217
rect 5008 3155 5018 3189
rect 5052 3155 5060 3189
rect 5008 3133 5060 3155
rect 5114 3205 5166 3217
rect 5114 3171 5122 3205
rect 5156 3171 5166 3205
rect 5114 3133 5166 3171
rect 5196 3133 5238 3217
rect 5268 3203 5334 3217
rect 5268 3169 5284 3203
rect 5318 3169 5334 3203
rect 5268 3133 5334 3169
rect 5364 3133 5406 3217
rect 5436 3133 5482 3217
rect 5512 3185 5606 3217
rect 5512 3151 5542 3185
rect 5576 3151 5606 3185
rect 5512 3133 5606 3151
rect 5556 3109 5606 3133
rect 5636 3178 5688 3217
rect 5636 3144 5646 3178
rect 5680 3144 5688 3178
rect 5636 3109 5688 3144
rect 5742 3179 5794 3217
rect 5742 3145 5750 3179
rect 5784 3145 5794 3179
rect 5742 3133 5794 3145
rect 5824 3205 5889 3217
rect 5824 3171 5845 3205
rect 5879 3171 5889 3205
rect 5824 3133 5889 3171
rect 5839 3087 5889 3133
rect 5919 3155 5971 3217
rect 5919 3121 5929 3155
rect 5963 3121 5971 3155
rect 5919 3087 5971 3121
rect 6375 3186 6427 3217
rect 6375 3152 6383 3186
rect 6417 3152 6427 3186
rect 6375 3107 6427 3152
rect 7005 3186 7057 3217
rect 7005 3152 7015 3186
rect 7049 3152 7057 3186
rect 7005 3107 7057 3152
rect 7203 3155 7255 3217
rect 7203 3121 7211 3155
rect 7245 3121 7255 3155
rect 7203 3087 7255 3121
rect 7285 3205 7357 3217
rect 7285 3171 7295 3205
rect 7329 3171 7357 3205
rect 7285 3133 7357 3171
rect 7411 3189 7463 3217
rect 7411 3155 7419 3189
rect 7453 3155 7463 3189
rect 7411 3133 7463 3155
rect 7493 3133 7554 3217
rect 7584 3209 7703 3217
rect 7584 3175 7637 3209
rect 7671 3175 7703 3209
rect 7584 3133 7703 3175
rect 7733 3145 7799 3217
rect 7829 3205 7908 3217
rect 7829 3171 7849 3205
rect 7883 3171 7908 3205
rect 7829 3145 7908 3171
rect 7938 3209 8007 3217
rect 7938 3175 7959 3209
rect 7993 3175 8007 3209
rect 7938 3145 8007 3175
rect 7733 3133 7783 3145
rect 7285 3087 7335 3133
rect 7953 3089 8007 3145
rect 8037 3205 8139 3217
rect 8037 3171 8071 3205
rect 8105 3171 8139 3205
rect 8037 3133 8139 3171
rect 8169 3133 8211 3217
rect 8241 3145 8377 3217
rect 8407 3203 8473 3217
rect 8407 3169 8417 3203
rect 8451 3169 8473 3203
rect 8407 3145 8473 3169
rect 8503 3203 8568 3217
rect 8503 3169 8524 3203
rect 8558 3169 8568 3203
rect 8503 3145 8568 3169
rect 8241 3133 8359 3145
rect 8037 3089 8087 3133
rect 8518 3133 8568 3145
rect 8598 3209 8703 3217
rect 8598 3175 8657 3209
rect 8691 3175 8703 3209
rect 8598 3133 8703 3175
rect 8771 3179 8823 3217
rect 8771 3145 8779 3179
rect 8813 3145 8823 3179
rect 8771 3133 8823 3145
rect 8853 3205 8907 3217
rect 8853 3171 8863 3205
rect 8897 3171 8907 3205
rect 8853 3133 8907 3171
rect 8937 3179 8989 3217
rect 8937 3145 8947 3179
rect 8981 3145 8989 3179
rect 8937 3133 8989 3145
rect 9043 3179 9095 3217
rect 9043 3145 9051 3179
rect 9085 3145 9095 3179
rect 9043 3107 9095 3145
rect 9305 3179 9357 3217
rect 9305 3145 9315 3179
rect 9349 3145 9357 3179
rect 9305 3107 9357 3145
rect 9411 3205 9464 3217
rect 9411 3171 9419 3205
rect 9453 3171 9464 3205
rect 9411 3133 9464 3171
rect 9494 3192 9550 3217
rect 9494 3158 9505 3192
rect 9539 3158 9550 3192
rect 9494 3133 9550 3158
rect 9580 3192 9636 3217
rect 9580 3158 9591 3192
rect 9625 3158 9636 3192
rect 9580 3133 9636 3158
rect 9666 3192 9722 3217
rect 9666 3158 9677 3192
rect 9711 3158 9722 3192
rect 9666 3133 9722 3158
rect 9752 3192 9808 3217
rect 9752 3158 9763 3192
rect 9797 3158 9808 3192
rect 9752 3133 9808 3158
rect 9838 3192 9894 3217
rect 9838 3158 9849 3192
rect 9883 3158 9894 3192
rect 9838 3133 9894 3158
rect 9924 3201 9980 3217
rect 9924 3167 9935 3201
rect 9969 3167 9980 3201
rect 9924 3133 9980 3167
rect 10010 3192 10066 3217
rect 10010 3158 10021 3192
rect 10055 3158 10066 3192
rect 10010 3133 10066 3158
rect 10096 3201 10152 3217
rect 10096 3167 10107 3201
rect 10141 3167 10152 3201
rect 10096 3133 10152 3167
rect 10182 3192 10238 3217
rect 10182 3158 10193 3192
rect 10227 3158 10238 3192
rect 10182 3133 10238 3158
rect 10268 3201 10324 3217
rect 10268 3167 10279 3201
rect 10313 3167 10324 3201
rect 10268 3133 10324 3167
rect 10354 3192 10410 3217
rect 10354 3158 10365 3192
rect 10399 3158 10410 3192
rect 10354 3133 10410 3158
rect 10440 3201 10495 3217
rect 10440 3167 10451 3201
rect 10485 3167 10495 3201
rect 10440 3133 10495 3167
rect 10525 3192 10581 3217
rect 10525 3158 10536 3192
rect 10570 3158 10581 3192
rect 10525 3133 10581 3158
rect 10611 3201 10667 3217
rect 10611 3167 10622 3201
rect 10656 3167 10667 3201
rect 10611 3133 10667 3167
rect 10697 3192 10753 3217
rect 10697 3158 10708 3192
rect 10742 3158 10753 3192
rect 10697 3133 10753 3158
rect 10783 3201 10839 3217
rect 10783 3167 10794 3201
rect 10828 3167 10839 3201
rect 10783 3133 10839 3167
rect 10869 3192 10925 3217
rect 10869 3158 10880 3192
rect 10914 3158 10925 3192
rect 10869 3133 10925 3158
rect 10955 3201 11011 3217
rect 10955 3167 10966 3201
rect 11000 3167 11011 3201
rect 10955 3133 11011 3167
rect 11041 3192 11097 3217
rect 11041 3158 11052 3192
rect 11086 3158 11097 3192
rect 11041 3133 11097 3158
rect 11127 3201 11180 3217
rect 11127 3167 11138 3201
rect 11172 3167 11180 3201
rect 11127 3133 11180 3167
rect 11711 3155 11763 3217
rect 11711 3121 11719 3155
rect 11753 3121 11763 3155
rect 11711 3087 11763 3121
rect 11793 3205 11865 3217
rect 11793 3171 11803 3205
rect 11837 3171 11865 3205
rect 11793 3133 11865 3171
rect 11919 3189 11971 3217
rect 11919 3155 11927 3189
rect 11961 3155 11971 3189
rect 11919 3133 11971 3155
rect 12001 3133 12062 3217
rect 12092 3209 12211 3217
rect 12092 3175 12145 3209
rect 12179 3175 12211 3209
rect 12092 3133 12211 3175
rect 12241 3145 12307 3217
rect 12337 3205 12416 3217
rect 12337 3171 12357 3205
rect 12391 3171 12416 3205
rect 12337 3145 12416 3171
rect 12446 3209 12515 3217
rect 12446 3175 12467 3209
rect 12501 3175 12515 3209
rect 12446 3145 12515 3175
rect 12241 3133 12291 3145
rect 11793 3087 11843 3133
rect 12461 3089 12515 3145
rect 12545 3205 12647 3217
rect 12545 3171 12579 3205
rect 12613 3171 12647 3205
rect 12545 3133 12647 3171
rect 12677 3133 12719 3217
rect 12749 3145 12885 3217
rect 12915 3203 12981 3217
rect 12915 3169 12925 3203
rect 12959 3169 12981 3203
rect 12915 3145 12981 3169
rect 13011 3203 13076 3217
rect 13011 3169 13032 3203
rect 13066 3169 13076 3203
rect 13011 3145 13076 3169
rect 12749 3133 12867 3145
rect 12545 3089 12595 3133
rect 13026 3133 13076 3145
rect 13106 3209 13211 3217
rect 13106 3175 13165 3209
rect 13199 3175 13211 3209
rect 13106 3133 13211 3175
rect 13279 3179 13331 3217
rect 13279 3145 13287 3179
rect 13321 3145 13331 3179
rect 13279 3133 13331 3145
rect 13361 3205 13415 3217
rect 13361 3171 13371 3205
rect 13405 3171 13415 3205
rect 13361 3133 13415 3171
rect 13445 3179 13497 3217
rect 13445 3145 13455 3179
rect 13489 3145 13497 3179
rect 13445 3133 13497 3145
rect 13551 3179 13603 3217
rect 13551 3145 13559 3179
rect 13593 3145 13603 3179
rect 13551 3107 13603 3145
rect 13813 3179 13865 3217
rect 13813 3145 13823 3179
rect 13857 3145 13865 3179
rect 13813 3107 13865 3145
rect 13919 3192 13971 3217
rect 13919 3158 13927 3192
rect 13961 3158 13971 3192
rect 13919 3133 13971 3158
rect 14001 3205 14066 3217
rect 14001 3171 14020 3205
rect 14054 3171 14066 3205
rect 14001 3133 14066 3171
rect 14016 3087 14066 3133
rect 14096 3175 14150 3217
rect 14096 3141 14106 3175
rect 14140 3141 14150 3175
rect 14096 3087 14150 3141
rect 14180 3201 14233 3217
rect 14180 3167 14190 3201
rect 14224 3167 14233 3201
rect 14180 3133 14233 3167
rect 14180 3099 14190 3133
rect 14224 3099 14233 3133
rect 14287 3186 14339 3217
rect 14287 3152 14295 3186
rect 14329 3152 14339 3186
rect 14287 3107 14339 3152
rect 15285 3186 15337 3217
rect 15285 3152 15295 3186
rect 15329 3152 15337 3186
rect 15285 3107 15337 3152
rect 15391 3186 15443 3217
rect 15391 3152 15399 3186
rect 15433 3152 15443 3186
rect 15391 3107 15443 3152
rect 16389 3186 16441 3217
rect 16389 3152 16399 3186
rect 16433 3152 16441 3186
rect 16389 3107 16441 3152
rect 14180 3087 14233 3099
rect 16679 3186 16731 3217
rect 16679 3152 16687 3186
rect 16721 3152 16731 3186
rect 16679 3107 16731 3152
rect 17677 3186 17729 3217
rect 17677 3152 17687 3186
rect 17721 3152 17729 3186
rect 17677 3107 17729 3152
rect 17783 3186 17835 3217
rect 17783 3152 17791 3186
rect 17825 3152 17835 3186
rect 17783 3107 17835 3152
rect 18413 3186 18465 3217
rect 18413 3152 18423 3186
rect 18457 3152 18465 3186
rect 18413 3107 18465 3152
rect 18611 3184 18663 3217
rect 18611 3150 18619 3184
rect 18653 3150 18663 3184
rect 18611 3107 18663 3150
rect 18781 3184 18833 3217
rect 18781 3150 18791 3184
rect 18825 3150 18833 3184
rect 18781 3107 18833 3150
rect 1131 2290 1183 2333
rect 1131 2256 1139 2290
rect 1173 2256 1183 2290
rect 1131 2223 1183 2256
rect 1301 2290 1353 2333
rect 1301 2256 1311 2290
rect 1345 2256 1353 2290
rect 1301 2223 1353 2256
rect 1407 2290 1459 2333
rect 1407 2256 1415 2290
rect 1449 2256 1459 2290
rect 1407 2223 1459 2256
rect 1577 2290 1629 2333
rect 1577 2256 1587 2290
rect 1621 2256 1629 2290
rect 1577 2223 1629 2256
rect 1683 2295 1735 2307
rect 1683 2261 1691 2295
rect 1725 2261 1735 2295
rect 1683 2223 1735 2261
rect 1765 2269 1819 2307
rect 1765 2235 1775 2269
rect 1809 2235 1819 2269
rect 1765 2223 1819 2235
rect 1849 2295 1901 2307
rect 1849 2261 1859 2295
rect 1893 2261 1901 2295
rect 1849 2223 1901 2261
rect 1969 2265 2074 2307
rect 1969 2231 1981 2265
rect 2015 2231 2074 2265
rect 1969 2223 2074 2231
rect 2104 2295 2154 2307
rect 2585 2307 2635 2351
rect 2313 2295 2431 2307
rect 2104 2271 2169 2295
rect 2104 2237 2114 2271
rect 2148 2237 2169 2271
rect 2104 2223 2169 2237
rect 2199 2271 2265 2295
rect 2199 2237 2221 2271
rect 2255 2237 2265 2271
rect 2199 2223 2265 2237
rect 2295 2223 2431 2295
rect 2461 2223 2503 2307
rect 2533 2269 2635 2307
rect 2533 2235 2567 2269
rect 2601 2235 2635 2269
rect 2533 2223 2635 2235
rect 2665 2295 2719 2351
rect 3337 2307 3387 2353
rect 2889 2295 2939 2307
rect 2665 2265 2734 2295
rect 2665 2231 2679 2265
rect 2713 2231 2734 2265
rect 2665 2223 2734 2231
rect 2764 2269 2843 2295
rect 2764 2235 2789 2269
rect 2823 2235 2843 2269
rect 2764 2223 2843 2235
rect 2873 2223 2939 2295
rect 2969 2265 3088 2307
rect 2969 2231 3001 2265
rect 3035 2231 3088 2265
rect 2969 2223 3088 2231
rect 3118 2223 3179 2307
rect 3209 2285 3261 2307
rect 3209 2251 3219 2285
rect 3253 2251 3261 2285
rect 3209 2223 3261 2251
rect 3315 2269 3387 2307
rect 3315 2235 3343 2269
rect 3377 2235 3387 2269
rect 3315 2223 3387 2235
rect 3417 2319 3469 2353
rect 3417 2285 3427 2319
rect 3461 2285 3469 2319
rect 3417 2223 3469 2285
rect 3799 2295 3851 2333
rect 3799 2261 3807 2295
rect 3841 2261 3851 2295
rect 3799 2223 3851 2261
rect 4061 2295 4113 2333
rect 4061 2261 4071 2295
rect 4105 2261 4113 2295
rect 4061 2223 4113 2261
rect 4259 2295 4311 2307
rect 4259 2261 4267 2295
rect 4301 2261 4311 2295
rect 4259 2223 4311 2261
rect 4341 2269 4395 2307
rect 4341 2235 4351 2269
rect 4385 2235 4395 2269
rect 4341 2223 4395 2235
rect 4425 2295 4477 2307
rect 4425 2261 4435 2295
rect 4469 2261 4477 2295
rect 4425 2223 4477 2261
rect 4545 2265 4650 2307
rect 4545 2231 4557 2265
rect 4591 2231 4650 2265
rect 4545 2223 4650 2231
rect 4680 2295 4730 2307
rect 5161 2307 5211 2351
rect 4889 2295 5007 2307
rect 4680 2271 4745 2295
rect 4680 2237 4690 2271
rect 4724 2237 4745 2271
rect 4680 2223 4745 2237
rect 4775 2271 4841 2295
rect 4775 2237 4797 2271
rect 4831 2237 4841 2271
rect 4775 2223 4841 2237
rect 4871 2223 5007 2295
rect 5037 2223 5079 2307
rect 5109 2269 5211 2307
rect 5109 2235 5143 2269
rect 5177 2235 5211 2269
rect 5109 2223 5211 2235
rect 5241 2295 5295 2351
rect 5913 2307 5963 2353
rect 5465 2295 5515 2307
rect 5241 2265 5310 2295
rect 5241 2231 5255 2265
rect 5289 2231 5310 2265
rect 5241 2223 5310 2231
rect 5340 2269 5419 2295
rect 5340 2235 5365 2269
rect 5399 2235 5419 2269
rect 5340 2223 5419 2235
rect 5449 2223 5515 2295
rect 5545 2265 5664 2307
rect 5545 2231 5577 2265
rect 5611 2231 5664 2265
rect 5545 2223 5664 2231
rect 5694 2223 5755 2307
rect 5785 2285 5837 2307
rect 5785 2251 5795 2285
rect 5829 2251 5837 2285
rect 5785 2223 5837 2251
rect 5891 2269 5963 2307
rect 5891 2235 5919 2269
rect 5953 2235 5963 2269
rect 5891 2223 5963 2235
rect 5993 2319 6045 2353
rect 5993 2285 6003 2319
rect 6037 2285 6045 2319
rect 5993 2223 6045 2285
rect 6375 2288 6427 2333
rect 6375 2254 6383 2288
rect 6417 2254 6427 2288
rect 6375 2223 6427 2254
rect 7373 2288 7425 2333
rect 7373 2254 7383 2288
rect 7417 2254 7425 2288
rect 7373 2223 7425 2254
rect 7479 2288 7531 2333
rect 7479 2254 7487 2288
rect 7521 2254 7531 2288
rect 7479 2223 7531 2254
rect 8477 2288 8529 2333
rect 8477 2254 8487 2288
rect 8521 2254 8529 2288
rect 8477 2223 8529 2254
rect 8583 2290 8635 2333
rect 8583 2256 8591 2290
rect 8625 2256 8635 2290
rect 8583 2223 8635 2256
rect 8753 2290 8805 2333
rect 8753 2256 8763 2290
rect 8797 2256 8805 2290
rect 8753 2223 8805 2256
rect 9135 2319 9187 2353
rect 9135 2285 9143 2319
rect 9177 2285 9187 2319
rect 9135 2223 9187 2285
rect 9217 2307 9267 2353
rect 9217 2269 9289 2307
rect 9217 2235 9227 2269
rect 9261 2235 9289 2269
rect 9217 2223 9289 2235
rect 9343 2285 9395 2307
rect 9343 2251 9351 2285
rect 9385 2251 9395 2285
rect 9343 2223 9395 2251
rect 9425 2223 9486 2307
rect 9516 2265 9635 2307
rect 9516 2231 9569 2265
rect 9603 2231 9635 2265
rect 9516 2223 9635 2231
rect 9665 2295 9715 2307
rect 9885 2295 9939 2351
rect 9665 2223 9731 2295
rect 9761 2269 9840 2295
rect 9761 2235 9781 2269
rect 9815 2235 9840 2269
rect 9761 2223 9840 2235
rect 9870 2265 9939 2295
rect 9870 2231 9891 2265
rect 9925 2231 9939 2265
rect 9870 2223 9939 2231
rect 9969 2307 10019 2351
rect 9969 2269 10071 2307
rect 9969 2235 10003 2269
rect 10037 2235 10071 2269
rect 9969 2223 10071 2235
rect 10101 2223 10143 2307
rect 10173 2295 10291 2307
rect 10450 2295 10500 2307
rect 10173 2223 10309 2295
rect 10339 2271 10405 2295
rect 10339 2237 10349 2271
rect 10383 2237 10405 2271
rect 10339 2223 10405 2237
rect 10435 2271 10500 2295
rect 10435 2237 10456 2271
rect 10490 2237 10500 2271
rect 10435 2223 10500 2237
rect 10530 2265 10635 2307
rect 10530 2231 10589 2265
rect 10623 2231 10635 2265
rect 10530 2223 10635 2231
rect 10703 2295 10755 2307
rect 10703 2261 10711 2295
rect 10745 2261 10755 2295
rect 10703 2223 10755 2261
rect 10785 2269 10839 2307
rect 10785 2235 10795 2269
rect 10829 2235 10839 2269
rect 10785 2223 10839 2235
rect 10869 2295 10921 2307
rect 10869 2261 10879 2295
rect 10913 2261 10921 2295
rect 10869 2223 10921 2261
rect 10975 2295 11027 2333
rect 10975 2261 10983 2295
rect 11017 2261 11027 2295
rect 10975 2223 11027 2261
rect 11237 2295 11289 2333
rect 11237 2261 11247 2295
rect 11281 2261 11289 2295
rect 11237 2223 11289 2261
rect 11527 2295 11579 2333
rect 11527 2261 11535 2295
rect 11569 2261 11579 2295
rect 11527 2223 11579 2261
rect 11789 2295 11841 2333
rect 11789 2261 11799 2295
rect 11833 2261 11841 2295
rect 11789 2223 11841 2261
rect 11987 2319 12039 2353
rect 11987 2285 11995 2319
rect 12029 2285 12039 2319
rect 11987 2223 12039 2285
rect 12069 2307 12119 2353
rect 12069 2269 12141 2307
rect 12069 2235 12079 2269
rect 12113 2235 12141 2269
rect 12069 2223 12141 2235
rect 12195 2285 12247 2307
rect 12195 2251 12203 2285
rect 12237 2251 12247 2285
rect 12195 2223 12247 2251
rect 12277 2223 12338 2307
rect 12368 2265 12487 2307
rect 12368 2231 12421 2265
rect 12455 2231 12487 2265
rect 12368 2223 12487 2231
rect 12517 2295 12567 2307
rect 12737 2295 12791 2351
rect 12517 2223 12583 2295
rect 12613 2269 12692 2295
rect 12613 2235 12633 2269
rect 12667 2235 12692 2269
rect 12613 2223 12692 2235
rect 12722 2265 12791 2295
rect 12722 2231 12743 2265
rect 12777 2231 12791 2265
rect 12722 2223 12791 2231
rect 12821 2307 12871 2351
rect 12821 2269 12923 2307
rect 12821 2235 12855 2269
rect 12889 2235 12923 2269
rect 12821 2223 12923 2235
rect 12953 2223 12995 2307
rect 13025 2295 13143 2307
rect 13302 2295 13352 2307
rect 13025 2223 13161 2295
rect 13191 2271 13257 2295
rect 13191 2237 13201 2271
rect 13235 2237 13257 2271
rect 13191 2223 13257 2237
rect 13287 2271 13352 2295
rect 13287 2237 13308 2271
rect 13342 2237 13352 2271
rect 13287 2223 13352 2237
rect 13382 2265 13487 2307
rect 13382 2231 13441 2265
rect 13475 2231 13487 2265
rect 13382 2223 13487 2231
rect 13555 2295 13607 2307
rect 13555 2261 13563 2295
rect 13597 2261 13607 2295
rect 13555 2223 13607 2261
rect 13637 2269 13691 2307
rect 13637 2235 13647 2269
rect 13681 2235 13691 2269
rect 13637 2223 13691 2235
rect 13721 2295 13773 2307
rect 13721 2261 13731 2295
rect 13765 2261 13773 2295
rect 13721 2223 13773 2261
rect 14287 2319 14339 2353
rect 14287 2285 14295 2319
rect 14329 2285 14339 2319
rect 14287 2223 14339 2285
rect 14369 2307 14419 2353
rect 14369 2269 14441 2307
rect 14369 2235 14379 2269
rect 14413 2235 14441 2269
rect 14369 2223 14441 2235
rect 14495 2285 14547 2307
rect 14495 2251 14503 2285
rect 14537 2251 14547 2285
rect 14495 2223 14547 2251
rect 14577 2223 14638 2307
rect 14668 2265 14787 2307
rect 14668 2231 14721 2265
rect 14755 2231 14787 2265
rect 14668 2223 14787 2231
rect 14817 2295 14867 2307
rect 15037 2295 15091 2351
rect 14817 2223 14883 2295
rect 14913 2269 14992 2295
rect 14913 2235 14933 2269
rect 14967 2235 14992 2269
rect 14913 2223 14992 2235
rect 15022 2265 15091 2295
rect 15022 2231 15043 2265
rect 15077 2231 15091 2265
rect 15022 2223 15091 2231
rect 15121 2307 15171 2351
rect 15121 2269 15223 2307
rect 15121 2235 15155 2269
rect 15189 2235 15223 2269
rect 15121 2223 15223 2235
rect 15253 2223 15295 2307
rect 15325 2295 15443 2307
rect 15602 2295 15652 2307
rect 15325 2223 15461 2295
rect 15491 2271 15557 2295
rect 15491 2237 15501 2271
rect 15535 2237 15557 2271
rect 15491 2223 15557 2237
rect 15587 2271 15652 2295
rect 15587 2237 15608 2271
rect 15642 2237 15652 2271
rect 15587 2223 15652 2237
rect 15682 2265 15787 2307
rect 15682 2231 15741 2265
rect 15775 2231 15787 2265
rect 15682 2223 15787 2231
rect 15855 2295 15907 2307
rect 15855 2261 15863 2295
rect 15897 2261 15907 2295
rect 15855 2223 15907 2261
rect 15937 2269 15991 2307
rect 15937 2235 15947 2269
rect 15981 2235 15991 2269
rect 15937 2223 15991 2235
rect 16021 2295 16073 2307
rect 16021 2261 16031 2295
rect 16065 2261 16073 2295
rect 16021 2223 16073 2261
rect 16127 2295 16179 2333
rect 16127 2261 16135 2295
rect 16169 2261 16179 2295
rect 16127 2223 16179 2261
rect 16389 2295 16441 2333
rect 16389 2261 16399 2295
rect 16433 2261 16441 2295
rect 16389 2223 16441 2261
rect 16679 2288 16731 2333
rect 16679 2254 16687 2288
rect 16721 2254 16731 2288
rect 16679 2223 16731 2254
rect 17309 2288 17361 2333
rect 17604 2307 17654 2353
rect 17309 2254 17319 2288
rect 17353 2254 17361 2288
rect 17309 2223 17361 2254
rect 17507 2282 17559 2307
rect 17507 2248 17515 2282
rect 17549 2248 17559 2282
rect 17507 2223 17559 2248
rect 17589 2269 17654 2307
rect 17589 2235 17608 2269
rect 17642 2235 17654 2269
rect 17589 2223 17654 2235
rect 17684 2299 17738 2353
rect 17684 2265 17694 2299
rect 17728 2265 17738 2299
rect 17684 2223 17738 2265
rect 17768 2341 17821 2353
rect 17768 2307 17778 2341
rect 17812 2307 17821 2341
rect 17768 2273 17821 2307
rect 17768 2239 17778 2273
rect 17812 2239 17821 2273
rect 17768 2223 17821 2239
rect 17875 2288 17927 2333
rect 17875 2254 17883 2288
rect 17917 2254 17927 2288
rect 17875 2223 17927 2254
rect 18505 2288 18557 2333
rect 18505 2254 18515 2288
rect 18549 2254 18557 2288
rect 18505 2223 18557 2254
rect 18611 2290 18663 2333
rect 18611 2256 18619 2290
rect 18653 2256 18663 2290
rect 18611 2223 18663 2256
rect 18781 2290 18833 2333
rect 18781 2256 18791 2290
rect 18825 2256 18833 2290
rect 18781 2223 18833 2256
<< pdiff >>
rect 1591 7301 1644 7319
rect 1131 7260 1183 7293
rect 1131 7226 1139 7260
rect 1173 7226 1183 7260
rect 1131 7165 1183 7226
rect 1131 7131 1139 7165
rect 1173 7131 1183 7165
rect 1131 7119 1183 7131
rect 1301 7260 1353 7293
rect 1301 7226 1311 7260
rect 1345 7226 1353 7260
rect 1301 7165 1353 7226
rect 1301 7131 1311 7165
rect 1345 7131 1353 7165
rect 1301 7119 1353 7131
rect 1591 7267 1600 7301
rect 1634 7267 1644 7301
rect 1591 7233 1644 7267
rect 1591 7199 1600 7233
rect 1634 7199 1644 7233
rect 1591 7165 1644 7199
rect 1591 7131 1600 7165
rect 1634 7131 1644 7165
rect 1591 7119 1644 7131
rect 1674 7270 1728 7319
rect 1674 7236 1684 7270
rect 1718 7236 1728 7270
rect 1674 7189 1728 7236
rect 1674 7155 1684 7189
rect 1718 7155 1728 7189
rect 1674 7119 1728 7155
rect 1758 7255 1808 7319
rect 1758 7241 1823 7255
rect 1758 7207 1770 7241
rect 1804 7207 1823 7241
rect 1758 7173 1823 7207
rect 1758 7139 1770 7173
rect 1804 7139 1823 7173
rect 1758 7127 1823 7139
rect 1853 7241 1905 7255
rect 1853 7207 1863 7241
rect 1897 7207 1905 7241
rect 1853 7173 1905 7207
rect 1853 7139 1863 7173
rect 1897 7139 1905 7173
rect 1853 7127 1905 7139
rect 1959 7165 2011 7293
rect 1959 7131 1967 7165
rect 2001 7131 2011 7165
rect 1758 7119 1808 7127
rect 1959 7119 2011 7131
rect 2957 7165 3009 7293
rect 2957 7131 2967 7165
rect 3001 7131 3009 7165
rect 2957 7119 3009 7131
rect 3063 7267 3115 7293
rect 3063 7233 3071 7267
rect 3105 7233 3115 7267
rect 3063 7165 3115 7233
rect 3063 7131 3071 7165
rect 3105 7131 3115 7165
rect 3063 7119 3115 7131
rect 3509 7267 3561 7293
rect 3509 7233 3519 7267
rect 3553 7233 3561 7267
rect 3509 7165 3561 7233
rect 3509 7131 3519 7165
rect 3553 7131 3561 7165
rect 3983 7301 4036 7319
rect 3983 7267 3992 7301
rect 4026 7267 4036 7301
rect 3983 7233 4036 7267
rect 3983 7199 3992 7233
rect 4026 7199 4036 7233
rect 3983 7165 4036 7199
rect 3509 7119 3561 7131
rect 3983 7131 3992 7165
rect 4026 7131 4036 7165
rect 3983 7119 4036 7131
rect 4066 7270 4120 7319
rect 4066 7236 4076 7270
rect 4110 7236 4120 7270
rect 4066 7189 4120 7236
rect 4066 7155 4076 7189
rect 4110 7155 4120 7189
rect 4066 7119 4120 7155
rect 4150 7255 4200 7319
rect 5639 7301 5692 7319
rect 4150 7241 4215 7255
rect 4150 7207 4162 7241
rect 4196 7207 4215 7241
rect 4150 7173 4215 7207
rect 4150 7139 4162 7173
rect 4196 7139 4215 7173
rect 4150 7127 4215 7139
rect 4245 7241 4297 7255
rect 4245 7207 4255 7241
rect 4289 7207 4297 7241
rect 4245 7173 4297 7207
rect 4245 7139 4255 7173
rect 4289 7139 4297 7173
rect 4245 7127 4297 7139
rect 4351 7165 4403 7293
rect 4351 7131 4359 7165
rect 4393 7131 4403 7165
rect 4150 7119 4200 7127
rect 4351 7119 4403 7131
rect 5349 7165 5401 7293
rect 5349 7131 5359 7165
rect 5393 7131 5401 7165
rect 5349 7119 5401 7131
rect 5639 7267 5648 7301
rect 5682 7267 5692 7301
rect 5639 7233 5692 7267
rect 5639 7199 5648 7233
rect 5682 7199 5692 7233
rect 5639 7165 5692 7199
rect 5639 7131 5648 7165
rect 5682 7131 5692 7165
rect 5639 7119 5692 7131
rect 5722 7270 5776 7319
rect 5722 7236 5732 7270
rect 5766 7236 5776 7270
rect 5722 7189 5776 7236
rect 5722 7155 5732 7189
rect 5766 7155 5776 7189
rect 5722 7119 5776 7155
rect 5806 7255 5856 7319
rect 6007 7260 6059 7293
rect 5806 7241 5871 7255
rect 5806 7207 5818 7241
rect 5852 7207 5871 7241
rect 5806 7173 5871 7207
rect 5806 7139 5818 7173
rect 5852 7139 5871 7173
rect 5806 7127 5871 7139
rect 5901 7241 5953 7255
rect 5901 7207 5911 7241
rect 5945 7207 5953 7241
rect 5901 7173 5953 7207
rect 5901 7139 5911 7173
rect 5945 7139 5953 7173
rect 5901 7127 5953 7139
rect 6007 7226 6015 7260
rect 6049 7226 6059 7260
rect 6007 7165 6059 7226
rect 6007 7131 6015 7165
rect 6049 7131 6059 7165
rect 5806 7119 5856 7127
rect 6007 7119 6059 7131
rect 6177 7260 6229 7293
rect 6177 7226 6187 7260
rect 6221 7226 6229 7260
rect 6177 7165 6229 7226
rect 6177 7131 6187 7165
rect 6221 7131 6229 7165
rect 7847 7301 7900 7319
rect 6375 7165 6427 7293
rect 6177 7119 6229 7131
rect 6375 7131 6383 7165
rect 6417 7131 6427 7165
rect 6375 7119 6427 7131
rect 7373 7165 7425 7293
rect 7373 7131 7383 7165
rect 7417 7131 7425 7165
rect 7373 7119 7425 7131
rect 7479 7267 7531 7293
rect 7479 7233 7487 7267
rect 7521 7233 7531 7267
rect 7479 7165 7531 7233
rect 7479 7131 7487 7165
rect 7521 7131 7531 7165
rect 7479 7119 7531 7131
rect 7741 7267 7793 7293
rect 7741 7233 7751 7267
rect 7785 7233 7793 7267
rect 7741 7165 7793 7233
rect 7741 7131 7751 7165
rect 7785 7131 7793 7165
rect 7741 7119 7793 7131
rect 7847 7267 7856 7301
rect 7890 7267 7900 7301
rect 7847 7233 7900 7267
rect 7847 7199 7856 7233
rect 7890 7199 7900 7233
rect 7847 7165 7900 7199
rect 7847 7131 7856 7165
rect 7890 7131 7900 7165
rect 7847 7119 7900 7131
rect 7930 7270 7984 7319
rect 7930 7236 7940 7270
rect 7974 7236 7984 7270
rect 7930 7189 7984 7236
rect 7930 7155 7940 7189
rect 7974 7155 7984 7189
rect 7930 7119 7984 7155
rect 8014 7255 8064 7319
rect 8215 7267 8267 7293
rect 8014 7241 8079 7255
rect 8014 7207 8026 7241
rect 8060 7207 8079 7241
rect 8014 7173 8079 7207
rect 8014 7139 8026 7173
rect 8060 7139 8079 7173
rect 8014 7127 8079 7139
rect 8109 7241 8161 7255
rect 8109 7207 8119 7241
rect 8153 7207 8161 7241
rect 8109 7173 8161 7207
rect 8109 7139 8119 7173
rect 8153 7139 8161 7173
rect 8109 7127 8161 7139
rect 8215 7233 8223 7267
rect 8257 7233 8267 7267
rect 8215 7165 8267 7233
rect 8215 7131 8223 7165
rect 8257 7131 8267 7165
rect 8014 7119 8064 7127
rect 8215 7119 8267 7131
rect 8661 7267 8713 7293
rect 8661 7233 8671 7267
rect 8705 7233 8713 7267
rect 8661 7165 8713 7233
rect 8661 7131 8671 7165
rect 8705 7131 8713 7165
rect 8951 7267 9003 7293
rect 8951 7233 8959 7267
rect 8993 7233 9003 7267
rect 8951 7165 9003 7233
rect 8661 7119 8713 7131
rect 8951 7131 8959 7165
rect 8993 7131 9003 7165
rect 8951 7119 9003 7131
rect 9397 7267 9449 7293
rect 9397 7233 9407 7267
rect 9441 7233 9449 7267
rect 9397 7165 9449 7233
rect 9397 7131 9407 7165
rect 9441 7131 9449 7165
rect 9397 7119 9449 7131
rect 9687 7267 9739 7293
rect 9687 7233 9695 7267
rect 9729 7233 9739 7267
rect 9687 7165 9739 7233
rect 9687 7131 9695 7165
rect 9729 7131 9739 7165
rect 9687 7119 9739 7131
rect 9949 7267 10001 7293
rect 9949 7233 9959 7267
rect 9993 7233 10001 7267
rect 9949 7165 10001 7233
rect 9949 7131 9959 7165
rect 9993 7131 10001 7165
rect 9949 7119 10001 7131
rect 10055 7284 10108 7319
rect 10055 7250 10063 7284
rect 10097 7250 10108 7284
rect 10055 7179 10108 7250
rect 10055 7145 10063 7179
rect 10097 7145 10108 7179
rect 10055 7119 10108 7145
rect 10138 7245 10203 7319
rect 10138 7211 10149 7245
rect 10183 7211 10203 7245
rect 10138 7177 10203 7211
rect 10138 7143 10149 7177
rect 10183 7143 10203 7177
rect 10138 7119 10203 7143
rect 10233 7179 10287 7319
rect 10233 7145 10243 7179
rect 10277 7145 10287 7179
rect 10233 7119 10287 7145
rect 10317 7174 10369 7319
rect 10317 7140 10327 7174
rect 10361 7140 10369 7174
rect 10317 7119 10369 7140
rect 10423 7267 10475 7293
rect 10423 7233 10431 7267
rect 10465 7233 10475 7267
rect 10423 7165 10475 7233
rect 10423 7131 10431 7165
rect 10465 7131 10475 7165
rect 10423 7119 10475 7131
rect 11053 7267 11105 7293
rect 11053 7233 11063 7267
rect 11097 7233 11105 7267
rect 11053 7165 11105 7233
rect 11053 7131 11063 7165
rect 11097 7131 11105 7165
rect 11053 7119 11105 7131
rect 11159 7260 11211 7293
rect 11159 7226 11167 7260
rect 11201 7226 11211 7260
rect 11159 7165 11211 7226
rect 11159 7131 11167 7165
rect 11201 7131 11211 7165
rect 11159 7119 11211 7131
rect 11329 7260 11381 7293
rect 11329 7226 11339 7260
rect 11373 7226 11381 7260
rect 11329 7165 11381 7226
rect 11329 7131 11339 7165
rect 11373 7131 11381 7165
rect 11527 7267 11579 7293
rect 11527 7233 11535 7267
rect 11569 7233 11579 7267
rect 11527 7165 11579 7233
rect 11329 7119 11381 7131
rect 11527 7131 11535 7165
rect 11569 7131 11579 7165
rect 11527 7119 11579 7131
rect 12157 7267 12209 7293
rect 12157 7233 12167 7267
rect 12201 7233 12209 7267
rect 12360 7255 12410 7319
rect 12157 7165 12209 7233
rect 12157 7131 12167 7165
rect 12201 7131 12209 7165
rect 12157 7119 12209 7131
rect 12263 7241 12315 7255
rect 12263 7207 12271 7241
rect 12305 7207 12315 7241
rect 12263 7173 12315 7207
rect 12263 7139 12271 7173
rect 12305 7139 12315 7173
rect 12263 7127 12315 7139
rect 12345 7241 12410 7255
rect 12345 7207 12364 7241
rect 12398 7207 12410 7241
rect 12345 7173 12410 7207
rect 12345 7139 12364 7173
rect 12398 7139 12410 7173
rect 12345 7127 12410 7139
rect 12360 7119 12410 7127
rect 12440 7270 12494 7319
rect 12440 7236 12450 7270
rect 12484 7236 12494 7270
rect 12440 7189 12494 7236
rect 12440 7155 12450 7189
rect 12484 7155 12494 7189
rect 12440 7119 12494 7155
rect 12524 7301 12577 7319
rect 12524 7267 12534 7301
rect 12568 7267 12577 7301
rect 12524 7233 12577 7267
rect 12524 7199 12534 7233
rect 12568 7199 12577 7233
rect 12524 7165 12577 7199
rect 12524 7131 12534 7165
rect 12568 7131 12577 7165
rect 12524 7119 12577 7131
rect 12631 7165 12683 7293
rect 12631 7131 12639 7165
rect 12673 7131 12683 7165
rect 12631 7119 12683 7131
rect 13629 7165 13681 7293
rect 13629 7131 13639 7165
rect 13673 7131 13681 7165
rect 13629 7119 13681 7131
rect 13735 7260 13787 7293
rect 13735 7226 13743 7260
rect 13777 7226 13787 7260
rect 13735 7165 13787 7226
rect 13735 7131 13743 7165
rect 13777 7131 13787 7165
rect 13735 7119 13787 7131
rect 13905 7260 13957 7293
rect 13905 7226 13915 7260
rect 13949 7226 13957 7260
rect 13905 7165 13957 7226
rect 13905 7131 13915 7165
rect 13949 7131 13957 7165
rect 14103 7267 14155 7293
rect 14103 7233 14111 7267
rect 14145 7233 14155 7267
rect 14103 7165 14155 7233
rect 13905 7119 13957 7131
rect 14103 7131 14111 7165
rect 14145 7131 14155 7165
rect 14103 7119 14155 7131
rect 14365 7267 14417 7293
rect 14365 7233 14375 7267
rect 14409 7233 14417 7267
rect 14568 7255 14618 7319
rect 14365 7165 14417 7233
rect 14365 7131 14375 7165
rect 14409 7131 14417 7165
rect 14365 7119 14417 7131
rect 14471 7241 14523 7255
rect 14471 7207 14479 7241
rect 14513 7207 14523 7241
rect 14471 7173 14523 7207
rect 14471 7139 14479 7173
rect 14513 7139 14523 7173
rect 14471 7127 14523 7139
rect 14553 7241 14618 7255
rect 14553 7207 14572 7241
rect 14606 7207 14618 7241
rect 14553 7173 14618 7207
rect 14553 7139 14572 7173
rect 14606 7139 14618 7173
rect 14553 7127 14618 7139
rect 14568 7119 14618 7127
rect 14648 7270 14702 7319
rect 14648 7236 14658 7270
rect 14692 7236 14702 7270
rect 14648 7189 14702 7236
rect 14648 7155 14658 7189
rect 14692 7155 14702 7189
rect 14648 7119 14702 7155
rect 14732 7301 14785 7319
rect 14732 7267 14742 7301
rect 14776 7267 14785 7301
rect 14732 7233 14785 7267
rect 14732 7199 14742 7233
rect 14776 7199 14785 7233
rect 14732 7165 14785 7199
rect 14732 7131 14742 7165
rect 14776 7131 14785 7165
rect 14732 7119 14785 7131
rect 14839 7165 14891 7293
rect 14839 7131 14847 7165
rect 14881 7131 14891 7165
rect 14839 7119 14891 7131
rect 15837 7165 15889 7293
rect 15837 7131 15847 7165
rect 15881 7131 15889 7165
rect 15837 7119 15889 7131
rect 15943 7267 15995 7293
rect 15943 7233 15951 7267
rect 15985 7233 15995 7267
rect 15943 7165 15995 7233
rect 15943 7131 15951 7165
rect 15985 7131 15995 7165
rect 15943 7119 15995 7131
rect 16389 7267 16441 7293
rect 16389 7233 16399 7267
rect 16433 7233 16441 7267
rect 16389 7165 16441 7233
rect 16389 7131 16399 7165
rect 16433 7131 16441 7165
rect 16960 7255 17010 7319
rect 16863 7241 16915 7255
rect 16863 7207 16871 7241
rect 16905 7207 16915 7241
rect 16863 7173 16915 7207
rect 16863 7139 16871 7173
rect 16905 7139 16915 7173
rect 16389 7119 16441 7131
rect 16863 7127 16915 7139
rect 16945 7241 17010 7255
rect 16945 7207 16964 7241
rect 16998 7207 17010 7241
rect 16945 7173 17010 7207
rect 16945 7139 16964 7173
rect 16998 7139 17010 7173
rect 16945 7127 17010 7139
rect 16960 7119 17010 7127
rect 17040 7270 17094 7319
rect 17040 7236 17050 7270
rect 17084 7236 17094 7270
rect 17040 7189 17094 7236
rect 17040 7155 17050 7189
rect 17084 7155 17094 7189
rect 17040 7119 17094 7155
rect 17124 7301 17177 7319
rect 17124 7267 17134 7301
rect 17168 7267 17177 7301
rect 17124 7233 17177 7267
rect 17124 7199 17134 7233
rect 17168 7199 17177 7233
rect 17124 7165 17177 7199
rect 17124 7131 17134 7165
rect 17168 7131 17177 7165
rect 17124 7119 17177 7131
rect 17231 7267 17283 7293
rect 17231 7233 17239 7267
rect 17273 7233 17283 7267
rect 17231 7165 17283 7233
rect 17231 7131 17239 7165
rect 17273 7131 17283 7165
rect 17231 7119 17283 7131
rect 17861 7267 17913 7293
rect 17861 7233 17871 7267
rect 17905 7233 17913 7267
rect 18156 7255 18206 7319
rect 17861 7165 17913 7233
rect 17861 7131 17871 7165
rect 17905 7131 17913 7165
rect 17861 7119 17913 7131
rect 18059 7241 18111 7255
rect 18059 7207 18067 7241
rect 18101 7207 18111 7241
rect 18059 7173 18111 7207
rect 18059 7139 18067 7173
rect 18101 7139 18111 7173
rect 18059 7127 18111 7139
rect 18141 7241 18206 7255
rect 18141 7207 18160 7241
rect 18194 7207 18206 7241
rect 18141 7173 18206 7207
rect 18141 7139 18160 7173
rect 18194 7139 18206 7173
rect 18141 7127 18206 7139
rect 18156 7119 18206 7127
rect 18236 7270 18290 7319
rect 18236 7236 18246 7270
rect 18280 7236 18290 7270
rect 18236 7189 18290 7236
rect 18236 7155 18246 7189
rect 18280 7155 18290 7189
rect 18236 7119 18290 7155
rect 18320 7301 18373 7319
rect 18320 7267 18330 7301
rect 18364 7267 18373 7301
rect 18320 7233 18373 7267
rect 18320 7199 18330 7233
rect 18364 7199 18373 7233
rect 18320 7165 18373 7199
rect 18320 7131 18330 7165
rect 18364 7131 18373 7165
rect 18320 7119 18373 7131
rect 18611 7260 18663 7293
rect 18611 7226 18619 7260
rect 18653 7226 18663 7260
rect 18611 7165 18663 7226
rect 18611 7131 18619 7165
rect 18653 7131 18663 7165
rect 18611 7119 18663 7131
rect 18781 7260 18833 7293
rect 18781 7226 18791 7260
rect 18825 7226 18833 7260
rect 18781 7165 18833 7226
rect 18781 7131 18791 7165
rect 18825 7131 18833 7165
rect 18781 7119 18833 7131
rect 1131 7013 1183 7025
rect 1131 6979 1139 7013
rect 1173 6979 1183 7013
rect 1131 6918 1183 6979
rect 1131 6884 1139 6918
rect 1173 6884 1183 6918
rect 1131 6851 1183 6884
rect 1301 7013 1353 7025
rect 1301 6979 1311 7013
rect 1345 6979 1353 7013
rect 1301 6918 1353 6979
rect 1301 6884 1311 6918
rect 1345 6884 1353 6918
rect 1301 6851 1353 6884
rect 1407 7013 1459 7025
rect 1407 6979 1415 7013
rect 1449 6979 1459 7013
rect 1407 6851 1459 6979
rect 2405 7013 2457 7025
rect 2405 6979 2415 7013
rect 2449 6979 2457 7013
rect 2405 6851 2457 6979
rect 2511 7013 2563 7025
rect 2511 6979 2519 7013
rect 2553 6979 2563 7013
rect 2511 6851 2563 6979
rect 3509 7013 3561 7025
rect 3509 6979 3519 7013
rect 3553 6979 3561 7013
rect 3799 7013 3851 7025
rect 3509 6851 3561 6979
rect 3799 6979 3807 7013
rect 3841 6979 3851 7013
rect 3799 6851 3851 6979
rect 4797 7013 4849 7025
rect 4797 6979 4807 7013
rect 4841 6979 4849 7013
rect 4797 6851 4849 6979
rect 4903 7013 4955 7025
rect 4903 6979 4911 7013
rect 4945 6979 4955 7013
rect 4903 6851 4955 6979
rect 5901 7013 5953 7025
rect 5901 6979 5911 7013
rect 5945 6979 5953 7013
rect 5901 6851 5953 6979
rect 6007 7013 6059 7025
rect 6007 6979 6015 7013
rect 6049 6979 6059 7013
rect 6007 6851 6059 6979
rect 7005 7013 7057 7025
rect 7005 6979 7015 7013
rect 7049 6979 7057 7013
rect 7005 6851 7057 6979
rect 7111 7013 7163 7025
rect 7111 6979 7119 7013
rect 7153 6979 7163 7013
rect 7111 6851 7163 6979
rect 8109 7013 8161 7025
rect 8109 6979 8119 7013
rect 8153 6979 8161 7013
rect 8109 6851 8161 6979
rect 8215 7013 8267 7025
rect 8215 6979 8223 7013
rect 8257 6979 8267 7013
rect 8215 6911 8267 6979
rect 8215 6877 8223 6911
rect 8257 6877 8267 6911
rect 8215 6851 8267 6877
rect 8661 7013 8713 7025
rect 8661 6979 8671 7013
rect 8705 6979 8713 7013
rect 8951 7013 9003 7025
rect 8661 6911 8713 6979
rect 8661 6877 8671 6911
rect 8705 6877 8713 6911
rect 8661 6851 8713 6877
rect 8951 6979 8959 7013
rect 8993 6979 9003 7013
rect 8951 6851 9003 6979
rect 9949 7013 10001 7025
rect 9949 6979 9959 7013
rect 9993 6979 10001 7013
rect 9949 6851 10001 6979
rect 10055 7013 10107 7025
rect 10055 6979 10063 7013
rect 10097 6979 10107 7013
rect 10055 6851 10107 6979
rect 11053 7013 11105 7025
rect 11053 6979 11063 7013
rect 11097 6979 11105 7013
rect 11053 6851 11105 6979
rect 11159 7013 11211 7025
rect 11159 6979 11167 7013
rect 11201 6979 11211 7013
rect 11159 6851 11211 6979
rect 12157 7013 12209 7025
rect 12157 6979 12167 7013
rect 12201 6979 12209 7013
rect 12157 6851 12209 6979
rect 12263 7013 12315 7025
rect 12263 6979 12271 7013
rect 12305 6979 12315 7013
rect 12263 6851 12315 6979
rect 13261 7013 13313 7025
rect 13261 6979 13271 7013
rect 13305 6979 13313 7013
rect 13261 6851 13313 6979
rect 13367 7013 13419 7025
rect 13367 6979 13375 7013
rect 13409 6979 13419 7013
rect 13367 6911 13419 6979
rect 13367 6877 13375 6911
rect 13409 6877 13419 6911
rect 13367 6851 13419 6877
rect 13813 7013 13865 7025
rect 13813 6979 13823 7013
rect 13857 6979 13865 7013
rect 14103 7013 14155 7025
rect 13813 6911 13865 6979
rect 13813 6877 13823 6911
rect 13857 6877 13865 6911
rect 13813 6851 13865 6877
rect 14103 6979 14111 7013
rect 14145 6979 14155 7013
rect 14103 6851 14155 6979
rect 15101 7013 15153 7025
rect 15101 6979 15111 7013
rect 15145 6979 15153 7013
rect 15101 6851 15153 6979
rect 15207 7013 15259 7025
rect 15207 6979 15215 7013
rect 15249 6979 15259 7013
rect 15207 6851 15259 6979
rect 16205 7013 16257 7025
rect 16205 6979 16215 7013
rect 16249 6979 16257 7013
rect 16205 6851 16257 6979
rect 16311 7013 16363 7025
rect 16311 6979 16319 7013
rect 16353 6979 16363 7013
rect 16311 6851 16363 6979
rect 17309 7013 17361 7025
rect 17309 6979 17319 7013
rect 17353 6979 17361 7013
rect 17309 6851 17361 6979
rect 17415 7013 17467 7025
rect 17415 6979 17423 7013
rect 17457 6979 17467 7013
rect 17415 6851 17467 6979
rect 18413 7013 18465 7025
rect 18413 6979 18423 7013
rect 18457 6979 18465 7013
rect 18413 6851 18465 6979
rect 18611 7013 18663 7025
rect 18611 6979 18619 7013
rect 18653 6979 18663 7013
rect 18611 6918 18663 6979
rect 18611 6884 18619 6918
rect 18653 6884 18663 6918
rect 18611 6851 18663 6884
rect 18781 7013 18833 7025
rect 18781 6979 18791 7013
rect 18825 6979 18833 7013
rect 18781 6918 18833 6979
rect 18781 6884 18791 6918
rect 18825 6884 18833 6918
rect 18781 6851 18833 6884
rect 1131 6172 1183 6205
rect 1131 6138 1139 6172
rect 1173 6138 1183 6172
rect 1131 6077 1183 6138
rect 1131 6043 1139 6077
rect 1173 6043 1183 6077
rect 1131 6031 1183 6043
rect 1301 6172 1353 6205
rect 1301 6138 1311 6172
rect 1345 6138 1353 6172
rect 1301 6077 1353 6138
rect 1301 6043 1311 6077
rect 1345 6043 1353 6077
rect 1301 6031 1353 6043
rect 1407 6077 1459 6205
rect 1407 6043 1415 6077
rect 1449 6043 1459 6077
rect 1407 6031 1459 6043
rect 2405 6077 2457 6205
rect 2405 6043 2415 6077
rect 2449 6043 2457 6077
rect 2405 6031 2457 6043
rect 2511 6077 2563 6205
rect 2511 6043 2519 6077
rect 2553 6043 2563 6077
rect 2511 6031 2563 6043
rect 3509 6077 3561 6205
rect 3509 6043 3519 6077
rect 3553 6043 3561 6077
rect 3509 6031 3561 6043
rect 3615 6077 3667 6205
rect 3615 6043 3623 6077
rect 3657 6043 3667 6077
rect 3615 6031 3667 6043
rect 4613 6077 4665 6205
rect 4613 6043 4623 6077
rect 4657 6043 4665 6077
rect 4613 6031 4665 6043
rect 4719 6077 4771 6205
rect 4719 6043 4727 6077
rect 4761 6043 4771 6077
rect 4719 6031 4771 6043
rect 5717 6077 5769 6205
rect 5717 6043 5727 6077
rect 5761 6043 5769 6077
rect 5717 6031 5769 6043
rect 5823 6179 5875 6205
rect 5823 6145 5831 6179
rect 5865 6145 5875 6179
rect 5823 6077 5875 6145
rect 5823 6043 5831 6077
rect 5865 6043 5875 6077
rect 5823 6031 5875 6043
rect 6085 6179 6137 6205
rect 6085 6145 6095 6179
rect 6129 6145 6137 6179
rect 6085 6077 6137 6145
rect 6085 6043 6095 6077
rect 6129 6043 6137 6077
rect 8072 6213 8124 6231
rect 6375 6077 6427 6205
rect 6085 6031 6137 6043
rect 6375 6043 6383 6077
rect 6417 6043 6427 6077
rect 6375 6031 6427 6043
rect 7373 6077 7425 6205
rect 7373 6043 7383 6077
rect 7417 6043 7425 6077
rect 7373 6031 7425 6043
rect 7479 6179 7531 6205
rect 7479 6145 7487 6179
rect 7521 6145 7531 6179
rect 7479 6077 7531 6145
rect 7479 6043 7487 6077
rect 7521 6043 7531 6077
rect 7479 6031 7531 6043
rect 7925 6179 7977 6205
rect 7925 6145 7935 6179
rect 7969 6145 7977 6179
rect 8072 6179 8080 6213
rect 8114 6179 8124 6213
rect 8072 6147 8124 6179
rect 8154 6147 8196 6231
rect 8226 6161 8293 6231
rect 8226 6147 8249 6161
rect 7925 6077 7977 6145
rect 8241 6127 8249 6147
rect 8283 6127 8293 6161
rect 7925 6043 7935 6077
rect 7969 6043 7977 6077
rect 7925 6031 7977 6043
rect 8241 6093 8293 6127
rect 8241 6059 8249 6093
rect 8283 6059 8293 6093
rect 8241 6031 8293 6059
rect 8323 6145 8391 6231
rect 8323 6111 8349 6145
rect 8383 6111 8391 6145
rect 8323 6077 8391 6111
rect 8323 6043 8349 6077
rect 8383 6043 8391 6077
rect 8323 6031 8391 6043
rect 8491 6077 8543 6205
rect 8491 6043 8499 6077
rect 8533 6043 8543 6077
rect 8491 6031 8543 6043
rect 9489 6077 9541 6205
rect 9489 6043 9499 6077
rect 9533 6043 9541 6077
rect 9489 6031 9541 6043
rect 9595 6077 9647 6205
rect 9595 6043 9603 6077
rect 9637 6043 9647 6077
rect 9595 6031 9647 6043
rect 10593 6077 10645 6205
rect 10593 6043 10603 6077
rect 10637 6043 10645 6077
rect 10593 6031 10645 6043
rect 10699 6179 10751 6205
rect 10699 6145 10707 6179
rect 10741 6145 10751 6179
rect 10699 6077 10751 6145
rect 10699 6043 10707 6077
rect 10741 6043 10751 6077
rect 10699 6031 10751 6043
rect 11329 6179 11381 6205
rect 11329 6145 11339 6179
rect 11373 6145 11381 6179
rect 11329 6077 11381 6145
rect 11329 6043 11339 6077
rect 11373 6043 11381 6077
rect 11527 6077 11579 6205
rect 11329 6031 11381 6043
rect 11527 6043 11535 6077
rect 11569 6043 11579 6077
rect 11527 6031 11579 6043
rect 12525 6077 12577 6205
rect 12525 6043 12535 6077
rect 12569 6043 12577 6077
rect 12525 6031 12577 6043
rect 12631 6077 12683 6205
rect 12631 6043 12639 6077
rect 12673 6043 12683 6077
rect 12631 6031 12683 6043
rect 13629 6077 13681 6205
rect 13629 6043 13639 6077
rect 13673 6043 13681 6077
rect 13629 6031 13681 6043
rect 13735 6077 13787 6205
rect 13735 6043 13743 6077
rect 13777 6043 13787 6077
rect 13735 6031 13787 6043
rect 14733 6077 14785 6205
rect 14733 6043 14743 6077
rect 14777 6043 14785 6077
rect 14733 6031 14785 6043
rect 14839 6077 14891 6205
rect 14839 6043 14847 6077
rect 14881 6043 14891 6077
rect 14839 6031 14891 6043
rect 15837 6077 15889 6205
rect 15837 6043 15847 6077
rect 15881 6043 15889 6077
rect 15837 6031 15889 6043
rect 15943 6179 15995 6205
rect 15943 6145 15951 6179
rect 15985 6145 15995 6179
rect 15943 6077 15995 6145
rect 15943 6043 15951 6077
rect 15985 6043 15995 6077
rect 15943 6031 15995 6043
rect 16389 6179 16441 6205
rect 16389 6145 16399 6179
rect 16433 6145 16441 6179
rect 16389 6077 16441 6145
rect 16389 6043 16399 6077
rect 16433 6043 16441 6077
rect 16679 6077 16731 6205
rect 16389 6031 16441 6043
rect 16679 6043 16687 6077
rect 16721 6043 16731 6077
rect 16679 6031 16731 6043
rect 17677 6077 17729 6205
rect 17677 6043 17687 6077
rect 17721 6043 17729 6077
rect 17677 6031 17729 6043
rect 17783 6179 17835 6205
rect 17783 6145 17791 6179
rect 17825 6145 17835 6179
rect 17783 6077 17835 6145
rect 17783 6043 17791 6077
rect 17825 6043 17835 6077
rect 17783 6031 17835 6043
rect 18413 6179 18465 6205
rect 18413 6145 18423 6179
rect 18457 6145 18465 6179
rect 18413 6077 18465 6145
rect 18413 6043 18423 6077
rect 18457 6043 18465 6077
rect 18413 6031 18465 6043
rect 18611 6172 18663 6205
rect 18611 6138 18619 6172
rect 18653 6138 18663 6172
rect 18611 6077 18663 6138
rect 18611 6043 18619 6077
rect 18653 6043 18663 6077
rect 18611 6031 18663 6043
rect 18781 6172 18833 6205
rect 18781 6138 18791 6172
rect 18825 6138 18833 6172
rect 18781 6077 18833 6138
rect 18781 6043 18791 6077
rect 18825 6043 18833 6077
rect 18781 6031 18833 6043
rect 1131 5925 1183 5937
rect 1131 5891 1139 5925
rect 1173 5891 1183 5925
rect 1131 5830 1183 5891
rect 1131 5796 1139 5830
rect 1173 5796 1183 5830
rect 1131 5763 1183 5796
rect 1301 5925 1353 5937
rect 1301 5891 1311 5925
rect 1345 5891 1353 5925
rect 1301 5830 1353 5891
rect 1301 5796 1311 5830
rect 1345 5796 1353 5830
rect 1301 5763 1353 5796
rect 1407 5925 1459 5937
rect 1407 5891 1415 5925
rect 1449 5891 1459 5925
rect 1407 5763 1459 5891
rect 2405 5925 2457 5937
rect 2405 5891 2415 5925
rect 2449 5891 2457 5925
rect 2405 5763 2457 5891
rect 2511 5925 2563 5937
rect 2511 5891 2519 5925
rect 2553 5891 2563 5925
rect 2511 5763 2563 5891
rect 3509 5925 3561 5937
rect 3509 5891 3519 5925
rect 3553 5891 3561 5925
rect 3799 5925 3851 5937
rect 3509 5763 3561 5891
rect 3799 5891 3807 5925
rect 3841 5891 3851 5925
rect 3799 5763 3851 5891
rect 4797 5925 4849 5937
rect 4797 5891 4807 5925
rect 4841 5891 4849 5925
rect 4797 5763 4849 5891
rect 4903 5925 4955 5937
rect 4903 5891 4911 5925
rect 4945 5891 4955 5925
rect 4903 5763 4955 5891
rect 5901 5925 5953 5937
rect 5901 5891 5911 5925
rect 5945 5891 5953 5925
rect 5901 5763 5953 5891
rect 6007 5925 6059 5937
rect 6007 5891 6015 5925
rect 6049 5891 6059 5925
rect 6007 5823 6059 5891
rect 6007 5789 6015 5823
rect 6049 5789 6059 5823
rect 6007 5763 6059 5789
rect 6637 5925 6689 5937
rect 6637 5891 6647 5925
rect 6681 5891 6689 5925
rect 6637 5823 6689 5891
rect 6637 5789 6647 5823
rect 6681 5789 6689 5823
rect 6637 5763 6689 5789
rect 6743 5917 6795 5937
rect 6743 5883 6751 5917
rect 6785 5883 6795 5917
rect 6743 5836 6795 5883
rect 6743 5802 6751 5836
rect 6785 5802 6795 5836
rect 6743 5779 6795 5802
rect 6825 5917 6883 5937
rect 6825 5883 6837 5917
rect 6871 5883 6883 5917
rect 6825 5849 6883 5883
rect 6825 5815 6837 5849
rect 6871 5815 6883 5849
rect 6825 5779 6883 5815
rect 6913 5917 6965 5937
rect 6913 5883 6923 5917
rect 6957 5883 6965 5917
rect 6913 5849 6965 5883
rect 6913 5815 6923 5849
rect 6957 5815 6965 5849
rect 6913 5779 6965 5815
rect 7019 5925 7071 5937
rect 7019 5891 7027 5925
rect 7061 5891 7071 5925
rect 7019 5823 7071 5891
rect 7019 5789 7027 5823
rect 7061 5789 7071 5823
rect 7019 5763 7071 5789
rect 7465 5925 7517 5937
rect 7465 5891 7475 5925
rect 7509 5891 7517 5925
rect 8211 5925 8263 5937
rect 8211 5898 8219 5925
rect 7465 5823 7517 5891
rect 7465 5789 7475 5823
rect 7509 5789 7517 5823
rect 7613 5865 7669 5898
rect 7613 5831 7625 5865
rect 7659 5831 7669 5865
rect 7613 5814 7669 5831
rect 7699 5865 7765 5898
rect 7699 5831 7711 5865
rect 7745 5831 7765 5865
rect 7699 5814 7765 5831
rect 7795 5814 7837 5898
rect 7867 5865 8051 5898
rect 7867 5831 7908 5865
rect 7942 5831 7983 5865
rect 8017 5831 8051 5865
rect 7867 5814 8051 5831
rect 8081 5814 8154 5898
rect 8184 5891 8219 5898
rect 8253 5891 8263 5925
rect 8184 5857 8263 5891
rect 8184 5823 8219 5857
rect 8253 5823 8263 5857
rect 8184 5814 8263 5823
rect 7465 5763 7517 5789
rect 8211 5789 8263 5814
rect 8211 5755 8219 5789
rect 8253 5755 8263 5789
rect 8211 5737 8263 5755
rect 8293 5925 8345 5937
rect 8293 5891 8303 5925
rect 8337 5891 8345 5925
rect 8293 5857 8345 5891
rect 8293 5823 8303 5857
rect 8337 5823 8345 5857
rect 8293 5789 8345 5823
rect 8293 5755 8303 5789
rect 8337 5755 8345 5789
rect 8399 5925 8451 5937
rect 8399 5891 8407 5925
rect 8441 5891 8451 5925
rect 8399 5823 8451 5891
rect 8399 5789 8407 5823
rect 8441 5789 8451 5823
rect 8399 5763 8451 5789
rect 8661 5925 8713 5937
rect 8661 5891 8671 5925
rect 8705 5891 8713 5925
rect 8951 5925 9003 5937
rect 8661 5823 8713 5891
rect 8661 5789 8671 5823
rect 8705 5789 8713 5823
rect 8661 5763 8713 5789
rect 8293 5737 8345 5755
rect 8951 5891 8959 5925
rect 8993 5891 9003 5925
rect 8951 5763 9003 5891
rect 9949 5925 10001 5937
rect 9949 5891 9959 5925
rect 9993 5891 10001 5925
rect 9949 5763 10001 5891
rect 10055 5925 10107 5937
rect 10055 5891 10063 5925
rect 10097 5891 10107 5925
rect 10055 5763 10107 5891
rect 11053 5925 11105 5937
rect 11053 5891 11063 5925
rect 11097 5891 11105 5925
rect 11053 5763 11105 5891
rect 11159 5925 11211 5937
rect 11159 5891 11167 5925
rect 11201 5891 11211 5925
rect 11159 5823 11211 5891
rect 11159 5789 11167 5823
rect 11201 5789 11211 5823
rect 11159 5763 11211 5789
rect 11421 5925 11473 5937
rect 11421 5891 11431 5925
rect 11465 5891 11473 5925
rect 11421 5823 11473 5891
rect 11737 5909 11789 5937
rect 11737 5875 11745 5909
rect 11779 5875 11789 5909
rect 11421 5789 11431 5823
rect 11465 5789 11473 5823
rect 11737 5841 11789 5875
rect 11737 5821 11745 5841
rect 11421 5763 11473 5789
rect 11568 5789 11620 5821
rect 11568 5755 11576 5789
rect 11610 5755 11620 5789
rect 11568 5737 11620 5755
rect 11650 5737 11692 5821
rect 11722 5807 11745 5821
rect 11779 5807 11789 5841
rect 11722 5737 11789 5807
rect 11819 5925 11887 5937
rect 11819 5891 11845 5925
rect 11879 5891 11887 5925
rect 11819 5857 11887 5891
rect 11819 5823 11845 5857
rect 11879 5823 11887 5857
rect 11819 5737 11887 5823
rect 11987 5925 12039 5937
rect 11987 5891 11995 5925
rect 12029 5891 12039 5925
rect 11987 5823 12039 5891
rect 11987 5789 11995 5823
rect 12029 5789 12039 5823
rect 11987 5763 12039 5789
rect 12617 5925 12669 5937
rect 12617 5891 12627 5925
rect 12661 5891 12669 5925
rect 12617 5823 12669 5891
rect 13025 5909 13077 5937
rect 13025 5875 13033 5909
rect 13067 5875 13077 5909
rect 12617 5789 12627 5823
rect 12661 5789 12669 5823
rect 13025 5841 13077 5875
rect 13025 5821 13033 5841
rect 12617 5763 12669 5789
rect 12856 5789 12908 5821
rect 12856 5755 12864 5789
rect 12898 5755 12908 5789
rect 12856 5737 12908 5755
rect 12938 5737 12980 5821
rect 13010 5807 13033 5821
rect 13067 5807 13077 5841
rect 13010 5737 13077 5807
rect 13107 5925 13175 5937
rect 13107 5891 13133 5925
rect 13167 5891 13175 5925
rect 13107 5857 13175 5891
rect 13107 5823 13133 5857
rect 13167 5823 13175 5857
rect 13107 5737 13175 5823
rect 13275 5925 13327 5937
rect 13275 5891 13283 5925
rect 13317 5891 13327 5925
rect 13275 5823 13327 5891
rect 13275 5789 13283 5823
rect 13317 5789 13327 5823
rect 13275 5763 13327 5789
rect 13905 5925 13957 5937
rect 13905 5891 13915 5925
rect 13949 5891 13957 5925
rect 14103 5925 14155 5937
rect 13905 5823 13957 5891
rect 13905 5789 13915 5823
rect 13949 5789 13957 5823
rect 13905 5763 13957 5789
rect 14103 5891 14111 5925
rect 14145 5891 14155 5925
rect 14103 5763 14155 5891
rect 15101 5925 15153 5937
rect 15101 5891 15111 5925
rect 15145 5891 15153 5925
rect 15101 5763 15153 5891
rect 15207 5925 15259 5937
rect 15207 5891 15215 5925
rect 15249 5891 15259 5925
rect 15207 5763 15259 5891
rect 16205 5925 16257 5937
rect 16205 5891 16215 5925
rect 16249 5891 16257 5925
rect 16205 5763 16257 5891
rect 16311 5925 16363 5937
rect 16311 5891 16319 5925
rect 16353 5891 16363 5925
rect 16311 5763 16363 5891
rect 17309 5925 17361 5937
rect 17309 5891 17319 5925
rect 17353 5891 17361 5925
rect 17309 5763 17361 5891
rect 17415 5925 17467 5937
rect 17415 5891 17423 5925
rect 17457 5891 17467 5925
rect 17415 5763 17467 5891
rect 18413 5925 18465 5937
rect 18413 5891 18423 5925
rect 18457 5891 18465 5925
rect 18413 5763 18465 5891
rect 18611 5925 18663 5937
rect 18611 5891 18619 5925
rect 18653 5891 18663 5925
rect 18611 5830 18663 5891
rect 18611 5796 18619 5830
rect 18653 5796 18663 5830
rect 18611 5763 18663 5796
rect 18781 5925 18833 5937
rect 18781 5891 18791 5925
rect 18825 5891 18833 5925
rect 18781 5830 18833 5891
rect 18781 5796 18791 5830
rect 18825 5796 18833 5830
rect 18781 5763 18833 5796
rect 1131 5084 1183 5117
rect 1131 5050 1139 5084
rect 1173 5050 1183 5084
rect 1131 4989 1183 5050
rect 1131 4955 1139 4989
rect 1173 4955 1183 4989
rect 1131 4943 1183 4955
rect 1301 5084 1353 5117
rect 1301 5050 1311 5084
rect 1345 5050 1353 5084
rect 1301 4989 1353 5050
rect 1301 4955 1311 4989
rect 1345 4955 1353 4989
rect 1301 4943 1353 4955
rect 1407 4989 1459 5117
rect 1407 4955 1415 4989
rect 1449 4955 1459 4989
rect 1407 4943 1459 4955
rect 2405 4989 2457 5117
rect 2405 4955 2415 4989
rect 2449 4955 2457 4989
rect 2405 4943 2457 4955
rect 2511 5084 2563 5117
rect 2511 5050 2519 5084
rect 2553 5050 2563 5084
rect 2511 4989 2563 5050
rect 2511 4955 2519 4989
rect 2553 4955 2563 4989
rect 2511 4943 2563 4955
rect 2681 5084 2733 5117
rect 2681 5050 2691 5084
rect 2725 5050 2733 5084
rect 2681 4989 2733 5050
rect 2681 4955 2691 4989
rect 2725 4955 2733 4989
rect 2681 4943 2733 4955
rect 2787 5065 2839 5077
rect 2787 5031 2795 5065
rect 2829 5031 2839 5065
rect 2787 4997 2839 5031
rect 2787 4963 2795 4997
rect 2829 4963 2839 4997
rect 2787 4949 2839 4963
rect 2869 5013 2923 5077
rect 2869 4979 2879 5013
rect 2913 4979 2923 5013
rect 2869 4949 2923 4979
rect 2953 5065 3005 5077
rect 2953 5031 2963 5065
rect 2997 5031 3005 5065
rect 2953 4997 3005 5031
rect 2953 4963 2963 4997
rect 2997 4963 3005 4997
rect 2953 4949 3005 4963
rect 3138 4989 3190 5027
rect 3138 4955 3146 4989
rect 3180 4955 3190 4989
rect 3138 4943 3190 4955
rect 3220 4997 3282 5027
rect 3220 4963 3230 4997
rect 3264 4963 3282 4997
rect 3220 4943 3282 4963
rect 3312 4991 3381 5027
rect 3312 4957 3323 4991
rect 3357 4957 3381 4991
rect 3312 4943 3381 4957
rect 3411 5015 3521 5027
rect 3411 4981 3477 5015
rect 3511 4981 3521 5015
rect 3411 4943 3521 4981
rect 3551 4999 3618 5027
rect 3551 4965 3574 4999
rect 3608 4965 3618 4999
rect 3551 4943 3618 4965
rect 3648 5015 3700 5027
rect 3648 4981 3658 5015
rect 3692 4981 3700 5015
rect 3648 4943 3700 4981
rect 3763 4989 3815 5111
rect 3763 4955 3771 4989
rect 3805 4955 3815 4989
rect 3763 4943 3815 4955
rect 3845 5027 3899 5111
rect 4441 5071 4491 5143
rect 4425 5057 4491 5071
rect 3845 4997 3914 5027
rect 3845 4963 3859 4997
rect 3893 4963 3914 4997
rect 3845 4943 3914 4963
rect 3944 4990 4000 5027
rect 3944 4956 3956 4990
rect 3990 4956 4000 4990
rect 3944 4943 4000 4956
rect 4030 4943 4084 5027
rect 4114 4989 4192 5027
rect 4114 4955 4148 4989
rect 4182 4955 4192 4989
rect 4114 4943 4192 4955
rect 4222 5015 4276 5027
rect 4222 4981 4232 5015
rect 4266 4981 4276 5015
rect 4222 4943 4276 4981
rect 4306 4989 4360 5027
rect 4306 4955 4318 4989
rect 4352 4955 4360 4989
rect 4306 4943 4360 4955
rect 4425 5023 4447 5057
rect 4481 5023 4491 5057
rect 4425 4989 4491 5023
rect 4425 4955 4447 4989
rect 4481 4955 4491 4989
rect 4425 4943 4491 4955
rect 4521 5093 4573 5143
rect 4521 5059 4531 5093
rect 4565 5059 4573 5093
rect 4521 5025 4573 5059
rect 4521 4991 4531 5025
rect 4565 4991 4573 5025
rect 4521 4943 4573 4991
rect 4627 4989 4679 5117
rect 4627 4955 4635 4989
rect 4669 4955 4679 4989
rect 4627 4943 4679 4955
rect 5625 4989 5677 5117
rect 5625 4955 5635 4989
rect 5669 4955 5677 4989
rect 5625 4943 5677 4955
rect 5731 5091 5783 5117
rect 5731 5057 5739 5091
rect 5773 5057 5783 5091
rect 5731 4989 5783 5057
rect 5731 4955 5739 4989
rect 5773 4955 5783 4989
rect 5731 4943 5783 4955
rect 6177 5091 6229 5117
rect 6177 5057 6187 5091
rect 6221 5057 6229 5091
rect 6177 4989 6229 5057
rect 6177 4955 6187 4989
rect 6221 4955 6229 4989
rect 6651 5125 6703 5143
rect 6375 5084 6427 5117
rect 6375 5050 6383 5084
rect 6417 5050 6427 5084
rect 6375 4989 6427 5050
rect 6177 4943 6229 4955
rect 6375 4955 6383 4989
rect 6417 4955 6427 4989
rect 6375 4943 6427 4955
rect 6545 5084 6597 5117
rect 6545 5050 6555 5084
rect 6589 5050 6597 5084
rect 6545 4989 6597 5050
rect 6545 4955 6555 4989
rect 6589 4955 6597 4989
rect 6545 4943 6597 4955
rect 6651 5091 6659 5125
rect 6693 5091 6703 5125
rect 6651 5057 6703 5091
rect 6651 5023 6659 5057
rect 6693 5023 6703 5057
rect 6651 4989 6703 5023
rect 6651 4955 6659 4989
rect 6693 4955 6703 4989
rect 6651 4943 6703 4955
rect 6733 5125 6785 5143
rect 6733 5091 6743 5125
rect 6777 5091 6785 5125
rect 6733 5066 6785 5091
rect 7479 5091 7531 5117
rect 6733 5057 6812 5066
rect 6733 5023 6743 5057
rect 6777 5023 6812 5057
rect 6733 4989 6812 5023
rect 6733 4955 6743 4989
rect 6777 4982 6812 4989
rect 6842 4982 6915 5066
rect 6945 5049 7129 5066
rect 6945 5015 6979 5049
rect 7013 5015 7054 5049
rect 7088 5015 7129 5049
rect 6945 4982 7129 5015
rect 7159 4982 7201 5066
rect 7231 5049 7297 5066
rect 7231 5015 7251 5049
rect 7285 5015 7297 5049
rect 7231 4982 7297 5015
rect 7327 5049 7383 5066
rect 7327 5015 7337 5049
rect 7371 5015 7383 5049
rect 7327 4982 7383 5015
rect 7479 5057 7487 5091
rect 7521 5057 7531 5091
rect 7479 4989 7531 5057
rect 6777 4955 6785 4982
rect 6733 4943 6785 4955
rect 7479 4955 7487 4989
rect 7521 4955 7531 4989
rect 7479 4943 7531 4955
rect 7741 5091 7793 5117
rect 7741 5057 7751 5091
rect 7785 5057 7793 5091
rect 7741 4989 7793 5057
rect 7741 4955 7751 4989
rect 7785 4955 7793 4989
rect 7741 4943 7793 4955
rect 7847 5065 7899 5077
rect 7847 5031 7855 5065
rect 7889 5031 7899 5065
rect 7847 4997 7899 5031
rect 7847 4963 7855 4997
rect 7889 4963 7899 4997
rect 7847 4949 7899 4963
rect 7929 5013 7983 5077
rect 7929 4979 7939 5013
rect 7973 4979 7983 5013
rect 7929 4949 7983 4979
rect 8013 5065 8065 5077
rect 8013 5031 8023 5065
rect 8057 5031 8065 5065
rect 8013 4997 8065 5031
rect 8013 4963 8023 4997
rect 8057 4963 8065 4997
rect 8013 4949 8065 4963
rect 8198 4989 8250 5027
rect 8198 4955 8206 4989
rect 8240 4955 8250 4989
rect 8198 4943 8250 4955
rect 8280 4997 8342 5027
rect 8280 4963 8290 4997
rect 8324 4963 8342 4997
rect 8280 4943 8342 4963
rect 8372 4991 8441 5027
rect 8372 4957 8383 4991
rect 8417 4957 8441 4991
rect 8372 4943 8441 4957
rect 8471 5015 8581 5027
rect 8471 4981 8537 5015
rect 8571 4981 8581 5015
rect 8471 4943 8581 4981
rect 8611 4999 8678 5027
rect 8611 4965 8634 4999
rect 8668 4965 8678 4999
rect 8611 4943 8678 4965
rect 8708 5015 8760 5027
rect 8708 4981 8718 5015
rect 8752 4981 8760 5015
rect 8708 4943 8760 4981
rect 8823 4989 8875 5111
rect 8823 4955 8831 4989
rect 8865 4955 8875 4989
rect 8823 4943 8875 4955
rect 8905 5027 8959 5111
rect 9501 5071 9551 5143
rect 9485 5057 9551 5071
rect 8905 4997 8974 5027
rect 8905 4963 8919 4997
rect 8953 4963 8974 4997
rect 8905 4943 8974 4963
rect 9004 4990 9060 5027
rect 9004 4956 9016 4990
rect 9050 4956 9060 4990
rect 9004 4943 9060 4956
rect 9090 4943 9144 5027
rect 9174 4989 9252 5027
rect 9174 4955 9208 4989
rect 9242 4955 9252 4989
rect 9174 4943 9252 4955
rect 9282 5015 9336 5027
rect 9282 4981 9292 5015
rect 9326 4981 9336 5015
rect 9282 4943 9336 4981
rect 9366 4989 9420 5027
rect 9366 4955 9378 4989
rect 9412 4955 9420 4989
rect 9366 4943 9420 4955
rect 9485 5023 9507 5057
rect 9541 5023 9551 5057
rect 9485 4989 9551 5023
rect 9485 4955 9507 4989
rect 9541 4955 9551 4989
rect 9485 4943 9551 4955
rect 9581 5093 9633 5143
rect 9581 5059 9591 5093
rect 9625 5059 9633 5093
rect 9581 5025 9633 5059
rect 9581 4991 9591 5025
rect 9625 4991 9633 5025
rect 9581 4943 9633 4991
rect 9687 5091 9739 5117
rect 9687 5057 9695 5091
rect 9729 5057 9739 5091
rect 9687 4989 9739 5057
rect 9687 4955 9695 4989
rect 9729 4955 9739 4989
rect 9687 4943 9739 4955
rect 9949 5091 10001 5117
rect 9949 5057 9959 5091
rect 9993 5057 10001 5091
rect 10695 5125 10747 5143
rect 10695 5091 10703 5125
rect 10737 5091 10747 5125
rect 10695 5066 10747 5091
rect 9949 4989 10001 5057
rect 9949 4955 9959 4989
rect 9993 4955 10001 4989
rect 10097 5049 10153 5066
rect 10097 5015 10109 5049
rect 10143 5015 10153 5049
rect 10097 4982 10153 5015
rect 10183 5049 10249 5066
rect 10183 5015 10195 5049
rect 10229 5015 10249 5049
rect 10183 4982 10249 5015
rect 10279 4982 10321 5066
rect 10351 5049 10535 5066
rect 10351 5015 10392 5049
rect 10426 5015 10467 5049
rect 10501 5015 10535 5049
rect 10351 4982 10535 5015
rect 10565 4982 10638 5066
rect 10668 5057 10747 5066
rect 10668 5023 10703 5057
rect 10737 5023 10747 5057
rect 10668 4989 10747 5023
rect 10668 4982 10703 4989
rect 9949 4943 10001 4955
rect 10695 4955 10703 4982
rect 10737 4955 10747 4989
rect 10695 4943 10747 4955
rect 10777 5125 10829 5143
rect 10777 5091 10787 5125
rect 10821 5091 10829 5125
rect 10777 5057 10829 5091
rect 10777 5023 10787 5057
rect 10821 5023 10829 5057
rect 10777 4989 10829 5023
rect 10777 4955 10787 4989
rect 10821 4955 10829 4989
rect 10777 4943 10829 4955
rect 10883 5091 10935 5117
rect 10883 5057 10891 5091
rect 10925 5057 10935 5091
rect 10883 4989 10935 5057
rect 10883 4955 10891 4989
rect 10925 4955 10935 4989
rect 10883 4943 10935 4955
rect 11329 5091 11381 5117
rect 11329 5057 11339 5091
rect 11373 5057 11381 5091
rect 11329 4989 11381 5057
rect 11329 4955 11339 4989
rect 11373 4955 11381 4989
rect 11711 5125 11763 5143
rect 11711 5091 11719 5125
rect 11753 5091 11763 5125
rect 11711 5057 11763 5091
rect 11711 5023 11719 5057
rect 11753 5023 11763 5057
rect 11711 4989 11763 5023
rect 11329 4943 11381 4955
rect 11711 4955 11719 4989
rect 11753 4955 11763 4989
rect 11711 4943 11763 4955
rect 11793 5125 11845 5143
rect 11793 5091 11803 5125
rect 11837 5091 11845 5125
rect 11793 5066 11845 5091
rect 12539 5091 12591 5117
rect 11793 5057 11872 5066
rect 11793 5023 11803 5057
rect 11837 5023 11872 5057
rect 11793 4989 11872 5023
rect 11793 4955 11803 4989
rect 11837 4982 11872 4989
rect 11902 4982 11975 5066
rect 12005 5049 12189 5066
rect 12005 5015 12039 5049
rect 12073 5015 12114 5049
rect 12148 5015 12189 5049
rect 12005 4982 12189 5015
rect 12219 4982 12261 5066
rect 12291 5049 12357 5066
rect 12291 5015 12311 5049
rect 12345 5015 12357 5049
rect 12291 4982 12357 5015
rect 12387 5049 12443 5066
rect 12387 5015 12397 5049
rect 12431 5015 12443 5049
rect 12387 4982 12443 5015
rect 12539 5057 12547 5091
rect 12581 5057 12591 5091
rect 12539 4989 12591 5057
rect 11837 4955 11845 4982
rect 11793 4943 11845 4955
rect 12539 4955 12547 4989
rect 12581 4955 12591 4989
rect 12539 4943 12591 4955
rect 12801 5091 12853 5117
rect 12801 5057 12811 5091
rect 12845 5057 12853 5091
rect 13547 5125 13599 5143
rect 13547 5091 13555 5125
rect 13589 5091 13599 5125
rect 13547 5066 13599 5091
rect 12801 4989 12853 5057
rect 12801 4955 12811 4989
rect 12845 4955 12853 4989
rect 12949 5049 13005 5066
rect 12949 5015 12961 5049
rect 12995 5015 13005 5049
rect 12949 4982 13005 5015
rect 13035 5049 13101 5066
rect 13035 5015 13047 5049
rect 13081 5015 13101 5049
rect 13035 4982 13101 5015
rect 13131 4982 13173 5066
rect 13203 5049 13387 5066
rect 13203 5015 13244 5049
rect 13278 5015 13319 5049
rect 13353 5015 13387 5049
rect 13203 4982 13387 5015
rect 13417 4982 13490 5066
rect 13520 5057 13599 5066
rect 13520 5023 13555 5057
rect 13589 5023 13599 5057
rect 13520 4989 13599 5023
rect 13520 4982 13555 4989
rect 12801 4943 12853 4955
rect 13547 4955 13555 4982
rect 13589 4955 13599 4989
rect 13547 4943 13599 4955
rect 13629 5125 13681 5143
rect 13629 5091 13639 5125
rect 13673 5091 13681 5125
rect 13629 5057 13681 5091
rect 13629 5023 13639 5057
rect 13673 5023 13681 5057
rect 13629 4989 13681 5023
rect 13629 4955 13639 4989
rect 13673 4955 13681 4989
rect 13629 4943 13681 4955
rect 13735 4989 13787 5117
rect 13735 4955 13743 4989
rect 13777 4955 13787 4989
rect 13735 4943 13787 4955
rect 14733 4989 14785 5117
rect 14733 4955 14743 4989
rect 14777 4955 14785 4989
rect 14733 4943 14785 4955
rect 14839 4989 14891 5117
rect 14839 4955 14847 4989
rect 14881 4955 14891 4989
rect 14839 4943 14891 4955
rect 15837 4989 15889 5117
rect 15837 4955 15847 4989
rect 15881 4955 15889 4989
rect 15837 4943 15889 4955
rect 15943 5091 15995 5117
rect 15943 5057 15951 5091
rect 15985 5057 15995 5091
rect 15943 4989 15995 5057
rect 15943 4955 15951 4989
rect 15985 4955 15995 4989
rect 15943 4943 15995 4955
rect 16389 5091 16441 5117
rect 16389 5057 16399 5091
rect 16433 5057 16441 5091
rect 16389 4989 16441 5057
rect 16389 4955 16399 4989
rect 16433 4955 16441 4989
rect 16679 4989 16731 5117
rect 16389 4943 16441 4955
rect 16679 4955 16687 4989
rect 16721 4955 16731 4989
rect 16679 4943 16731 4955
rect 17677 4989 17729 5117
rect 17677 4955 17687 4989
rect 17721 4955 17729 4989
rect 17677 4943 17729 4955
rect 17783 5091 17835 5117
rect 17783 5057 17791 5091
rect 17825 5057 17835 5091
rect 17783 4989 17835 5057
rect 17783 4955 17791 4989
rect 17825 4955 17835 4989
rect 17783 4943 17835 4955
rect 18413 5091 18465 5117
rect 18413 5057 18423 5091
rect 18457 5057 18465 5091
rect 18413 4989 18465 5057
rect 18413 4955 18423 4989
rect 18457 4955 18465 4989
rect 18413 4943 18465 4955
rect 18611 5084 18663 5117
rect 18611 5050 18619 5084
rect 18653 5050 18663 5084
rect 18611 4989 18663 5050
rect 18611 4955 18619 4989
rect 18653 4955 18663 4989
rect 18611 4943 18663 4955
rect 18781 5084 18833 5117
rect 18781 5050 18791 5084
rect 18825 5050 18833 5084
rect 18781 4989 18833 5050
rect 18781 4955 18791 4989
rect 18825 4955 18833 4989
rect 18781 4943 18833 4955
rect 1131 4837 1183 4849
rect 1131 4803 1139 4837
rect 1173 4803 1183 4837
rect 1131 4742 1183 4803
rect 1131 4708 1139 4742
rect 1173 4708 1183 4742
rect 1131 4675 1183 4708
rect 1301 4837 1353 4849
rect 1301 4803 1311 4837
rect 1345 4803 1353 4837
rect 1301 4742 1353 4803
rect 1301 4708 1311 4742
rect 1345 4708 1353 4742
rect 1301 4675 1353 4708
rect 1407 4837 1459 4849
rect 1407 4803 1415 4837
rect 1449 4803 1459 4837
rect 1407 4735 1459 4803
rect 1407 4701 1415 4735
rect 1449 4701 1459 4735
rect 1407 4675 1459 4701
rect 2037 4837 2089 4849
rect 2037 4803 2047 4837
rect 2081 4803 2089 4837
rect 2037 4735 2089 4803
rect 2037 4701 2047 4735
rect 2081 4701 2089 4735
rect 2037 4675 2089 4701
rect 2143 4837 2195 4849
rect 2143 4803 2151 4837
rect 2185 4803 2195 4837
rect 2143 4742 2195 4803
rect 2143 4708 2151 4742
rect 2185 4708 2195 4742
rect 2143 4675 2195 4708
rect 2313 4837 2365 4849
rect 2313 4803 2323 4837
rect 2357 4803 2365 4837
rect 2313 4742 2365 4803
rect 2313 4708 2323 4742
rect 2357 4708 2365 4742
rect 2313 4675 2365 4708
rect 2438 4811 2490 4849
rect 2438 4777 2446 4811
rect 2480 4777 2490 4811
rect 2438 4649 2490 4777
rect 2520 4837 2585 4849
rect 2520 4803 2536 4837
rect 2570 4803 2585 4837
rect 2520 4765 2585 4803
rect 2685 4811 2737 4849
rect 2685 4777 2695 4811
rect 2729 4777 2737 4811
rect 2685 4765 2737 4777
rect 2791 4811 2843 4849
rect 2791 4777 2799 4811
rect 2833 4777 2843 4811
rect 2791 4765 2843 4777
rect 2943 4837 2997 4849
rect 2943 4803 2953 4837
rect 2987 4803 2997 4837
rect 2943 4765 2997 4803
rect 3027 4811 3079 4849
rect 3027 4777 3037 4811
rect 3071 4777 3079 4811
rect 3027 4765 3079 4777
rect 3155 4837 3207 4849
rect 3155 4803 3163 4837
rect 3197 4803 3207 4837
rect 2520 4649 2570 4765
rect 3155 4735 3207 4803
rect 3155 4701 3163 4735
rect 3197 4701 3207 4735
rect 3155 4675 3207 4701
rect 3601 4837 3653 4849
rect 3601 4803 3611 4837
rect 3645 4803 3653 4837
rect 3601 4735 3653 4803
rect 3601 4701 3611 4735
rect 3645 4701 3653 4735
rect 3601 4675 3653 4701
rect 3984 4823 4044 4849
rect 3984 4789 3999 4823
rect 4033 4789 4044 4823
rect 3984 4755 4044 4789
rect 3984 4721 3999 4755
rect 4033 4721 4044 4755
rect 3984 4649 4044 4721
rect 4074 4829 4130 4849
rect 4074 4795 4085 4829
rect 4119 4795 4130 4829
rect 4074 4761 4130 4795
rect 4074 4727 4085 4761
rect 4119 4727 4130 4761
rect 4074 4693 4130 4727
rect 4074 4659 4085 4693
rect 4119 4659 4130 4693
rect 4074 4649 4130 4659
rect 4160 4837 4216 4849
rect 4160 4803 4171 4837
rect 4205 4803 4216 4837
rect 4160 4649 4216 4803
rect 4246 4802 4302 4849
rect 4246 4768 4257 4802
rect 4291 4768 4302 4802
rect 4246 4649 4302 4768
rect 4332 4837 4398 4849
rect 4332 4803 4353 4837
rect 4387 4803 4398 4837
rect 4332 4769 4398 4803
rect 4332 4735 4353 4769
rect 4387 4735 4398 4769
rect 4332 4649 4398 4735
rect 4428 4829 4481 4849
rect 4428 4795 4439 4829
rect 4473 4795 4481 4829
rect 4428 4707 4481 4795
rect 4428 4673 4439 4707
rect 4473 4673 4481 4707
rect 4535 4837 4587 4849
rect 4535 4803 4543 4837
rect 4577 4803 4587 4837
rect 4535 4735 4587 4803
rect 4535 4701 4543 4735
rect 4577 4701 4587 4735
rect 4535 4675 4587 4701
rect 4797 4837 4849 4849
rect 4797 4803 4807 4837
rect 4841 4803 4849 4837
rect 4797 4735 4849 4803
rect 4797 4701 4807 4735
rect 4841 4701 4849 4735
rect 4797 4675 4849 4701
rect 5087 4837 5139 4849
rect 5087 4803 5095 4837
rect 5129 4803 5139 4837
rect 5087 4735 5139 4803
rect 5087 4701 5095 4735
rect 5129 4701 5139 4735
rect 5087 4675 5139 4701
rect 5717 4837 5769 4849
rect 5717 4803 5727 4837
rect 5761 4803 5769 4837
rect 5717 4735 5769 4803
rect 5717 4701 5727 4735
rect 5761 4701 5769 4735
rect 5717 4675 5769 4701
rect 6053 4837 6121 4849
rect 6053 4803 6061 4837
rect 6095 4803 6121 4837
rect 6053 4769 6121 4803
rect 6053 4735 6061 4769
rect 6095 4735 6121 4769
rect 4428 4649 4481 4673
rect 6053 4649 6121 4735
rect 6151 4821 6203 4849
rect 6151 4787 6161 4821
rect 6195 4787 6203 4821
rect 6151 4753 6203 4787
rect 6467 4837 6519 4849
rect 6467 4803 6475 4837
rect 6509 4803 6519 4837
rect 6151 4719 6161 4753
rect 6195 4733 6203 4753
rect 6467 4735 6519 4803
rect 6195 4719 6218 4733
rect 6151 4649 6218 4719
rect 6248 4649 6290 4733
rect 6320 4701 6372 4733
rect 6320 4667 6330 4701
rect 6364 4667 6372 4701
rect 6467 4701 6475 4735
rect 6509 4701 6519 4735
rect 6467 4675 6519 4701
rect 6729 4837 6781 4849
rect 6729 4803 6739 4837
rect 6773 4803 6781 4837
rect 6729 4735 6781 4803
rect 7045 4821 7097 4849
rect 7045 4787 7053 4821
rect 7087 4787 7097 4821
rect 6729 4701 6739 4735
rect 6773 4701 6781 4735
rect 7045 4753 7097 4787
rect 7045 4733 7053 4753
rect 6729 4675 6781 4701
rect 6876 4701 6928 4733
rect 6320 4649 6372 4667
rect 6876 4667 6884 4701
rect 6918 4667 6928 4701
rect 6876 4649 6928 4667
rect 6958 4649 7000 4733
rect 7030 4719 7053 4733
rect 7087 4719 7097 4753
rect 7030 4649 7097 4719
rect 7127 4837 7195 4849
rect 7127 4803 7153 4837
rect 7187 4803 7195 4837
rect 7127 4769 7195 4803
rect 7127 4735 7153 4769
rect 7187 4735 7195 4769
rect 7127 4649 7195 4735
rect 7295 4837 7347 4849
rect 7295 4803 7303 4837
rect 7337 4803 7347 4837
rect 7295 4735 7347 4803
rect 7295 4701 7303 4735
rect 7337 4701 7347 4735
rect 7295 4675 7347 4701
rect 7741 4837 7793 4849
rect 7741 4803 7751 4837
rect 7785 4803 7793 4837
rect 7741 4735 7793 4803
rect 7741 4701 7751 4735
rect 7785 4701 7793 4735
rect 7741 4675 7793 4701
rect 7847 4837 7899 4849
rect 7847 4803 7855 4837
rect 7889 4803 7899 4837
rect 7847 4769 7899 4803
rect 7847 4735 7855 4769
rect 7889 4735 7899 4769
rect 7847 4701 7899 4735
rect 7847 4667 7855 4701
rect 7889 4667 7899 4701
rect 7847 4649 7899 4667
rect 7929 4837 7981 4849
rect 7929 4803 7939 4837
rect 7973 4810 7981 4837
rect 7973 4803 8008 4810
rect 7929 4769 8008 4803
rect 7929 4735 7939 4769
rect 7973 4735 8008 4769
rect 7929 4726 8008 4735
rect 8038 4726 8111 4810
rect 8141 4777 8325 4810
rect 8141 4743 8175 4777
rect 8209 4743 8250 4777
rect 8284 4743 8325 4777
rect 8141 4726 8325 4743
rect 8355 4726 8397 4810
rect 8427 4777 8493 4810
rect 8427 4743 8447 4777
rect 8481 4743 8493 4777
rect 8427 4726 8493 4743
rect 8523 4777 8579 4810
rect 8523 4743 8533 4777
rect 8567 4743 8579 4777
rect 8523 4726 8579 4743
rect 7929 4701 7981 4726
rect 7929 4667 7939 4701
rect 7973 4667 7981 4701
rect 7929 4649 7981 4667
rect 9345 4821 9397 4849
rect 9345 4787 9353 4821
rect 9387 4787 9397 4821
rect 9345 4753 9397 4787
rect 9345 4733 9353 4753
rect 9176 4701 9228 4733
rect 9176 4667 9184 4701
rect 9218 4667 9228 4701
rect 9176 4649 9228 4667
rect 9258 4649 9300 4733
rect 9330 4719 9353 4733
rect 9387 4719 9397 4753
rect 9330 4649 9397 4719
rect 9427 4837 9495 4849
rect 9427 4803 9453 4837
rect 9487 4803 9495 4837
rect 9427 4769 9495 4803
rect 9427 4735 9453 4769
rect 9487 4735 9495 4769
rect 9427 4649 9495 4735
rect 9595 4837 9647 4849
rect 9595 4803 9603 4837
rect 9637 4803 9647 4837
rect 9595 4735 9647 4803
rect 9595 4701 9603 4735
rect 9637 4701 9647 4735
rect 9595 4675 9647 4701
rect 9857 4837 9909 4849
rect 9857 4803 9867 4837
rect 9901 4803 9909 4837
rect 9857 4735 9909 4803
rect 9857 4701 9867 4735
rect 9901 4701 9909 4735
rect 9857 4675 9909 4701
rect 10147 4837 10199 4849
rect 10147 4803 10155 4837
rect 10189 4803 10199 4837
rect 10147 4735 10199 4803
rect 10147 4701 10155 4735
rect 10189 4701 10199 4735
rect 10147 4675 10199 4701
rect 10409 4837 10461 4849
rect 10409 4803 10419 4837
rect 10453 4803 10461 4837
rect 10409 4735 10461 4803
rect 10725 4821 10777 4849
rect 10725 4787 10733 4821
rect 10767 4787 10777 4821
rect 10409 4701 10419 4735
rect 10453 4701 10461 4735
rect 10725 4753 10777 4787
rect 10725 4733 10733 4753
rect 10409 4675 10461 4701
rect 10556 4701 10608 4733
rect 10556 4667 10564 4701
rect 10598 4667 10608 4701
rect 10556 4649 10608 4667
rect 10638 4649 10680 4733
rect 10710 4719 10733 4733
rect 10767 4719 10777 4753
rect 10710 4649 10777 4719
rect 10807 4837 10875 4849
rect 10807 4803 10833 4837
rect 10867 4803 10875 4837
rect 10807 4769 10875 4803
rect 10807 4735 10833 4769
rect 10867 4735 10875 4769
rect 10807 4649 10875 4735
rect 10975 4837 11027 4849
rect 10975 4803 10983 4837
rect 11017 4803 11027 4837
rect 10975 4735 11027 4803
rect 10975 4701 10983 4735
rect 11017 4701 11027 4735
rect 10975 4675 11027 4701
rect 11237 4837 11289 4849
rect 11237 4803 11247 4837
rect 11281 4803 11289 4837
rect 11237 4735 11289 4803
rect 11237 4701 11247 4735
rect 11281 4701 11289 4735
rect 11237 4675 11289 4701
rect 11343 4829 11395 4849
rect 11343 4795 11351 4829
rect 11385 4795 11395 4829
rect 11343 4761 11395 4795
rect 11343 4727 11351 4761
rect 11385 4727 11395 4761
rect 11343 4691 11395 4727
rect 11425 4829 11483 4849
rect 11425 4795 11437 4829
rect 11471 4795 11483 4829
rect 11425 4761 11483 4795
rect 11425 4727 11437 4761
rect 11471 4727 11483 4761
rect 11425 4691 11483 4727
rect 11513 4829 11565 4849
rect 11513 4795 11523 4829
rect 11557 4795 11565 4829
rect 11513 4748 11565 4795
rect 11513 4714 11523 4748
rect 11557 4714 11565 4748
rect 11513 4691 11565 4714
rect 11619 4837 11671 4849
rect 11619 4803 11627 4837
rect 11661 4803 11671 4837
rect 11619 4735 11671 4803
rect 11619 4701 11627 4735
rect 11661 4701 11671 4735
rect 11619 4675 11671 4701
rect 11881 4837 11933 4849
rect 11881 4803 11891 4837
rect 11925 4803 11933 4837
rect 12627 4837 12679 4849
rect 12627 4810 12635 4837
rect 11881 4735 11933 4803
rect 11881 4701 11891 4735
rect 11925 4701 11933 4735
rect 12029 4777 12085 4810
rect 12029 4743 12041 4777
rect 12075 4743 12085 4777
rect 12029 4726 12085 4743
rect 12115 4777 12181 4810
rect 12115 4743 12127 4777
rect 12161 4743 12181 4777
rect 12115 4726 12181 4743
rect 12211 4726 12253 4810
rect 12283 4777 12467 4810
rect 12283 4743 12324 4777
rect 12358 4743 12399 4777
rect 12433 4743 12467 4777
rect 12283 4726 12467 4743
rect 12497 4726 12570 4810
rect 12600 4803 12635 4810
rect 12669 4803 12679 4837
rect 12600 4769 12679 4803
rect 12600 4735 12635 4769
rect 12669 4735 12679 4769
rect 12600 4726 12679 4735
rect 11881 4675 11933 4701
rect 12627 4701 12679 4726
rect 12627 4667 12635 4701
rect 12669 4667 12679 4701
rect 12627 4649 12679 4667
rect 12709 4837 12761 4849
rect 12709 4803 12719 4837
rect 12753 4803 12761 4837
rect 12709 4769 12761 4803
rect 12709 4735 12719 4769
rect 12753 4735 12761 4769
rect 12709 4701 12761 4735
rect 12709 4667 12719 4701
rect 12753 4667 12761 4701
rect 12815 4837 12867 4849
rect 12815 4803 12823 4837
rect 12857 4803 12867 4837
rect 12815 4735 12867 4803
rect 12815 4701 12823 4735
rect 12857 4701 12867 4735
rect 12815 4675 12867 4701
rect 13077 4837 13129 4849
rect 13077 4803 13087 4837
rect 13121 4803 13129 4837
rect 13077 4735 13129 4803
rect 13077 4701 13087 4735
rect 13121 4701 13129 4735
rect 13077 4675 13129 4701
rect 13183 4829 13235 4849
rect 13183 4795 13191 4829
rect 13225 4795 13235 4829
rect 13183 4748 13235 4795
rect 13183 4714 13191 4748
rect 13225 4714 13235 4748
rect 13183 4691 13235 4714
rect 13265 4829 13323 4849
rect 13265 4795 13277 4829
rect 13311 4795 13323 4829
rect 13265 4761 13323 4795
rect 13265 4727 13277 4761
rect 13311 4727 13323 4761
rect 13265 4691 13323 4727
rect 13353 4829 13405 4849
rect 13353 4795 13363 4829
rect 13397 4795 13405 4829
rect 13353 4761 13405 4795
rect 13353 4727 13363 4761
rect 13397 4727 13405 4761
rect 13353 4691 13405 4727
rect 13459 4837 13511 4849
rect 13459 4803 13467 4837
rect 13501 4803 13511 4837
rect 13459 4735 13511 4803
rect 13459 4701 13467 4735
rect 13501 4701 13511 4735
rect 12709 4649 12761 4667
rect 13459 4675 13511 4701
rect 13905 4837 13957 4849
rect 13905 4803 13915 4837
rect 13949 4803 13957 4837
rect 14103 4837 14155 4849
rect 13905 4735 13957 4803
rect 13905 4701 13915 4735
rect 13949 4701 13957 4735
rect 13905 4675 13957 4701
rect 14103 4803 14111 4837
rect 14145 4803 14155 4837
rect 14103 4675 14155 4803
rect 15101 4837 15153 4849
rect 15101 4803 15111 4837
rect 15145 4803 15153 4837
rect 15101 4675 15153 4803
rect 15417 4821 15469 4849
rect 15417 4787 15425 4821
rect 15459 4787 15469 4821
rect 15417 4753 15469 4787
rect 15417 4733 15425 4753
rect 15248 4701 15300 4733
rect 15248 4667 15256 4701
rect 15290 4667 15300 4701
rect 15248 4649 15300 4667
rect 15330 4649 15372 4733
rect 15402 4719 15425 4733
rect 15459 4719 15469 4753
rect 15402 4649 15469 4719
rect 15499 4837 15567 4849
rect 15499 4803 15525 4837
rect 15559 4803 15567 4837
rect 15499 4769 15567 4803
rect 15499 4735 15525 4769
rect 15559 4735 15567 4769
rect 15499 4649 15567 4735
rect 15667 4837 15719 4849
rect 15667 4803 15675 4837
rect 15709 4803 15719 4837
rect 15667 4735 15719 4803
rect 15667 4701 15675 4735
rect 15709 4701 15719 4735
rect 15667 4675 15719 4701
rect 15929 4837 15981 4849
rect 15929 4803 15939 4837
rect 15973 4803 15981 4837
rect 15929 4735 15981 4803
rect 15929 4701 15939 4735
rect 15973 4701 15981 4735
rect 15929 4675 15981 4701
rect 16035 4829 16087 4849
rect 16035 4795 16043 4829
rect 16077 4795 16087 4829
rect 16035 4748 16087 4795
rect 16035 4714 16043 4748
rect 16077 4714 16087 4748
rect 16035 4691 16087 4714
rect 16117 4829 16175 4849
rect 16117 4795 16129 4829
rect 16163 4795 16175 4829
rect 16117 4761 16175 4795
rect 16117 4727 16129 4761
rect 16163 4727 16175 4761
rect 16117 4691 16175 4727
rect 16205 4829 16257 4849
rect 16205 4795 16215 4829
rect 16249 4795 16257 4829
rect 16205 4761 16257 4795
rect 16205 4727 16215 4761
rect 16249 4727 16257 4761
rect 16205 4691 16257 4727
rect 16311 4837 16363 4849
rect 16311 4803 16319 4837
rect 16353 4803 16363 4837
rect 16311 4735 16363 4803
rect 16311 4701 16319 4735
rect 16353 4701 16363 4735
rect 16311 4675 16363 4701
rect 16573 4837 16625 4849
rect 16573 4803 16583 4837
rect 16617 4803 16625 4837
rect 16573 4735 16625 4803
rect 16573 4701 16583 4735
rect 16617 4701 16625 4735
rect 16573 4675 16625 4701
rect 16679 4829 16731 4849
rect 16679 4795 16687 4829
rect 16721 4795 16731 4829
rect 16679 4748 16731 4795
rect 16679 4714 16687 4748
rect 16721 4714 16731 4748
rect 16679 4691 16731 4714
rect 16761 4829 16819 4849
rect 16761 4795 16773 4829
rect 16807 4795 16819 4829
rect 16761 4761 16819 4795
rect 16761 4727 16773 4761
rect 16807 4727 16819 4761
rect 16761 4691 16819 4727
rect 16849 4829 16901 4849
rect 16849 4795 16859 4829
rect 16893 4795 16901 4829
rect 16849 4761 16901 4795
rect 16849 4727 16859 4761
rect 16893 4727 16901 4761
rect 16849 4691 16901 4727
rect 16955 4837 17007 4849
rect 16955 4803 16963 4837
rect 16997 4803 17007 4837
rect 16955 4675 17007 4803
rect 17953 4837 18005 4849
rect 17953 4803 17963 4837
rect 17997 4803 18005 4837
rect 17953 4675 18005 4803
rect 18059 4837 18111 4849
rect 18059 4803 18067 4837
rect 18101 4803 18111 4837
rect 18059 4735 18111 4803
rect 18059 4701 18067 4735
rect 18101 4701 18111 4735
rect 18059 4675 18111 4701
rect 18505 4837 18557 4849
rect 18505 4803 18515 4837
rect 18549 4803 18557 4837
rect 18505 4735 18557 4803
rect 18505 4701 18515 4735
rect 18549 4701 18557 4735
rect 18505 4675 18557 4701
rect 18611 4837 18663 4849
rect 18611 4803 18619 4837
rect 18653 4803 18663 4837
rect 18611 4742 18663 4803
rect 18611 4708 18619 4742
rect 18653 4708 18663 4742
rect 18611 4675 18663 4708
rect 18781 4837 18833 4849
rect 18781 4803 18791 4837
rect 18825 4803 18833 4837
rect 18781 4742 18833 4803
rect 18781 4708 18791 4742
rect 18825 4708 18833 4742
rect 18781 4675 18833 4708
rect 1131 3996 1183 4029
rect 1131 3962 1139 3996
rect 1173 3962 1183 3996
rect 1131 3901 1183 3962
rect 1131 3867 1139 3901
rect 1173 3867 1183 3901
rect 1131 3855 1183 3867
rect 1301 3996 1353 4029
rect 1301 3962 1311 3996
rect 1345 3962 1353 3996
rect 1301 3901 1353 3962
rect 1301 3867 1311 3901
rect 1345 3867 1353 3901
rect 1301 3855 1353 3867
rect 1407 4003 1459 4029
rect 1407 3969 1415 4003
rect 1449 3969 1459 4003
rect 1407 3901 1459 3969
rect 1407 3867 1415 3901
rect 1449 3867 1459 3901
rect 1407 3855 1459 3867
rect 2037 4003 2089 4029
rect 2037 3969 2047 4003
rect 2081 3969 2089 4003
rect 2037 3901 2089 3969
rect 2037 3867 2047 3901
rect 2081 3867 2089 3901
rect 2037 3855 2089 3867
rect 2235 3977 2287 4013
rect 2235 3943 2243 3977
rect 2277 3943 2287 3977
rect 2235 3909 2287 3943
rect 2235 3875 2243 3909
rect 2277 3875 2287 3909
rect 2235 3855 2287 3875
rect 2317 3977 2375 4013
rect 2317 3943 2329 3977
rect 2363 3943 2375 3977
rect 2317 3909 2375 3943
rect 2317 3875 2329 3909
rect 2363 3875 2375 3909
rect 2317 3855 2375 3875
rect 2405 3990 2457 4013
rect 2405 3956 2415 3990
rect 2449 3956 2457 3990
rect 2405 3909 2457 3956
rect 2405 3875 2415 3909
rect 2449 3875 2457 3909
rect 2405 3855 2457 3875
rect 2511 4003 2563 4029
rect 2511 3969 2519 4003
rect 2553 3969 2563 4003
rect 2511 3901 2563 3969
rect 2511 3867 2519 3901
rect 2553 3867 2563 3901
rect 2511 3855 2563 3867
rect 2773 4003 2825 4029
rect 2773 3969 2783 4003
rect 2817 3969 2825 4003
rect 2773 3901 2825 3969
rect 2773 3867 2783 3901
rect 2817 3867 2825 3901
rect 2773 3855 2825 3867
rect 2879 3977 2931 3989
rect 2879 3943 2887 3977
rect 2921 3943 2931 3977
rect 2879 3909 2931 3943
rect 2879 3875 2887 3909
rect 2921 3875 2931 3909
rect 2879 3861 2931 3875
rect 2961 3925 3015 3989
rect 2961 3891 2971 3925
rect 3005 3891 3015 3925
rect 2961 3861 3015 3891
rect 3045 3977 3097 3989
rect 3045 3943 3055 3977
rect 3089 3943 3097 3977
rect 3045 3909 3097 3943
rect 3045 3875 3055 3909
rect 3089 3875 3097 3909
rect 3045 3861 3097 3875
rect 3230 3901 3282 3939
rect 3230 3867 3238 3901
rect 3272 3867 3282 3901
rect 3230 3855 3282 3867
rect 3312 3909 3374 3939
rect 3312 3875 3322 3909
rect 3356 3875 3374 3909
rect 3312 3855 3374 3875
rect 3404 3903 3473 3939
rect 3404 3869 3415 3903
rect 3449 3869 3473 3903
rect 3404 3855 3473 3869
rect 3503 3927 3613 3939
rect 3503 3893 3569 3927
rect 3603 3893 3613 3927
rect 3503 3855 3613 3893
rect 3643 3911 3710 3939
rect 3643 3877 3666 3911
rect 3700 3877 3710 3911
rect 3643 3855 3710 3877
rect 3740 3927 3792 3939
rect 3740 3893 3750 3927
rect 3784 3893 3792 3927
rect 3740 3855 3792 3893
rect 3855 3901 3907 4023
rect 3855 3867 3863 3901
rect 3897 3867 3907 3901
rect 3855 3855 3907 3867
rect 3937 3939 3991 4023
rect 4533 3983 4583 4055
rect 4517 3969 4583 3983
rect 3937 3909 4006 3939
rect 3937 3875 3951 3909
rect 3985 3875 4006 3909
rect 3937 3855 4006 3875
rect 4036 3902 4092 3939
rect 4036 3868 4048 3902
rect 4082 3868 4092 3902
rect 4036 3855 4092 3868
rect 4122 3855 4176 3939
rect 4206 3901 4284 3939
rect 4206 3867 4240 3901
rect 4274 3867 4284 3901
rect 4206 3855 4284 3867
rect 4314 3927 4368 3939
rect 4314 3893 4324 3927
rect 4358 3893 4368 3927
rect 4314 3855 4368 3893
rect 4398 3901 4452 3939
rect 4398 3867 4410 3901
rect 4444 3867 4452 3901
rect 4398 3855 4452 3867
rect 4517 3935 4539 3969
rect 4573 3935 4583 3969
rect 4517 3901 4583 3935
rect 4517 3867 4539 3901
rect 4573 3867 4583 3901
rect 4517 3855 4583 3867
rect 4613 4005 4665 4055
rect 4613 3971 4623 4005
rect 4657 3971 4665 4005
rect 4613 3937 4665 3971
rect 4613 3903 4623 3937
rect 4657 3903 4665 3937
rect 4613 3855 4665 3903
rect 4719 4003 4771 4029
rect 4719 3969 4727 4003
rect 4761 3969 4771 4003
rect 4719 3901 4771 3969
rect 4719 3867 4727 3901
rect 4761 3867 4771 3901
rect 4719 3855 4771 3867
rect 4981 4003 5033 4029
rect 4981 3969 4991 4003
rect 5025 3969 5033 4003
rect 4981 3901 5033 3969
rect 4981 3867 4991 3901
rect 5025 3867 5033 3901
rect 4981 3855 5033 3867
rect 5363 4003 5415 4029
rect 5363 3969 5371 4003
rect 5405 3969 5415 4003
rect 5363 3901 5415 3969
rect 5363 3867 5371 3901
rect 5405 3867 5415 3901
rect 5363 3855 5415 3867
rect 5993 4003 6045 4029
rect 5993 3969 6003 4003
rect 6037 3969 6045 4003
rect 5993 3901 6045 3969
rect 5993 3867 6003 3901
rect 6037 3867 6045 3901
rect 6375 3996 6427 4029
rect 6375 3962 6383 3996
rect 6417 3962 6427 3996
rect 6375 3901 6427 3962
rect 5993 3855 6045 3867
rect 6375 3867 6383 3901
rect 6417 3867 6427 3901
rect 6375 3855 6427 3867
rect 6545 3996 6597 4029
rect 6545 3962 6555 3996
rect 6589 3962 6597 3996
rect 6545 3901 6597 3962
rect 6545 3867 6555 3901
rect 6589 3867 6597 3901
rect 6545 3855 6597 3867
rect 6651 3990 6703 4013
rect 6651 3956 6659 3990
rect 6693 3956 6703 3990
rect 6651 3909 6703 3956
rect 6651 3875 6659 3909
rect 6693 3875 6703 3909
rect 6651 3855 6703 3875
rect 6733 3977 6791 4013
rect 6733 3943 6745 3977
rect 6779 3943 6791 3977
rect 6733 3909 6791 3943
rect 6733 3875 6745 3909
rect 6779 3875 6791 3909
rect 6733 3855 6791 3875
rect 6821 3977 6873 4013
rect 6821 3943 6831 3977
rect 6865 3943 6873 3977
rect 6821 3909 6873 3943
rect 6821 3875 6831 3909
rect 6865 3875 6873 3909
rect 6821 3855 6873 3875
rect 6927 4003 6979 4029
rect 6927 3969 6935 4003
rect 6969 3969 6979 4003
rect 6927 3901 6979 3969
rect 6927 3867 6935 3901
rect 6969 3867 6979 3901
rect 6927 3855 6979 3867
rect 7557 4003 7609 4029
rect 7557 3969 7567 4003
rect 7601 3969 7609 4003
rect 8303 4037 8355 4055
rect 8303 4003 8311 4037
rect 8345 4003 8355 4037
rect 8303 3978 8355 4003
rect 7557 3901 7609 3969
rect 7557 3867 7567 3901
rect 7601 3867 7609 3901
rect 7705 3961 7761 3978
rect 7705 3927 7717 3961
rect 7751 3927 7761 3961
rect 7705 3894 7761 3927
rect 7791 3961 7857 3978
rect 7791 3927 7803 3961
rect 7837 3927 7857 3961
rect 7791 3894 7857 3927
rect 7887 3894 7929 3978
rect 7959 3961 8143 3978
rect 7959 3927 8000 3961
rect 8034 3927 8075 3961
rect 8109 3927 8143 3961
rect 7959 3894 8143 3927
rect 8173 3894 8246 3978
rect 8276 3969 8355 3978
rect 8276 3935 8311 3969
rect 8345 3935 8355 3969
rect 8276 3901 8355 3935
rect 8276 3894 8311 3901
rect 7557 3855 7609 3867
rect 8303 3867 8311 3894
rect 8345 3867 8355 3901
rect 8303 3855 8355 3867
rect 8385 4037 8437 4055
rect 8385 4003 8395 4037
rect 8429 4003 8437 4037
rect 8385 3969 8437 4003
rect 8385 3935 8395 3969
rect 8429 3935 8437 3969
rect 8385 3901 8437 3935
rect 8385 3867 8395 3901
rect 8429 3867 8437 3901
rect 8385 3855 8437 3867
rect 8491 4003 8543 4029
rect 8491 3969 8499 4003
rect 8533 3969 8543 4003
rect 8491 3901 8543 3969
rect 8491 3867 8499 3901
rect 8533 3867 8543 3901
rect 8491 3855 8543 3867
rect 8753 4003 8805 4029
rect 8753 3969 8763 4003
rect 8797 3969 8805 4003
rect 8753 3901 8805 3969
rect 8753 3867 8763 3901
rect 8797 3867 8805 3901
rect 8753 3855 8805 3867
rect 8951 3969 9004 4055
rect 8951 3935 8959 3969
rect 8993 3935 9004 3969
rect 8951 3901 9004 3935
rect 8951 3867 8959 3901
rect 8993 3867 9004 3901
rect 8951 3855 9004 3867
rect 9034 3977 9090 4055
rect 9034 3943 9045 3977
rect 9079 3943 9090 3977
rect 9034 3909 9090 3943
rect 9034 3875 9045 3909
rect 9079 3875 9090 3909
rect 9034 3855 9090 3875
rect 9120 3969 9176 4055
rect 9120 3935 9131 3969
rect 9165 3935 9176 3969
rect 9120 3901 9176 3935
rect 9120 3867 9131 3901
rect 9165 3867 9176 3901
rect 9120 3855 9176 3867
rect 9206 3985 9262 4055
rect 9206 3951 9217 3985
rect 9251 3951 9262 3985
rect 9206 3917 9262 3951
rect 9206 3883 9217 3917
rect 9251 3883 9262 3917
rect 9206 3855 9262 3883
rect 9292 3969 9348 4055
rect 9292 3935 9303 3969
rect 9337 3935 9348 3969
rect 9292 3901 9348 3935
rect 9292 3867 9303 3901
rect 9337 3867 9348 3901
rect 9292 3855 9348 3867
rect 9378 4031 9434 4055
rect 9378 3997 9389 4031
rect 9423 3997 9434 4031
rect 9378 3945 9434 3997
rect 9378 3911 9389 3945
rect 9423 3911 9434 3945
rect 9378 3855 9434 3911
rect 9464 3925 9520 4055
rect 9464 3891 9475 3925
rect 9509 3891 9520 3925
rect 9464 3855 9520 3891
rect 9550 4031 9606 4055
rect 9550 3997 9561 4031
rect 9595 3997 9606 4031
rect 9550 3945 9606 3997
rect 9550 3911 9561 3945
rect 9595 3911 9606 3945
rect 9550 3855 9606 3911
rect 9636 3925 9692 4055
rect 9636 3891 9647 3925
rect 9681 3891 9692 3925
rect 9636 3855 9692 3891
rect 9722 4031 9778 4055
rect 9722 3997 9733 4031
rect 9767 3997 9778 4031
rect 9722 3945 9778 3997
rect 9722 3911 9733 3945
rect 9767 3911 9778 3945
rect 9722 3855 9778 3911
rect 9808 3925 9864 4055
rect 9808 3891 9819 3925
rect 9853 3891 9864 3925
rect 9808 3855 9864 3891
rect 9894 4031 9950 4055
rect 9894 3997 9905 4031
rect 9939 3997 9950 4031
rect 9894 3945 9950 3997
rect 9894 3911 9905 3945
rect 9939 3911 9950 3945
rect 9894 3855 9950 3911
rect 9980 3925 10035 4055
rect 9980 3891 9991 3925
rect 10025 3891 10035 3925
rect 9980 3855 10035 3891
rect 10065 4031 10121 4055
rect 10065 3997 10076 4031
rect 10110 3997 10121 4031
rect 10065 3945 10121 3997
rect 10065 3911 10076 3945
rect 10110 3911 10121 3945
rect 10065 3855 10121 3911
rect 10151 3925 10207 4055
rect 10151 3891 10162 3925
rect 10196 3891 10207 3925
rect 10151 3855 10207 3891
rect 10237 4031 10293 4055
rect 10237 3997 10248 4031
rect 10282 3997 10293 4031
rect 10237 3945 10293 3997
rect 10237 3911 10248 3945
rect 10282 3911 10293 3945
rect 10237 3855 10293 3911
rect 10323 3925 10379 4055
rect 10323 3891 10334 3925
rect 10368 3891 10379 3925
rect 10323 3855 10379 3891
rect 10409 4031 10465 4055
rect 10409 3997 10420 4031
rect 10454 3997 10465 4031
rect 10409 3945 10465 3997
rect 10409 3911 10420 3945
rect 10454 3911 10465 3945
rect 10409 3855 10465 3911
rect 10495 3925 10551 4055
rect 10495 3891 10506 3925
rect 10540 3891 10551 3925
rect 10495 3855 10551 3891
rect 10581 4031 10637 4055
rect 10581 3997 10592 4031
rect 10626 3997 10637 4031
rect 10581 3945 10637 3997
rect 10581 3911 10592 3945
rect 10626 3911 10637 3945
rect 10581 3855 10637 3911
rect 10667 3925 10720 4055
rect 10667 3891 10678 3925
rect 10712 3891 10720 3925
rect 10667 3855 10720 3891
rect 10791 4003 10843 4029
rect 10791 3969 10799 4003
rect 10833 3969 10843 4003
rect 10791 3901 10843 3969
rect 10791 3867 10799 3901
rect 10833 3867 10843 3901
rect 10791 3855 10843 3867
rect 11237 4003 11289 4029
rect 11237 3969 11247 4003
rect 11281 3969 11289 4003
rect 11237 3901 11289 3969
rect 11237 3867 11247 3901
rect 11281 3867 11289 3901
rect 11711 4005 11763 4055
rect 11711 3971 11719 4005
rect 11753 3971 11763 4005
rect 11711 3937 11763 3971
rect 11711 3903 11719 3937
rect 11753 3903 11763 3937
rect 11237 3855 11289 3867
rect 11711 3855 11763 3903
rect 11793 3983 11843 4055
rect 11793 3969 11859 3983
rect 11793 3935 11803 3969
rect 11837 3935 11859 3969
rect 12385 3939 12439 4023
rect 11793 3901 11859 3935
rect 11793 3867 11803 3901
rect 11837 3867 11859 3901
rect 11793 3855 11859 3867
rect 11924 3901 11978 3939
rect 11924 3867 11932 3901
rect 11966 3867 11978 3901
rect 11924 3855 11978 3867
rect 12008 3927 12062 3939
rect 12008 3893 12018 3927
rect 12052 3893 12062 3927
rect 12008 3855 12062 3893
rect 12092 3901 12170 3939
rect 12092 3867 12102 3901
rect 12136 3867 12170 3901
rect 12092 3855 12170 3867
rect 12200 3855 12254 3939
rect 12284 3902 12340 3939
rect 12284 3868 12294 3902
rect 12328 3868 12340 3902
rect 12284 3855 12340 3868
rect 12370 3909 12439 3939
rect 12370 3875 12391 3909
rect 12425 3875 12439 3909
rect 12370 3855 12439 3875
rect 12469 3901 12521 4023
rect 13551 4003 13603 4029
rect 13279 3977 13331 3989
rect 13279 3943 13287 3977
rect 13321 3943 13331 3977
rect 12469 3867 12479 3901
rect 12513 3867 12521 3901
rect 12469 3855 12521 3867
rect 12584 3927 12636 3939
rect 12584 3893 12592 3927
rect 12626 3893 12636 3927
rect 12584 3855 12636 3893
rect 12666 3911 12733 3939
rect 12666 3877 12676 3911
rect 12710 3877 12733 3911
rect 12666 3855 12733 3877
rect 12763 3927 12873 3939
rect 12763 3893 12773 3927
rect 12807 3893 12873 3927
rect 12763 3855 12873 3893
rect 12903 3903 12972 3939
rect 12903 3869 12927 3903
rect 12961 3869 12972 3903
rect 12903 3855 12972 3869
rect 13002 3909 13064 3939
rect 13002 3875 13020 3909
rect 13054 3875 13064 3909
rect 13002 3855 13064 3875
rect 13094 3901 13146 3939
rect 13094 3867 13104 3901
rect 13138 3867 13146 3901
rect 13094 3855 13146 3867
rect 13279 3909 13331 3943
rect 13279 3875 13287 3909
rect 13321 3875 13331 3909
rect 13279 3861 13331 3875
rect 13361 3925 13415 3989
rect 13361 3891 13371 3925
rect 13405 3891 13415 3925
rect 13361 3861 13415 3891
rect 13445 3977 13497 3989
rect 13445 3943 13455 3977
rect 13489 3943 13497 3977
rect 13445 3909 13497 3943
rect 13445 3875 13455 3909
rect 13489 3875 13497 3909
rect 13445 3861 13497 3875
rect 13551 3969 13559 4003
rect 13593 3969 13603 4003
rect 13551 3901 13603 3969
rect 13551 3867 13559 3901
rect 13593 3867 13603 3901
rect 13551 3855 13603 3867
rect 13813 4003 13865 4029
rect 13813 3969 13823 4003
rect 13857 3969 13865 4003
rect 13813 3901 13865 3969
rect 13813 3867 13823 3901
rect 13857 3867 13865 3901
rect 13813 3855 13865 3867
rect 13919 3977 13971 3989
rect 13919 3943 13927 3977
rect 13961 3943 13971 3977
rect 13919 3909 13971 3943
rect 13919 3875 13927 3909
rect 13961 3875 13971 3909
rect 13919 3861 13971 3875
rect 14001 3925 14055 3989
rect 14001 3891 14011 3925
rect 14045 3891 14055 3925
rect 14001 3861 14055 3891
rect 14085 3977 14137 3989
rect 14085 3943 14095 3977
rect 14129 3943 14137 3977
rect 14085 3909 14137 3943
rect 14085 3875 14095 3909
rect 14129 3875 14137 3909
rect 14085 3861 14137 3875
rect 14270 3901 14322 3939
rect 14270 3867 14278 3901
rect 14312 3867 14322 3901
rect 14270 3855 14322 3867
rect 14352 3909 14414 3939
rect 14352 3875 14362 3909
rect 14396 3875 14414 3909
rect 14352 3855 14414 3875
rect 14444 3903 14513 3939
rect 14444 3869 14455 3903
rect 14489 3869 14513 3903
rect 14444 3855 14513 3869
rect 14543 3927 14653 3939
rect 14543 3893 14609 3927
rect 14643 3893 14653 3927
rect 14543 3855 14653 3893
rect 14683 3911 14750 3939
rect 14683 3877 14706 3911
rect 14740 3877 14750 3911
rect 14683 3855 14750 3877
rect 14780 3927 14832 3939
rect 14780 3893 14790 3927
rect 14824 3893 14832 3927
rect 14780 3855 14832 3893
rect 14895 3901 14947 4023
rect 14895 3867 14903 3901
rect 14937 3867 14947 3901
rect 14895 3855 14947 3867
rect 14977 3939 15031 4023
rect 15573 3983 15623 4055
rect 15557 3969 15623 3983
rect 14977 3909 15046 3939
rect 14977 3875 14991 3909
rect 15025 3875 15046 3909
rect 14977 3855 15046 3875
rect 15076 3902 15132 3939
rect 15076 3868 15088 3902
rect 15122 3868 15132 3902
rect 15076 3855 15132 3868
rect 15162 3855 15216 3939
rect 15246 3901 15324 3939
rect 15246 3867 15280 3901
rect 15314 3867 15324 3901
rect 15246 3855 15324 3867
rect 15354 3927 15408 3939
rect 15354 3893 15364 3927
rect 15398 3893 15408 3927
rect 15354 3855 15408 3893
rect 15438 3901 15492 3939
rect 15438 3867 15450 3901
rect 15484 3867 15492 3901
rect 15438 3855 15492 3867
rect 15557 3935 15579 3969
rect 15613 3935 15623 3969
rect 15557 3901 15623 3935
rect 15557 3867 15579 3901
rect 15613 3867 15623 3901
rect 15557 3855 15623 3867
rect 15653 4005 15705 4055
rect 15653 3971 15663 4005
rect 15697 3971 15705 4005
rect 15653 3937 15705 3971
rect 15653 3903 15663 3937
rect 15697 3903 15705 3937
rect 15653 3855 15705 3903
rect 15759 4003 15811 4029
rect 15759 3969 15767 4003
rect 15801 3969 15811 4003
rect 15759 3901 15811 3969
rect 15759 3867 15767 3901
rect 15801 3867 15811 3901
rect 15759 3855 15811 3867
rect 16389 4003 16441 4029
rect 16389 3969 16399 4003
rect 16433 3969 16441 4003
rect 16389 3901 16441 3969
rect 16389 3867 16399 3901
rect 16433 3867 16441 3901
rect 16679 3901 16731 4029
rect 16389 3855 16441 3867
rect 16679 3867 16687 3901
rect 16721 3867 16731 3901
rect 16679 3855 16731 3867
rect 17677 3901 17729 4029
rect 17677 3867 17687 3901
rect 17721 3867 17729 3901
rect 17677 3855 17729 3867
rect 17783 4003 17835 4029
rect 17783 3969 17791 4003
rect 17825 3969 17835 4003
rect 17783 3901 17835 3969
rect 17783 3867 17791 3901
rect 17825 3867 17835 3901
rect 17783 3855 17835 3867
rect 18413 4003 18465 4029
rect 18413 3969 18423 4003
rect 18457 3969 18465 4003
rect 18413 3901 18465 3969
rect 18413 3867 18423 3901
rect 18457 3867 18465 3901
rect 18413 3855 18465 3867
rect 18611 3996 18663 4029
rect 18611 3962 18619 3996
rect 18653 3962 18663 3996
rect 18611 3901 18663 3962
rect 18611 3867 18619 3901
rect 18653 3867 18663 3901
rect 18611 3855 18663 3867
rect 18781 3996 18833 4029
rect 18781 3962 18791 3996
rect 18825 3962 18833 3996
rect 18781 3901 18833 3962
rect 18781 3867 18791 3901
rect 18825 3867 18833 3901
rect 18781 3855 18833 3867
rect 1131 3749 1183 3761
rect 1131 3715 1139 3749
rect 1173 3715 1183 3749
rect 1131 3654 1183 3715
rect 1131 3620 1139 3654
rect 1173 3620 1183 3654
rect 1131 3587 1183 3620
rect 1301 3749 1353 3761
rect 1301 3715 1311 3749
rect 1345 3715 1353 3749
rect 1301 3654 1353 3715
rect 1301 3620 1311 3654
rect 1345 3620 1353 3654
rect 1301 3587 1353 3620
rect 1407 3749 1459 3761
rect 1407 3715 1415 3749
rect 1449 3715 1459 3749
rect 1407 3654 1459 3715
rect 1407 3620 1415 3654
rect 1449 3620 1459 3654
rect 1407 3587 1459 3620
rect 1577 3749 1629 3761
rect 1577 3715 1587 3749
rect 1621 3715 1629 3749
rect 1577 3654 1629 3715
rect 1577 3620 1587 3654
rect 1621 3620 1629 3654
rect 1683 3741 1735 3755
rect 1683 3707 1691 3741
rect 1725 3707 1735 3741
rect 1683 3673 1735 3707
rect 1683 3639 1691 3673
rect 1725 3639 1735 3673
rect 1683 3627 1735 3639
rect 1765 3725 1819 3755
rect 1765 3691 1775 3725
rect 1809 3691 1819 3725
rect 1765 3627 1819 3691
rect 1849 3741 1901 3755
rect 1849 3707 1859 3741
rect 1893 3707 1901 3741
rect 1849 3673 1901 3707
rect 2034 3749 2086 3761
rect 2034 3715 2042 3749
rect 2076 3715 2086 3749
rect 2034 3677 2086 3715
rect 2116 3741 2178 3761
rect 2116 3707 2126 3741
rect 2160 3707 2178 3741
rect 2116 3677 2178 3707
rect 2208 3747 2277 3761
rect 2208 3713 2219 3747
rect 2253 3713 2277 3747
rect 2208 3677 2277 3713
rect 2307 3723 2417 3761
rect 2307 3689 2373 3723
rect 2407 3689 2417 3723
rect 2307 3677 2417 3689
rect 2447 3739 2514 3761
rect 2447 3705 2470 3739
rect 2504 3705 2514 3739
rect 2447 3677 2514 3705
rect 2544 3723 2596 3761
rect 2544 3689 2554 3723
rect 2588 3689 2596 3723
rect 2544 3677 2596 3689
rect 2659 3749 2711 3761
rect 2659 3715 2667 3749
rect 2701 3715 2711 3749
rect 1849 3639 1859 3673
rect 1893 3639 1901 3673
rect 1849 3627 1901 3639
rect 1577 3587 1629 3620
rect 2659 3593 2711 3715
rect 2741 3741 2810 3761
rect 2741 3707 2755 3741
rect 2789 3707 2810 3741
rect 2741 3677 2810 3707
rect 2840 3748 2896 3761
rect 2840 3714 2852 3748
rect 2886 3714 2896 3748
rect 2840 3677 2896 3714
rect 2926 3677 2980 3761
rect 3010 3749 3088 3761
rect 3010 3715 3044 3749
rect 3078 3715 3088 3749
rect 3010 3677 3088 3715
rect 3118 3723 3172 3761
rect 3118 3689 3128 3723
rect 3162 3689 3172 3723
rect 3118 3677 3172 3689
rect 3202 3749 3256 3761
rect 3202 3715 3214 3749
rect 3248 3715 3256 3749
rect 3202 3677 3256 3715
rect 3321 3749 3387 3761
rect 3321 3715 3343 3749
rect 3377 3715 3387 3749
rect 3321 3681 3387 3715
rect 2741 3593 2795 3677
rect 3321 3647 3343 3681
rect 3377 3647 3387 3681
rect 3321 3633 3387 3647
rect 3337 3561 3387 3633
rect 3417 3713 3469 3761
rect 3799 3749 3851 3761
rect 3417 3679 3427 3713
rect 3461 3679 3469 3713
rect 3417 3645 3469 3679
rect 3417 3611 3427 3645
rect 3461 3611 3469 3645
rect 3417 3561 3469 3611
rect 3799 3715 3807 3749
rect 3841 3715 3851 3749
rect 3799 3647 3851 3715
rect 3799 3613 3807 3647
rect 3841 3613 3851 3647
rect 3799 3587 3851 3613
rect 4429 3749 4481 3761
rect 4429 3715 4439 3749
rect 4473 3715 4481 3749
rect 4429 3647 4481 3715
rect 4429 3613 4439 3647
rect 4473 3613 4481 3647
rect 4429 3587 4481 3613
rect 4552 3725 4605 3761
rect 4552 3691 4560 3725
rect 4594 3691 4605 3725
rect 4552 3561 4605 3691
rect 4635 3705 4691 3761
rect 4635 3671 4646 3705
rect 4680 3671 4691 3705
rect 4635 3619 4691 3671
rect 4635 3585 4646 3619
rect 4680 3585 4691 3619
rect 4635 3561 4691 3585
rect 4721 3725 4777 3761
rect 4721 3691 4732 3725
rect 4766 3691 4777 3725
rect 4721 3561 4777 3691
rect 4807 3705 4863 3761
rect 4807 3671 4818 3705
rect 4852 3671 4863 3705
rect 4807 3619 4863 3671
rect 4807 3585 4818 3619
rect 4852 3585 4863 3619
rect 4807 3561 4863 3585
rect 4893 3725 4949 3761
rect 4893 3691 4904 3725
rect 4938 3691 4949 3725
rect 4893 3561 4949 3691
rect 4979 3705 5035 3761
rect 4979 3671 4990 3705
rect 5024 3671 5035 3705
rect 4979 3619 5035 3671
rect 4979 3585 4990 3619
rect 5024 3585 5035 3619
rect 4979 3561 5035 3585
rect 5065 3725 5121 3761
rect 5065 3691 5076 3725
rect 5110 3691 5121 3725
rect 5065 3561 5121 3691
rect 5151 3705 5207 3761
rect 5151 3671 5162 3705
rect 5196 3671 5207 3705
rect 5151 3619 5207 3671
rect 5151 3585 5162 3619
rect 5196 3585 5207 3619
rect 5151 3561 5207 3585
rect 5237 3725 5292 3761
rect 5237 3691 5247 3725
rect 5281 3691 5292 3725
rect 5237 3561 5292 3691
rect 5322 3705 5378 3761
rect 5322 3671 5333 3705
rect 5367 3671 5378 3705
rect 5322 3619 5378 3671
rect 5322 3585 5333 3619
rect 5367 3585 5378 3619
rect 5322 3561 5378 3585
rect 5408 3725 5464 3761
rect 5408 3691 5419 3725
rect 5453 3691 5464 3725
rect 5408 3561 5464 3691
rect 5494 3705 5550 3761
rect 5494 3671 5505 3705
rect 5539 3671 5550 3705
rect 5494 3619 5550 3671
rect 5494 3585 5505 3619
rect 5539 3585 5550 3619
rect 5494 3561 5550 3585
rect 5580 3725 5636 3761
rect 5580 3691 5591 3725
rect 5625 3691 5636 3725
rect 5580 3561 5636 3691
rect 5666 3705 5722 3761
rect 5666 3671 5677 3705
rect 5711 3671 5722 3705
rect 5666 3619 5722 3671
rect 5666 3585 5677 3619
rect 5711 3585 5722 3619
rect 5666 3561 5722 3585
rect 5752 3725 5808 3761
rect 5752 3691 5763 3725
rect 5797 3691 5808 3725
rect 5752 3561 5808 3691
rect 5838 3705 5894 3761
rect 5838 3671 5849 3705
rect 5883 3671 5894 3705
rect 5838 3619 5894 3671
rect 5838 3585 5849 3619
rect 5883 3585 5894 3619
rect 5838 3561 5894 3585
rect 5924 3749 5980 3761
rect 5924 3715 5935 3749
rect 5969 3715 5980 3749
rect 5924 3681 5980 3715
rect 5924 3647 5935 3681
rect 5969 3647 5980 3681
rect 5924 3561 5980 3647
rect 6010 3733 6066 3761
rect 6010 3699 6021 3733
rect 6055 3699 6066 3733
rect 6010 3665 6066 3699
rect 6010 3631 6021 3665
rect 6055 3631 6066 3665
rect 6010 3561 6066 3631
rect 6096 3749 6152 3761
rect 6096 3715 6107 3749
rect 6141 3715 6152 3749
rect 6096 3681 6152 3715
rect 6096 3647 6107 3681
rect 6141 3647 6152 3681
rect 6096 3561 6152 3647
rect 6182 3741 6238 3761
rect 6182 3707 6193 3741
rect 6227 3707 6238 3741
rect 6182 3673 6238 3707
rect 6182 3639 6193 3673
rect 6227 3639 6238 3673
rect 6182 3561 6238 3639
rect 6268 3749 6321 3761
rect 6268 3715 6279 3749
rect 6313 3715 6321 3749
rect 6268 3681 6321 3715
rect 6268 3647 6279 3681
rect 6313 3647 6321 3681
rect 6268 3561 6321 3647
rect 6375 3749 6427 3761
rect 6375 3715 6383 3749
rect 6417 3715 6427 3749
rect 6375 3647 6427 3715
rect 6375 3613 6383 3647
rect 6417 3613 6427 3647
rect 6375 3587 6427 3613
rect 6637 3749 6689 3761
rect 6637 3715 6647 3749
rect 6681 3715 6689 3749
rect 6637 3647 6689 3715
rect 6637 3613 6647 3647
rect 6681 3613 6689 3647
rect 6743 3741 6795 3755
rect 6743 3707 6751 3741
rect 6785 3707 6795 3741
rect 6743 3673 6795 3707
rect 6743 3639 6751 3673
rect 6785 3639 6795 3673
rect 6743 3627 6795 3639
rect 6825 3725 6879 3755
rect 6825 3691 6835 3725
rect 6869 3691 6879 3725
rect 6825 3627 6879 3691
rect 6909 3741 6961 3755
rect 6909 3707 6919 3741
rect 6953 3707 6961 3741
rect 6909 3673 6961 3707
rect 7094 3749 7146 3761
rect 7094 3715 7102 3749
rect 7136 3715 7146 3749
rect 7094 3677 7146 3715
rect 7176 3741 7238 3761
rect 7176 3707 7186 3741
rect 7220 3707 7238 3741
rect 7176 3677 7238 3707
rect 7268 3747 7337 3761
rect 7268 3713 7279 3747
rect 7313 3713 7337 3747
rect 7268 3677 7337 3713
rect 7367 3723 7477 3761
rect 7367 3689 7433 3723
rect 7467 3689 7477 3723
rect 7367 3677 7477 3689
rect 7507 3739 7574 3761
rect 7507 3705 7530 3739
rect 7564 3705 7574 3739
rect 7507 3677 7574 3705
rect 7604 3723 7656 3761
rect 7604 3689 7614 3723
rect 7648 3689 7656 3723
rect 7604 3677 7656 3689
rect 7719 3749 7771 3761
rect 7719 3715 7727 3749
rect 7761 3715 7771 3749
rect 6909 3639 6919 3673
rect 6953 3639 6961 3673
rect 6909 3627 6961 3639
rect 6637 3587 6689 3613
rect 7719 3593 7771 3715
rect 7801 3741 7870 3761
rect 7801 3707 7815 3741
rect 7849 3707 7870 3741
rect 7801 3677 7870 3707
rect 7900 3748 7956 3761
rect 7900 3714 7912 3748
rect 7946 3714 7956 3748
rect 7900 3677 7956 3714
rect 7986 3677 8040 3761
rect 8070 3749 8148 3761
rect 8070 3715 8104 3749
rect 8138 3715 8148 3749
rect 8070 3677 8148 3715
rect 8178 3723 8232 3761
rect 8178 3689 8188 3723
rect 8222 3689 8232 3723
rect 8178 3677 8232 3689
rect 8262 3749 8316 3761
rect 8262 3715 8274 3749
rect 8308 3715 8316 3749
rect 8262 3677 8316 3715
rect 8381 3749 8447 3761
rect 8381 3715 8403 3749
rect 8437 3715 8447 3749
rect 8381 3681 8447 3715
rect 7801 3593 7855 3677
rect 8381 3647 8403 3681
rect 8437 3647 8447 3681
rect 8381 3633 8447 3647
rect 8397 3561 8447 3633
rect 8477 3713 8529 3761
rect 8477 3679 8487 3713
rect 8521 3679 8529 3713
rect 8477 3645 8529 3679
rect 8477 3611 8487 3645
rect 8521 3611 8529 3645
rect 8477 3561 8529 3611
rect 8583 3749 8635 3761
rect 8583 3715 8591 3749
rect 8625 3715 8635 3749
rect 8583 3654 8635 3715
rect 8583 3620 8591 3654
rect 8625 3620 8635 3654
rect 8583 3587 8635 3620
rect 8753 3749 8805 3761
rect 9232 3753 9282 3761
rect 8753 3715 8763 3749
rect 8797 3715 8805 3749
rect 8753 3654 8805 3715
rect 8753 3620 8763 3654
rect 8797 3620 8805 3654
rect 8753 3587 8805 3620
rect 9135 3741 9187 3753
rect 9135 3707 9143 3741
rect 9177 3707 9187 3741
rect 9135 3673 9187 3707
rect 9135 3639 9143 3673
rect 9177 3639 9187 3673
rect 9135 3625 9187 3639
rect 9217 3741 9282 3753
rect 9217 3707 9236 3741
rect 9270 3707 9282 3741
rect 9217 3673 9282 3707
rect 9217 3639 9236 3673
rect 9270 3639 9282 3673
rect 9217 3625 9282 3639
rect 9232 3561 9282 3625
rect 9312 3725 9366 3761
rect 9312 3691 9322 3725
rect 9356 3691 9366 3725
rect 9312 3644 9366 3691
rect 9312 3610 9322 3644
rect 9356 3610 9366 3644
rect 9312 3561 9366 3610
rect 9396 3749 9449 3761
rect 9396 3715 9406 3749
rect 9440 3715 9449 3749
rect 9396 3681 9449 3715
rect 9396 3647 9406 3681
rect 9440 3647 9449 3681
rect 9396 3613 9449 3647
rect 9396 3579 9406 3613
rect 9440 3579 9449 3613
rect 9503 3749 9555 3761
rect 9503 3715 9511 3749
rect 9545 3715 9555 3749
rect 9503 3647 9555 3715
rect 9503 3613 9511 3647
rect 9545 3613 9555 3647
rect 9503 3587 9555 3613
rect 9949 3749 10001 3761
rect 9949 3715 9959 3749
rect 9993 3715 10001 3749
rect 9949 3647 10001 3715
rect 9949 3613 9959 3647
rect 9993 3613 10001 3647
rect 9949 3587 10001 3613
rect 10055 3741 10107 3761
rect 10055 3707 10063 3741
rect 10097 3707 10107 3741
rect 10055 3660 10107 3707
rect 10055 3626 10063 3660
rect 10097 3626 10107 3660
rect 10055 3603 10107 3626
rect 10137 3741 10195 3761
rect 10137 3707 10149 3741
rect 10183 3707 10195 3741
rect 10137 3673 10195 3707
rect 10137 3639 10149 3673
rect 10183 3639 10195 3673
rect 10137 3603 10195 3639
rect 10225 3741 10277 3761
rect 10225 3707 10235 3741
rect 10269 3707 10277 3741
rect 10225 3673 10277 3707
rect 10225 3639 10235 3673
rect 10269 3639 10277 3673
rect 10225 3603 10277 3639
rect 10331 3749 10383 3761
rect 10331 3715 10339 3749
rect 10373 3715 10383 3749
rect 10331 3647 10383 3715
rect 10331 3613 10339 3647
rect 10373 3613 10383 3647
rect 9396 3561 9449 3579
rect 10331 3587 10383 3613
rect 10777 3749 10829 3761
rect 10777 3715 10787 3749
rect 10821 3715 10829 3749
rect 10777 3647 10829 3715
rect 10777 3613 10787 3647
rect 10821 3613 10829 3647
rect 10777 3587 10829 3613
rect 10975 3741 11027 3761
rect 10975 3707 10983 3741
rect 11017 3707 11027 3741
rect 10975 3673 11027 3707
rect 10975 3639 10983 3673
rect 11017 3639 11027 3673
rect 10975 3603 11027 3639
rect 11057 3741 11115 3761
rect 11057 3707 11069 3741
rect 11103 3707 11115 3741
rect 11057 3673 11115 3707
rect 11057 3639 11069 3673
rect 11103 3639 11115 3673
rect 11057 3603 11115 3639
rect 11145 3741 11197 3761
rect 11145 3707 11155 3741
rect 11189 3707 11197 3741
rect 11145 3660 11197 3707
rect 11145 3626 11155 3660
rect 11189 3626 11197 3660
rect 11145 3603 11197 3626
rect 11251 3749 11303 3761
rect 11251 3715 11259 3749
rect 11293 3715 11303 3749
rect 11251 3647 11303 3715
rect 11251 3613 11259 3647
rect 11293 3613 11303 3647
rect 11251 3587 11303 3613
rect 11881 3749 11933 3761
rect 11881 3715 11891 3749
rect 11925 3715 11933 3749
rect 11881 3647 11933 3715
rect 11881 3613 11891 3647
rect 11925 3613 11933 3647
rect 11881 3587 11933 3613
rect 11987 3713 12039 3761
rect 11987 3679 11995 3713
rect 12029 3679 12039 3713
rect 11987 3645 12039 3679
rect 11987 3611 11995 3645
rect 12029 3611 12039 3645
rect 11987 3561 12039 3611
rect 12069 3749 12135 3761
rect 12069 3715 12079 3749
rect 12113 3715 12135 3749
rect 12069 3681 12135 3715
rect 12069 3647 12079 3681
rect 12113 3647 12135 3681
rect 12200 3749 12254 3761
rect 12200 3715 12208 3749
rect 12242 3715 12254 3749
rect 12200 3677 12254 3715
rect 12284 3723 12338 3761
rect 12284 3689 12294 3723
rect 12328 3689 12338 3723
rect 12284 3677 12338 3689
rect 12368 3749 12446 3761
rect 12368 3715 12378 3749
rect 12412 3715 12446 3749
rect 12368 3677 12446 3715
rect 12476 3677 12530 3761
rect 12560 3748 12616 3761
rect 12560 3714 12570 3748
rect 12604 3714 12616 3748
rect 12560 3677 12616 3714
rect 12646 3741 12715 3761
rect 12646 3707 12667 3741
rect 12701 3707 12715 3741
rect 12646 3677 12715 3707
rect 12069 3633 12135 3647
rect 12069 3561 12119 3633
rect 12661 3593 12715 3677
rect 12745 3749 12797 3761
rect 12745 3715 12755 3749
rect 12789 3715 12797 3749
rect 12745 3593 12797 3715
rect 12860 3723 12912 3761
rect 12860 3689 12868 3723
rect 12902 3689 12912 3723
rect 12860 3677 12912 3689
rect 12942 3739 13009 3761
rect 12942 3705 12952 3739
rect 12986 3705 13009 3739
rect 12942 3677 13009 3705
rect 13039 3723 13149 3761
rect 13039 3689 13049 3723
rect 13083 3689 13149 3723
rect 13039 3677 13149 3689
rect 13179 3747 13248 3761
rect 13179 3713 13203 3747
rect 13237 3713 13248 3747
rect 13179 3677 13248 3713
rect 13278 3741 13340 3761
rect 13278 3707 13296 3741
rect 13330 3707 13340 3741
rect 13278 3677 13340 3707
rect 13370 3749 13422 3761
rect 13370 3715 13380 3749
rect 13414 3715 13422 3749
rect 13370 3677 13422 3715
rect 13555 3741 13607 3755
rect 13555 3707 13563 3741
rect 13597 3707 13607 3741
rect 13555 3673 13607 3707
rect 13555 3639 13563 3673
rect 13597 3639 13607 3673
rect 13555 3627 13607 3639
rect 13637 3725 13691 3755
rect 13637 3691 13647 3725
rect 13681 3691 13691 3725
rect 13637 3627 13691 3691
rect 13721 3741 13773 3755
rect 14103 3749 14155 3761
rect 13721 3707 13731 3741
rect 13765 3707 13773 3741
rect 13721 3673 13773 3707
rect 13721 3639 13731 3673
rect 13765 3639 13773 3673
rect 13721 3627 13773 3639
rect 14103 3715 14111 3749
rect 14145 3715 14155 3749
rect 14103 3587 14155 3715
rect 15101 3749 15153 3761
rect 15101 3715 15111 3749
rect 15145 3715 15153 3749
rect 15101 3587 15153 3715
rect 15207 3749 15259 3761
rect 15207 3715 15215 3749
rect 15249 3715 15259 3749
rect 15207 3587 15259 3715
rect 16205 3749 16257 3761
rect 16205 3715 16215 3749
rect 16249 3715 16257 3749
rect 16205 3587 16257 3715
rect 16311 3749 16363 3761
rect 16311 3715 16319 3749
rect 16353 3715 16363 3749
rect 16311 3587 16363 3715
rect 17309 3749 17361 3761
rect 17309 3715 17319 3749
rect 17353 3715 17361 3749
rect 17309 3587 17361 3715
rect 17415 3749 17467 3761
rect 17415 3715 17423 3749
rect 17457 3715 17467 3749
rect 17415 3587 17467 3715
rect 18413 3749 18465 3761
rect 18413 3715 18423 3749
rect 18457 3715 18465 3749
rect 18413 3587 18465 3715
rect 18611 3749 18663 3761
rect 18611 3715 18619 3749
rect 18653 3715 18663 3749
rect 18611 3654 18663 3715
rect 18611 3620 18619 3654
rect 18653 3620 18663 3654
rect 18611 3587 18663 3620
rect 18781 3749 18833 3761
rect 18781 3715 18791 3749
rect 18825 3715 18833 3749
rect 18781 3654 18833 3715
rect 18781 3620 18791 3654
rect 18825 3620 18833 3654
rect 18781 3587 18833 3620
rect 1131 2908 1183 2941
rect 1131 2874 1139 2908
rect 1173 2874 1183 2908
rect 1131 2813 1183 2874
rect 1131 2779 1139 2813
rect 1173 2779 1183 2813
rect 1131 2767 1183 2779
rect 1301 2908 1353 2941
rect 1301 2874 1311 2908
rect 1345 2874 1353 2908
rect 1301 2813 1353 2874
rect 1301 2779 1311 2813
rect 1345 2779 1353 2813
rect 1301 2767 1353 2779
rect 1407 2915 1459 2941
rect 1407 2881 1415 2915
rect 1449 2881 1459 2915
rect 1407 2813 1459 2881
rect 1407 2779 1415 2813
rect 1449 2779 1459 2813
rect 1407 2767 1459 2779
rect 1853 2915 1905 2941
rect 1853 2881 1863 2915
rect 1897 2881 1905 2915
rect 1853 2813 1905 2881
rect 1853 2779 1863 2813
rect 1897 2779 1905 2813
rect 1853 2767 1905 2779
rect 1959 2917 2011 2967
rect 1959 2883 1967 2917
rect 2001 2883 2011 2917
rect 1959 2849 2011 2883
rect 1959 2815 1967 2849
rect 2001 2815 2011 2849
rect 1959 2767 2011 2815
rect 2041 2895 2091 2967
rect 2041 2881 2107 2895
rect 2041 2847 2051 2881
rect 2085 2847 2107 2881
rect 2633 2851 2687 2935
rect 2041 2813 2107 2847
rect 2041 2779 2051 2813
rect 2085 2779 2107 2813
rect 2041 2767 2107 2779
rect 2172 2813 2226 2851
rect 2172 2779 2180 2813
rect 2214 2779 2226 2813
rect 2172 2767 2226 2779
rect 2256 2839 2310 2851
rect 2256 2805 2266 2839
rect 2300 2805 2310 2839
rect 2256 2767 2310 2805
rect 2340 2813 2418 2851
rect 2340 2779 2350 2813
rect 2384 2779 2418 2813
rect 2340 2767 2418 2779
rect 2448 2767 2502 2851
rect 2532 2814 2588 2851
rect 2532 2780 2542 2814
rect 2576 2780 2588 2814
rect 2532 2767 2588 2780
rect 2618 2821 2687 2851
rect 2618 2787 2639 2821
rect 2673 2787 2687 2821
rect 2618 2767 2687 2787
rect 2717 2813 2769 2935
rect 3799 2915 3851 2941
rect 3527 2889 3579 2901
rect 3527 2855 3535 2889
rect 3569 2855 3579 2889
rect 2717 2779 2727 2813
rect 2761 2779 2769 2813
rect 2717 2767 2769 2779
rect 2832 2839 2884 2851
rect 2832 2805 2840 2839
rect 2874 2805 2884 2839
rect 2832 2767 2884 2805
rect 2914 2823 2981 2851
rect 2914 2789 2924 2823
rect 2958 2789 2981 2823
rect 2914 2767 2981 2789
rect 3011 2839 3121 2851
rect 3011 2805 3021 2839
rect 3055 2805 3121 2839
rect 3011 2767 3121 2805
rect 3151 2815 3220 2851
rect 3151 2781 3175 2815
rect 3209 2781 3220 2815
rect 3151 2767 3220 2781
rect 3250 2821 3312 2851
rect 3250 2787 3268 2821
rect 3302 2787 3312 2821
rect 3250 2767 3312 2787
rect 3342 2813 3394 2851
rect 3342 2779 3352 2813
rect 3386 2779 3394 2813
rect 3342 2767 3394 2779
rect 3527 2821 3579 2855
rect 3527 2787 3535 2821
rect 3569 2787 3579 2821
rect 3527 2773 3579 2787
rect 3609 2837 3663 2901
rect 3609 2803 3619 2837
rect 3653 2803 3663 2837
rect 3609 2773 3663 2803
rect 3693 2889 3745 2901
rect 3693 2855 3703 2889
rect 3737 2855 3745 2889
rect 3693 2821 3745 2855
rect 3693 2787 3703 2821
rect 3737 2787 3745 2821
rect 3693 2773 3745 2787
rect 3799 2881 3807 2915
rect 3841 2881 3851 2915
rect 3799 2813 3851 2881
rect 3799 2779 3807 2813
rect 3841 2779 3851 2813
rect 3799 2767 3851 2779
rect 4061 2915 4113 2941
rect 4061 2881 4071 2915
rect 4105 2881 4113 2915
rect 4061 2813 4113 2881
rect 4061 2779 4071 2813
rect 4105 2779 4113 2813
rect 4061 2767 4113 2779
rect 4167 2889 4219 2901
rect 4167 2855 4175 2889
rect 4209 2855 4219 2889
rect 4167 2821 4219 2855
rect 4167 2787 4175 2821
rect 4209 2787 4219 2821
rect 4167 2773 4219 2787
rect 4249 2837 4303 2901
rect 4249 2803 4259 2837
rect 4293 2803 4303 2837
rect 4249 2773 4303 2803
rect 4333 2889 4385 2901
rect 4333 2855 4343 2889
rect 4377 2855 4385 2889
rect 4333 2821 4385 2855
rect 4333 2787 4343 2821
rect 4377 2787 4385 2821
rect 4333 2773 4385 2787
rect 4439 2837 4491 2935
rect 4439 2803 4447 2837
rect 4481 2803 4491 2837
rect 4439 2767 4491 2803
rect 4521 2889 4573 2935
rect 4521 2855 4531 2889
rect 4565 2855 4573 2889
rect 4521 2851 4573 2855
rect 5555 2851 5606 2935
rect 4521 2821 4588 2851
rect 4521 2787 4531 2821
rect 4565 2787 4588 2821
rect 4521 2767 4588 2787
rect 4618 2814 4672 2851
rect 4618 2780 4628 2814
rect 4662 2780 4672 2814
rect 4618 2767 4672 2780
rect 4702 2767 4792 2851
rect 4822 2813 4898 2851
rect 4822 2779 4842 2813
rect 4876 2779 4898 2813
rect 4822 2767 4898 2779
rect 4928 2839 4982 2851
rect 4928 2805 4938 2839
rect 4972 2805 4982 2839
rect 4928 2767 4982 2805
rect 5012 2813 5066 2851
rect 5012 2779 5022 2813
rect 5056 2779 5066 2813
rect 5012 2767 5066 2779
rect 5096 2767 5142 2851
rect 5172 2815 5250 2851
rect 5172 2781 5182 2815
rect 5216 2781 5250 2815
rect 5172 2767 5250 2781
rect 5280 2767 5322 2851
rect 5352 2813 5404 2851
rect 5352 2779 5362 2813
rect 5396 2779 5404 2813
rect 5352 2767 5404 2779
rect 5458 2839 5510 2851
rect 5458 2805 5466 2839
rect 5500 2805 5510 2839
rect 5458 2767 5510 2805
rect 5540 2839 5606 2851
rect 5540 2805 5562 2839
rect 5596 2805 5606 2839
rect 5540 2767 5606 2805
rect 5636 2907 5688 2935
rect 5636 2873 5646 2907
rect 5680 2873 5688 2907
rect 5839 2895 5889 2967
rect 5636 2839 5688 2873
rect 5636 2805 5646 2839
rect 5680 2805 5688 2839
rect 5636 2767 5688 2805
rect 5742 2881 5794 2895
rect 5742 2847 5750 2881
rect 5784 2847 5794 2881
rect 5742 2813 5794 2847
rect 5742 2779 5750 2813
rect 5784 2779 5794 2813
rect 5742 2767 5794 2779
rect 5824 2881 5889 2895
rect 5824 2847 5845 2881
rect 5879 2847 5889 2881
rect 5824 2813 5889 2847
rect 5824 2779 5845 2813
rect 5879 2779 5889 2813
rect 5824 2767 5889 2779
rect 5919 2917 5971 2967
rect 5919 2883 5929 2917
rect 5963 2883 5971 2917
rect 5919 2849 5971 2883
rect 5919 2815 5929 2849
rect 5963 2815 5971 2849
rect 5919 2767 5971 2815
rect 6375 2915 6427 2941
rect 6375 2881 6383 2915
rect 6417 2881 6427 2915
rect 6375 2813 6427 2881
rect 6375 2779 6383 2813
rect 6417 2779 6427 2813
rect 6375 2767 6427 2779
rect 7005 2915 7057 2941
rect 7005 2881 7015 2915
rect 7049 2881 7057 2915
rect 7005 2813 7057 2881
rect 7005 2779 7015 2813
rect 7049 2779 7057 2813
rect 7005 2767 7057 2779
rect 7203 2917 7255 2967
rect 7203 2883 7211 2917
rect 7245 2883 7255 2917
rect 7203 2849 7255 2883
rect 7203 2815 7211 2849
rect 7245 2815 7255 2849
rect 7203 2767 7255 2815
rect 7285 2895 7335 2967
rect 7285 2881 7351 2895
rect 7285 2847 7295 2881
rect 7329 2847 7351 2881
rect 7877 2851 7931 2935
rect 7285 2813 7351 2847
rect 7285 2779 7295 2813
rect 7329 2779 7351 2813
rect 7285 2767 7351 2779
rect 7416 2813 7470 2851
rect 7416 2779 7424 2813
rect 7458 2779 7470 2813
rect 7416 2767 7470 2779
rect 7500 2839 7554 2851
rect 7500 2805 7510 2839
rect 7544 2805 7554 2839
rect 7500 2767 7554 2805
rect 7584 2813 7662 2851
rect 7584 2779 7594 2813
rect 7628 2779 7662 2813
rect 7584 2767 7662 2779
rect 7692 2767 7746 2851
rect 7776 2814 7832 2851
rect 7776 2780 7786 2814
rect 7820 2780 7832 2814
rect 7776 2767 7832 2780
rect 7862 2821 7931 2851
rect 7862 2787 7883 2821
rect 7917 2787 7931 2821
rect 7862 2767 7931 2787
rect 7961 2813 8013 2935
rect 9043 2915 9095 2941
rect 8771 2889 8823 2901
rect 8771 2855 8779 2889
rect 8813 2855 8823 2889
rect 7961 2779 7971 2813
rect 8005 2779 8013 2813
rect 7961 2767 8013 2779
rect 8076 2839 8128 2851
rect 8076 2805 8084 2839
rect 8118 2805 8128 2839
rect 8076 2767 8128 2805
rect 8158 2823 8225 2851
rect 8158 2789 8168 2823
rect 8202 2789 8225 2823
rect 8158 2767 8225 2789
rect 8255 2839 8365 2851
rect 8255 2805 8265 2839
rect 8299 2805 8365 2839
rect 8255 2767 8365 2805
rect 8395 2815 8464 2851
rect 8395 2781 8419 2815
rect 8453 2781 8464 2815
rect 8395 2767 8464 2781
rect 8494 2821 8556 2851
rect 8494 2787 8512 2821
rect 8546 2787 8556 2821
rect 8494 2767 8556 2787
rect 8586 2813 8638 2851
rect 8586 2779 8596 2813
rect 8630 2779 8638 2813
rect 8586 2767 8638 2779
rect 8771 2821 8823 2855
rect 8771 2787 8779 2821
rect 8813 2787 8823 2821
rect 8771 2773 8823 2787
rect 8853 2837 8907 2901
rect 8853 2803 8863 2837
rect 8897 2803 8907 2837
rect 8853 2773 8907 2803
rect 8937 2889 8989 2901
rect 8937 2855 8947 2889
rect 8981 2855 8989 2889
rect 8937 2821 8989 2855
rect 8937 2787 8947 2821
rect 8981 2787 8989 2821
rect 8937 2773 8989 2787
rect 9043 2881 9051 2915
rect 9085 2881 9095 2915
rect 9043 2813 9095 2881
rect 9043 2779 9051 2813
rect 9085 2779 9095 2813
rect 9043 2767 9095 2779
rect 9305 2915 9357 2941
rect 9305 2881 9315 2915
rect 9349 2881 9357 2915
rect 9305 2813 9357 2881
rect 9305 2779 9315 2813
rect 9349 2779 9357 2813
rect 9305 2767 9357 2779
rect 9411 2881 9464 2967
rect 9411 2847 9419 2881
rect 9453 2847 9464 2881
rect 9411 2813 9464 2847
rect 9411 2779 9419 2813
rect 9453 2779 9464 2813
rect 9411 2767 9464 2779
rect 9494 2889 9550 2967
rect 9494 2855 9505 2889
rect 9539 2855 9550 2889
rect 9494 2821 9550 2855
rect 9494 2787 9505 2821
rect 9539 2787 9550 2821
rect 9494 2767 9550 2787
rect 9580 2881 9636 2967
rect 9580 2847 9591 2881
rect 9625 2847 9636 2881
rect 9580 2813 9636 2847
rect 9580 2779 9591 2813
rect 9625 2779 9636 2813
rect 9580 2767 9636 2779
rect 9666 2897 9722 2967
rect 9666 2863 9677 2897
rect 9711 2863 9722 2897
rect 9666 2829 9722 2863
rect 9666 2795 9677 2829
rect 9711 2795 9722 2829
rect 9666 2767 9722 2795
rect 9752 2881 9808 2967
rect 9752 2847 9763 2881
rect 9797 2847 9808 2881
rect 9752 2813 9808 2847
rect 9752 2779 9763 2813
rect 9797 2779 9808 2813
rect 9752 2767 9808 2779
rect 9838 2943 9894 2967
rect 9838 2909 9849 2943
rect 9883 2909 9894 2943
rect 9838 2857 9894 2909
rect 9838 2823 9849 2857
rect 9883 2823 9894 2857
rect 9838 2767 9894 2823
rect 9924 2837 9980 2967
rect 9924 2803 9935 2837
rect 9969 2803 9980 2837
rect 9924 2767 9980 2803
rect 10010 2943 10066 2967
rect 10010 2909 10021 2943
rect 10055 2909 10066 2943
rect 10010 2857 10066 2909
rect 10010 2823 10021 2857
rect 10055 2823 10066 2857
rect 10010 2767 10066 2823
rect 10096 2837 10152 2967
rect 10096 2803 10107 2837
rect 10141 2803 10152 2837
rect 10096 2767 10152 2803
rect 10182 2943 10238 2967
rect 10182 2909 10193 2943
rect 10227 2909 10238 2943
rect 10182 2857 10238 2909
rect 10182 2823 10193 2857
rect 10227 2823 10238 2857
rect 10182 2767 10238 2823
rect 10268 2837 10324 2967
rect 10268 2803 10279 2837
rect 10313 2803 10324 2837
rect 10268 2767 10324 2803
rect 10354 2943 10410 2967
rect 10354 2909 10365 2943
rect 10399 2909 10410 2943
rect 10354 2857 10410 2909
rect 10354 2823 10365 2857
rect 10399 2823 10410 2857
rect 10354 2767 10410 2823
rect 10440 2837 10495 2967
rect 10440 2803 10451 2837
rect 10485 2803 10495 2837
rect 10440 2767 10495 2803
rect 10525 2943 10581 2967
rect 10525 2909 10536 2943
rect 10570 2909 10581 2943
rect 10525 2857 10581 2909
rect 10525 2823 10536 2857
rect 10570 2823 10581 2857
rect 10525 2767 10581 2823
rect 10611 2837 10667 2967
rect 10611 2803 10622 2837
rect 10656 2803 10667 2837
rect 10611 2767 10667 2803
rect 10697 2943 10753 2967
rect 10697 2909 10708 2943
rect 10742 2909 10753 2943
rect 10697 2857 10753 2909
rect 10697 2823 10708 2857
rect 10742 2823 10753 2857
rect 10697 2767 10753 2823
rect 10783 2837 10839 2967
rect 10783 2803 10794 2837
rect 10828 2803 10839 2837
rect 10783 2767 10839 2803
rect 10869 2943 10925 2967
rect 10869 2909 10880 2943
rect 10914 2909 10925 2943
rect 10869 2857 10925 2909
rect 10869 2823 10880 2857
rect 10914 2823 10925 2857
rect 10869 2767 10925 2823
rect 10955 2837 11011 2967
rect 10955 2803 10966 2837
rect 11000 2803 11011 2837
rect 10955 2767 11011 2803
rect 11041 2943 11097 2967
rect 11041 2909 11052 2943
rect 11086 2909 11097 2943
rect 11041 2857 11097 2909
rect 11041 2823 11052 2857
rect 11086 2823 11097 2857
rect 11041 2767 11097 2823
rect 11127 2837 11180 2967
rect 11127 2803 11138 2837
rect 11172 2803 11180 2837
rect 11127 2767 11180 2803
rect 11711 2917 11763 2967
rect 11711 2883 11719 2917
rect 11753 2883 11763 2917
rect 11711 2849 11763 2883
rect 11711 2815 11719 2849
rect 11753 2815 11763 2849
rect 11711 2767 11763 2815
rect 11793 2895 11843 2967
rect 11793 2881 11859 2895
rect 11793 2847 11803 2881
rect 11837 2847 11859 2881
rect 12385 2851 12439 2935
rect 11793 2813 11859 2847
rect 11793 2779 11803 2813
rect 11837 2779 11859 2813
rect 11793 2767 11859 2779
rect 11924 2813 11978 2851
rect 11924 2779 11932 2813
rect 11966 2779 11978 2813
rect 11924 2767 11978 2779
rect 12008 2839 12062 2851
rect 12008 2805 12018 2839
rect 12052 2805 12062 2839
rect 12008 2767 12062 2805
rect 12092 2813 12170 2851
rect 12092 2779 12102 2813
rect 12136 2779 12170 2813
rect 12092 2767 12170 2779
rect 12200 2767 12254 2851
rect 12284 2814 12340 2851
rect 12284 2780 12294 2814
rect 12328 2780 12340 2814
rect 12284 2767 12340 2780
rect 12370 2821 12439 2851
rect 12370 2787 12391 2821
rect 12425 2787 12439 2821
rect 12370 2767 12439 2787
rect 12469 2813 12521 2935
rect 13551 2915 13603 2941
rect 13279 2889 13331 2901
rect 13279 2855 13287 2889
rect 13321 2855 13331 2889
rect 12469 2779 12479 2813
rect 12513 2779 12521 2813
rect 12469 2767 12521 2779
rect 12584 2839 12636 2851
rect 12584 2805 12592 2839
rect 12626 2805 12636 2839
rect 12584 2767 12636 2805
rect 12666 2823 12733 2851
rect 12666 2789 12676 2823
rect 12710 2789 12733 2823
rect 12666 2767 12733 2789
rect 12763 2839 12873 2851
rect 12763 2805 12773 2839
rect 12807 2805 12873 2839
rect 12763 2767 12873 2805
rect 12903 2815 12972 2851
rect 12903 2781 12927 2815
rect 12961 2781 12972 2815
rect 12903 2767 12972 2781
rect 13002 2821 13064 2851
rect 13002 2787 13020 2821
rect 13054 2787 13064 2821
rect 13002 2767 13064 2787
rect 13094 2813 13146 2851
rect 13094 2779 13104 2813
rect 13138 2779 13146 2813
rect 13094 2767 13146 2779
rect 13279 2821 13331 2855
rect 13279 2787 13287 2821
rect 13321 2787 13331 2821
rect 13279 2773 13331 2787
rect 13361 2837 13415 2901
rect 13361 2803 13371 2837
rect 13405 2803 13415 2837
rect 13361 2773 13415 2803
rect 13445 2889 13497 2901
rect 13445 2855 13455 2889
rect 13489 2855 13497 2889
rect 13445 2821 13497 2855
rect 13445 2787 13455 2821
rect 13489 2787 13497 2821
rect 13445 2773 13497 2787
rect 13551 2881 13559 2915
rect 13593 2881 13603 2915
rect 13551 2813 13603 2881
rect 13551 2779 13559 2813
rect 13593 2779 13603 2813
rect 13551 2767 13603 2779
rect 13813 2915 13865 2941
rect 13813 2881 13823 2915
rect 13857 2881 13865 2915
rect 14016 2903 14066 2967
rect 13813 2813 13865 2881
rect 13813 2779 13823 2813
rect 13857 2779 13865 2813
rect 13813 2767 13865 2779
rect 13919 2889 13971 2903
rect 13919 2855 13927 2889
rect 13961 2855 13971 2889
rect 13919 2821 13971 2855
rect 13919 2787 13927 2821
rect 13961 2787 13971 2821
rect 13919 2775 13971 2787
rect 14001 2889 14066 2903
rect 14001 2855 14020 2889
rect 14054 2855 14066 2889
rect 14001 2821 14066 2855
rect 14001 2787 14020 2821
rect 14054 2787 14066 2821
rect 14001 2775 14066 2787
rect 14016 2767 14066 2775
rect 14096 2918 14150 2967
rect 14096 2884 14106 2918
rect 14140 2884 14150 2918
rect 14096 2837 14150 2884
rect 14096 2803 14106 2837
rect 14140 2803 14150 2837
rect 14096 2767 14150 2803
rect 14180 2949 14233 2967
rect 14180 2915 14190 2949
rect 14224 2915 14233 2949
rect 14180 2881 14233 2915
rect 14180 2847 14190 2881
rect 14224 2847 14233 2881
rect 14180 2813 14233 2847
rect 14180 2779 14190 2813
rect 14224 2779 14233 2813
rect 14180 2767 14233 2779
rect 14287 2813 14339 2941
rect 14287 2779 14295 2813
rect 14329 2779 14339 2813
rect 14287 2767 14339 2779
rect 15285 2813 15337 2941
rect 15285 2779 15295 2813
rect 15329 2779 15337 2813
rect 15285 2767 15337 2779
rect 15391 2813 15443 2941
rect 15391 2779 15399 2813
rect 15433 2779 15443 2813
rect 15391 2767 15443 2779
rect 16389 2813 16441 2941
rect 16389 2779 16399 2813
rect 16433 2779 16441 2813
rect 16679 2813 16731 2941
rect 16389 2767 16441 2779
rect 16679 2779 16687 2813
rect 16721 2779 16731 2813
rect 16679 2767 16731 2779
rect 17677 2813 17729 2941
rect 17677 2779 17687 2813
rect 17721 2779 17729 2813
rect 17677 2767 17729 2779
rect 17783 2915 17835 2941
rect 17783 2881 17791 2915
rect 17825 2881 17835 2915
rect 17783 2813 17835 2881
rect 17783 2779 17791 2813
rect 17825 2779 17835 2813
rect 17783 2767 17835 2779
rect 18413 2915 18465 2941
rect 18413 2881 18423 2915
rect 18457 2881 18465 2915
rect 18413 2813 18465 2881
rect 18413 2779 18423 2813
rect 18457 2779 18465 2813
rect 18413 2767 18465 2779
rect 18611 2908 18663 2941
rect 18611 2874 18619 2908
rect 18653 2874 18663 2908
rect 18611 2813 18663 2874
rect 18611 2779 18619 2813
rect 18653 2779 18663 2813
rect 18611 2767 18663 2779
rect 18781 2908 18833 2941
rect 18781 2874 18791 2908
rect 18825 2874 18833 2908
rect 18781 2813 18833 2874
rect 18781 2779 18791 2813
rect 18825 2779 18833 2813
rect 18781 2767 18833 2779
rect 1131 2661 1183 2673
rect 1131 2627 1139 2661
rect 1173 2627 1183 2661
rect 1131 2566 1183 2627
rect 1131 2532 1139 2566
rect 1173 2532 1183 2566
rect 1131 2499 1183 2532
rect 1301 2661 1353 2673
rect 1301 2627 1311 2661
rect 1345 2627 1353 2661
rect 1301 2566 1353 2627
rect 1301 2532 1311 2566
rect 1345 2532 1353 2566
rect 1301 2499 1353 2532
rect 1407 2661 1459 2673
rect 1407 2627 1415 2661
rect 1449 2627 1459 2661
rect 1407 2566 1459 2627
rect 1407 2532 1415 2566
rect 1449 2532 1459 2566
rect 1407 2499 1459 2532
rect 1577 2661 1629 2673
rect 1577 2627 1587 2661
rect 1621 2627 1629 2661
rect 1577 2566 1629 2627
rect 1577 2532 1587 2566
rect 1621 2532 1629 2566
rect 1683 2653 1735 2667
rect 1683 2619 1691 2653
rect 1725 2619 1735 2653
rect 1683 2585 1735 2619
rect 1683 2551 1691 2585
rect 1725 2551 1735 2585
rect 1683 2539 1735 2551
rect 1765 2637 1819 2667
rect 1765 2603 1775 2637
rect 1809 2603 1819 2637
rect 1765 2539 1819 2603
rect 1849 2653 1901 2667
rect 1849 2619 1859 2653
rect 1893 2619 1901 2653
rect 1849 2585 1901 2619
rect 2034 2661 2086 2673
rect 2034 2627 2042 2661
rect 2076 2627 2086 2661
rect 2034 2589 2086 2627
rect 2116 2653 2178 2673
rect 2116 2619 2126 2653
rect 2160 2619 2178 2653
rect 2116 2589 2178 2619
rect 2208 2659 2277 2673
rect 2208 2625 2219 2659
rect 2253 2625 2277 2659
rect 2208 2589 2277 2625
rect 2307 2635 2417 2673
rect 2307 2601 2373 2635
rect 2407 2601 2417 2635
rect 2307 2589 2417 2601
rect 2447 2651 2514 2673
rect 2447 2617 2470 2651
rect 2504 2617 2514 2651
rect 2447 2589 2514 2617
rect 2544 2635 2596 2673
rect 2544 2601 2554 2635
rect 2588 2601 2596 2635
rect 2544 2589 2596 2601
rect 2659 2661 2711 2673
rect 2659 2627 2667 2661
rect 2701 2627 2711 2661
rect 1849 2551 1859 2585
rect 1893 2551 1901 2585
rect 1849 2539 1901 2551
rect 1577 2499 1629 2532
rect 2659 2505 2711 2627
rect 2741 2653 2810 2673
rect 2741 2619 2755 2653
rect 2789 2619 2810 2653
rect 2741 2589 2810 2619
rect 2840 2660 2896 2673
rect 2840 2626 2852 2660
rect 2886 2626 2896 2660
rect 2840 2589 2896 2626
rect 2926 2589 2980 2673
rect 3010 2661 3088 2673
rect 3010 2627 3044 2661
rect 3078 2627 3088 2661
rect 3010 2589 3088 2627
rect 3118 2635 3172 2673
rect 3118 2601 3128 2635
rect 3162 2601 3172 2635
rect 3118 2589 3172 2601
rect 3202 2661 3256 2673
rect 3202 2627 3214 2661
rect 3248 2627 3256 2661
rect 3202 2589 3256 2627
rect 3321 2661 3387 2673
rect 3321 2627 3343 2661
rect 3377 2627 3387 2661
rect 3321 2593 3387 2627
rect 2741 2505 2795 2589
rect 3321 2559 3343 2593
rect 3377 2559 3387 2593
rect 3321 2545 3387 2559
rect 3337 2473 3387 2545
rect 3417 2625 3469 2673
rect 3799 2661 3851 2673
rect 3417 2591 3427 2625
rect 3461 2591 3469 2625
rect 3417 2557 3469 2591
rect 3417 2523 3427 2557
rect 3461 2523 3469 2557
rect 3417 2473 3469 2523
rect 3799 2627 3807 2661
rect 3841 2627 3851 2661
rect 3799 2559 3851 2627
rect 3799 2525 3807 2559
rect 3841 2525 3851 2559
rect 3799 2499 3851 2525
rect 4061 2661 4113 2673
rect 4061 2627 4071 2661
rect 4105 2627 4113 2661
rect 4061 2559 4113 2627
rect 4061 2525 4071 2559
rect 4105 2525 4113 2559
rect 4259 2653 4311 2667
rect 4259 2619 4267 2653
rect 4301 2619 4311 2653
rect 4259 2585 4311 2619
rect 4259 2551 4267 2585
rect 4301 2551 4311 2585
rect 4259 2539 4311 2551
rect 4341 2637 4395 2667
rect 4341 2603 4351 2637
rect 4385 2603 4395 2637
rect 4341 2539 4395 2603
rect 4425 2653 4477 2667
rect 4425 2619 4435 2653
rect 4469 2619 4477 2653
rect 4425 2585 4477 2619
rect 4610 2661 4662 2673
rect 4610 2627 4618 2661
rect 4652 2627 4662 2661
rect 4610 2589 4662 2627
rect 4692 2653 4754 2673
rect 4692 2619 4702 2653
rect 4736 2619 4754 2653
rect 4692 2589 4754 2619
rect 4784 2659 4853 2673
rect 4784 2625 4795 2659
rect 4829 2625 4853 2659
rect 4784 2589 4853 2625
rect 4883 2635 4993 2673
rect 4883 2601 4949 2635
rect 4983 2601 4993 2635
rect 4883 2589 4993 2601
rect 5023 2651 5090 2673
rect 5023 2617 5046 2651
rect 5080 2617 5090 2651
rect 5023 2589 5090 2617
rect 5120 2635 5172 2673
rect 5120 2601 5130 2635
rect 5164 2601 5172 2635
rect 5120 2589 5172 2601
rect 5235 2661 5287 2673
rect 5235 2627 5243 2661
rect 5277 2627 5287 2661
rect 4425 2551 4435 2585
rect 4469 2551 4477 2585
rect 4425 2539 4477 2551
rect 4061 2499 4113 2525
rect 5235 2505 5287 2627
rect 5317 2653 5386 2673
rect 5317 2619 5331 2653
rect 5365 2619 5386 2653
rect 5317 2589 5386 2619
rect 5416 2660 5472 2673
rect 5416 2626 5428 2660
rect 5462 2626 5472 2660
rect 5416 2589 5472 2626
rect 5502 2589 5556 2673
rect 5586 2661 5664 2673
rect 5586 2627 5620 2661
rect 5654 2627 5664 2661
rect 5586 2589 5664 2627
rect 5694 2635 5748 2673
rect 5694 2601 5704 2635
rect 5738 2601 5748 2635
rect 5694 2589 5748 2601
rect 5778 2661 5832 2673
rect 5778 2627 5790 2661
rect 5824 2627 5832 2661
rect 5778 2589 5832 2627
rect 5897 2661 5963 2673
rect 5897 2627 5919 2661
rect 5953 2627 5963 2661
rect 5897 2593 5963 2627
rect 5317 2505 5371 2589
rect 5897 2559 5919 2593
rect 5953 2559 5963 2593
rect 5897 2545 5963 2559
rect 5913 2473 5963 2545
rect 5993 2625 6045 2673
rect 6375 2661 6427 2673
rect 5993 2591 6003 2625
rect 6037 2591 6045 2625
rect 5993 2557 6045 2591
rect 5993 2523 6003 2557
rect 6037 2523 6045 2557
rect 5993 2473 6045 2523
rect 6375 2627 6383 2661
rect 6417 2627 6427 2661
rect 6375 2499 6427 2627
rect 7373 2661 7425 2673
rect 7373 2627 7383 2661
rect 7417 2627 7425 2661
rect 7373 2499 7425 2627
rect 7479 2661 7531 2673
rect 7479 2627 7487 2661
rect 7521 2627 7531 2661
rect 7479 2499 7531 2627
rect 8477 2661 8529 2673
rect 8477 2627 8487 2661
rect 8521 2627 8529 2661
rect 8477 2499 8529 2627
rect 8583 2661 8635 2673
rect 8583 2627 8591 2661
rect 8625 2627 8635 2661
rect 8583 2566 8635 2627
rect 8583 2532 8591 2566
rect 8625 2532 8635 2566
rect 8583 2499 8635 2532
rect 8753 2661 8805 2673
rect 8753 2627 8763 2661
rect 8797 2627 8805 2661
rect 8753 2566 8805 2627
rect 8753 2532 8763 2566
rect 8797 2532 8805 2566
rect 8753 2499 8805 2532
rect 9135 2625 9187 2673
rect 9135 2591 9143 2625
rect 9177 2591 9187 2625
rect 9135 2557 9187 2591
rect 9135 2523 9143 2557
rect 9177 2523 9187 2557
rect 9135 2473 9187 2523
rect 9217 2661 9283 2673
rect 9217 2627 9227 2661
rect 9261 2627 9283 2661
rect 9217 2593 9283 2627
rect 9217 2559 9227 2593
rect 9261 2559 9283 2593
rect 9348 2661 9402 2673
rect 9348 2627 9356 2661
rect 9390 2627 9402 2661
rect 9348 2589 9402 2627
rect 9432 2635 9486 2673
rect 9432 2601 9442 2635
rect 9476 2601 9486 2635
rect 9432 2589 9486 2601
rect 9516 2661 9594 2673
rect 9516 2627 9526 2661
rect 9560 2627 9594 2661
rect 9516 2589 9594 2627
rect 9624 2589 9678 2673
rect 9708 2660 9764 2673
rect 9708 2626 9718 2660
rect 9752 2626 9764 2660
rect 9708 2589 9764 2626
rect 9794 2653 9863 2673
rect 9794 2619 9815 2653
rect 9849 2619 9863 2653
rect 9794 2589 9863 2619
rect 9217 2545 9283 2559
rect 9217 2473 9267 2545
rect 9809 2505 9863 2589
rect 9893 2661 9945 2673
rect 9893 2627 9903 2661
rect 9937 2627 9945 2661
rect 9893 2505 9945 2627
rect 10008 2635 10060 2673
rect 10008 2601 10016 2635
rect 10050 2601 10060 2635
rect 10008 2589 10060 2601
rect 10090 2651 10157 2673
rect 10090 2617 10100 2651
rect 10134 2617 10157 2651
rect 10090 2589 10157 2617
rect 10187 2635 10297 2673
rect 10187 2601 10197 2635
rect 10231 2601 10297 2635
rect 10187 2589 10297 2601
rect 10327 2659 10396 2673
rect 10327 2625 10351 2659
rect 10385 2625 10396 2659
rect 10327 2589 10396 2625
rect 10426 2653 10488 2673
rect 10426 2619 10444 2653
rect 10478 2619 10488 2653
rect 10426 2589 10488 2619
rect 10518 2661 10570 2673
rect 10518 2627 10528 2661
rect 10562 2627 10570 2661
rect 10518 2589 10570 2627
rect 10703 2653 10755 2667
rect 10703 2619 10711 2653
rect 10745 2619 10755 2653
rect 10703 2585 10755 2619
rect 10703 2551 10711 2585
rect 10745 2551 10755 2585
rect 10703 2539 10755 2551
rect 10785 2637 10839 2667
rect 10785 2603 10795 2637
rect 10829 2603 10839 2637
rect 10785 2539 10839 2603
rect 10869 2653 10921 2667
rect 10869 2619 10879 2653
rect 10913 2619 10921 2653
rect 10869 2585 10921 2619
rect 10869 2551 10879 2585
rect 10913 2551 10921 2585
rect 10869 2539 10921 2551
rect 10975 2661 11027 2673
rect 10975 2627 10983 2661
rect 11017 2627 11027 2661
rect 10975 2559 11027 2627
rect 10975 2525 10983 2559
rect 11017 2525 11027 2559
rect 10975 2499 11027 2525
rect 11237 2661 11289 2673
rect 11237 2627 11247 2661
rect 11281 2627 11289 2661
rect 11527 2661 11579 2673
rect 11237 2559 11289 2627
rect 11237 2525 11247 2559
rect 11281 2525 11289 2559
rect 11237 2499 11289 2525
rect 11527 2627 11535 2661
rect 11569 2627 11579 2661
rect 11527 2559 11579 2627
rect 11527 2525 11535 2559
rect 11569 2525 11579 2559
rect 11527 2499 11579 2525
rect 11789 2661 11841 2673
rect 11789 2627 11799 2661
rect 11833 2627 11841 2661
rect 11789 2559 11841 2627
rect 11789 2525 11799 2559
rect 11833 2525 11841 2559
rect 11789 2499 11841 2525
rect 11987 2625 12039 2673
rect 11987 2591 11995 2625
rect 12029 2591 12039 2625
rect 11987 2557 12039 2591
rect 11987 2523 11995 2557
rect 12029 2523 12039 2557
rect 11987 2473 12039 2523
rect 12069 2661 12135 2673
rect 12069 2627 12079 2661
rect 12113 2627 12135 2661
rect 12069 2593 12135 2627
rect 12069 2559 12079 2593
rect 12113 2559 12135 2593
rect 12200 2661 12254 2673
rect 12200 2627 12208 2661
rect 12242 2627 12254 2661
rect 12200 2589 12254 2627
rect 12284 2635 12338 2673
rect 12284 2601 12294 2635
rect 12328 2601 12338 2635
rect 12284 2589 12338 2601
rect 12368 2661 12446 2673
rect 12368 2627 12378 2661
rect 12412 2627 12446 2661
rect 12368 2589 12446 2627
rect 12476 2589 12530 2673
rect 12560 2660 12616 2673
rect 12560 2626 12570 2660
rect 12604 2626 12616 2660
rect 12560 2589 12616 2626
rect 12646 2653 12715 2673
rect 12646 2619 12667 2653
rect 12701 2619 12715 2653
rect 12646 2589 12715 2619
rect 12069 2545 12135 2559
rect 12069 2473 12119 2545
rect 12661 2505 12715 2589
rect 12745 2661 12797 2673
rect 12745 2627 12755 2661
rect 12789 2627 12797 2661
rect 12745 2505 12797 2627
rect 12860 2635 12912 2673
rect 12860 2601 12868 2635
rect 12902 2601 12912 2635
rect 12860 2589 12912 2601
rect 12942 2651 13009 2673
rect 12942 2617 12952 2651
rect 12986 2617 13009 2651
rect 12942 2589 13009 2617
rect 13039 2635 13149 2673
rect 13039 2601 13049 2635
rect 13083 2601 13149 2635
rect 13039 2589 13149 2601
rect 13179 2659 13248 2673
rect 13179 2625 13203 2659
rect 13237 2625 13248 2659
rect 13179 2589 13248 2625
rect 13278 2653 13340 2673
rect 13278 2619 13296 2653
rect 13330 2619 13340 2653
rect 13278 2589 13340 2619
rect 13370 2661 13422 2673
rect 13370 2627 13380 2661
rect 13414 2627 13422 2661
rect 13370 2589 13422 2627
rect 13555 2653 13607 2667
rect 13555 2619 13563 2653
rect 13597 2619 13607 2653
rect 13555 2585 13607 2619
rect 13555 2551 13563 2585
rect 13597 2551 13607 2585
rect 13555 2539 13607 2551
rect 13637 2637 13691 2667
rect 13637 2603 13647 2637
rect 13681 2603 13691 2637
rect 13637 2539 13691 2603
rect 13721 2653 13773 2667
rect 13721 2619 13731 2653
rect 13765 2619 13773 2653
rect 13721 2585 13773 2619
rect 13721 2551 13731 2585
rect 13765 2551 13773 2585
rect 13721 2539 13773 2551
rect 14287 2625 14339 2673
rect 14287 2591 14295 2625
rect 14329 2591 14339 2625
rect 14287 2557 14339 2591
rect 14287 2523 14295 2557
rect 14329 2523 14339 2557
rect 14287 2473 14339 2523
rect 14369 2661 14435 2673
rect 14369 2627 14379 2661
rect 14413 2627 14435 2661
rect 14369 2593 14435 2627
rect 14369 2559 14379 2593
rect 14413 2559 14435 2593
rect 14500 2661 14554 2673
rect 14500 2627 14508 2661
rect 14542 2627 14554 2661
rect 14500 2589 14554 2627
rect 14584 2635 14638 2673
rect 14584 2601 14594 2635
rect 14628 2601 14638 2635
rect 14584 2589 14638 2601
rect 14668 2661 14746 2673
rect 14668 2627 14678 2661
rect 14712 2627 14746 2661
rect 14668 2589 14746 2627
rect 14776 2589 14830 2673
rect 14860 2660 14916 2673
rect 14860 2626 14870 2660
rect 14904 2626 14916 2660
rect 14860 2589 14916 2626
rect 14946 2653 15015 2673
rect 14946 2619 14967 2653
rect 15001 2619 15015 2653
rect 14946 2589 15015 2619
rect 14369 2545 14435 2559
rect 14369 2473 14419 2545
rect 14961 2505 15015 2589
rect 15045 2661 15097 2673
rect 15045 2627 15055 2661
rect 15089 2627 15097 2661
rect 15045 2505 15097 2627
rect 15160 2635 15212 2673
rect 15160 2601 15168 2635
rect 15202 2601 15212 2635
rect 15160 2589 15212 2601
rect 15242 2651 15309 2673
rect 15242 2617 15252 2651
rect 15286 2617 15309 2651
rect 15242 2589 15309 2617
rect 15339 2635 15449 2673
rect 15339 2601 15349 2635
rect 15383 2601 15449 2635
rect 15339 2589 15449 2601
rect 15479 2659 15548 2673
rect 15479 2625 15503 2659
rect 15537 2625 15548 2659
rect 15479 2589 15548 2625
rect 15578 2653 15640 2673
rect 15578 2619 15596 2653
rect 15630 2619 15640 2653
rect 15578 2589 15640 2619
rect 15670 2661 15722 2673
rect 15670 2627 15680 2661
rect 15714 2627 15722 2661
rect 15670 2589 15722 2627
rect 15855 2653 15907 2667
rect 15855 2619 15863 2653
rect 15897 2619 15907 2653
rect 15855 2585 15907 2619
rect 15855 2551 15863 2585
rect 15897 2551 15907 2585
rect 15855 2539 15907 2551
rect 15937 2637 15991 2667
rect 15937 2603 15947 2637
rect 15981 2603 15991 2637
rect 15937 2539 15991 2603
rect 16021 2653 16073 2667
rect 16021 2619 16031 2653
rect 16065 2619 16073 2653
rect 16021 2585 16073 2619
rect 16021 2551 16031 2585
rect 16065 2551 16073 2585
rect 16021 2539 16073 2551
rect 16127 2661 16179 2673
rect 16127 2627 16135 2661
rect 16169 2627 16179 2661
rect 16127 2559 16179 2627
rect 16127 2525 16135 2559
rect 16169 2525 16179 2559
rect 16127 2499 16179 2525
rect 16389 2661 16441 2673
rect 16389 2627 16399 2661
rect 16433 2627 16441 2661
rect 16679 2661 16731 2673
rect 16389 2559 16441 2627
rect 16389 2525 16399 2559
rect 16433 2525 16441 2559
rect 16389 2499 16441 2525
rect 16679 2627 16687 2661
rect 16721 2627 16731 2661
rect 16679 2559 16731 2627
rect 16679 2525 16687 2559
rect 16721 2525 16731 2559
rect 16679 2499 16731 2525
rect 17309 2661 17361 2673
rect 17604 2665 17654 2673
rect 17309 2627 17319 2661
rect 17353 2627 17361 2661
rect 17309 2559 17361 2627
rect 17309 2525 17319 2559
rect 17353 2525 17361 2559
rect 17507 2653 17559 2665
rect 17507 2619 17515 2653
rect 17549 2619 17559 2653
rect 17507 2585 17559 2619
rect 17507 2551 17515 2585
rect 17549 2551 17559 2585
rect 17507 2537 17559 2551
rect 17589 2653 17654 2665
rect 17589 2619 17608 2653
rect 17642 2619 17654 2653
rect 17589 2585 17654 2619
rect 17589 2551 17608 2585
rect 17642 2551 17654 2585
rect 17589 2537 17654 2551
rect 17309 2499 17361 2525
rect 17604 2473 17654 2537
rect 17684 2637 17738 2673
rect 17684 2603 17694 2637
rect 17728 2603 17738 2637
rect 17684 2556 17738 2603
rect 17684 2522 17694 2556
rect 17728 2522 17738 2556
rect 17684 2473 17738 2522
rect 17768 2661 17821 2673
rect 17768 2627 17778 2661
rect 17812 2627 17821 2661
rect 17768 2593 17821 2627
rect 17768 2559 17778 2593
rect 17812 2559 17821 2593
rect 17768 2525 17821 2559
rect 17768 2491 17778 2525
rect 17812 2491 17821 2525
rect 17875 2661 17927 2673
rect 17875 2627 17883 2661
rect 17917 2627 17927 2661
rect 17875 2559 17927 2627
rect 17875 2525 17883 2559
rect 17917 2525 17927 2559
rect 17875 2499 17927 2525
rect 18505 2661 18557 2673
rect 18505 2627 18515 2661
rect 18549 2627 18557 2661
rect 18505 2559 18557 2627
rect 18505 2525 18515 2559
rect 18549 2525 18557 2559
rect 18505 2499 18557 2525
rect 18611 2661 18663 2673
rect 18611 2627 18619 2661
rect 18653 2627 18663 2661
rect 18611 2566 18663 2627
rect 18611 2532 18619 2566
rect 18653 2532 18663 2566
rect 18611 2499 18663 2532
rect 18781 2661 18833 2673
rect 18781 2627 18791 2661
rect 18825 2627 18833 2661
rect 18781 2566 18833 2627
rect 18781 2532 18791 2566
rect 18825 2532 18833 2566
rect 18781 2499 18833 2532
rect 17768 2473 17821 2491
<< ndiffc >>
rect 1139 7502 1173 7536
rect 1311 7502 1345 7536
rect 1600 7519 1634 7553
rect 1600 7451 1634 7485
rect 1684 7493 1718 7527
rect 1770 7523 1804 7557
rect 1863 7510 1897 7544
rect 1967 7504 2001 7538
rect 2967 7504 3001 7538
rect 3071 7504 3105 7538
rect 3519 7504 3553 7538
rect 3992 7519 4026 7553
rect 3992 7451 4026 7485
rect 4076 7493 4110 7527
rect 4162 7523 4196 7557
rect 4255 7510 4289 7544
rect 4359 7504 4393 7538
rect 5359 7504 5393 7538
rect 5648 7519 5682 7553
rect 5648 7451 5682 7485
rect 5732 7493 5766 7527
rect 5818 7523 5852 7557
rect 5911 7510 5945 7544
rect 6015 7502 6049 7536
rect 6187 7502 6221 7536
rect 6383 7504 6417 7538
rect 7383 7504 7417 7538
rect 7487 7497 7521 7531
rect 7751 7497 7785 7531
rect 7856 7519 7890 7553
rect 7856 7451 7890 7485
rect 7940 7493 7974 7527
rect 8026 7523 8060 7557
rect 8119 7510 8153 7544
rect 8223 7504 8257 7538
rect 8671 7504 8705 7538
rect 8959 7504 8993 7538
rect 9407 7504 9441 7538
rect 9695 7497 9729 7531
rect 9959 7497 9993 7531
rect 10063 7515 10097 7549
rect 10149 7519 10183 7553
rect 10243 7515 10277 7549
rect 10327 7519 10361 7553
rect 10431 7504 10465 7538
rect 11063 7504 11097 7538
rect 11167 7502 11201 7536
rect 11339 7502 11373 7536
rect 11535 7504 11569 7538
rect 12167 7504 12201 7538
rect 12271 7510 12305 7544
rect 12364 7523 12398 7557
rect 12450 7493 12484 7527
rect 12534 7519 12568 7553
rect 12534 7451 12568 7485
rect 12639 7504 12673 7538
rect 13639 7504 13673 7538
rect 13743 7502 13777 7536
rect 13915 7502 13949 7536
rect 14111 7497 14145 7531
rect 14375 7497 14409 7531
rect 14479 7510 14513 7544
rect 14572 7523 14606 7557
rect 14658 7493 14692 7527
rect 14742 7519 14776 7553
rect 14742 7451 14776 7485
rect 14847 7504 14881 7538
rect 15847 7504 15881 7538
rect 15951 7504 15985 7538
rect 16399 7504 16433 7538
rect 16871 7510 16905 7544
rect 16964 7523 16998 7557
rect 17050 7493 17084 7527
rect 17134 7519 17168 7553
rect 17134 7451 17168 7485
rect 17239 7504 17273 7538
rect 17871 7504 17905 7538
rect 18067 7510 18101 7544
rect 18160 7523 18194 7557
rect 18246 7493 18280 7527
rect 18330 7519 18364 7553
rect 18330 7451 18364 7485
rect 18619 7502 18653 7536
rect 18791 7502 18825 7536
rect 1139 6608 1173 6642
rect 1311 6608 1345 6642
rect 1415 6606 1449 6640
rect 2415 6606 2449 6640
rect 2519 6606 2553 6640
rect 3519 6606 3553 6640
rect 3807 6606 3841 6640
rect 4807 6606 4841 6640
rect 4911 6606 4945 6640
rect 5911 6606 5945 6640
rect 6015 6606 6049 6640
rect 7015 6606 7049 6640
rect 7119 6606 7153 6640
rect 8119 6606 8153 6640
rect 8223 6606 8257 6640
rect 8671 6606 8705 6640
rect 8959 6606 8993 6640
rect 9959 6606 9993 6640
rect 10063 6606 10097 6640
rect 11063 6606 11097 6640
rect 11167 6606 11201 6640
rect 12167 6606 12201 6640
rect 12271 6606 12305 6640
rect 13271 6606 13305 6640
rect 13375 6606 13409 6640
rect 13823 6606 13857 6640
rect 14111 6606 14145 6640
rect 15111 6606 15145 6640
rect 15215 6606 15249 6640
rect 16215 6606 16249 6640
rect 16319 6606 16353 6640
rect 17319 6606 17353 6640
rect 17423 6606 17457 6640
rect 18423 6606 18457 6640
rect 18619 6608 18653 6642
rect 18791 6608 18825 6642
rect 1139 6414 1173 6448
rect 1311 6414 1345 6448
rect 1415 6416 1449 6450
rect 2415 6416 2449 6450
rect 2519 6416 2553 6450
rect 3519 6416 3553 6450
rect 3623 6416 3657 6450
rect 4623 6416 4657 6450
rect 4727 6416 4761 6450
rect 5727 6416 5761 6450
rect 5831 6409 5865 6443
rect 6095 6409 6129 6443
rect 6383 6416 6417 6450
rect 7383 6416 7417 6450
rect 7487 6416 7521 6450
rect 7935 6416 7969 6450
rect 8068 6425 8102 6459
rect 8152 6425 8186 6459
rect 8248 6425 8282 6459
rect 8333 6433 8367 6467
rect 8333 6365 8367 6399
rect 8499 6416 8533 6450
rect 9499 6416 9533 6450
rect 9603 6416 9637 6450
rect 10603 6416 10637 6450
rect 10707 6416 10741 6450
rect 11339 6416 11373 6450
rect 11535 6416 11569 6450
rect 12535 6416 12569 6450
rect 12639 6416 12673 6450
rect 13639 6416 13673 6450
rect 13743 6416 13777 6450
rect 14743 6416 14777 6450
rect 14847 6416 14881 6450
rect 15847 6416 15881 6450
rect 15951 6416 15985 6450
rect 16399 6416 16433 6450
rect 16687 6416 16721 6450
rect 17687 6416 17721 6450
rect 17791 6416 17825 6450
rect 18423 6416 18457 6450
rect 18619 6414 18653 6448
rect 18791 6414 18825 6448
rect 1139 5520 1173 5554
rect 1311 5520 1345 5554
rect 1415 5518 1449 5552
rect 2415 5518 2449 5552
rect 2519 5518 2553 5552
rect 3519 5518 3553 5552
rect 3807 5518 3841 5552
rect 4807 5518 4841 5552
rect 4911 5518 4945 5552
rect 5911 5518 5945 5552
rect 6015 5518 6049 5552
rect 6647 5518 6681 5552
rect 6751 5529 6785 5563
rect 6837 5499 6871 5533
rect 6923 5512 6957 5546
rect 7027 5518 7061 5552
rect 7475 5518 7509 5552
rect 7625 5514 7659 5548
rect 7709 5514 7743 5548
rect 7777 5514 7811 5548
rect 8012 5514 8046 5548
rect 8219 5499 8253 5533
rect 8303 5518 8337 5552
rect 8407 5525 8441 5559
rect 8671 5525 8705 5559
rect 8959 5518 8993 5552
rect 9959 5518 9993 5552
rect 10063 5518 10097 5552
rect 11063 5518 11097 5552
rect 11167 5525 11201 5559
rect 11431 5525 11465 5559
rect 11564 5509 11598 5543
rect 11648 5509 11682 5543
rect 11744 5509 11778 5543
rect 11829 5569 11863 5603
rect 11829 5501 11863 5535
rect 11995 5518 12029 5552
rect 12627 5518 12661 5552
rect 12852 5509 12886 5543
rect 12936 5509 12970 5543
rect 13032 5509 13066 5543
rect 13117 5569 13151 5603
rect 13117 5501 13151 5535
rect 13283 5518 13317 5552
rect 13915 5518 13949 5552
rect 14111 5518 14145 5552
rect 15111 5518 15145 5552
rect 15215 5518 15249 5552
rect 16215 5518 16249 5552
rect 16319 5518 16353 5552
rect 17319 5518 17353 5552
rect 17423 5518 17457 5552
rect 18423 5518 18457 5552
rect 18619 5520 18653 5554
rect 18791 5520 18825 5554
rect 1139 5326 1173 5360
rect 1311 5326 1345 5360
rect 1415 5328 1449 5362
rect 2415 5328 2449 5362
rect 2519 5326 2553 5360
rect 2691 5326 2725 5360
rect 2795 5321 2829 5355
rect 2879 5347 2913 5381
rect 2963 5321 2997 5355
rect 3085 5351 3119 5385
rect 3218 5345 3252 5379
rect 3325 5345 3359 5379
rect 3671 5347 3705 5381
rect 3783 5351 3817 5385
rect 3893 5347 3927 5381
rect 4105 5351 4139 5385
rect 4323 5331 4357 5365
rect 4447 5347 4481 5381
rect 4531 5297 4565 5331
rect 4635 5328 4669 5362
rect 5635 5328 5669 5362
rect 5739 5328 5773 5362
rect 6187 5328 6221 5362
rect 6383 5326 6417 5360
rect 6555 5326 6589 5360
rect 6659 5328 6693 5362
rect 6743 5347 6777 5381
rect 6950 5332 6984 5366
rect 7185 5332 7219 5366
rect 7253 5332 7287 5366
rect 7337 5332 7371 5366
rect 7487 5321 7521 5355
rect 7751 5321 7785 5355
rect 7855 5321 7889 5355
rect 7939 5347 7973 5381
rect 8023 5321 8057 5355
rect 8145 5351 8179 5385
rect 8278 5345 8312 5379
rect 8385 5345 8419 5379
rect 8731 5347 8765 5381
rect 8843 5351 8877 5385
rect 8953 5347 8987 5381
rect 9165 5351 9199 5385
rect 9383 5331 9417 5365
rect 9507 5347 9541 5381
rect 9591 5297 9625 5331
rect 9695 5321 9729 5355
rect 9959 5321 9993 5355
rect 10109 5332 10143 5366
rect 10193 5332 10227 5366
rect 10261 5332 10295 5366
rect 10496 5332 10530 5366
rect 10703 5347 10737 5381
rect 10787 5328 10821 5362
rect 10891 5328 10925 5362
rect 11339 5328 11373 5362
rect 11719 5328 11753 5362
rect 11803 5347 11837 5381
rect 12010 5332 12044 5366
rect 12245 5332 12279 5366
rect 12313 5332 12347 5366
rect 12397 5332 12431 5366
rect 12547 5321 12581 5355
rect 12811 5321 12845 5355
rect 12961 5332 12995 5366
rect 13045 5332 13079 5366
rect 13113 5332 13147 5366
rect 13348 5332 13382 5366
rect 13555 5347 13589 5381
rect 13639 5328 13673 5362
rect 13743 5328 13777 5362
rect 14743 5328 14777 5362
rect 14847 5328 14881 5362
rect 15847 5328 15881 5362
rect 15951 5328 15985 5362
rect 16399 5328 16433 5362
rect 16687 5328 16721 5362
rect 17687 5328 17721 5362
rect 17791 5328 17825 5362
rect 18423 5328 18457 5362
rect 18619 5326 18653 5360
rect 18791 5326 18825 5360
rect 1139 4432 1173 4466
rect 1311 4432 1345 4466
rect 1415 4430 1449 4464
rect 2047 4430 2081 4464
rect 2151 4432 2185 4466
rect 2323 4432 2357 4466
rect 2446 4437 2480 4471
rect 2536 4411 2570 4445
rect 2695 4437 2729 4471
rect 2799 4437 2833 4471
rect 2953 4411 2987 4445
rect 3037 4437 3071 4471
rect 3163 4430 3197 4464
rect 3611 4430 3645 4464
rect 3998 4415 4032 4449
rect 4084 4437 4118 4471
rect 4170 4415 4204 4449
rect 4256 4437 4290 4471
rect 4353 4415 4387 4449
rect 4439 4419 4473 4453
rect 4543 4437 4577 4471
rect 4807 4437 4841 4471
rect 5095 4430 5129 4464
rect 5727 4430 5761 4464
rect 6077 4481 6111 4515
rect 6077 4413 6111 4447
rect 6162 4421 6196 4455
rect 6258 4421 6292 4455
rect 6342 4421 6376 4455
rect 6475 4437 6509 4471
rect 6739 4437 6773 4471
rect 6872 4421 6906 4455
rect 6956 4421 6990 4455
rect 7052 4421 7086 4455
rect 7137 4481 7171 4515
rect 7137 4413 7171 4447
rect 7303 4430 7337 4464
rect 7751 4430 7785 4464
rect 7855 4430 7889 4464
rect 7939 4411 7973 4445
rect 8146 4426 8180 4460
rect 8381 4426 8415 4460
rect 8449 4426 8483 4460
rect 8533 4426 8567 4460
rect 9172 4421 9206 4455
rect 9256 4421 9290 4455
rect 9352 4421 9386 4455
rect 9437 4481 9471 4515
rect 9437 4413 9471 4447
rect 9603 4437 9637 4471
rect 9867 4437 9901 4471
rect 10155 4437 10189 4471
rect 10419 4437 10453 4471
rect 10552 4421 10586 4455
rect 10636 4421 10670 4455
rect 10732 4421 10766 4455
rect 10817 4481 10851 4515
rect 10817 4413 10851 4447
rect 10983 4437 11017 4471
rect 11247 4437 11281 4471
rect 11351 4424 11385 4458
rect 11437 4411 11471 4445
rect 11523 4441 11557 4475
rect 11627 4437 11661 4471
rect 11891 4437 11925 4471
rect 12041 4426 12075 4460
rect 12125 4426 12159 4460
rect 12193 4426 12227 4460
rect 12428 4426 12462 4460
rect 12635 4411 12669 4445
rect 12719 4430 12753 4464
rect 12823 4437 12857 4471
rect 13087 4437 13121 4471
rect 13191 4441 13225 4475
rect 13277 4411 13311 4445
rect 13363 4424 13397 4458
rect 13467 4430 13501 4464
rect 13915 4430 13949 4464
rect 14111 4430 14145 4464
rect 15111 4430 15145 4464
rect 15244 4421 15278 4455
rect 15328 4421 15362 4455
rect 15424 4421 15458 4455
rect 15509 4481 15543 4515
rect 15509 4413 15543 4447
rect 15675 4437 15709 4471
rect 15939 4437 15973 4471
rect 16043 4441 16077 4475
rect 16129 4411 16163 4445
rect 16215 4424 16249 4458
rect 16319 4437 16353 4471
rect 16583 4437 16617 4471
rect 16687 4441 16721 4475
rect 16773 4411 16807 4445
rect 16859 4424 16893 4458
rect 16963 4430 16997 4464
rect 17963 4430 17997 4464
rect 18067 4430 18101 4464
rect 18515 4430 18549 4464
rect 18619 4432 18653 4466
rect 18791 4432 18825 4466
rect 1139 4238 1173 4272
rect 1311 4238 1345 4272
rect 1415 4240 1449 4274
rect 2047 4240 2081 4274
rect 2243 4246 2277 4280
rect 2329 4259 2363 4293
rect 2415 4229 2449 4263
rect 2519 4233 2553 4267
rect 2783 4233 2817 4267
rect 2887 4233 2921 4267
rect 2971 4259 3005 4293
rect 3055 4233 3089 4267
rect 3177 4263 3211 4297
rect 3310 4257 3344 4291
rect 3417 4257 3451 4291
rect 3763 4259 3797 4293
rect 3875 4263 3909 4297
rect 3985 4259 4019 4293
rect 4197 4263 4231 4297
rect 4415 4243 4449 4277
rect 4539 4259 4573 4293
rect 4623 4209 4657 4243
rect 4727 4233 4761 4267
rect 4991 4233 5025 4267
rect 5371 4240 5405 4274
rect 6003 4240 6037 4274
rect 6383 4238 6417 4272
rect 6555 4238 6589 4272
rect 6659 4229 6693 4263
rect 6745 4259 6779 4293
rect 6831 4246 6865 4280
rect 6935 4240 6969 4274
rect 7567 4240 7601 4274
rect 7717 4244 7751 4278
rect 7801 4244 7835 4278
rect 7869 4244 7903 4278
rect 8104 4244 8138 4278
rect 8311 4259 8345 4293
rect 8395 4240 8429 4274
rect 8499 4233 8533 4267
rect 8763 4233 8797 4267
rect 8959 4259 8993 4293
rect 9045 4246 9079 4280
rect 9131 4246 9165 4280
rect 9217 4246 9251 4280
rect 9303 4246 9337 4280
rect 9389 4246 9423 4280
rect 9475 4255 9509 4289
rect 9561 4246 9595 4280
rect 9647 4255 9681 4289
rect 9733 4246 9767 4280
rect 9819 4255 9853 4289
rect 9905 4246 9939 4280
rect 9991 4255 10025 4289
rect 10076 4246 10110 4280
rect 10162 4255 10196 4289
rect 10248 4246 10282 4280
rect 10334 4255 10368 4289
rect 10420 4246 10454 4280
rect 10506 4255 10540 4289
rect 10592 4246 10626 4280
rect 10678 4255 10712 4289
rect 10799 4240 10833 4274
rect 11247 4240 11281 4274
rect 11719 4209 11753 4243
rect 11803 4259 11837 4293
rect 11927 4243 11961 4277
rect 12145 4263 12179 4297
rect 12357 4259 12391 4293
rect 12467 4263 12501 4297
rect 12579 4259 12613 4293
rect 12925 4257 12959 4291
rect 13032 4257 13066 4291
rect 13165 4263 13199 4297
rect 13287 4233 13321 4267
rect 13371 4259 13405 4293
rect 13455 4233 13489 4267
rect 13559 4233 13593 4267
rect 13823 4233 13857 4267
rect 13927 4233 13961 4267
rect 14011 4259 14045 4293
rect 14095 4233 14129 4267
rect 14217 4263 14251 4297
rect 14350 4257 14384 4291
rect 14457 4257 14491 4291
rect 14803 4259 14837 4293
rect 14915 4263 14949 4297
rect 15025 4259 15059 4293
rect 15237 4263 15271 4297
rect 15455 4243 15489 4277
rect 15579 4259 15613 4293
rect 15663 4209 15697 4243
rect 15767 4240 15801 4274
rect 16399 4240 16433 4274
rect 16687 4240 16721 4274
rect 17687 4240 17721 4274
rect 17791 4240 17825 4274
rect 18423 4240 18457 4274
rect 18619 4238 18653 4272
rect 18791 4238 18825 4272
rect 1139 3344 1173 3378
rect 1311 3344 1345 3378
rect 1415 3344 1449 3378
rect 1587 3344 1621 3378
rect 1691 3349 1725 3383
rect 1775 3323 1809 3357
rect 1859 3349 1893 3383
rect 1981 3319 2015 3353
rect 2114 3325 2148 3359
rect 2221 3325 2255 3359
rect 2567 3323 2601 3357
rect 2679 3319 2713 3353
rect 2789 3323 2823 3357
rect 3001 3319 3035 3353
rect 3219 3339 3253 3373
rect 3343 3323 3377 3357
rect 3427 3373 3461 3407
rect 3807 3342 3841 3376
rect 4439 3342 4473 3376
rect 4560 3327 4594 3361
rect 4646 3336 4680 3370
rect 4732 3327 4766 3361
rect 4818 3336 4852 3370
rect 4904 3327 4938 3361
rect 4990 3336 5024 3370
rect 5076 3327 5110 3361
rect 5162 3336 5196 3370
rect 5247 3327 5281 3361
rect 5333 3336 5367 3370
rect 5419 3327 5453 3361
rect 5505 3336 5539 3370
rect 5591 3327 5625 3361
rect 5677 3336 5711 3370
rect 5763 3327 5797 3361
rect 5849 3336 5883 3370
rect 5935 3336 5969 3370
rect 6021 3336 6055 3370
rect 6107 3336 6141 3370
rect 6193 3336 6227 3370
rect 6279 3323 6313 3357
rect 6383 3349 6417 3383
rect 6647 3349 6681 3383
rect 6751 3349 6785 3383
rect 6835 3323 6869 3357
rect 6919 3349 6953 3383
rect 7041 3319 7075 3353
rect 7174 3325 7208 3359
rect 7281 3325 7315 3359
rect 7627 3323 7661 3357
rect 7739 3319 7773 3353
rect 7849 3323 7883 3357
rect 8061 3319 8095 3353
rect 8279 3339 8313 3373
rect 8403 3323 8437 3357
rect 8487 3373 8521 3407
rect 8591 3344 8625 3378
rect 8763 3344 8797 3378
rect 9143 3336 9177 3370
rect 9236 3323 9270 3357
rect 9322 3353 9356 3387
rect 9406 3395 9440 3429
rect 9406 3327 9440 3361
rect 9511 3342 9545 3376
rect 9959 3342 9993 3376
rect 10063 3353 10097 3387
rect 10149 3323 10183 3357
rect 10235 3336 10269 3370
rect 10339 3342 10373 3376
rect 10787 3342 10821 3376
rect 10983 3336 11017 3370
rect 11069 3323 11103 3357
rect 11155 3353 11189 3387
rect 11259 3342 11293 3376
rect 11891 3342 11925 3376
rect 11995 3373 12029 3407
rect 12079 3323 12113 3357
rect 12203 3339 12237 3373
rect 12421 3319 12455 3353
rect 12633 3323 12667 3357
rect 12743 3319 12777 3353
rect 12855 3323 12889 3357
rect 13201 3325 13235 3359
rect 13308 3325 13342 3359
rect 13441 3319 13475 3353
rect 13563 3349 13597 3383
rect 13647 3323 13681 3357
rect 13731 3349 13765 3383
rect 14111 3342 14145 3376
rect 15111 3342 15145 3376
rect 15215 3342 15249 3376
rect 16215 3342 16249 3376
rect 16319 3342 16353 3376
rect 17319 3342 17353 3376
rect 17423 3342 17457 3376
rect 18423 3342 18457 3376
rect 18619 3344 18653 3378
rect 18791 3344 18825 3378
rect 1139 3150 1173 3184
rect 1311 3150 1345 3184
rect 1415 3152 1449 3186
rect 1863 3152 1897 3186
rect 1967 3121 2001 3155
rect 2051 3171 2085 3205
rect 2175 3155 2209 3189
rect 2393 3175 2427 3209
rect 2605 3171 2639 3205
rect 2715 3175 2749 3209
rect 2827 3171 2861 3205
rect 3173 3169 3207 3203
rect 3280 3169 3314 3203
rect 3413 3175 3447 3209
rect 3535 3145 3569 3179
rect 3619 3171 3653 3205
rect 3703 3145 3737 3179
rect 3807 3145 3841 3179
rect 4071 3145 4105 3179
rect 4175 3145 4209 3179
rect 4259 3171 4293 3205
rect 4343 3145 4377 3179
rect 4447 3171 4481 3205
rect 4531 3153 4565 3187
rect 4641 3171 4675 3205
rect 4862 3175 4896 3209
rect 5018 3155 5052 3189
rect 5122 3171 5156 3205
rect 5284 3169 5318 3203
rect 5542 3151 5576 3185
rect 5646 3144 5680 3178
rect 5750 3145 5784 3179
rect 5845 3171 5879 3205
rect 5929 3121 5963 3155
rect 6383 3152 6417 3186
rect 7015 3152 7049 3186
rect 7211 3121 7245 3155
rect 7295 3171 7329 3205
rect 7419 3155 7453 3189
rect 7637 3175 7671 3209
rect 7849 3171 7883 3205
rect 7959 3175 7993 3209
rect 8071 3171 8105 3205
rect 8417 3169 8451 3203
rect 8524 3169 8558 3203
rect 8657 3175 8691 3209
rect 8779 3145 8813 3179
rect 8863 3171 8897 3205
rect 8947 3145 8981 3179
rect 9051 3145 9085 3179
rect 9315 3145 9349 3179
rect 9419 3171 9453 3205
rect 9505 3158 9539 3192
rect 9591 3158 9625 3192
rect 9677 3158 9711 3192
rect 9763 3158 9797 3192
rect 9849 3158 9883 3192
rect 9935 3167 9969 3201
rect 10021 3158 10055 3192
rect 10107 3167 10141 3201
rect 10193 3158 10227 3192
rect 10279 3167 10313 3201
rect 10365 3158 10399 3192
rect 10451 3167 10485 3201
rect 10536 3158 10570 3192
rect 10622 3167 10656 3201
rect 10708 3158 10742 3192
rect 10794 3167 10828 3201
rect 10880 3158 10914 3192
rect 10966 3167 11000 3201
rect 11052 3158 11086 3192
rect 11138 3167 11172 3201
rect 11719 3121 11753 3155
rect 11803 3171 11837 3205
rect 11927 3155 11961 3189
rect 12145 3175 12179 3209
rect 12357 3171 12391 3205
rect 12467 3175 12501 3209
rect 12579 3171 12613 3205
rect 12925 3169 12959 3203
rect 13032 3169 13066 3203
rect 13165 3175 13199 3209
rect 13287 3145 13321 3179
rect 13371 3171 13405 3205
rect 13455 3145 13489 3179
rect 13559 3145 13593 3179
rect 13823 3145 13857 3179
rect 13927 3158 13961 3192
rect 14020 3171 14054 3205
rect 14106 3141 14140 3175
rect 14190 3167 14224 3201
rect 14190 3099 14224 3133
rect 14295 3152 14329 3186
rect 15295 3152 15329 3186
rect 15399 3152 15433 3186
rect 16399 3152 16433 3186
rect 16687 3152 16721 3186
rect 17687 3152 17721 3186
rect 17791 3152 17825 3186
rect 18423 3152 18457 3186
rect 18619 3150 18653 3184
rect 18791 3150 18825 3184
rect 1139 2256 1173 2290
rect 1311 2256 1345 2290
rect 1415 2256 1449 2290
rect 1587 2256 1621 2290
rect 1691 2261 1725 2295
rect 1775 2235 1809 2269
rect 1859 2261 1893 2295
rect 1981 2231 2015 2265
rect 2114 2237 2148 2271
rect 2221 2237 2255 2271
rect 2567 2235 2601 2269
rect 2679 2231 2713 2265
rect 2789 2235 2823 2269
rect 3001 2231 3035 2265
rect 3219 2251 3253 2285
rect 3343 2235 3377 2269
rect 3427 2285 3461 2319
rect 3807 2261 3841 2295
rect 4071 2261 4105 2295
rect 4267 2261 4301 2295
rect 4351 2235 4385 2269
rect 4435 2261 4469 2295
rect 4557 2231 4591 2265
rect 4690 2237 4724 2271
rect 4797 2237 4831 2271
rect 5143 2235 5177 2269
rect 5255 2231 5289 2265
rect 5365 2235 5399 2269
rect 5577 2231 5611 2265
rect 5795 2251 5829 2285
rect 5919 2235 5953 2269
rect 6003 2285 6037 2319
rect 6383 2254 6417 2288
rect 7383 2254 7417 2288
rect 7487 2254 7521 2288
rect 8487 2254 8521 2288
rect 8591 2256 8625 2290
rect 8763 2256 8797 2290
rect 9143 2285 9177 2319
rect 9227 2235 9261 2269
rect 9351 2251 9385 2285
rect 9569 2231 9603 2265
rect 9781 2235 9815 2269
rect 9891 2231 9925 2265
rect 10003 2235 10037 2269
rect 10349 2237 10383 2271
rect 10456 2237 10490 2271
rect 10589 2231 10623 2265
rect 10711 2261 10745 2295
rect 10795 2235 10829 2269
rect 10879 2261 10913 2295
rect 10983 2261 11017 2295
rect 11247 2261 11281 2295
rect 11535 2261 11569 2295
rect 11799 2261 11833 2295
rect 11995 2285 12029 2319
rect 12079 2235 12113 2269
rect 12203 2251 12237 2285
rect 12421 2231 12455 2265
rect 12633 2235 12667 2269
rect 12743 2231 12777 2265
rect 12855 2235 12889 2269
rect 13201 2237 13235 2271
rect 13308 2237 13342 2271
rect 13441 2231 13475 2265
rect 13563 2261 13597 2295
rect 13647 2235 13681 2269
rect 13731 2261 13765 2295
rect 14295 2285 14329 2319
rect 14379 2235 14413 2269
rect 14503 2251 14537 2285
rect 14721 2231 14755 2265
rect 14933 2235 14967 2269
rect 15043 2231 15077 2265
rect 15155 2235 15189 2269
rect 15501 2237 15535 2271
rect 15608 2237 15642 2271
rect 15741 2231 15775 2265
rect 15863 2261 15897 2295
rect 15947 2235 15981 2269
rect 16031 2261 16065 2295
rect 16135 2261 16169 2295
rect 16399 2261 16433 2295
rect 16687 2254 16721 2288
rect 17319 2254 17353 2288
rect 17515 2248 17549 2282
rect 17608 2235 17642 2269
rect 17694 2265 17728 2299
rect 17778 2307 17812 2341
rect 17778 2239 17812 2273
rect 17883 2254 17917 2288
rect 18515 2254 18549 2288
rect 18619 2256 18653 2290
rect 18791 2256 18825 2290
<< pdiffc >>
rect 1139 7226 1173 7260
rect 1139 7131 1173 7165
rect 1311 7226 1345 7260
rect 1311 7131 1345 7165
rect 1600 7267 1634 7301
rect 1600 7199 1634 7233
rect 1600 7131 1634 7165
rect 1684 7236 1718 7270
rect 1684 7155 1718 7189
rect 1770 7207 1804 7241
rect 1770 7139 1804 7173
rect 1863 7207 1897 7241
rect 1863 7139 1897 7173
rect 1967 7131 2001 7165
rect 2967 7131 3001 7165
rect 3071 7233 3105 7267
rect 3071 7131 3105 7165
rect 3519 7233 3553 7267
rect 3519 7131 3553 7165
rect 3992 7267 4026 7301
rect 3992 7199 4026 7233
rect 3992 7131 4026 7165
rect 4076 7236 4110 7270
rect 4076 7155 4110 7189
rect 4162 7207 4196 7241
rect 4162 7139 4196 7173
rect 4255 7207 4289 7241
rect 4255 7139 4289 7173
rect 4359 7131 4393 7165
rect 5359 7131 5393 7165
rect 5648 7267 5682 7301
rect 5648 7199 5682 7233
rect 5648 7131 5682 7165
rect 5732 7236 5766 7270
rect 5732 7155 5766 7189
rect 5818 7207 5852 7241
rect 5818 7139 5852 7173
rect 5911 7207 5945 7241
rect 5911 7139 5945 7173
rect 6015 7226 6049 7260
rect 6015 7131 6049 7165
rect 6187 7226 6221 7260
rect 6187 7131 6221 7165
rect 6383 7131 6417 7165
rect 7383 7131 7417 7165
rect 7487 7233 7521 7267
rect 7487 7131 7521 7165
rect 7751 7233 7785 7267
rect 7751 7131 7785 7165
rect 7856 7267 7890 7301
rect 7856 7199 7890 7233
rect 7856 7131 7890 7165
rect 7940 7236 7974 7270
rect 7940 7155 7974 7189
rect 8026 7207 8060 7241
rect 8026 7139 8060 7173
rect 8119 7207 8153 7241
rect 8119 7139 8153 7173
rect 8223 7233 8257 7267
rect 8223 7131 8257 7165
rect 8671 7233 8705 7267
rect 8671 7131 8705 7165
rect 8959 7233 8993 7267
rect 8959 7131 8993 7165
rect 9407 7233 9441 7267
rect 9407 7131 9441 7165
rect 9695 7233 9729 7267
rect 9695 7131 9729 7165
rect 9959 7233 9993 7267
rect 9959 7131 9993 7165
rect 10063 7250 10097 7284
rect 10063 7145 10097 7179
rect 10149 7211 10183 7245
rect 10149 7143 10183 7177
rect 10243 7145 10277 7179
rect 10327 7140 10361 7174
rect 10431 7233 10465 7267
rect 10431 7131 10465 7165
rect 11063 7233 11097 7267
rect 11063 7131 11097 7165
rect 11167 7226 11201 7260
rect 11167 7131 11201 7165
rect 11339 7226 11373 7260
rect 11339 7131 11373 7165
rect 11535 7233 11569 7267
rect 11535 7131 11569 7165
rect 12167 7233 12201 7267
rect 12167 7131 12201 7165
rect 12271 7207 12305 7241
rect 12271 7139 12305 7173
rect 12364 7207 12398 7241
rect 12364 7139 12398 7173
rect 12450 7236 12484 7270
rect 12450 7155 12484 7189
rect 12534 7267 12568 7301
rect 12534 7199 12568 7233
rect 12534 7131 12568 7165
rect 12639 7131 12673 7165
rect 13639 7131 13673 7165
rect 13743 7226 13777 7260
rect 13743 7131 13777 7165
rect 13915 7226 13949 7260
rect 13915 7131 13949 7165
rect 14111 7233 14145 7267
rect 14111 7131 14145 7165
rect 14375 7233 14409 7267
rect 14375 7131 14409 7165
rect 14479 7207 14513 7241
rect 14479 7139 14513 7173
rect 14572 7207 14606 7241
rect 14572 7139 14606 7173
rect 14658 7236 14692 7270
rect 14658 7155 14692 7189
rect 14742 7267 14776 7301
rect 14742 7199 14776 7233
rect 14742 7131 14776 7165
rect 14847 7131 14881 7165
rect 15847 7131 15881 7165
rect 15951 7233 15985 7267
rect 15951 7131 15985 7165
rect 16399 7233 16433 7267
rect 16399 7131 16433 7165
rect 16871 7207 16905 7241
rect 16871 7139 16905 7173
rect 16964 7207 16998 7241
rect 16964 7139 16998 7173
rect 17050 7236 17084 7270
rect 17050 7155 17084 7189
rect 17134 7267 17168 7301
rect 17134 7199 17168 7233
rect 17134 7131 17168 7165
rect 17239 7233 17273 7267
rect 17239 7131 17273 7165
rect 17871 7233 17905 7267
rect 17871 7131 17905 7165
rect 18067 7207 18101 7241
rect 18067 7139 18101 7173
rect 18160 7207 18194 7241
rect 18160 7139 18194 7173
rect 18246 7236 18280 7270
rect 18246 7155 18280 7189
rect 18330 7267 18364 7301
rect 18330 7199 18364 7233
rect 18330 7131 18364 7165
rect 18619 7226 18653 7260
rect 18619 7131 18653 7165
rect 18791 7226 18825 7260
rect 18791 7131 18825 7165
rect 1139 6979 1173 7013
rect 1139 6884 1173 6918
rect 1311 6979 1345 7013
rect 1311 6884 1345 6918
rect 1415 6979 1449 7013
rect 2415 6979 2449 7013
rect 2519 6979 2553 7013
rect 3519 6979 3553 7013
rect 3807 6979 3841 7013
rect 4807 6979 4841 7013
rect 4911 6979 4945 7013
rect 5911 6979 5945 7013
rect 6015 6979 6049 7013
rect 7015 6979 7049 7013
rect 7119 6979 7153 7013
rect 8119 6979 8153 7013
rect 8223 6979 8257 7013
rect 8223 6877 8257 6911
rect 8671 6979 8705 7013
rect 8671 6877 8705 6911
rect 8959 6979 8993 7013
rect 9959 6979 9993 7013
rect 10063 6979 10097 7013
rect 11063 6979 11097 7013
rect 11167 6979 11201 7013
rect 12167 6979 12201 7013
rect 12271 6979 12305 7013
rect 13271 6979 13305 7013
rect 13375 6979 13409 7013
rect 13375 6877 13409 6911
rect 13823 6979 13857 7013
rect 13823 6877 13857 6911
rect 14111 6979 14145 7013
rect 15111 6979 15145 7013
rect 15215 6979 15249 7013
rect 16215 6979 16249 7013
rect 16319 6979 16353 7013
rect 17319 6979 17353 7013
rect 17423 6979 17457 7013
rect 18423 6979 18457 7013
rect 18619 6979 18653 7013
rect 18619 6884 18653 6918
rect 18791 6979 18825 7013
rect 18791 6884 18825 6918
rect 1139 6138 1173 6172
rect 1139 6043 1173 6077
rect 1311 6138 1345 6172
rect 1311 6043 1345 6077
rect 1415 6043 1449 6077
rect 2415 6043 2449 6077
rect 2519 6043 2553 6077
rect 3519 6043 3553 6077
rect 3623 6043 3657 6077
rect 4623 6043 4657 6077
rect 4727 6043 4761 6077
rect 5727 6043 5761 6077
rect 5831 6145 5865 6179
rect 5831 6043 5865 6077
rect 6095 6145 6129 6179
rect 6095 6043 6129 6077
rect 6383 6043 6417 6077
rect 7383 6043 7417 6077
rect 7487 6145 7521 6179
rect 7487 6043 7521 6077
rect 7935 6145 7969 6179
rect 8080 6179 8114 6213
rect 8249 6127 8283 6161
rect 7935 6043 7969 6077
rect 8249 6059 8283 6093
rect 8349 6111 8383 6145
rect 8349 6043 8383 6077
rect 8499 6043 8533 6077
rect 9499 6043 9533 6077
rect 9603 6043 9637 6077
rect 10603 6043 10637 6077
rect 10707 6145 10741 6179
rect 10707 6043 10741 6077
rect 11339 6145 11373 6179
rect 11339 6043 11373 6077
rect 11535 6043 11569 6077
rect 12535 6043 12569 6077
rect 12639 6043 12673 6077
rect 13639 6043 13673 6077
rect 13743 6043 13777 6077
rect 14743 6043 14777 6077
rect 14847 6043 14881 6077
rect 15847 6043 15881 6077
rect 15951 6145 15985 6179
rect 15951 6043 15985 6077
rect 16399 6145 16433 6179
rect 16399 6043 16433 6077
rect 16687 6043 16721 6077
rect 17687 6043 17721 6077
rect 17791 6145 17825 6179
rect 17791 6043 17825 6077
rect 18423 6145 18457 6179
rect 18423 6043 18457 6077
rect 18619 6138 18653 6172
rect 18619 6043 18653 6077
rect 18791 6138 18825 6172
rect 18791 6043 18825 6077
rect 1139 5891 1173 5925
rect 1139 5796 1173 5830
rect 1311 5891 1345 5925
rect 1311 5796 1345 5830
rect 1415 5891 1449 5925
rect 2415 5891 2449 5925
rect 2519 5891 2553 5925
rect 3519 5891 3553 5925
rect 3807 5891 3841 5925
rect 4807 5891 4841 5925
rect 4911 5891 4945 5925
rect 5911 5891 5945 5925
rect 6015 5891 6049 5925
rect 6015 5789 6049 5823
rect 6647 5891 6681 5925
rect 6647 5789 6681 5823
rect 6751 5883 6785 5917
rect 6751 5802 6785 5836
rect 6837 5883 6871 5917
rect 6837 5815 6871 5849
rect 6923 5883 6957 5917
rect 6923 5815 6957 5849
rect 7027 5891 7061 5925
rect 7027 5789 7061 5823
rect 7475 5891 7509 5925
rect 7475 5789 7509 5823
rect 7625 5831 7659 5865
rect 7711 5831 7745 5865
rect 7908 5831 7942 5865
rect 7983 5831 8017 5865
rect 8219 5891 8253 5925
rect 8219 5823 8253 5857
rect 8219 5755 8253 5789
rect 8303 5891 8337 5925
rect 8303 5823 8337 5857
rect 8303 5755 8337 5789
rect 8407 5891 8441 5925
rect 8407 5789 8441 5823
rect 8671 5891 8705 5925
rect 8671 5789 8705 5823
rect 8959 5891 8993 5925
rect 9959 5891 9993 5925
rect 10063 5891 10097 5925
rect 11063 5891 11097 5925
rect 11167 5891 11201 5925
rect 11167 5789 11201 5823
rect 11431 5891 11465 5925
rect 11745 5875 11779 5909
rect 11431 5789 11465 5823
rect 11576 5755 11610 5789
rect 11745 5807 11779 5841
rect 11845 5891 11879 5925
rect 11845 5823 11879 5857
rect 11995 5891 12029 5925
rect 11995 5789 12029 5823
rect 12627 5891 12661 5925
rect 13033 5875 13067 5909
rect 12627 5789 12661 5823
rect 12864 5755 12898 5789
rect 13033 5807 13067 5841
rect 13133 5891 13167 5925
rect 13133 5823 13167 5857
rect 13283 5891 13317 5925
rect 13283 5789 13317 5823
rect 13915 5891 13949 5925
rect 13915 5789 13949 5823
rect 14111 5891 14145 5925
rect 15111 5891 15145 5925
rect 15215 5891 15249 5925
rect 16215 5891 16249 5925
rect 16319 5891 16353 5925
rect 17319 5891 17353 5925
rect 17423 5891 17457 5925
rect 18423 5891 18457 5925
rect 18619 5891 18653 5925
rect 18619 5796 18653 5830
rect 18791 5891 18825 5925
rect 18791 5796 18825 5830
rect 1139 5050 1173 5084
rect 1139 4955 1173 4989
rect 1311 5050 1345 5084
rect 1311 4955 1345 4989
rect 1415 4955 1449 4989
rect 2415 4955 2449 4989
rect 2519 5050 2553 5084
rect 2519 4955 2553 4989
rect 2691 5050 2725 5084
rect 2691 4955 2725 4989
rect 2795 5031 2829 5065
rect 2795 4963 2829 4997
rect 2879 4979 2913 5013
rect 2963 5031 2997 5065
rect 2963 4963 2997 4997
rect 3146 4955 3180 4989
rect 3230 4963 3264 4997
rect 3323 4957 3357 4991
rect 3477 4981 3511 5015
rect 3574 4965 3608 4999
rect 3658 4981 3692 5015
rect 3771 4955 3805 4989
rect 3859 4963 3893 4997
rect 3956 4956 3990 4990
rect 4148 4955 4182 4989
rect 4232 4981 4266 5015
rect 4318 4955 4352 4989
rect 4447 5023 4481 5057
rect 4447 4955 4481 4989
rect 4531 5059 4565 5093
rect 4531 4991 4565 5025
rect 4635 4955 4669 4989
rect 5635 4955 5669 4989
rect 5739 5057 5773 5091
rect 5739 4955 5773 4989
rect 6187 5057 6221 5091
rect 6187 4955 6221 4989
rect 6383 5050 6417 5084
rect 6383 4955 6417 4989
rect 6555 5050 6589 5084
rect 6555 4955 6589 4989
rect 6659 5091 6693 5125
rect 6659 5023 6693 5057
rect 6659 4955 6693 4989
rect 6743 5091 6777 5125
rect 6743 5023 6777 5057
rect 6743 4955 6777 4989
rect 6979 5015 7013 5049
rect 7054 5015 7088 5049
rect 7251 5015 7285 5049
rect 7337 5015 7371 5049
rect 7487 5057 7521 5091
rect 7487 4955 7521 4989
rect 7751 5057 7785 5091
rect 7751 4955 7785 4989
rect 7855 5031 7889 5065
rect 7855 4963 7889 4997
rect 7939 4979 7973 5013
rect 8023 5031 8057 5065
rect 8023 4963 8057 4997
rect 8206 4955 8240 4989
rect 8290 4963 8324 4997
rect 8383 4957 8417 4991
rect 8537 4981 8571 5015
rect 8634 4965 8668 4999
rect 8718 4981 8752 5015
rect 8831 4955 8865 4989
rect 8919 4963 8953 4997
rect 9016 4956 9050 4990
rect 9208 4955 9242 4989
rect 9292 4981 9326 5015
rect 9378 4955 9412 4989
rect 9507 5023 9541 5057
rect 9507 4955 9541 4989
rect 9591 5059 9625 5093
rect 9591 4991 9625 5025
rect 9695 5057 9729 5091
rect 9695 4955 9729 4989
rect 9959 5057 9993 5091
rect 10703 5091 10737 5125
rect 9959 4955 9993 4989
rect 10109 5015 10143 5049
rect 10195 5015 10229 5049
rect 10392 5015 10426 5049
rect 10467 5015 10501 5049
rect 10703 5023 10737 5057
rect 10703 4955 10737 4989
rect 10787 5091 10821 5125
rect 10787 5023 10821 5057
rect 10787 4955 10821 4989
rect 10891 5057 10925 5091
rect 10891 4955 10925 4989
rect 11339 5057 11373 5091
rect 11339 4955 11373 4989
rect 11719 5091 11753 5125
rect 11719 5023 11753 5057
rect 11719 4955 11753 4989
rect 11803 5091 11837 5125
rect 11803 5023 11837 5057
rect 11803 4955 11837 4989
rect 12039 5015 12073 5049
rect 12114 5015 12148 5049
rect 12311 5015 12345 5049
rect 12397 5015 12431 5049
rect 12547 5057 12581 5091
rect 12547 4955 12581 4989
rect 12811 5057 12845 5091
rect 13555 5091 13589 5125
rect 12811 4955 12845 4989
rect 12961 5015 12995 5049
rect 13047 5015 13081 5049
rect 13244 5015 13278 5049
rect 13319 5015 13353 5049
rect 13555 5023 13589 5057
rect 13555 4955 13589 4989
rect 13639 5091 13673 5125
rect 13639 5023 13673 5057
rect 13639 4955 13673 4989
rect 13743 4955 13777 4989
rect 14743 4955 14777 4989
rect 14847 4955 14881 4989
rect 15847 4955 15881 4989
rect 15951 5057 15985 5091
rect 15951 4955 15985 4989
rect 16399 5057 16433 5091
rect 16399 4955 16433 4989
rect 16687 4955 16721 4989
rect 17687 4955 17721 4989
rect 17791 5057 17825 5091
rect 17791 4955 17825 4989
rect 18423 5057 18457 5091
rect 18423 4955 18457 4989
rect 18619 5050 18653 5084
rect 18619 4955 18653 4989
rect 18791 5050 18825 5084
rect 18791 4955 18825 4989
rect 1139 4803 1173 4837
rect 1139 4708 1173 4742
rect 1311 4803 1345 4837
rect 1311 4708 1345 4742
rect 1415 4803 1449 4837
rect 1415 4701 1449 4735
rect 2047 4803 2081 4837
rect 2047 4701 2081 4735
rect 2151 4803 2185 4837
rect 2151 4708 2185 4742
rect 2323 4803 2357 4837
rect 2323 4708 2357 4742
rect 2446 4777 2480 4811
rect 2536 4803 2570 4837
rect 2695 4777 2729 4811
rect 2799 4777 2833 4811
rect 2953 4803 2987 4837
rect 3037 4777 3071 4811
rect 3163 4803 3197 4837
rect 3163 4701 3197 4735
rect 3611 4803 3645 4837
rect 3611 4701 3645 4735
rect 3999 4789 4033 4823
rect 3999 4721 4033 4755
rect 4085 4795 4119 4829
rect 4085 4727 4119 4761
rect 4085 4659 4119 4693
rect 4171 4803 4205 4837
rect 4257 4768 4291 4802
rect 4353 4803 4387 4837
rect 4353 4735 4387 4769
rect 4439 4795 4473 4829
rect 4439 4673 4473 4707
rect 4543 4803 4577 4837
rect 4543 4701 4577 4735
rect 4807 4803 4841 4837
rect 4807 4701 4841 4735
rect 5095 4803 5129 4837
rect 5095 4701 5129 4735
rect 5727 4803 5761 4837
rect 5727 4701 5761 4735
rect 6061 4803 6095 4837
rect 6061 4735 6095 4769
rect 6161 4787 6195 4821
rect 6475 4803 6509 4837
rect 6161 4719 6195 4753
rect 6330 4667 6364 4701
rect 6475 4701 6509 4735
rect 6739 4803 6773 4837
rect 7053 4787 7087 4821
rect 6739 4701 6773 4735
rect 6884 4667 6918 4701
rect 7053 4719 7087 4753
rect 7153 4803 7187 4837
rect 7153 4735 7187 4769
rect 7303 4803 7337 4837
rect 7303 4701 7337 4735
rect 7751 4803 7785 4837
rect 7751 4701 7785 4735
rect 7855 4803 7889 4837
rect 7855 4735 7889 4769
rect 7855 4667 7889 4701
rect 7939 4803 7973 4837
rect 7939 4735 7973 4769
rect 8175 4743 8209 4777
rect 8250 4743 8284 4777
rect 8447 4743 8481 4777
rect 8533 4743 8567 4777
rect 7939 4667 7973 4701
rect 9353 4787 9387 4821
rect 9184 4667 9218 4701
rect 9353 4719 9387 4753
rect 9453 4803 9487 4837
rect 9453 4735 9487 4769
rect 9603 4803 9637 4837
rect 9603 4701 9637 4735
rect 9867 4803 9901 4837
rect 9867 4701 9901 4735
rect 10155 4803 10189 4837
rect 10155 4701 10189 4735
rect 10419 4803 10453 4837
rect 10733 4787 10767 4821
rect 10419 4701 10453 4735
rect 10564 4667 10598 4701
rect 10733 4719 10767 4753
rect 10833 4803 10867 4837
rect 10833 4735 10867 4769
rect 10983 4803 11017 4837
rect 10983 4701 11017 4735
rect 11247 4803 11281 4837
rect 11247 4701 11281 4735
rect 11351 4795 11385 4829
rect 11351 4727 11385 4761
rect 11437 4795 11471 4829
rect 11437 4727 11471 4761
rect 11523 4795 11557 4829
rect 11523 4714 11557 4748
rect 11627 4803 11661 4837
rect 11627 4701 11661 4735
rect 11891 4803 11925 4837
rect 11891 4701 11925 4735
rect 12041 4743 12075 4777
rect 12127 4743 12161 4777
rect 12324 4743 12358 4777
rect 12399 4743 12433 4777
rect 12635 4803 12669 4837
rect 12635 4735 12669 4769
rect 12635 4667 12669 4701
rect 12719 4803 12753 4837
rect 12719 4735 12753 4769
rect 12719 4667 12753 4701
rect 12823 4803 12857 4837
rect 12823 4701 12857 4735
rect 13087 4803 13121 4837
rect 13087 4701 13121 4735
rect 13191 4795 13225 4829
rect 13191 4714 13225 4748
rect 13277 4795 13311 4829
rect 13277 4727 13311 4761
rect 13363 4795 13397 4829
rect 13363 4727 13397 4761
rect 13467 4803 13501 4837
rect 13467 4701 13501 4735
rect 13915 4803 13949 4837
rect 13915 4701 13949 4735
rect 14111 4803 14145 4837
rect 15111 4803 15145 4837
rect 15425 4787 15459 4821
rect 15256 4667 15290 4701
rect 15425 4719 15459 4753
rect 15525 4803 15559 4837
rect 15525 4735 15559 4769
rect 15675 4803 15709 4837
rect 15675 4701 15709 4735
rect 15939 4803 15973 4837
rect 15939 4701 15973 4735
rect 16043 4795 16077 4829
rect 16043 4714 16077 4748
rect 16129 4795 16163 4829
rect 16129 4727 16163 4761
rect 16215 4795 16249 4829
rect 16215 4727 16249 4761
rect 16319 4803 16353 4837
rect 16319 4701 16353 4735
rect 16583 4803 16617 4837
rect 16583 4701 16617 4735
rect 16687 4795 16721 4829
rect 16687 4714 16721 4748
rect 16773 4795 16807 4829
rect 16773 4727 16807 4761
rect 16859 4795 16893 4829
rect 16859 4727 16893 4761
rect 16963 4803 16997 4837
rect 17963 4803 17997 4837
rect 18067 4803 18101 4837
rect 18067 4701 18101 4735
rect 18515 4803 18549 4837
rect 18515 4701 18549 4735
rect 18619 4803 18653 4837
rect 18619 4708 18653 4742
rect 18791 4803 18825 4837
rect 18791 4708 18825 4742
rect 1139 3962 1173 3996
rect 1139 3867 1173 3901
rect 1311 3962 1345 3996
rect 1311 3867 1345 3901
rect 1415 3969 1449 4003
rect 1415 3867 1449 3901
rect 2047 3969 2081 4003
rect 2047 3867 2081 3901
rect 2243 3943 2277 3977
rect 2243 3875 2277 3909
rect 2329 3943 2363 3977
rect 2329 3875 2363 3909
rect 2415 3956 2449 3990
rect 2415 3875 2449 3909
rect 2519 3969 2553 4003
rect 2519 3867 2553 3901
rect 2783 3969 2817 4003
rect 2783 3867 2817 3901
rect 2887 3943 2921 3977
rect 2887 3875 2921 3909
rect 2971 3891 3005 3925
rect 3055 3943 3089 3977
rect 3055 3875 3089 3909
rect 3238 3867 3272 3901
rect 3322 3875 3356 3909
rect 3415 3869 3449 3903
rect 3569 3893 3603 3927
rect 3666 3877 3700 3911
rect 3750 3893 3784 3927
rect 3863 3867 3897 3901
rect 3951 3875 3985 3909
rect 4048 3868 4082 3902
rect 4240 3867 4274 3901
rect 4324 3893 4358 3927
rect 4410 3867 4444 3901
rect 4539 3935 4573 3969
rect 4539 3867 4573 3901
rect 4623 3971 4657 4005
rect 4623 3903 4657 3937
rect 4727 3969 4761 4003
rect 4727 3867 4761 3901
rect 4991 3969 5025 4003
rect 4991 3867 5025 3901
rect 5371 3969 5405 4003
rect 5371 3867 5405 3901
rect 6003 3969 6037 4003
rect 6003 3867 6037 3901
rect 6383 3962 6417 3996
rect 6383 3867 6417 3901
rect 6555 3962 6589 3996
rect 6555 3867 6589 3901
rect 6659 3956 6693 3990
rect 6659 3875 6693 3909
rect 6745 3943 6779 3977
rect 6745 3875 6779 3909
rect 6831 3943 6865 3977
rect 6831 3875 6865 3909
rect 6935 3969 6969 4003
rect 6935 3867 6969 3901
rect 7567 3969 7601 4003
rect 8311 4003 8345 4037
rect 7567 3867 7601 3901
rect 7717 3927 7751 3961
rect 7803 3927 7837 3961
rect 8000 3927 8034 3961
rect 8075 3927 8109 3961
rect 8311 3935 8345 3969
rect 8311 3867 8345 3901
rect 8395 4003 8429 4037
rect 8395 3935 8429 3969
rect 8395 3867 8429 3901
rect 8499 3969 8533 4003
rect 8499 3867 8533 3901
rect 8763 3969 8797 4003
rect 8763 3867 8797 3901
rect 8959 3935 8993 3969
rect 8959 3867 8993 3901
rect 9045 3943 9079 3977
rect 9045 3875 9079 3909
rect 9131 3935 9165 3969
rect 9131 3867 9165 3901
rect 9217 3951 9251 3985
rect 9217 3883 9251 3917
rect 9303 3935 9337 3969
rect 9303 3867 9337 3901
rect 9389 3997 9423 4031
rect 9389 3911 9423 3945
rect 9475 3891 9509 3925
rect 9561 3997 9595 4031
rect 9561 3911 9595 3945
rect 9647 3891 9681 3925
rect 9733 3997 9767 4031
rect 9733 3911 9767 3945
rect 9819 3891 9853 3925
rect 9905 3997 9939 4031
rect 9905 3911 9939 3945
rect 9991 3891 10025 3925
rect 10076 3997 10110 4031
rect 10076 3911 10110 3945
rect 10162 3891 10196 3925
rect 10248 3997 10282 4031
rect 10248 3911 10282 3945
rect 10334 3891 10368 3925
rect 10420 3997 10454 4031
rect 10420 3911 10454 3945
rect 10506 3891 10540 3925
rect 10592 3997 10626 4031
rect 10592 3911 10626 3945
rect 10678 3891 10712 3925
rect 10799 3969 10833 4003
rect 10799 3867 10833 3901
rect 11247 3969 11281 4003
rect 11247 3867 11281 3901
rect 11719 3971 11753 4005
rect 11719 3903 11753 3937
rect 11803 3935 11837 3969
rect 11803 3867 11837 3901
rect 11932 3867 11966 3901
rect 12018 3893 12052 3927
rect 12102 3867 12136 3901
rect 12294 3868 12328 3902
rect 12391 3875 12425 3909
rect 13287 3943 13321 3977
rect 12479 3867 12513 3901
rect 12592 3893 12626 3927
rect 12676 3877 12710 3911
rect 12773 3893 12807 3927
rect 12927 3869 12961 3903
rect 13020 3875 13054 3909
rect 13104 3867 13138 3901
rect 13287 3875 13321 3909
rect 13371 3891 13405 3925
rect 13455 3943 13489 3977
rect 13455 3875 13489 3909
rect 13559 3969 13593 4003
rect 13559 3867 13593 3901
rect 13823 3969 13857 4003
rect 13823 3867 13857 3901
rect 13927 3943 13961 3977
rect 13927 3875 13961 3909
rect 14011 3891 14045 3925
rect 14095 3943 14129 3977
rect 14095 3875 14129 3909
rect 14278 3867 14312 3901
rect 14362 3875 14396 3909
rect 14455 3869 14489 3903
rect 14609 3893 14643 3927
rect 14706 3877 14740 3911
rect 14790 3893 14824 3927
rect 14903 3867 14937 3901
rect 14991 3875 15025 3909
rect 15088 3868 15122 3902
rect 15280 3867 15314 3901
rect 15364 3893 15398 3927
rect 15450 3867 15484 3901
rect 15579 3935 15613 3969
rect 15579 3867 15613 3901
rect 15663 3971 15697 4005
rect 15663 3903 15697 3937
rect 15767 3969 15801 4003
rect 15767 3867 15801 3901
rect 16399 3969 16433 4003
rect 16399 3867 16433 3901
rect 16687 3867 16721 3901
rect 17687 3867 17721 3901
rect 17791 3969 17825 4003
rect 17791 3867 17825 3901
rect 18423 3969 18457 4003
rect 18423 3867 18457 3901
rect 18619 3962 18653 3996
rect 18619 3867 18653 3901
rect 18791 3962 18825 3996
rect 18791 3867 18825 3901
rect 1139 3715 1173 3749
rect 1139 3620 1173 3654
rect 1311 3715 1345 3749
rect 1311 3620 1345 3654
rect 1415 3715 1449 3749
rect 1415 3620 1449 3654
rect 1587 3715 1621 3749
rect 1587 3620 1621 3654
rect 1691 3707 1725 3741
rect 1691 3639 1725 3673
rect 1775 3691 1809 3725
rect 1859 3707 1893 3741
rect 2042 3715 2076 3749
rect 2126 3707 2160 3741
rect 2219 3713 2253 3747
rect 2373 3689 2407 3723
rect 2470 3705 2504 3739
rect 2554 3689 2588 3723
rect 2667 3715 2701 3749
rect 1859 3639 1893 3673
rect 2755 3707 2789 3741
rect 2852 3714 2886 3748
rect 3044 3715 3078 3749
rect 3128 3689 3162 3723
rect 3214 3715 3248 3749
rect 3343 3715 3377 3749
rect 3343 3647 3377 3681
rect 3427 3679 3461 3713
rect 3427 3611 3461 3645
rect 3807 3715 3841 3749
rect 3807 3613 3841 3647
rect 4439 3715 4473 3749
rect 4439 3613 4473 3647
rect 4560 3691 4594 3725
rect 4646 3671 4680 3705
rect 4646 3585 4680 3619
rect 4732 3691 4766 3725
rect 4818 3671 4852 3705
rect 4818 3585 4852 3619
rect 4904 3691 4938 3725
rect 4990 3671 5024 3705
rect 4990 3585 5024 3619
rect 5076 3691 5110 3725
rect 5162 3671 5196 3705
rect 5162 3585 5196 3619
rect 5247 3691 5281 3725
rect 5333 3671 5367 3705
rect 5333 3585 5367 3619
rect 5419 3691 5453 3725
rect 5505 3671 5539 3705
rect 5505 3585 5539 3619
rect 5591 3691 5625 3725
rect 5677 3671 5711 3705
rect 5677 3585 5711 3619
rect 5763 3691 5797 3725
rect 5849 3671 5883 3705
rect 5849 3585 5883 3619
rect 5935 3715 5969 3749
rect 5935 3647 5969 3681
rect 6021 3699 6055 3733
rect 6021 3631 6055 3665
rect 6107 3715 6141 3749
rect 6107 3647 6141 3681
rect 6193 3707 6227 3741
rect 6193 3639 6227 3673
rect 6279 3715 6313 3749
rect 6279 3647 6313 3681
rect 6383 3715 6417 3749
rect 6383 3613 6417 3647
rect 6647 3715 6681 3749
rect 6647 3613 6681 3647
rect 6751 3707 6785 3741
rect 6751 3639 6785 3673
rect 6835 3691 6869 3725
rect 6919 3707 6953 3741
rect 7102 3715 7136 3749
rect 7186 3707 7220 3741
rect 7279 3713 7313 3747
rect 7433 3689 7467 3723
rect 7530 3705 7564 3739
rect 7614 3689 7648 3723
rect 7727 3715 7761 3749
rect 6919 3639 6953 3673
rect 7815 3707 7849 3741
rect 7912 3714 7946 3748
rect 8104 3715 8138 3749
rect 8188 3689 8222 3723
rect 8274 3715 8308 3749
rect 8403 3715 8437 3749
rect 8403 3647 8437 3681
rect 8487 3679 8521 3713
rect 8487 3611 8521 3645
rect 8591 3715 8625 3749
rect 8591 3620 8625 3654
rect 8763 3715 8797 3749
rect 8763 3620 8797 3654
rect 9143 3707 9177 3741
rect 9143 3639 9177 3673
rect 9236 3707 9270 3741
rect 9236 3639 9270 3673
rect 9322 3691 9356 3725
rect 9322 3610 9356 3644
rect 9406 3715 9440 3749
rect 9406 3647 9440 3681
rect 9406 3579 9440 3613
rect 9511 3715 9545 3749
rect 9511 3613 9545 3647
rect 9959 3715 9993 3749
rect 9959 3613 9993 3647
rect 10063 3707 10097 3741
rect 10063 3626 10097 3660
rect 10149 3707 10183 3741
rect 10149 3639 10183 3673
rect 10235 3707 10269 3741
rect 10235 3639 10269 3673
rect 10339 3715 10373 3749
rect 10339 3613 10373 3647
rect 10787 3715 10821 3749
rect 10787 3613 10821 3647
rect 10983 3707 11017 3741
rect 10983 3639 11017 3673
rect 11069 3707 11103 3741
rect 11069 3639 11103 3673
rect 11155 3707 11189 3741
rect 11155 3626 11189 3660
rect 11259 3715 11293 3749
rect 11259 3613 11293 3647
rect 11891 3715 11925 3749
rect 11891 3613 11925 3647
rect 11995 3679 12029 3713
rect 11995 3611 12029 3645
rect 12079 3715 12113 3749
rect 12079 3647 12113 3681
rect 12208 3715 12242 3749
rect 12294 3689 12328 3723
rect 12378 3715 12412 3749
rect 12570 3714 12604 3748
rect 12667 3707 12701 3741
rect 12755 3715 12789 3749
rect 12868 3689 12902 3723
rect 12952 3705 12986 3739
rect 13049 3689 13083 3723
rect 13203 3713 13237 3747
rect 13296 3707 13330 3741
rect 13380 3715 13414 3749
rect 13563 3707 13597 3741
rect 13563 3639 13597 3673
rect 13647 3691 13681 3725
rect 13731 3707 13765 3741
rect 13731 3639 13765 3673
rect 14111 3715 14145 3749
rect 15111 3715 15145 3749
rect 15215 3715 15249 3749
rect 16215 3715 16249 3749
rect 16319 3715 16353 3749
rect 17319 3715 17353 3749
rect 17423 3715 17457 3749
rect 18423 3715 18457 3749
rect 18619 3715 18653 3749
rect 18619 3620 18653 3654
rect 18791 3715 18825 3749
rect 18791 3620 18825 3654
rect 1139 2874 1173 2908
rect 1139 2779 1173 2813
rect 1311 2874 1345 2908
rect 1311 2779 1345 2813
rect 1415 2881 1449 2915
rect 1415 2779 1449 2813
rect 1863 2881 1897 2915
rect 1863 2779 1897 2813
rect 1967 2883 2001 2917
rect 1967 2815 2001 2849
rect 2051 2847 2085 2881
rect 2051 2779 2085 2813
rect 2180 2779 2214 2813
rect 2266 2805 2300 2839
rect 2350 2779 2384 2813
rect 2542 2780 2576 2814
rect 2639 2787 2673 2821
rect 3535 2855 3569 2889
rect 2727 2779 2761 2813
rect 2840 2805 2874 2839
rect 2924 2789 2958 2823
rect 3021 2805 3055 2839
rect 3175 2781 3209 2815
rect 3268 2787 3302 2821
rect 3352 2779 3386 2813
rect 3535 2787 3569 2821
rect 3619 2803 3653 2837
rect 3703 2855 3737 2889
rect 3703 2787 3737 2821
rect 3807 2881 3841 2915
rect 3807 2779 3841 2813
rect 4071 2881 4105 2915
rect 4071 2779 4105 2813
rect 4175 2855 4209 2889
rect 4175 2787 4209 2821
rect 4259 2803 4293 2837
rect 4343 2855 4377 2889
rect 4343 2787 4377 2821
rect 4447 2803 4481 2837
rect 4531 2855 4565 2889
rect 4531 2787 4565 2821
rect 4628 2780 4662 2814
rect 4842 2779 4876 2813
rect 4938 2805 4972 2839
rect 5022 2779 5056 2813
rect 5182 2781 5216 2815
rect 5362 2779 5396 2813
rect 5466 2805 5500 2839
rect 5562 2805 5596 2839
rect 5646 2873 5680 2907
rect 5646 2805 5680 2839
rect 5750 2847 5784 2881
rect 5750 2779 5784 2813
rect 5845 2847 5879 2881
rect 5845 2779 5879 2813
rect 5929 2883 5963 2917
rect 5929 2815 5963 2849
rect 6383 2881 6417 2915
rect 6383 2779 6417 2813
rect 7015 2881 7049 2915
rect 7015 2779 7049 2813
rect 7211 2883 7245 2917
rect 7211 2815 7245 2849
rect 7295 2847 7329 2881
rect 7295 2779 7329 2813
rect 7424 2779 7458 2813
rect 7510 2805 7544 2839
rect 7594 2779 7628 2813
rect 7786 2780 7820 2814
rect 7883 2787 7917 2821
rect 8779 2855 8813 2889
rect 7971 2779 8005 2813
rect 8084 2805 8118 2839
rect 8168 2789 8202 2823
rect 8265 2805 8299 2839
rect 8419 2781 8453 2815
rect 8512 2787 8546 2821
rect 8596 2779 8630 2813
rect 8779 2787 8813 2821
rect 8863 2803 8897 2837
rect 8947 2855 8981 2889
rect 8947 2787 8981 2821
rect 9051 2881 9085 2915
rect 9051 2779 9085 2813
rect 9315 2881 9349 2915
rect 9315 2779 9349 2813
rect 9419 2847 9453 2881
rect 9419 2779 9453 2813
rect 9505 2855 9539 2889
rect 9505 2787 9539 2821
rect 9591 2847 9625 2881
rect 9591 2779 9625 2813
rect 9677 2863 9711 2897
rect 9677 2795 9711 2829
rect 9763 2847 9797 2881
rect 9763 2779 9797 2813
rect 9849 2909 9883 2943
rect 9849 2823 9883 2857
rect 9935 2803 9969 2837
rect 10021 2909 10055 2943
rect 10021 2823 10055 2857
rect 10107 2803 10141 2837
rect 10193 2909 10227 2943
rect 10193 2823 10227 2857
rect 10279 2803 10313 2837
rect 10365 2909 10399 2943
rect 10365 2823 10399 2857
rect 10451 2803 10485 2837
rect 10536 2909 10570 2943
rect 10536 2823 10570 2857
rect 10622 2803 10656 2837
rect 10708 2909 10742 2943
rect 10708 2823 10742 2857
rect 10794 2803 10828 2837
rect 10880 2909 10914 2943
rect 10880 2823 10914 2857
rect 10966 2803 11000 2837
rect 11052 2909 11086 2943
rect 11052 2823 11086 2857
rect 11138 2803 11172 2837
rect 11719 2883 11753 2917
rect 11719 2815 11753 2849
rect 11803 2847 11837 2881
rect 11803 2779 11837 2813
rect 11932 2779 11966 2813
rect 12018 2805 12052 2839
rect 12102 2779 12136 2813
rect 12294 2780 12328 2814
rect 12391 2787 12425 2821
rect 13287 2855 13321 2889
rect 12479 2779 12513 2813
rect 12592 2805 12626 2839
rect 12676 2789 12710 2823
rect 12773 2805 12807 2839
rect 12927 2781 12961 2815
rect 13020 2787 13054 2821
rect 13104 2779 13138 2813
rect 13287 2787 13321 2821
rect 13371 2803 13405 2837
rect 13455 2855 13489 2889
rect 13455 2787 13489 2821
rect 13559 2881 13593 2915
rect 13559 2779 13593 2813
rect 13823 2881 13857 2915
rect 13823 2779 13857 2813
rect 13927 2855 13961 2889
rect 13927 2787 13961 2821
rect 14020 2855 14054 2889
rect 14020 2787 14054 2821
rect 14106 2884 14140 2918
rect 14106 2803 14140 2837
rect 14190 2915 14224 2949
rect 14190 2847 14224 2881
rect 14190 2779 14224 2813
rect 14295 2779 14329 2813
rect 15295 2779 15329 2813
rect 15399 2779 15433 2813
rect 16399 2779 16433 2813
rect 16687 2779 16721 2813
rect 17687 2779 17721 2813
rect 17791 2881 17825 2915
rect 17791 2779 17825 2813
rect 18423 2881 18457 2915
rect 18423 2779 18457 2813
rect 18619 2874 18653 2908
rect 18619 2779 18653 2813
rect 18791 2874 18825 2908
rect 18791 2779 18825 2813
rect 1139 2627 1173 2661
rect 1139 2532 1173 2566
rect 1311 2627 1345 2661
rect 1311 2532 1345 2566
rect 1415 2627 1449 2661
rect 1415 2532 1449 2566
rect 1587 2627 1621 2661
rect 1587 2532 1621 2566
rect 1691 2619 1725 2653
rect 1691 2551 1725 2585
rect 1775 2603 1809 2637
rect 1859 2619 1893 2653
rect 2042 2627 2076 2661
rect 2126 2619 2160 2653
rect 2219 2625 2253 2659
rect 2373 2601 2407 2635
rect 2470 2617 2504 2651
rect 2554 2601 2588 2635
rect 2667 2627 2701 2661
rect 1859 2551 1893 2585
rect 2755 2619 2789 2653
rect 2852 2626 2886 2660
rect 3044 2627 3078 2661
rect 3128 2601 3162 2635
rect 3214 2627 3248 2661
rect 3343 2627 3377 2661
rect 3343 2559 3377 2593
rect 3427 2591 3461 2625
rect 3427 2523 3461 2557
rect 3807 2627 3841 2661
rect 3807 2525 3841 2559
rect 4071 2627 4105 2661
rect 4071 2525 4105 2559
rect 4267 2619 4301 2653
rect 4267 2551 4301 2585
rect 4351 2603 4385 2637
rect 4435 2619 4469 2653
rect 4618 2627 4652 2661
rect 4702 2619 4736 2653
rect 4795 2625 4829 2659
rect 4949 2601 4983 2635
rect 5046 2617 5080 2651
rect 5130 2601 5164 2635
rect 5243 2627 5277 2661
rect 4435 2551 4469 2585
rect 5331 2619 5365 2653
rect 5428 2626 5462 2660
rect 5620 2627 5654 2661
rect 5704 2601 5738 2635
rect 5790 2627 5824 2661
rect 5919 2627 5953 2661
rect 5919 2559 5953 2593
rect 6003 2591 6037 2625
rect 6003 2523 6037 2557
rect 6383 2627 6417 2661
rect 7383 2627 7417 2661
rect 7487 2627 7521 2661
rect 8487 2627 8521 2661
rect 8591 2627 8625 2661
rect 8591 2532 8625 2566
rect 8763 2627 8797 2661
rect 8763 2532 8797 2566
rect 9143 2591 9177 2625
rect 9143 2523 9177 2557
rect 9227 2627 9261 2661
rect 9227 2559 9261 2593
rect 9356 2627 9390 2661
rect 9442 2601 9476 2635
rect 9526 2627 9560 2661
rect 9718 2626 9752 2660
rect 9815 2619 9849 2653
rect 9903 2627 9937 2661
rect 10016 2601 10050 2635
rect 10100 2617 10134 2651
rect 10197 2601 10231 2635
rect 10351 2625 10385 2659
rect 10444 2619 10478 2653
rect 10528 2627 10562 2661
rect 10711 2619 10745 2653
rect 10711 2551 10745 2585
rect 10795 2603 10829 2637
rect 10879 2619 10913 2653
rect 10879 2551 10913 2585
rect 10983 2627 11017 2661
rect 10983 2525 11017 2559
rect 11247 2627 11281 2661
rect 11247 2525 11281 2559
rect 11535 2627 11569 2661
rect 11535 2525 11569 2559
rect 11799 2627 11833 2661
rect 11799 2525 11833 2559
rect 11995 2591 12029 2625
rect 11995 2523 12029 2557
rect 12079 2627 12113 2661
rect 12079 2559 12113 2593
rect 12208 2627 12242 2661
rect 12294 2601 12328 2635
rect 12378 2627 12412 2661
rect 12570 2626 12604 2660
rect 12667 2619 12701 2653
rect 12755 2627 12789 2661
rect 12868 2601 12902 2635
rect 12952 2617 12986 2651
rect 13049 2601 13083 2635
rect 13203 2625 13237 2659
rect 13296 2619 13330 2653
rect 13380 2627 13414 2661
rect 13563 2619 13597 2653
rect 13563 2551 13597 2585
rect 13647 2603 13681 2637
rect 13731 2619 13765 2653
rect 13731 2551 13765 2585
rect 14295 2591 14329 2625
rect 14295 2523 14329 2557
rect 14379 2627 14413 2661
rect 14379 2559 14413 2593
rect 14508 2627 14542 2661
rect 14594 2601 14628 2635
rect 14678 2627 14712 2661
rect 14870 2626 14904 2660
rect 14967 2619 15001 2653
rect 15055 2627 15089 2661
rect 15168 2601 15202 2635
rect 15252 2617 15286 2651
rect 15349 2601 15383 2635
rect 15503 2625 15537 2659
rect 15596 2619 15630 2653
rect 15680 2627 15714 2661
rect 15863 2619 15897 2653
rect 15863 2551 15897 2585
rect 15947 2603 15981 2637
rect 16031 2619 16065 2653
rect 16031 2551 16065 2585
rect 16135 2627 16169 2661
rect 16135 2525 16169 2559
rect 16399 2627 16433 2661
rect 16399 2525 16433 2559
rect 16687 2627 16721 2661
rect 16687 2525 16721 2559
rect 17319 2627 17353 2661
rect 17319 2525 17353 2559
rect 17515 2619 17549 2653
rect 17515 2551 17549 2585
rect 17608 2619 17642 2653
rect 17608 2551 17642 2585
rect 17694 2603 17728 2637
rect 17694 2522 17728 2556
rect 17778 2627 17812 2661
rect 17778 2559 17812 2593
rect 17778 2491 17812 2525
rect 17883 2627 17917 2661
rect 17883 2525 17917 2559
rect 18515 2627 18549 2661
rect 18515 2525 18549 2559
rect 18619 2627 18653 2661
rect 18619 2532 18653 2566
rect 18791 2627 18825 2661
rect 18791 2532 18825 2566
<< psubdiff >>
rect 3709 7505 3743 7552
rect 3709 7447 3743 7471
rect 6285 7505 6319 7552
rect 6285 7447 6319 7471
rect 8861 7505 8895 7552
rect 8861 7447 8895 7471
rect 11437 7505 11471 7552
rect 11437 7447 11471 7471
rect 14013 7505 14047 7552
rect 14013 7447 14047 7471
rect 16589 7505 16623 7552
rect 16589 7447 16623 7471
rect 3709 6673 3743 6697
rect 3709 6592 3743 6639
rect 8861 6673 8895 6697
rect 8861 6592 8895 6639
rect 14013 6673 14047 6697
rect 14013 6592 14047 6639
rect 6285 6417 6319 6464
rect 6285 6359 6319 6383
rect 11437 6417 11471 6464
rect 11437 6359 11471 6383
rect 16589 6417 16623 6464
rect 16589 6359 16623 6383
rect 3709 5585 3743 5609
rect 3709 5504 3743 5551
rect 8861 5585 8895 5609
rect 8861 5504 8895 5551
rect 14013 5585 14047 5609
rect 14013 5504 14047 5551
rect 6285 5329 6319 5376
rect 6285 5271 6319 5295
rect 11437 5329 11471 5376
rect 11437 5271 11471 5295
rect 16589 5329 16623 5376
rect 16589 5271 16623 5295
rect 3709 4497 3743 4521
rect 3709 4416 3743 4463
rect 8861 4497 8895 4521
rect 8861 4416 8895 4463
rect 14013 4497 14047 4521
rect 14013 4416 14047 4463
rect 6285 4241 6319 4288
rect 6285 4183 6319 4207
rect 11437 4241 11471 4288
rect 11437 4183 11471 4207
rect 16589 4241 16623 4288
rect 16589 4183 16623 4207
rect 3709 3409 3743 3433
rect 3709 3328 3743 3375
rect 8861 3409 8895 3433
rect 8861 3328 8895 3375
rect 14013 3409 14047 3433
rect 14013 3328 14047 3375
rect 6285 3153 6319 3200
rect 6285 3095 6319 3119
rect 11437 3153 11471 3200
rect 11437 3095 11471 3119
rect 16589 3153 16623 3200
rect 16589 3095 16623 3119
rect 3709 2321 3743 2345
rect 3709 2240 3743 2287
rect 6285 2321 6319 2345
rect 6285 2240 6319 2287
rect 8861 2321 8895 2345
rect 8861 2240 8895 2287
rect 11437 2321 11471 2345
rect 11437 2240 11471 2287
rect 14013 2321 14047 2345
rect 14013 2240 14047 2287
rect 16589 2321 16623 2345
rect 16589 2240 16623 2287
<< nsubdiff >>
rect 3709 7287 3743 7311
rect 3709 7194 3743 7253
rect 3709 7136 3743 7160
rect 6285 7287 6319 7311
rect 6285 7194 6319 7253
rect 6285 7136 6319 7160
rect 8861 7287 8895 7311
rect 8861 7194 8895 7253
rect 8861 7136 8895 7160
rect 11437 7287 11471 7311
rect 11437 7194 11471 7253
rect 11437 7136 11471 7160
rect 14013 7287 14047 7311
rect 14013 7194 14047 7253
rect 14013 7136 14047 7160
rect 16589 7287 16623 7311
rect 16589 7194 16623 7253
rect 16589 7136 16623 7160
rect 3709 6984 3743 7008
rect 3709 6891 3743 6950
rect 3709 6833 3743 6857
rect 8861 6984 8895 7008
rect 8861 6891 8895 6950
rect 8861 6833 8895 6857
rect 14013 6984 14047 7008
rect 14013 6891 14047 6950
rect 14013 6833 14047 6857
rect 6285 6199 6319 6223
rect 6285 6106 6319 6165
rect 6285 6048 6319 6072
rect 11437 6199 11471 6223
rect 11437 6106 11471 6165
rect 11437 6048 11471 6072
rect 16589 6199 16623 6223
rect 16589 6106 16623 6165
rect 16589 6048 16623 6072
rect 3709 5896 3743 5920
rect 3709 5803 3743 5862
rect 3709 5745 3743 5769
rect 8861 5896 8895 5920
rect 8861 5803 8895 5862
rect 8861 5745 8895 5769
rect 14013 5896 14047 5920
rect 14013 5803 14047 5862
rect 14013 5745 14047 5769
rect 6285 5111 6319 5135
rect 6285 5018 6319 5077
rect 6285 4960 6319 4984
rect 11437 5111 11471 5135
rect 11437 5018 11471 5077
rect 11437 4960 11471 4984
rect 16589 5111 16623 5135
rect 16589 5018 16623 5077
rect 16589 4960 16623 4984
rect 3709 4808 3743 4832
rect 3709 4715 3743 4774
rect 3709 4657 3743 4681
rect 8861 4808 8895 4832
rect 8861 4715 8895 4774
rect 8861 4657 8895 4681
rect 14013 4808 14047 4832
rect 14013 4715 14047 4774
rect 14013 4657 14047 4681
rect 6285 4023 6319 4047
rect 6285 3930 6319 3989
rect 6285 3872 6319 3896
rect 11437 4023 11471 4047
rect 11437 3930 11471 3989
rect 11437 3872 11471 3896
rect 16589 4023 16623 4047
rect 16589 3930 16623 3989
rect 16589 3872 16623 3896
rect 3709 3720 3743 3744
rect 3709 3627 3743 3686
rect 3709 3569 3743 3593
rect 8861 3720 8895 3744
rect 8861 3627 8895 3686
rect 8861 3569 8895 3593
rect 14013 3720 14047 3744
rect 14013 3627 14047 3686
rect 14013 3569 14047 3593
rect 6285 2935 6319 2959
rect 6285 2842 6319 2901
rect 6285 2784 6319 2808
rect 11437 2935 11471 2959
rect 11437 2842 11471 2901
rect 11437 2784 11471 2808
rect 16589 2935 16623 2959
rect 16589 2842 16623 2901
rect 16589 2784 16623 2808
rect 3709 2632 3743 2656
rect 3709 2539 3743 2598
rect 3709 2481 3743 2505
rect 6285 2632 6319 2656
rect 6285 2539 6319 2598
rect 6285 2481 6319 2505
rect 8861 2632 8895 2656
rect 8861 2539 8895 2598
rect 8861 2481 8895 2505
rect 11437 2632 11471 2656
rect 11437 2539 11471 2598
rect 11437 2481 11471 2505
rect 14013 2632 14047 2656
rect 14013 2539 14047 2598
rect 14013 2481 14047 2505
rect 16589 2632 16623 2656
rect 16589 2539 16623 2598
rect 16589 2481 16623 2505
<< psubdiffcont >>
rect 3709 7471 3743 7505
rect 6285 7471 6319 7505
rect 8861 7471 8895 7505
rect 11437 7471 11471 7505
rect 14013 7471 14047 7505
rect 16589 7471 16623 7505
rect 3709 6639 3743 6673
rect 8861 6639 8895 6673
rect 14013 6639 14047 6673
rect 6285 6383 6319 6417
rect 11437 6383 11471 6417
rect 16589 6383 16623 6417
rect 3709 5551 3743 5585
rect 8861 5551 8895 5585
rect 14013 5551 14047 5585
rect 6285 5295 6319 5329
rect 11437 5295 11471 5329
rect 16589 5295 16623 5329
rect 3709 4463 3743 4497
rect 8861 4463 8895 4497
rect 14013 4463 14047 4497
rect 6285 4207 6319 4241
rect 11437 4207 11471 4241
rect 16589 4207 16623 4241
rect 3709 3375 3743 3409
rect 8861 3375 8895 3409
rect 14013 3375 14047 3409
rect 6285 3119 6319 3153
rect 11437 3119 11471 3153
rect 16589 3119 16623 3153
rect 3709 2287 3743 2321
rect 6285 2287 6319 2321
rect 8861 2287 8895 2321
rect 11437 2287 11471 2321
rect 14013 2287 14047 2321
rect 16589 2287 16623 2321
<< nsubdiffcont >>
rect 3709 7253 3743 7287
rect 3709 7160 3743 7194
rect 6285 7253 6319 7287
rect 6285 7160 6319 7194
rect 8861 7253 8895 7287
rect 8861 7160 8895 7194
rect 11437 7253 11471 7287
rect 11437 7160 11471 7194
rect 14013 7253 14047 7287
rect 14013 7160 14047 7194
rect 16589 7253 16623 7287
rect 16589 7160 16623 7194
rect 3709 6950 3743 6984
rect 3709 6857 3743 6891
rect 8861 6950 8895 6984
rect 8861 6857 8895 6891
rect 14013 6950 14047 6984
rect 14013 6857 14047 6891
rect 6285 6165 6319 6199
rect 6285 6072 6319 6106
rect 11437 6165 11471 6199
rect 11437 6072 11471 6106
rect 16589 6165 16623 6199
rect 16589 6072 16623 6106
rect 3709 5862 3743 5896
rect 3709 5769 3743 5803
rect 8861 5862 8895 5896
rect 8861 5769 8895 5803
rect 14013 5862 14047 5896
rect 14013 5769 14047 5803
rect 6285 5077 6319 5111
rect 6285 4984 6319 5018
rect 11437 5077 11471 5111
rect 11437 4984 11471 5018
rect 16589 5077 16623 5111
rect 16589 4984 16623 5018
rect 3709 4774 3743 4808
rect 3709 4681 3743 4715
rect 8861 4774 8895 4808
rect 8861 4681 8895 4715
rect 14013 4774 14047 4808
rect 14013 4681 14047 4715
rect 6285 3989 6319 4023
rect 6285 3896 6319 3930
rect 11437 3989 11471 4023
rect 11437 3896 11471 3930
rect 16589 3989 16623 4023
rect 16589 3896 16623 3930
rect 3709 3686 3743 3720
rect 3709 3593 3743 3627
rect 8861 3686 8895 3720
rect 8861 3593 8895 3627
rect 14013 3686 14047 3720
rect 14013 3593 14047 3627
rect 6285 2901 6319 2935
rect 6285 2808 6319 2842
rect 11437 2901 11471 2935
rect 11437 2808 11471 2842
rect 16589 2901 16623 2935
rect 16589 2808 16623 2842
rect 3709 2598 3743 2632
rect 3709 2505 3743 2539
rect 6285 2598 6319 2632
rect 6285 2505 6319 2539
rect 8861 2598 8895 2632
rect 8861 2505 8895 2539
rect 11437 2598 11471 2632
rect 11437 2505 11471 2539
rect 14013 2598 14047 2632
rect 14013 2505 14047 2539
rect 16589 2598 16623 2632
rect 16589 2505 16623 2539
<< poly >>
rect 1183 7569 1301 7595
rect 1644 7569 1674 7595
rect 1728 7569 1758 7595
rect 1823 7569 1853 7595
rect 2011 7569 2957 7595
rect 3115 7569 3509 7595
rect 4036 7569 4066 7595
rect 4120 7569 4150 7595
rect 4215 7569 4245 7595
rect 4403 7569 5349 7595
rect 5692 7569 5722 7595
rect 5776 7569 5806 7595
rect 5871 7569 5901 7595
rect 6059 7569 6177 7595
rect 6427 7569 7373 7595
rect 7531 7569 7741 7595
rect 7900 7569 7930 7595
rect 7984 7569 8014 7595
rect 8079 7569 8109 7595
rect 8267 7569 8661 7595
rect 9003 7569 9397 7595
rect 1183 7433 1301 7459
rect 1263 7431 1301 7433
rect 1263 7415 1329 7431
rect 1155 7375 1221 7391
rect 1155 7341 1171 7375
rect 1205 7341 1221 7375
rect 1263 7381 1279 7415
rect 1313 7381 1329 7415
rect 1263 7365 1329 7381
rect 1644 7417 1674 7439
rect 1728 7417 1758 7439
rect 1823 7417 1853 7485
rect 2011 7433 2957 7459
rect 3115 7433 3509 7459
rect 1644 7401 1781 7417
rect 1644 7367 1737 7401
rect 1771 7367 1781 7401
rect 1155 7325 1221 7341
rect 1183 7323 1221 7325
rect 1644 7351 1781 7367
rect 1823 7401 1905 7417
rect 1823 7367 1861 7401
rect 1895 7367 1905 7401
rect 2503 7411 2957 7433
rect 1823 7351 1905 7367
rect 2011 7375 2461 7391
rect 1183 7293 1301 7323
rect 1644 7319 1674 7351
rect 1728 7319 1758 7351
rect 1823 7255 1853 7351
rect 2011 7341 2283 7375
rect 2317 7341 2461 7375
rect 2503 7377 2647 7411
rect 2681 7377 2957 7411
rect 3333 7411 3509 7433
rect 2503 7361 2957 7377
rect 3115 7375 3291 7391
rect 2011 7319 2461 7341
rect 3115 7341 3131 7375
rect 3165 7341 3241 7375
rect 3275 7341 3291 7375
rect 3333 7377 3349 7411
rect 3383 7377 3459 7411
rect 3493 7377 3509 7411
rect 3333 7361 3509 7377
rect 4036 7417 4066 7439
rect 4120 7417 4150 7439
rect 4215 7417 4245 7485
rect 4403 7433 5349 7459
rect 4036 7401 4173 7417
rect 4036 7367 4129 7401
rect 4163 7367 4173 7401
rect 3115 7319 3291 7341
rect 4036 7351 4173 7367
rect 4215 7401 4297 7417
rect 4215 7367 4253 7401
rect 4287 7367 4297 7401
rect 4895 7411 5349 7433
rect 4215 7351 4297 7367
rect 4403 7375 4853 7391
rect 4036 7319 4066 7351
rect 4120 7319 4150 7351
rect 2011 7293 2957 7319
rect 3115 7293 3509 7319
rect 1183 7093 1301 7119
rect 1644 7093 1674 7119
rect 1728 7093 1758 7119
rect 1823 7101 1853 7127
rect 4215 7255 4245 7351
rect 4403 7341 4675 7375
rect 4709 7341 4853 7375
rect 4895 7377 5039 7411
rect 5073 7377 5349 7411
rect 4895 7361 5349 7377
rect 5692 7417 5722 7439
rect 5776 7417 5806 7439
rect 5871 7417 5901 7485
rect 6059 7433 6177 7459
rect 6427 7433 7373 7459
rect 7531 7433 7741 7459
rect 6139 7431 6177 7433
rect 5692 7401 5829 7417
rect 5692 7367 5785 7401
rect 5819 7367 5829 7401
rect 4403 7319 4853 7341
rect 5692 7351 5829 7367
rect 5871 7401 5953 7417
rect 5871 7367 5909 7401
rect 5943 7367 5953 7401
rect 6139 7415 6205 7431
rect 5871 7351 5953 7367
rect 6031 7375 6097 7391
rect 5692 7319 5722 7351
rect 5776 7319 5806 7351
rect 4403 7293 5349 7319
rect 2011 7093 2957 7119
rect 3115 7093 3509 7119
rect 4036 7093 4066 7119
rect 4120 7093 4150 7119
rect 4215 7101 4245 7127
rect 5871 7255 5901 7351
rect 6031 7341 6047 7375
rect 6081 7341 6097 7375
rect 6139 7381 6155 7415
rect 6189 7381 6205 7415
rect 6919 7411 7373 7433
rect 6139 7365 6205 7381
rect 6427 7375 6877 7391
rect 6031 7325 6097 7341
rect 6059 7323 6097 7325
rect 6427 7341 6699 7375
rect 6733 7341 6877 7375
rect 6919 7377 7063 7411
rect 7097 7377 7373 7411
rect 7657 7427 7741 7433
rect 7657 7411 7799 7427
rect 6919 7361 7373 7377
rect 7473 7375 7615 7391
rect 6059 7293 6177 7323
rect 6427 7319 6877 7341
rect 7473 7341 7489 7375
rect 7523 7341 7615 7375
rect 7657 7377 7749 7411
rect 7783 7377 7799 7411
rect 7657 7361 7799 7377
rect 7900 7417 7930 7439
rect 7984 7417 8014 7439
rect 8079 7417 8109 7485
rect 8267 7433 8661 7459
rect 9739 7569 9949 7595
rect 10108 7569 10138 7595
rect 10203 7569 10233 7595
rect 10287 7569 10317 7595
rect 10475 7569 11053 7595
rect 11211 7569 11329 7595
rect 11579 7569 12157 7595
rect 12315 7569 12345 7595
rect 12410 7569 12440 7595
rect 12494 7569 12524 7595
rect 12683 7569 13629 7595
rect 13787 7569 13905 7595
rect 14155 7569 14365 7595
rect 14523 7569 14553 7595
rect 14618 7569 14648 7595
rect 14702 7569 14732 7595
rect 14891 7569 15837 7595
rect 15995 7569 16389 7595
rect 16915 7569 16945 7595
rect 17010 7569 17040 7595
rect 17094 7569 17124 7595
rect 17283 7569 17861 7595
rect 18111 7569 18141 7595
rect 18206 7569 18236 7595
rect 18290 7569 18320 7595
rect 18663 7569 18781 7595
rect 9003 7433 9397 7459
rect 9739 7433 9949 7459
rect 7900 7401 8037 7417
rect 7900 7367 7993 7401
rect 8027 7367 8037 7401
rect 7473 7325 7615 7341
rect 7531 7319 7615 7325
rect 7900 7351 8037 7367
rect 8079 7401 8161 7417
rect 8079 7367 8117 7401
rect 8151 7367 8161 7401
rect 8485 7411 8661 7433
rect 8079 7351 8161 7367
rect 8267 7375 8443 7391
rect 7900 7319 7930 7351
rect 7984 7319 8014 7351
rect 4403 7093 5349 7119
rect 5692 7093 5722 7119
rect 5776 7093 5806 7119
rect 5871 7101 5901 7127
rect 6427 7293 7373 7319
rect 7531 7293 7741 7319
rect 8079 7255 8109 7351
rect 8267 7341 8283 7375
rect 8317 7341 8393 7375
rect 8427 7341 8443 7375
rect 8485 7377 8501 7411
rect 8535 7377 8611 7411
rect 8645 7377 8661 7411
rect 9221 7411 9397 7433
rect 8485 7361 8661 7377
rect 9003 7375 9179 7391
rect 8267 7319 8443 7341
rect 9003 7341 9019 7375
rect 9053 7341 9129 7375
rect 9163 7341 9179 7375
rect 9221 7377 9237 7411
rect 9271 7377 9347 7411
rect 9381 7377 9397 7411
rect 9865 7427 9949 7433
rect 10108 7436 10138 7485
rect 10203 7467 10233 7485
rect 10287 7467 10317 7485
rect 9865 7411 10007 7427
rect 10108 7421 10161 7436
rect 9221 7361 9397 7377
rect 9681 7375 9823 7391
rect 9003 7319 9179 7341
rect 9681 7341 9697 7375
rect 9731 7341 9823 7375
rect 9865 7377 9957 7411
rect 9991 7377 10007 7411
rect 9865 7361 10007 7377
rect 10097 7401 10161 7421
rect 10097 7367 10117 7401
rect 10151 7367 10161 7401
rect 9681 7325 9823 7341
rect 10097 7337 10161 7367
rect 10203 7401 10317 7467
rect 10475 7433 11053 7459
rect 11211 7433 11329 7459
rect 11579 7433 12157 7459
rect 10203 7367 10221 7401
rect 10255 7367 10317 7401
rect 10781 7411 11053 7433
rect 10203 7337 10317 7367
rect 9739 7319 9823 7325
rect 10108 7319 10138 7337
rect 10203 7319 10233 7337
rect 10287 7319 10317 7337
rect 10475 7375 10739 7391
rect 10475 7341 10491 7375
rect 10525 7341 10590 7375
rect 10624 7341 10689 7375
rect 10723 7341 10739 7375
rect 10781 7377 10797 7411
rect 10831 7377 10900 7411
rect 10934 7377 11003 7411
rect 11037 7377 11053 7411
rect 11291 7431 11329 7433
rect 11291 7415 11357 7431
rect 10781 7361 11053 7377
rect 11183 7375 11249 7391
rect 10475 7319 10739 7341
rect 11183 7341 11199 7375
rect 11233 7341 11249 7375
rect 11291 7381 11307 7415
rect 11341 7381 11357 7415
rect 11885 7411 12157 7433
rect 12315 7417 12345 7485
rect 12410 7417 12440 7439
rect 12494 7417 12524 7439
rect 12683 7433 13629 7459
rect 13787 7433 13905 7459
rect 14155 7433 14365 7459
rect 11291 7365 11357 7381
rect 11579 7375 11843 7391
rect 11183 7325 11249 7341
rect 11211 7323 11249 7325
rect 11579 7341 11595 7375
rect 11629 7341 11694 7375
rect 11728 7341 11793 7375
rect 11827 7341 11843 7375
rect 11885 7377 11901 7411
rect 11935 7377 12004 7411
rect 12038 7377 12107 7411
rect 12141 7377 12157 7411
rect 11885 7361 12157 7377
rect 12263 7401 12345 7417
rect 12263 7367 12273 7401
rect 12307 7367 12345 7401
rect 12263 7351 12345 7367
rect 12387 7401 12524 7417
rect 12387 7367 12397 7401
rect 12431 7367 12524 7401
rect 13175 7411 13629 7433
rect 12387 7351 12524 7367
rect 8267 7293 8661 7319
rect 6059 7093 6177 7119
rect 6427 7093 7373 7119
rect 7531 7093 7741 7119
rect 7900 7093 7930 7119
rect 7984 7093 8014 7119
rect 8079 7101 8109 7127
rect 9003 7293 9397 7319
rect 9739 7293 9949 7319
rect 10475 7293 11053 7319
rect 11211 7293 11329 7323
rect 11579 7319 11843 7341
rect 11579 7293 12157 7319
rect 12315 7255 12345 7351
rect 12410 7319 12440 7351
rect 12494 7319 12524 7351
rect 12683 7375 13133 7391
rect 12683 7341 12955 7375
rect 12989 7341 13133 7375
rect 13175 7377 13319 7411
rect 13353 7377 13629 7411
rect 13867 7431 13905 7433
rect 13867 7415 13933 7431
rect 13175 7361 13629 7377
rect 13759 7375 13825 7391
rect 12683 7319 13133 7341
rect 13759 7341 13775 7375
rect 13809 7341 13825 7375
rect 13867 7381 13883 7415
rect 13917 7381 13933 7415
rect 14281 7427 14365 7433
rect 14281 7411 14423 7427
rect 14523 7417 14553 7485
rect 14618 7417 14648 7439
rect 14702 7417 14732 7439
rect 14891 7433 15837 7459
rect 15995 7433 16389 7459
rect 13867 7365 13933 7381
rect 14097 7375 14239 7391
rect 13759 7325 13825 7341
rect 14097 7341 14113 7375
rect 14147 7341 14239 7375
rect 14281 7377 14373 7411
rect 14407 7377 14423 7411
rect 14281 7361 14423 7377
rect 14471 7401 14553 7417
rect 14471 7367 14481 7401
rect 14515 7367 14553 7401
rect 14471 7351 14553 7367
rect 14595 7401 14732 7417
rect 14595 7367 14605 7401
rect 14639 7367 14732 7401
rect 15383 7411 15837 7433
rect 14595 7351 14732 7367
rect 14097 7325 14239 7341
rect 13787 7323 13825 7325
rect 8267 7093 8661 7119
rect 9003 7093 9397 7119
rect 9739 7093 9949 7119
rect 10108 7093 10138 7119
rect 10203 7093 10233 7119
rect 10287 7093 10317 7119
rect 10475 7093 11053 7119
rect 11211 7093 11329 7119
rect 11579 7093 12157 7119
rect 12315 7101 12345 7127
rect 12683 7293 13629 7319
rect 13787 7293 13905 7323
rect 14155 7319 14239 7325
rect 14155 7293 14365 7319
rect 14523 7255 14553 7351
rect 14618 7319 14648 7351
rect 14702 7319 14732 7351
rect 14891 7375 15341 7391
rect 14891 7341 15163 7375
rect 15197 7341 15341 7375
rect 15383 7377 15527 7411
rect 15561 7377 15837 7411
rect 16213 7411 16389 7433
rect 16915 7417 16945 7485
rect 17010 7417 17040 7439
rect 17094 7417 17124 7439
rect 17283 7433 17861 7459
rect 15383 7361 15837 7377
rect 15995 7375 16171 7391
rect 14891 7319 15341 7341
rect 15995 7341 16011 7375
rect 16045 7341 16121 7375
rect 16155 7341 16171 7375
rect 16213 7377 16229 7411
rect 16263 7377 16339 7411
rect 16373 7377 16389 7411
rect 16213 7361 16389 7377
rect 16863 7401 16945 7417
rect 16863 7367 16873 7401
rect 16907 7367 16945 7401
rect 16863 7351 16945 7367
rect 16987 7401 17124 7417
rect 16987 7367 16997 7401
rect 17031 7367 17124 7401
rect 17589 7411 17861 7433
rect 18111 7417 18141 7485
rect 18206 7417 18236 7439
rect 18290 7417 18320 7439
rect 18663 7433 18781 7459
rect 18663 7431 18701 7433
rect 16987 7351 17124 7367
rect 15995 7319 16171 7341
rect 12410 7093 12440 7119
rect 12494 7093 12524 7119
rect 12683 7093 13629 7119
rect 13787 7093 13905 7119
rect 14155 7093 14365 7119
rect 14523 7101 14553 7127
rect 14891 7293 15837 7319
rect 15995 7293 16389 7319
rect 16915 7255 16945 7351
rect 17010 7319 17040 7351
rect 17094 7319 17124 7351
rect 17283 7375 17547 7391
rect 17283 7341 17299 7375
rect 17333 7341 17398 7375
rect 17432 7341 17497 7375
rect 17531 7341 17547 7375
rect 17589 7377 17605 7411
rect 17639 7377 17708 7411
rect 17742 7377 17811 7411
rect 17845 7377 17861 7411
rect 17589 7361 17861 7377
rect 18059 7401 18141 7417
rect 18059 7367 18069 7401
rect 18103 7367 18141 7401
rect 18059 7351 18141 7367
rect 18183 7401 18320 7417
rect 18183 7367 18193 7401
rect 18227 7367 18320 7401
rect 18183 7351 18320 7367
rect 18635 7415 18701 7431
rect 18635 7381 18651 7415
rect 18685 7381 18701 7415
rect 18635 7365 18701 7381
rect 18743 7375 18809 7391
rect 17283 7319 17547 7341
rect 14618 7093 14648 7119
rect 14702 7093 14732 7119
rect 14891 7093 15837 7119
rect 15995 7093 16389 7119
rect 16915 7101 16945 7127
rect 17283 7293 17861 7319
rect 18111 7255 18141 7351
rect 18206 7319 18236 7351
rect 18290 7319 18320 7351
rect 18743 7341 18759 7375
rect 18793 7341 18809 7375
rect 18743 7325 18809 7341
rect 18743 7323 18781 7325
rect 17010 7093 17040 7119
rect 17094 7093 17124 7119
rect 17283 7093 17861 7119
rect 18111 7101 18141 7127
rect 18663 7293 18781 7323
rect 18206 7093 18236 7119
rect 18290 7093 18320 7119
rect 18663 7093 18781 7119
rect 1183 7025 1301 7051
rect 1459 7025 2405 7051
rect 2563 7025 3509 7051
rect 3851 7025 4797 7051
rect 4955 7025 5901 7051
rect 6059 7025 7005 7051
rect 7163 7025 8109 7051
rect 8267 7025 8661 7051
rect 9003 7025 9949 7051
rect 10107 7025 11053 7051
rect 11211 7025 12157 7051
rect 12315 7025 13261 7051
rect 13419 7025 13813 7051
rect 14155 7025 15101 7051
rect 15259 7025 16205 7051
rect 16363 7025 17309 7051
rect 17467 7025 18413 7051
rect 18663 7025 18781 7051
rect 1183 6821 1301 6851
rect 1459 6825 2405 6851
rect 2563 6825 3509 6851
rect 3851 6825 4797 6851
rect 4955 6825 5901 6851
rect 6059 6825 7005 6851
rect 7163 6825 8109 6851
rect 8267 6825 8661 6851
rect 9003 6825 9949 6851
rect 10107 6825 11053 6851
rect 11211 6825 12157 6851
rect 12315 6825 13261 6851
rect 13419 6825 13813 6851
rect 14155 6825 15101 6851
rect 15259 6825 16205 6851
rect 16363 6825 17309 6851
rect 17467 6825 18413 6851
rect 1183 6819 1221 6821
rect 1155 6803 1221 6819
rect 1155 6769 1171 6803
rect 1205 6769 1221 6803
rect 1459 6803 1909 6825
rect 1155 6753 1221 6769
rect 1263 6763 1329 6779
rect 1263 6729 1279 6763
rect 1313 6729 1329 6763
rect 1459 6769 1731 6803
rect 1765 6769 1909 6803
rect 2563 6803 3013 6825
rect 1459 6753 1909 6769
rect 1951 6767 2405 6783
rect 1263 6713 1329 6729
rect 1951 6733 2095 6767
rect 2129 6733 2405 6767
rect 2563 6769 2835 6803
rect 2869 6769 3013 6803
rect 3851 6803 4301 6825
rect 2563 6753 3013 6769
rect 3055 6767 3509 6783
rect 1263 6711 1301 6713
rect 1951 6711 2405 6733
rect 3055 6733 3199 6767
rect 3233 6733 3509 6767
rect 3851 6769 4123 6803
rect 4157 6769 4301 6803
rect 4955 6803 5405 6825
rect 3851 6753 4301 6769
rect 4343 6767 4797 6783
rect 3055 6711 3509 6733
rect 4343 6733 4487 6767
rect 4521 6733 4797 6767
rect 4955 6769 5227 6803
rect 5261 6769 5405 6803
rect 6059 6803 6509 6825
rect 4955 6753 5405 6769
rect 5447 6767 5901 6783
rect 4343 6711 4797 6733
rect 5447 6733 5591 6767
rect 5625 6733 5901 6767
rect 6059 6769 6331 6803
rect 6365 6769 6509 6803
rect 7163 6803 7613 6825
rect 6059 6753 6509 6769
rect 6551 6767 7005 6783
rect 5447 6711 5901 6733
rect 6551 6733 6695 6767
rect 6729 6733 7005 6767
rect 7163 6769 7435 6803
rect 7469 6769 7613 6803
rect 8267 6803 8443 6825
rect 7163 6753 7613 6769
rect 7655 6767 8109 6783
rect 6551 6711 7005 6733
rect 7655 6733 7799 6767
rect 7833 6733 8109 6767
rect 8267 6769 8283 6803
rect 8317 6769 8393 6803
rect 8427 6769 8443 6803
rect 9003 6803 9453 6825
rect 8267 6753 8443 6769
rect 8485 6767 8661 6783
rect 7655 6711 8109 6733
rect 8485 6733 8501 6767
rect 8535 6733 8611 6767
rect 8645 6733 8661 6767
rect 9003 6769 9275 6803
rect 9309 6769 9453 6803
rect 10107 6803 10557 6825
rect 9003 6753 9453 6769
rect 9495 6767 9949 6783
rect 8485 6711 8661 6733
rect 9495 6733 9639 6767
rect 9673 6733 9949 6767
rect 10107 6769 10379 6803
rect 10413 6769 10557 6803
rect 11211 6803 11661 6825
rect 10107 6753 10557 6769
rect 10599 6767 11053 6783
rect 9495 6711 9949 6733
rect 10599 6733 10743 6767
rect 10777 6733 11053 6767
rect 11211 6769 11483 6803
rect 11517 6769 11661 6803
rect 12315 6803 12765 6825
rect 11211 6753 11661 6769
rect 11703 6767 12157 6783
rect 10599 6711 11053 6733
rect 11703 6733 11847 6767
rect 11881 6733 12157 6767
rect 12315 6769 12587 6803
rect 12621 6769 12765 6803
rect 13419 6803 13595 6825
rect 12315 6753 12765 6769
rect 12807 6767 13261 6783
rect 11703 6711 12157 6733
rect 12807 6733 12951 6767
rect 12985 6733 13261 6767
rect 13419 6769 13435 6803
rect 13469 6769 13545 6803
rect 13579 6769 13595 6803
rect 14155 6803 14605 6825
rect 13419 6753 13595 6769
rect 13637 6767 13813 6783
rect 12807 6711 13261 6733
rect 13637 6733 13653 6767
rect 13687 6733 13763 6767
rect 13797 6733 13813 6767
rect 14155 6769 14427 6803
rect 14461 6769 14605 6803
rect 15259 6803 15709 6825
rect 14155 6753 14605 6769
rect 14647 6767 15101 6783
rect 13637 6711 13813 6733
rect 14647 6733 14791 6767
rect 14825 6733 15101 6767
rect 15259 6769 15531 6803
rect 15565 6769 15709 6803
rect 16363 6803 16813 6825
rect 15259 6753 15709 6769
rect 15751 6767 16205 6783
rect 14647 6711 15101 6733
rect 15751 6733 15895 6767
rect 15929 6733 16205 6767
rect 16363 6769 16635 6803
rect 16669 6769 16813 6803
rect 17467 6803 17917 6825
rect 18663 6821 18781 6851
rect 16363 6753 16813 6769
rect 16855 6767 17309 6783
rect 15751 6711 16205 6733
rect 16855 6733 16999 6767
rect 17033 6733 17309 6767
rect 17467 6769 17739 6803
rect 17773 6769 17917 6803
rect 18743 6819 18781 6821
rect 18743 6803 18809 6819
rect 17467 6753 17917 6769
rect 17959 6767 18413 6783
rect 16855 6711 17309 6733
rect 17959 6733 18103 6767
rect 18137 6733 18413 6767
rect 17959 6711 18413 6733
rect 18635 6763 18701 6779
rect 18635 6729 18651 6763
rect 18685 6729 18701 6763
rect 18743 6769 18759 6803
rect 18793 6769 18809 6803
rect 18743 6753 18809 6769
rect 18635 6713 18701 6729
rect 1183 6685 1301 6711
rect 1459 6685 2405 6711
rect 2563 6685 3509 6711
rect 3851 6685 4797 6711
rect 4955 6685 5901 6711
rect 6059 6685 7005 6711
rect 7163 6685 8109 6711
rect 8267 6685 8661 6711
rect 9003 6685 9949 6711
rect 10107 6685 11053 6711
rect 11211 6685 12157 6711
rect 12315 6685 13261 6711
rect 13419 6685 13813 6711
rect 14155 6685 15101 6711
rect 15259 6685 16205 6711
rect 16363 6685 17309 6711
rect 17467 6685 18413 6711
rect 18663 6711 18701 6713
rect 18663 6685 18781 6711
rect 1183 6549 1301 6575
rect 1459 6549 2405 6575
rect 2563 6549 3509 6575
rect 3851 6549 4797 6575
rect 4955 6549 5901 6575
rect 6059 6549 7005 6575
rect 7163 6549 8109 6575
rect 8267 6549 8661 6575
rect 9003 6549 9949 6575
rect 10107 6549 11053 6575
rect 11211 6549 12157 6575
rect 12315 6549 13261 6575
rect 13419 6549 13813 6575
rect 14155 6549 15101 6575
rect 15259 6549 16205 6575
rect 16363 6549 17309 6575
rect 17467 6549 18413 6575
rect 18663 6549 18781 6575
rect 1183 6481 1301 6507
rect 1459 6481 2405 6507
rect 2563 6481 3509 6507
rect 3667 6481 4613 6507
rect 4771 6481 5717 6507
rect 5875 6481 6085 6507
rect 6427 6481 7373 6507
rect 7531 6481 7925 6507
rect 8112 6481 8142 6507
rect 8196 6481 8226 6507
rect 8293 6481 8323 6507
rect 8543 6481 9489 6507
rect 9647 6481 10593 6507
rect 10751 6481 11329 6507
rect 11579 6481 12525 6507
rect 12683 6481 13629 6507
rect 13787 6481 14733 6507
rect 14891 6481 15837 6507
rect 15995 6481 16389 6507
rect 16731 6481 17677 6507
rect 17835 6481 18413 6507
rect 18663 6481 18781 6507
rect 1183 6345 1301 6371
rect 1459 6345 2405 6371
rect 2563 6345 3509 6371
rect 3667 6345 4613 6371
rect 4771 6345 5717 6371
rect 5875 6345 6085 6371
rect 6427 6345 7373 6371
rect 7531 6345 7925 6371
rect 1263 6343 1301 6345
rect 1263 6327 1329 6343
rect 1155 6287 1221 6303
rect 1155 6253 1171 6287
rect 1205 6253 1221 6287
rect 1263 6293 1279 6327
rect 1313 6293 1329 6327
rect 1951 6323 2405 6345
rect 1263 6277 1329 6293
rect 1459 6287 1909 6303
rect 1155 6237 1221 6253
rect 1183 6235 1221 6237
rect 1459 6253 1731 6287
rect 1765 6253 1909 6287
rect 1951 6289 2095 6323
rect 2129 6289 2405 6323
rect 3055 6323 3509 6345
rect 1951 6273 2405 6289
rect 2563 6287 3013 6303
rect 1183 6205 1301 6235
rect 1459 6231 1909 6253
rect 2563 6253 2835 6287
rect 2869 6253 3013 6287
rect 3055 6289 3199 6323
rect 3233 6289 3509 6323
rect 4159 6323 4613 6345
rect 3055 6273 3509 6289
rect 3667 6287 4117 6303
rect 2563 6231 3013 6253
rect 3667 6253 3939 6287
rect 3973 6253 4117 6287
rect 4159 6289 4303 6323
rect 4337 6289 4613 6323
rect 5263 6323 5717 6345
rect 4159 6273 4613 6289
rect 4771 6287 5221 6303
rect 3667 6231 4117 6253
rect 4771 6253 5043 6287
rect 5077 6253 5221 6287
rect 5263 6289 5407 6323
rect 5441 6289 5717 6323
rect 6001 6339 6085 6345
rect 6001 6323 6143 6339
rect 5263 6273 5717 6289
rect 5817 6287 5959 6303
rect 4771 6231 5221 6253
rect 5817 6253 5833 6287
rect 5867 6253 5959 6287
rect 6001 6289 6093 6323
rect 6127 6289 6143 6323
rect 6919 6323 7373 6345
rect 6001 6273 6143 6289
rect 6427 6287 6877 6303
rect 5817 6237 5959 6253
rect 5875 6231 5959 6237
rect 6427 6253 6699 6287
rect 6733 6253 6877 6287
rect 6919 6289 7063 6323
rect 7097 6289 7373 6323
rect 7749 6323 7925 6345
rect 8112 6329 8142 6397
rect 8196 6329 8226 6397
rect 8293 6329 8323 6351
rect 8543 6345 9489 6371
rect 9647 6345 10593 6371
rect 10751 6345 11329 6371
rect 11579 6345 12525 6371
rect 12683 6345 13629 6371
rect 13787 6345 14733 6371
rect 14891 6345 15837 6371
rect 15995 6345 16389 6371
rect 16731 6345 17677 6371
rect 17835 6345 18413 6371
rect 6919 6273 7373 6289
rect 7531 6287 7707 6303
rect 6427 6231 6877 6253
rect 7531 6253 7547 6287
rect 7581 6253 7657 6287
rect 7691 6253 7707 6287
rect 7749 6289 7765 6323
rect 7799 6289 7875 6323
rect 7909 6289 7925 6323
rect 7749 6273 7925 6289
rect 8054 6313 8154 6329
rect 8054 6279 8070 6313
rect 8104 6279 8154 6313
rect 8054 6263 8154 6279
rect 7531 6231 7707 6253
rect 8124 6231 8154 6263
rect 8196 6313 8250 6329
rect 8196 6279 8206 6313
rect 8240 6279 8250 6313
rect 8196 6263 8250 6279
rect 8293 6313 8359 6329
rect 8293 6279 8309 6313
rect 8343 6279 8359 6313
rect 9035 6323 9489 6345
rect 8293 6263 8359 6279
rect 8543 6287 8993 6303
rect 8196 6231 8226 6263
rect 8293 6231 8323 6263
rect 8543 6253 8815 6287
rect 8849 6253 8993 6287
rect 9035 6289 9179 6323
rect 9213 6289 9489 6323
rect 10139 6323 10593 6345
rect 9035 6273 9489 6289
rect 9647 6287 10097 6303
rect 8543 6231 8993 6253
rect 9647 6253 9919 6287
rect 9953 6253 10097 6287
rect 10139 6289 10283 6323
rect 10317 6289 10593 6323
rect 11057 6323 11329 6345
rect 10139 6273 10593 6289
rect 10751 6287 11015 6303
rect 9647 6231 10097 6253
rect 10751 6253 10767 6287
rect 10801 6253 10866 6287
rect 10900 6253 10965 6287
rect 10999 6253 11015 6287
rect 11057 6289 11073 6323
rect 11107 6289 11176 6323
rect 11210 6289 11279 6323
rect 11313 6289 11329 6323
rect 12071 6323 12525 6345
rect 11057 6273 11329 6289
rect 11579 6287 12029 6303
rect 10751 6231 11015 6253
rect 11579 6253 11851 6287
rect 11885 6253 12029 6287
rect 12071 6289 12215 6323
rect 12249 6289 12525 6323
rect 13175 6323 13629 6345
rect 12071 6273 12525 6289
rect 12683 6287 13133 6303
rect 11579 6231 12029 6253
rect 12683 6253 12955 6287
rect 12989 6253 13133 6287
rect 13175 6289 13319 6323
rect 13353 6289 13629 6323
rect 14279 6323 14733 6345
rect 13175 6273 13629 6289
rect 13787 6287 14237 6303
rect 12683 6231 13133 6253
rect 13787 6253 14059 6287
rect 14093 6253 14237 6287
rect 14279 6289 14423 6323
rect 14457 6289 14733 6323
rect 15383 6323 15837 6345
rect 14279 6273 14733 6289
rect 14891 6287 15341 6303
rect 13787 6231 14237 6253
rect 14891 6253 15163 6287
rect 15197 6253 15341 6287
rect 15383 6289 15527 6323
rect 15561 6289 15837 6323
rect 16213 6323 16389 6345
rect 15383 6273 15837 6289
rect 15995 6287 16171 6303
rect 14891 6231 15341 6253
rect 15995 6253 16011 6287
rect 16045 6253 16121 6287
rect 16155 6253 16171 6287
rect 16213 6289 16229 6323
rect 16263 6289 16339 6323
rect 16373 6289 16389 6323
rect 17223 6323 17677 6345
rect 16213 6273 16389 6289
rect 16731 6287 17181 6303
rect 15995 6231 16171 6253
rect 16731 6253 17003 6287
rect 17037 6253 17181 6287
rect 17223 6289 17367 6323
rect 17401 6289 17677 6323
rect 18141 6323 18413 6345
rect 18663 6345 18781 6371
rect 18663 6343 18701 6345
rect 17223 6273 17677 6289
rect 17835 6287 18099 6303
rect 16731 6231 17181 6253
rect 17835 6253 17851 6287
rect 17885 6253 17950 6287
rect 17984 6253 18049 6287
rect 18083 6253 18099 6287
rect 18141 6289 18157 6323
rect 18191 6289 18260 6323
rect 18294 6289 18363 6323
rect 18397 6289 18413 6323
rect 18141 6273 18413 6289
rect 18635 6327 18701 6343
rect 18635 6293 18651 6327
rect 18685 6293 18701 6327
rect 18635 6277 18701 6293
rect 18743 6287 18809 6303
rect 17835 6231 18099 6253
rect 18743 6253 18759 6287
rect 18793 6253 18809 6287
rect 18743 6237 18809 6253
rect 18743 6235 18781 6237
rect 1459 6205 2405 6231
rect 2563 6205 3509 6231
rect 3667 6205 4613 6231
rect 4771 6205 5717 6231
rect 5875 6205 6085 6231
rect 6427 6205 7373 6231
rect 7531 6205 7925 6231
rect 8124 6121 8154 6147
rect 8196 6121 8226 6147
rect 8543 6205 9489 6231
rect 9647 6205 10593 6231
rect 10751 6205 11329 6231
rect 11579 6205 12525 6231
rect 12683 6205 13629 6231
rect 13787 6205 14733 6231
rect 14891 6205 15837 6231
rect 15995 6205 16389 6231
rect 16731 6205 17677 6231
rect 17835 6205 18413 6231
rect 18663 6205 18781 6235
rect 1183 6005 1301 6031
rect 1459 6005 2405 6031
rect 2563 6005 3509 6031
rect 3667 6005 4613 6031
rect 4771 6005 5717 6031
rect 5875 6005 6085 6031
rect 6427 6005 7373 6031
rect 7531 6005 7925 6031
rect 8293 6005 8323 6031
rect 8543 6005 9489 6031
rect 9647 6005 10593 6031
rect 10751 6005 11329 6031
rect 11579 6005 12525 6031
rect 12683 6005 13629 6031
rect 13787 6005 14733 6031
rect 14891 6005 15837 6031
rect 15995 6005 16389 6031
rect 16731 6005 17677 6031
rect 17835 6005 18413 6031
rect 18663 6005 18781 6031
rect 1183 5937 1301 5963
rect 1459 5937 2405 5963
rect 2563 5937 3509 5963
rect 3851 5937 4797 5963
rect 4955 5937 5901 5963
rect 6059 5937 6637 5963
rect 6795 5937 6825 5963
rect 6883 5937 6913 5963
rect 7071 5937 7465 5963
rect 8263 5937 8293 5963
rect 8451 5937 8661 5963
rect 9003 5937 9949 5963
rect 10107 5937 11053 5963
rect 11211 5937 11421 5963
rect 11789 5937 11819 5963
rect 12039 5937 12617 5963
rect 13077 5937 13107 5963
rect 13327 5937 13905 5963
rect 14155 5937 15101 5963
rect 15259 5937 16205 5963
rect 16363 5937 17309 5963
rect 17467 5937 18413 5963
rect 18663 5937 18781 5963
rect 1183 5733 1301 5763
rect 1459 5737 2405 5763
rect 2563 5737 3509 5763
rect 3851 5737 4797 5763
rect 4955 5737 5901 5763
rect 6059 5737 6637 5763
rect 1183 5731 1221 5733
rect 1155 5715 1221 5731
rect 1155 5681 1171 5715
rect 1205 5681 1221 5715
rect 1459 5715 1909 5737
rect 1155 5665 1221 5681
rect 1263 5675 1329 5691
rect 1263 5641 1279 5675
rect 1313 5641 1329 5675
rect 1459 5681 1731 5715
rect 1765 5681 1909 5715
rect 2563 5715 3013 5737
rect 1459 5665 1909 5681
rect 1951 5679 2405 5695
rect 1263 5625 1329 5641
rect 1951 5645 2095 5679
rect 2129 5645 2405 5679
rect 2563 5681 2835 5715
rect 2869 5681 3013 5715
rect 3851 5715 4301 5737
rect 2563 5665 3013 5681
rect 3055 5679 3509 5695
rect 1263 5623 1301 5625
rect 1951 5623 2405 5645
rect 3055 5645 3199 5679
rect 3233 5645 3509 5679
rect 3851 5681 4123 5715
rect 4157 5681 4301 5715
rect 4955 5715 5405 5737
rect 3851 5665 4301 5681
rect 4343 5679 4797 5695
rect 3055 5623 3509 5645
rect 4343 5645 4487 5679
rect 4521 5645 4797 5679
rect 4955 5681 5227 5715
rect 5261 5681 5405 5715
rect 6059 5715 6323 5737
rect 6795 5718 6825 5779
rect 6883 5764 6913 5779
rect 6883 5740 6919 5764
rect 7669 5898 7699 5924
rect 7765 5898 7795 5924
rect 7837 5898 7867 5924
rect 8051 5898 8081 5924
rect 8154 5898 8184 5924
rect 7669 5782 7699 5814
rect 7669 5766 7723 5782
rect 4955 5665 5405 5681
rect 5447 5679 5901 5695
rect 4343 5623 4797 5645
rect 5447 5645 5591 5679
rect 5625 5645 5901 5679
rect 6059 5681 6075 5715
rect 6109 5681 6174 5715
rect 6208 5681 6273 5715
rect 6307 5681 6323 5715
rect 6791 5702 6845 5718
rect 6059 5665 6323 5681
rect 6365 5679 6637 5695
rect 5447 5623 5901 5645
rect 6365 5645 6381 5679
rect 6415 5645 6484 5679
rect 6518 5645 6587 5679
rect 6621 5645 6637 5679
rect 6791 5668 6801 5702
rect 6835 5668 6845 5702
rect 6791 5652 6845 5668
rect 6889 5705 6919 5740
rect 7071 5737 7465 5763
rect 7071 5715 7247 5737
rect 6889 5689 6965 5705
rect 6889 5655 6921 5689
rect 6955 5655 6965 5689
rect 7071 5681 7087 5715
rect 7121 5681 7197 5715
rect 7231 5681 7247 5715
rect 7669 5732 7679 5766
rect 7713 5732 7723 5766
rect 7669 5716 7723 5732
rect 7071 5665 7247 5681
rect 7289 5679 7465 5695
rect 6365 5623 6637 5645
rect 1183 5597 1301 5623
rect 1459 5597 2405 5623
rect 2563 5597 3509 5623
rect 3851 5597 4797 5623
rect 4955 5597 5901 5623
rect 6059 5597 6637 5623
rect 6795 5591 6825 5652
rect 6889 5639 6965 5655
rect 7289 5645 7305 5679
rect 7339 5645 7415 5679
rect 7449 5645 7465 5679
rect 6889 5630 6919 5639
rect 6883 5606 6919 5630
rect 7289 5623 7465 5645
rect 6883 5591 6913 5606
rect 7071 5597 7465 5623
rect 7669 5571 7699 5716
rect 7765 5663 7795 5814
rect 7837 5782 7867 5814
rect 8051 5799 8081 5814
rect 7837 5766 7891 5782
rect 7837 5732 7847 5766
rect 7881 5732 7891 5766
rect 7837 5716 7891 5732
rect 7933 5769 8081 5799
rect 7933 5669 7963 5769
rect 8154 5705 8184 5814
rect 8451 5737 8661 5763
rect 11620 5821 11650 5847
rect 11692 5821 11722 5847
rect 9003 5737 9949 5763
rect 10107 5737 11053 5763
rect 11211 5737 11421 5763
rect 12908 5821 12938 5847
rect 12980 5821 13010 5847
rect 12039 5737 12617 5763
rect 13327 5737 13905 5763
rect 14155 5737 15101 5763
rect 15259 5737 16205 5763
rect 16363 5737 17309 5763
rect 17467 5737 18413 5763
rect 8263 5705 8293 5737
rect 8451 5731 8535 5737
rect 8393 5715 8535 5731
rect 8146 5689 8200 5705
rect 7741 5653 7807 5663
rect 7741 5619 7757 5653
rect 7791 5639 7807 5653
rect 7909 5653 7963 5669
rect 7791 5619 7867 5639
rect 7741 5609 7867 5619
rect 7837 5571 7867 5609
rect 7909 5619 7919 5653
rect 7953 5619 7963 5653
rect 7909 5603 7963 5619
rect 8005 5653 8088 5669
rect 8005 5619 8015 5653
rect 8049 5619 8088 5653
rect 8146 5655 8156 5689
rect 8190 5655 8200 5689
rect 8146 5639 8200 5655
rect 8242 5689 8296 5705
rect 8242 5655 8252 5689
rect 8286 5655 8296 5689
rect 8393 5681 8409 5715
rect 8443 5681 8535 5715
rect 9003 5715 9453 5737
rect 8393 5665 8535 5681
rect 8577 5679 8719 5695
rect 8242 5639 8296 5655
rect 8577 5645 8669 5679
rect 8703 5645 8719 5679
rect 9003 5681 9275 5715
rect 9309 5681 9453 5715
rect 10107 5715 10557 5737
rect 11211 5731 11295 5737
rect 9003 5665 9453 5681
rect 9495 5679 9949 5695
rect 8005 5603 8088 5619
rect 7933 5571 7963 5603
rect 8058 5571 8088 5603
rect 8154 5571 8184 5639
rect 8263 5617 8293 5639
rect 8577 5629 8719 5645
rect 9495 5645 9639 5679
rect 9673 5645 9949 5679
rect 10107 5681 10379 5715
rect 10413 5681 10557 5715
rect 11153 5715 11295 5731
rect 10107 5665 10557 5681
rect 10599 5679 11053 5695
rect 8577 5623 8661 5629
rect 9495 5623 9949 5645
rect 10599 5645 10743 5679
rect 10777 5645 11053 5679
rect 11153 5681 11169 5715
rect 11203 5681 11295 5715
rect 11620 5705 11650 5737
rect 11153 5665 11295 5681
rect 11337 5679 11479 5695
rect 10599 5623 11053 5645
rect 11337 5645 11429 5679
rect 11463 5645 11479 5679
rect 11337 5629 11479 5645
rect 11550 5689 11650 5705
rect 11550 5655 11566 5689
rect 11600 5655 11650 5689
rect 11550 5639 11650 5655
rect 11692 5705 11722 5737
rect 11789 5705 11819 5737
rect 12039 5715 12303 5737
rect 11692 5689 11746 5705
rect 11692 5655 11702 5689
rect 11736 5655 11746 5689
rect 11692 5639 11746 5655
rect 11789 5689 11855 5705
rect 11789 5655 11805 5689
rect 11839 5655 11855 5689
rect 12039 5681 12055 5715
rect 12089 5681 12154 5715
rect 12188 5681 12253 5715
rect 12287 5681 12303 5715
rect 12908 5705 12938 5737
rect 12039 5665 12303 5681
rect 12345 5679 12617 5695
rect 11789 5639 11855 5655
rect 12345 5645 12361 5679
rect 12395 5645 12464 5679
rect 12498 5645 12567 5679
rect 12601 5645 12617 5679
rect 11337 5623 11421 5629
rect 8451 5597 8661 5623
rect 9003 5597 9949 5623
rect 10107 5597 11053 5623
rect 11211 5597 11421 5623
rect 11608 5571 11638 5639
rect 11692 5571 11722 5639
rect 11789 5617 11819 5639
rect 12345 5623 12617 5645
rect 12838 5689 12938 5705
rect 12838 5655 12854 5689
rect 12888 5655 12938 5689
rect 12838 5639 12938 5655
rect 12980 5705 13010 5737
rect 13077 5705 13107 5737
rect 13327 5715 13591 5737
rect 12980 5689 13034 5705
rect 12980 5655 12990 5689
rect 13024 5655 13034 5689
rect 12980 5639 13034 5655
rect 13077 5689 13143 5705
rect 13077 5655 13093 5689
rect 13127 5655 13143 5689
rect 13327 5681 13343 5715
rect 13377 5681 13442 5715
rect 13476 5681 13541 5715
rect 13575 5681 13591 5715
rect 14155 5715 14605 5737
rect 13327 5665 13591 5681
rect 13633 5679 13905 5695
rect 13077 5639 13143 5655
rect 13633 5645 13649 5679
rect 13683 5645 13752 5679
rect 13786 5645 13855 5679
rect 13889 5645 13905 5679
rect 14155 5681 14427 5715
rect 14461 5681 14605 5715
rect 15259 5715 15709 5737
rect 14155 5665 14605 5681
rect 14647 5679 15101 5695
rect 12039 5597 12617 5623
rect 12896 5571 12926 5639
rect 12980 5571 13010 5639
rect 13077 5617 13107 5639
rect 13633 5623 13905 5645
rect 14647 5645 14791 5679
rect 14825 5645 15101 5679
rect 15259 5681 15531 5715
rect 15565 5681 15709 5715
rect 16363 5715 16813 5737
rect 15259 5665 15709 5681
rect 15751 5679 16205 5695
rect 14647 5623 15101 5645
rect 15751 5645 15895 5679
rect 15929 5645 16205 5679
rect 16363 5681 16635 5715
rect 16669 5681 16813 5715
rect 17467 5715 17917 5737
rect 18663 5733 18781 5763
rect 16363 5665 16813 5681
rect 16855 5679 17309 5695
rect 15751 5623 16205 5645
rect 16855 5645 16999 5679
rect 17033 5645 17309 5679
rect 17467 5681 17739 5715
rect 17773 5681 17917 5715
rect 18743 5731 18781 5733
rect 18743 5715 18809 5731
rect 17467 5665 17917 5681
rect 17959 5679 18413 5695
rect 16855 5623 17309 5645
rect 17959 5645 18103 5679
rect 18137 5645 18413 5679
rect 17959 5623 18413 5645
rect 18635 5675 18701 5691
rect 18635 5641 18651 5675
rect 18685 5641 18701 5675
rect 18743 5681 18759 5715
rect 18793 5681 18809 5715
rect 18743 5665 18809 5681
rect 18635 5625 18701 5641
rect 13327 5597 13905 5623
rect 14155 5597 15101 5623
rect 15259 5597 16205 5623
rect 16363 5597 17309 5623
rect 17467 5597 18413 5623
rect 18663 5623 18701 5625
rect 18663 5597 18781 5623
rect 1183 5461 1301 5487
rect 1459 5461 2405 5487
rect 2563 5461 3509 5487
rect 3851 5461 4797 5487
rect 4955 5461 5901 5487
rect 6059 5461 6637 5487
rect 6795 5461 6825 5487
rect 6883 5461 6913 5487
rect 7071 5461 7465 5487
rect 7669 5461 7699 5487
rect 7837 5461 7867 5487
rect 7933 5461 7963 5487
rect 8058 5461 8088 5487
rect 8154 5461 8184 5487
rect 8263 5461 8293 5487
rect 8451 5461 8661 5487
rect 9003 5461 9949 5487
rect 10107 5461 11053 5487
rect 11211 5461 11421 5487
rect 11608 5461 11638 5487
rect 11692 5461 11722 5487
rect 11789 5461 11819 5487
rect 12039 5461 12617 5487
rect 12896 5461 12926 5487
rect 12980 5461 13010 5487
rect 13077 5461 13107 5487
rect 13327 5461 13905 5487
rect 14155 5461 15101 5487
rect 15259 5461 16205 5487
rect 16363 5461 17309 5487
rect 17467 5461 18413 5487
rect 18663 5461 18781 5487
rect 1183 5393 1301 5419
rect 1459 5393 2405 5419
rect 2563 5393 2681 5419
rect 2839 5393 2869 5419
rect 2923 5393 2953 5419
rect 3178 5393 3208 5419
rect 3273 5393 3303 5419
rect 3369 5393 3399 5419
rect 3535 5393 3565 5419
rect 3607 5393 3637 5419
rect 3739 5393 3769 5419
rect 3838 5393 3868 5419
rect 3947 5393 3977 5419
rect 4043 5393 4073 5419
rect 4192 5393 4222 5419
rect 4283 5393 4313 5419
rect 4491 5393 4521 5419
rect 4679 5393 5625 5419
rect 5783 5393 6177 5419
rect 6427 5393 6545 5419
rect 6703 5393 6733 5419
rect 6812 5393 6842 5419
rect 6908 5393 6938 5419
rect 7033 5393 7063 5419
rect 7129 5393 7159 5419
rect 7297 5393 7327 5419
rect 7531 5393 7741 5419
rect 7899 5393 7929 5419
rect 7983 5393 8013 5419
rect 8238 5393 8268 5419
rect 8333 5393 8363 5419
rect 8429 5393 8459 5419
rect 8595 5393 8625 5419
rect 8667 5393 8697 5419
rect 8799 5393 8829 5419
rect 8898 5393 8928 5419
rect 9007 5393 9037 5419
rect 9103 5393 9133 5419
rect 9252 5393 9282 5419
rect 9343 5393 9373 5419
rect 9551 5393 9581 5419
rect 9739 5393 9949 5419
rect 10153 5393 10183 5419
rect 10321 5393 10351 5419
rect 10417 5393 10447 5419
rect 10542 5393 10572 5419
rect 10638 5393 10668 5419
rect 10747 5393 10777 5419
rect 10935 5393 11329 5419
rect 11763 5393 11793 5419
rect 11872 5393 11902 5419
rect 11968 5393 11998 5419
rect 12093 5393 12123 5419
rect 12189 5393 12219 5419
rect 12357 5393 12387 5419
rect 12591 5393 12801 5419
rect 13005 5393 13035 5419
rect 13173 5393 13203 5419
rect 13269 5393 13299 5419
rect 13394 5393 13424 5419
rect 13490 5393 13520 5419
rect 13599 5393 13629 5419
rect 13787 5393 14733 5419
rect 14891 5393 15837 5419
rect 15995 5393 16389 5419
rect 16731 5393 17677 5419
rect 17835 5393 18413 5419
rect 18663 5393 18781 5419
rect 2839 5294 2869 5309
rect 1183 5257 1301 5283
rect 1459 5257 2405 5283
rect 2563 5257 2681 5283
rect 1263 5255 1301 5257
rect 1263 5239 1329 5255
rect 1155 5199 1221 5215
rect 1155 5165 1171 5199
rect 1205 5165 1221 5199
rect 1263 5205 1279 5239
rect 1313 5205 1329 5239
rect 1951 5235 2405 5257
rect 1263 5189 1329 5205
rect 1459 5199 1909 5215
rect 1155 5149 1221 5165
rect 1183 5147 1221 5149
rect 1459 5165 1731 5199
rect 1765 5165 1909 5199
rect 1951 5201 2095 5235
rect 2129 5201 2405 5235
rect 2643 5255 2681 5257
rect 2806 5264 2869 5294
rect 2643 5239 2709 5255
rect 2806 5241 2836 5264
rect 1951 5185 2405 5201
rect 2535 5199 2601 5215
rect 1183 5117 1301 5147
rect 1459 5143 1909 5165
rect 2535 5165 2551 5199
rect 2585 5165 2601 5199
rect 2643 5205 2659 5239
rect 2693 5205 2709 5239
rect 2643 5189 2709 5205
rect 2782 5225 2836 5241
rect 2782 5191 2792 5225
rect 2826 5191 2836 5225
rect 2923 5220 2953 5309
rect 2782 5175 2836 5191
rect 2535 5149 2601 5165
rect 2563 5147 2601 5149
rect 1459 5117 2405 5143
rect 2563 5117 2681 5147
rect 2806 5122 2836 5175
rect 2878 5210 2953 5220
rect 2878 5176 2894 5210
rect 2928 5176 2953 5210
rect 3178 5180 3208 5309
rect 3273 5287 3303 5321
rect 3369 5287 3399 5321
rect 3250 5271 3304 5287
rect 3250 5237 3260 5271
rect 3294 5237 3304 5271
rect 3250 5221 3304 5237
rect 3346 5277 3412 5287
rect 3346 5243 3362 5277
rect 3396 5243 3412 5277
rect 3346 5233 3412 5243
rect 2878 5166 2953 5176
rect 2806 5092 2869 5122
rect 2839 5077 2869 5092
rect 2923 5077 2953 5166
rect 3091 5164 3208 5180
rect 3091 5130 3101 5164
rect 3135 5144 3208 5164
rect 3273 5191 3304 5221
rect 3273 5161 3411 5191
rect 3135 5130 3220 5144
rect 3091 5114 3220 5130
rect 3190 5027 3220 5114
rect 3266 5109 3332 5119
rect 3266 5075 3282 5109
rect 3316 5075 3332 5109
rect 3266 5065 3332 5075
rect 3282 5027 3312 5065
rect 3381 5027 3411 5161
rect 3535 5151 3565 5309
rect 3607 5287 3637 5309
rect 3607 5271 3661 5287
rect 3607 5237 3617 5271
rect 3651 5237 3661 5271
rect 3838 5299 3868 5321
rect 3838 5283 3905 5299
rect 3739 5239 3769 5265
rect 3607 5221 3661 5237
rect 3703 5223 3769 5239
rect 3838 5249 3861 5283
rect 3895 5249 3905 5283
rect 3838 5233 3905 5249
rect 3947 5251 3977 5321
rect 4043 5277 4073 5309
rect 4043 5261 4145 5277
rect 3947 5235 4001 5251
rect 4043 5247 4101 5261
rect 3521 5135 3576 5151
rect 3521 5101 3531 5135
rect 3565 5101 3576 5135
rect 3521 5085 3576 5101
rect 3521 5027 3551 5085
rect 3618 5027 3648 5221
rect 3703 5189 3713 5223
rect 3747 5189 3769 5223
rect 3947 5203 3957 5235
rect 3935 5201 3957 5203
rect 3991 5201 4001 5235
rect 3935 5191 4001 5201
rect 3703 5173 3769 5189
rect 3739 5156 3769 5173
rect 3914 5185 4001 5191
rect 4084 5227 4101 5247
rect 4135 5227 4145 5261
rect 4192 5249 4222 5309
rect 4084 5211 4145 5227
rect 4187 5233 4241 5249
rect 3914 5173 3977 5185
rect 3914 5161 3964 5173
rect 3739 5126 3845 5156
rect 3815 5111 3845 5126
rect 1183 4917 1301 4943
rect 1459 4917 2405 4943
rect 2563 4917 2681 4943
rect 2839 4923 2869 4949
rect 2923 4923 2953 4949
rect 3914 5027 3944 5161
rect 3986 5109 4040 5125
rect 3986 5075 3996 5109
rect 4030 5075 4040 5109
rect 3986 5059 4040 5075
rect 4000 5027 4030 5059
rect 4084 5027 4114 5211
rect 4187 5199 4197 5233
rect 4231 5199 4241 5233
rect 4187 5183 4241 5199
rect 4192 5027 4222 5183
rect 4283 5141 4313 5309
rect 4491 5241 4521 5263
rect 4679 5257 5625 5283
rect 5783 5257 6177 5283
rect 6427 5257 6545 5283
rect 4462 5225 4521 5241
rect 4462 5191 4472 5225
rect 4506 5191 4521 5225
rect 5171 5235 5625 5257
rect 4462 5175 4521 5191
rect 4491 5143 4521 5175
rect 4679 5199 5129 5215
rect 4679 5165 4951 5199
rect 4985 5165 5129 5199
rect 5171 5201 5315 5235
rect 5349 5201 5625 5235
rect 6001 5235 6177 5257
rect 5171 5185 5625 5201
rect 5783 5199 5959 5215
rect 4679 5143 5129 5165
rect 5783 5165 5799 5199
rect 5833 5165 5909 5199
rect 5943 5165 5959 5199
rect 6001 5201 6017 5235
rect 6051 5201 6127 5235
rect 6161 5201 6177 5235
rect 6507 5255 6545 5257
rect 6507 5239 6573 5255
rect 6703 5241 6733 5263
rect 6812 5241 6842 5309
rect 6908 5277 6938 5309
rect 7033 5277 7063 5309
rect 6908 5261 6991 5277
rect 6001 5185 6177 5201
rect 6399 5199 6465 5215
rect 5783 5143 5959 5165
rect 6399 5165 6415 5199
rect 6449 5165 6465 5199
rect 6507 5205 6523 5239
rect 6557 5205 6573 5239
rect 6507 5189 6573 5205
rect 6700 5225 6754 5241
rect 6700 5191 6710 5225
rect 6744 5191 6754 5225
rect 6700 5175 6754 5191
rect 6796 5225 6850 5241
rect 6796 5191 6806 5225
rect 6840 5191 6850 5225
rect 6908 5227 6947 5261
rect 6981 5227 6991 5261
rect 6908 5211 6991 5227
rect 7033 5261 7087 5277
rect 7033 5227 7043 5261
rect 7077 5227 7087 5261
rect 7129 5271 7159 5309
rect 7129 5261 7255 5271
rect 7129 5241 7205 5261
rect 7033 5211 7087 5227
rect 7189 5227 7205 5241
rect 7239 5227 7255 5261
rect 7189 5217 7255 5227
rect 6796 5175 6850 5191
rect 6399 5149 6465 5165
rect 6427 5147 6465 5149
rect 4264 5125 4318 5141
rect 4264 5091 4274 5125
rect 4308 5091 4318 5125
rect 4264 5075 4318 5091
rect 4276 5027 4306 5075
rect 4679 5117 5625 5143
rect 5783 5117 6177 5143
rect 6427 5117 6545 5147
rect 6703 5143 6733 5175
rect 6812 5066 6842 5175
rect 7033 5111 7063 5211
rect 6915 5081 7063 5111
rect 7105 5148 7159 5164
rect 7105 5114 7115 5148
rect 7149 5114 7159 5148
rect 7105 5098 7159 5114
rect 6915 5066 6945 5081
rect 7129 5066 7159 5098
rect 7201 5066 7231 5217
rect 7297 5164 7327 5309
rect 7899 5294 7929 5309
rect 7531 5257 7741 5283
rect 7657 5251 7741 5257
rect 7866 5264 7929 5294
rect 7657 5235 7799 5251
rect 7866 5241 7896 5264
rect 7273 5148 7327 5164
rect 7473 5199 7615 5215
rect 7473 5165 7489 5199
rect 7523 5165 7615 5199
rect 7657 5201 7749 5235
rect 7783 5201 7799 5235
rect 7657 5185 7799 5201
rect 7842 5225 7896 5241
rect 7842 5191 7852 5225
rect 7886 5191 7896 5225
rect 7983 5220 8013 5309
rect 7842 5175 7896 5191
rect 7473 5149 7615 5165
rect 7273 5114 7283 5148
rect 7317 5114 7327 5148
rect 7531 5143 7615 5149
rect 7531 5117 7741 5143
rect 7866 5122 7896 5175
rect 7938 5210 8013 5220
rect 7938 5176 7954 5210
rect 7988 5176 8013 5210
rect 8238 5180 8268 5309
rect 8333 5287 8363 5321
rect 8429 5287 8459 5321
rect 8310 5271 8364 5287
rect 8310 5237 8320 5271
rect 8354 5237 8364 5271
rect 8310 5221 8364 5237
rect 8406 5277 8472 5287
rect 8406 5243 8422 5277
rect 8456 5243 8472 5277
rect 8406 5233 8472 5243
rect 7938 5166 8013 5176
rect 7273 5098 7327 5114
rect 7297 5066 7327 5098
rect 6812 4956 6842 4982
rect 6915 4956 6945 4982
rect 7129 4956 7159 4982
rect 7201 4956 7231 4982
rect 7297 4956 7327 4982
rect 7866 5092 7929 5122
rect 7899 5077 7929 5092
rect 7983 5077 8013 5166
rect 8151 5164 8268 5180
rect 8151 5130 8161 5164
rect 8195 5144 8268 5164
rect 8333 5191 8364 5221
rect 8333 5161 8471 5191
rect 8195 5130 8280 5144
rect 8151 5114 8280 5130
rect 8250 5027 8280 5114
rect 8326 5109 8392 5119
rect 8326 5075 8342 5109
rect 8376 5075 8392 5109
rect 8326 5065 8392 5075
rect 8342 5027 8372 5065
rect 8441 5027 8471 5161
rect 8595 5151 8625 5309
rect 8667 5287 8697 5309
rect 8667 5271 8721 5287
rect 8667 5237 8677 5271
rect 8711 5237 8721 5271
rect 8898 5299 8928 5321
rect 8898 5283 8965 5299
rect 8799 5239 8829 5265
rect 8667 5221 8721 5237
rect 8763 5223 8829 5239
rect 8898 5249 8921 5283
rect 8955 5249 8965 5283
rect 8898 5233 8965 5249
rect 9007 5251 9037 5321
rect 9103 5277 9133 5309
rect 9103 5261 9205 5277
rect 9007 5235 9061 5251
rect 9103 5247 9161 5261
rect 8581 5135 8636 5151
rect 8581 5101 8591 5135
rect 8625 5101 8636 5135
rect 8581 5085 8636 5101
rect 8581 5027 8611 5085
rect 8678 5027 8708 5221
rect 8763 5189 8773 5223
rect 8807 5189 8829 5223
rect 9007 5203 9017 5235
rect 8995 5201 9017 5203
rect 9051 5201 9061 5235
rect 8995 5191 9061 5201
rect 8763 5173 8829 5189
rect 8799 5156 8829 5173
rect 8974 5185 9061 5191
rect 9144 5227 9161 5247
rect 9195 5227 9205 5261
rect 9252 5249 9282 5309
rect 9144 5211 9205 5227
rect 9247 5233 9301 5249
rect 8974 5173 9037 5185
rect 8974 5161 9024 5173
rect 8799 5126 8905 5156
rect 8875 5111 8905 5126
rect 3190 4917 3220 4943
rect 3282 4917 3312 4943
rect 3381 4917 3411 4943
rect 3521 4917 3551 4943
rect 3618 4917 3648 4943
rect 3815 4917 3845 4943
rect 3914 4917 3944 4943
rect 4000 4917 4030 4943
rect 4084 4917 4114 4943
rect 4192 4917 4222 4943
rect 4276 4917 4306 4943
rect 4491 4917 4521 4943
rect 4679 4917 5625 4943
rect 5783 4917 6177 4943
rect 6427 4917 6545 4943
rect 6703 4917 6733 4943
rect 7531 4917 7741 4943
rect 7899 4923 7929 4949
rect 7983 4923 8013 4949
rect 8974 5027 9004 5161
rect 9046 5109 9100 5125
rect 9046 5075 9056 5109
rect 9090 5075 9100 5109
rect 9046 5059 9100 5075
rect 9060 5027 9090 5059
rect 9144 5027 9174 5211
rect 9247 5199 9257 5233
rect 9291 5199 9301 5233
rect 9247 5183 9301 5199
rect 9252 5027 9282 5183
rect 9343 5141 9373 5309
rect 9551 5241 9581 5263
rect 9739 5257 9949 5283
rect 9522 5225 9581 5241
rect 9522 5191 9532 5225
rect 9566 5191 9581 5225
rect 9865 5251 9949 5257
rect 9865 5235 10007 5251
rect 9522 5175 9581 5191
rect 9551 5143 9581 5175
rect 9681 5199 9823 5215
rect 9681 5165 9697 5199
rect 9731 5165 9823 5199
rect 9865 5201 9957 5235
rect 9991 5201 10007 5235
rect 9865 5185 10007 5201
rect 9681 5149 9823 5165
rect 9739 5143 9823 5149
rect 10153 5164 10183 5309
rect 10321 5271 10351 5309
rect 10417 5277 10447 5309
rect 10542 5277 10572 5309
rect 10225 5261 10351 5271
rect 10225 5227 10241 5261
rect 10275 5241 10351 5261
rect 10393 5261 10447 5277
rect 10275 5227 10291 5241
rect 10225 5217 10291 5227
rect 10393 5227 10403 5261
rect 10437 5227 10447 5261
rect 10153 5148 10207 5164
rect 9324 5125 9378 5141
rect 9324 5091 9334 5125
rect 9368 5091 9378 5125
rect 9324 5075 9378 5091
rect 9336 5027 9366 5075
rect 9739 5117 9949 5143
rect 10153 5114 10163 5148
rect 10197 5114 10207 5148
rect 10153 5098 10207 5114
rect 10153 5066 10183 5098
rect 10249 5066 10279 5217
rect 10393 5211 10447 5227
rect 10489 5261 10572 5277
rect 10489 5227 10499 5261
rect 10533 5227 10572 5261
rect 10638 5241 10668 5309
rect 10747 5241 10777 5263
rect 10935 5257 11329 5283
rect 10489 5211 10572 5227
rect 10630 5225 10684 5241
rect 10321 5148 10375 5164
rect 10321 5114 10331 5148
rect 10365 5114 10375 5148
rect 10321 5098 10375 5114
rect 10417 5111 10447 5211
rect 10630 5191 10640 5225
rect 10674 5191 10684 5225
rect 10630 5175 10684 5191
rect 10726 5225 10780 5241
rect 10726 5191 10736 5225
rect 10770 5191 10780 5225
rect 11153 5235 11329 5257
rect 11763 5241 11793 5263
rect 11872 5241 11902 5309
rect 11968 5277 11998 5309
rect 12093 5277 12123 5309
rect 11968 5261 12051 5277
rect 10726 5175 10780 5191
rect 10935 5199 11111 5215
rect 10321 5066 10351 5098
rect 10417 5081 10565 5111
rect 10535 5066 10565 5081
rect 10638 5066 10668 5175
rect 10747 5143 10777 5175
rect 10935 5165 10951 5199
rect 10985 5165 11061 5199
rect 11095 5165 11111 5199
rect 11153 5201 11169 5235
rect 11203 5201 11279 5235
rect 11313 5201 11329 5235
rect 11153 5185 11329 5201
rect 11760 5225 11814 5241
rect 11760 5191 11770 5225
rect 11804 5191 11814 5225
rect 11760 5175 11814 5191
rect 11856 5225 11910 5241
rect 11856 5191 11866 5225
rect 11900 5191 11910 5225
rect 11968 5227 12007 5261
rect 12041 5227 12051 5261
rect 11968 5211 12051 5227
rect 12093 5261 12147 5277
rect 12093 5227 12103 5261
rect 12137 5227 12147 5261
rect 12189 5271 12219 5309
rect 12189 5261 12315 5271
rect 12189 5241 12265 5261
rect 12093 5211 12147 5227
rect 12249 5227 12265 5241
rect 12299 5227 12315 5261
rect 12249 5217 12315 5227
rect 11856 5175 11910 5191
rect 10935 5143 11111 5165
rect 11763 5143 11793 5175
rect 10153 4956 10183 4982
rect 10249 4956 10279 4982
rect 10321 4956 10351 4982
rect 10535 4956 10565 4982
rect 10638 4956 10668 4982
rect 10935 5117 11329 5143
rect 11872 5066 11902 5175
rect 12093 5111 12123 5211
rect 11975 5081 12123 5111
rect 12165 5148 12219 5164
rect 12165 5114 12175 5148
rect 12209 5114 12219 5148
rect 12165 5098 12219 5114
rect 11975 5066 12005 5081
rect 12189 5066 12219 5098
rect 12261 5066 12291 5217
rect 12357 5164 12387 5309
rect 12591 5257 12801 5283
rect 12717 5251 12801 5257
rect 12717 5235 12859 5251
rect 12333 5148 12387 5164
rect 12533 5199 12675 5215
rect 12533 5165 12549 5199
rect 12583 5165 12675 5199
rect 12717 5201 12809 5235
rect 12843 5201 12859 5235
rect 12717 5185 12859 5201
rect 12533 5149 12675 5165
rect 12333 5114 12343 5148
rect 12377 5114 12387 5148
rect 12591 5143 12675 5149
rect 13005 5164 13035 5309
rect 13173 5271 13203 5309
rect 13269 5277 13299 5309
rect 13394 5277 13424 5309
rect 13077 5261 13203 5271
rect 13077 5227 13093 5261
rect 13127 5241 13203 5261
rect 13245 5261 13299 5277
rect 13127 5227 13143 5241
rect 13077 5217 13143 5227
rect 13245 5227 13255 5261
rect 13289 5227 13299 5261
rect 13005 5148 13059 5164
rect 12591 5117 12801 5143
rect 12333 5098 12387 5114
rect 12357 5066 12387 5098
rect 11872 4956 11902 4982
rect 11975 4956 12005 4982
rect 12189 4956 12219 4982
rect 12261 4956 12291 4982
rect 12357 4956 12387 4982
rect 13005 5114 13015 5148
rect 13049 5114 13059 5148
rect 13005 5098 13059 5114
rect 13005 5066 13035 5098
rect 13101 5066 13131 5217
rect 13245 5211 13299 5227
rect 13341 5261 13424 5277
rect 13341 5227 13351 5261
rect 13385 5227 13424 5261
rect 13490 5241 13520 5309
rect 13599 5241 13629 5263
rect 13787 5257 14733 5283
rect 14891 5257 15837 5283
rect 15995 5257 16389 5283
rect 16731 5257 17677 5283
rect 17835 5257 18413 5283
rect 13341 5211 13424 5227
rect 13482 5225 13536 5241
rect 13173 5148 13227 5164
rect 13173 5114 13183 5148
rect 13217 5114 13227 5148
rect 13173 5098 13227 5114
rect 13269 5111 13299 5211
rect 13482 5191 13492 5225
rect 13526 5191 13536 5225
rect 13482 5175 13536 5191
rect 13578 5225 13632 5241
rect 13578 5191 13588 5225
rect 13622 5191 13632 5225
rect 14279 5235 14733 5257
rect 13578 5175 13632 5191
rect 13787 5199 14237 5215
rect 13173 5066 13203 5098
rect 13269 5081 13417 5111
rect 13387 5066 13417 5081
rect 13490 5066 13520 5175
rect 13599 5143 13629 5175
rect 13787 5165 14059 5199
rect 14093 5165 14237 5199
rect 14279 5201 14423 5235
rect 14457 5201 14733 5235
rect 15383 5235 15837 5257
rect 14279 5185 14733 5201
rect 14891 5199 15341 5215
rect 13787 5143 14237 5165
rect 14891 5165 15163 5199
rect 15197 5165 15341 5199
rect 15383 5201 15527 5235
rect 15561 5201 15837 5235
rect 16213 5235 16389 5257
rect 15383 5185 15837 5201
rect 15995 5199 16171 5215
rect 14891 5143 15341 5165
rect 15995 5165 16011 5199
rect 16045 5165 16121 5199
rect 16155 5165 16171 5199
rect 16213 5201 16229 5235
rect 16263 5201 16339 5235
rect 16373 5201 16389 5235
rect 17223 5235 17677 5257
rect 16213 5185 16389 5201
rect 16731 5199 17181 5215
rect 15995 5143 16171 5165
rect 16731 5165 17003 5199
rect 17037 5165 17181 5199
rect 17223 5201 17367 5235
rect 17401 5201 17677 5235
rect 18141 5235 18413 5257
rect 18663 5257 18781 5283
rect 18663 5255 18701 5257
rect 17223 5185 17677 5201
rect 17835 5199 18099 5215
rect 16731 5143 17181 5165
rect 17835 5165 17851 5199
rect 17885 5165 17950 5199
rect 17984 5165 18049 5199
rect 18083 5165 18099 5199
rect 18141 5201 18157 5235
rect 18191 5201 18260 5235
rect 18294 5201 18363 5235
rect 18397 5201 18413 5235
rect 18141 5185 18413 5201
rect 18635 5239 18701 5255
rect 18635 5205 18651 5239
rect 18685 5205 18701 5239
rect 18635 5189 18701 5205
rect 18743 5199 18809 5215
rect 17835 5143 18099 5165
rect 18743 5165 18759 5199
rect 18793 5165 18809 5199
rect 18743 5149 18809 5165
rect 18743 5147 18781 5149
rect 13005 4956 13035 4982
rect 13101 4956 13131 4982
rect 13173 4956 13203 4982
rect 13387 4956 13417 4982
rect 13490 4956 13520 4982
rect 13787 5117 14733 5143
rect 14891 5117 15837 5143
rect 15995 5117 16389 5143
rect 16731 5117 17677 5143
rect 17835 5117 18413 5143
rect 18663 5117 18781 5147
rect 8250 4917 8280 4943
rect 8342 4917 8372 4943
rect 8441 4917 8471 4943
rect 8581 4917 8611 4943
rect 8678 4917 8708 4943
rect 8875 4917 8905 4943
rect 8974 4917 9004 4943
rect 9060 4917 9090 4943
rect 9144 4917 9174 4943
rect 9252 4917 9282 4943
rect 9336 4917 9366 4943
rect 9551 4917 9581 4943
rect 9739 4917 9949 4943
rect 10747 4917 10777 4943
rect 10935 4917 11329 4943
rect 11763 4917 11793 4943
rect 12591 4917 12801 4943
rect 13599 4917 13629 4943
rect 13787 4917 14733 4943
rect 14891 4917 15837 4943
rect 15995 4917 16389 4943
rect 16731 4917 17677 4943
rect 17835 4917 18413 4943
rect 18663 4917 18781 4943
rect 1183 4849 1301 4875
rect 1459 4849 2037 4875
rect 2195 4849 2313 4875
rect 2490 4849 2520 4875
rect 2585 4849 2685 4875
rect 2843 4849 2943 4875
rect 2997 4849 3027 4875
rect 3207 4849 3601 4875
rect 4044 4849 4074 4875
rect 4130 4849 4160 4875
rect 4216 4849 4246 4875
rect 4302 4849 4332 4875
rect 4398 4849 4428 4875
rect 4587 4849 4797 4875
rect 5139 4849 5717 4875
rect 6121 4849 6151 4875
rect 6519 4849 6729 4875
rect 7097 4849 7127 4875
rect 7347 4849 7741 4875
rect 7899 4849 7929 4875
rect 9397 4849 9427 4875
rect 9647 4849 9857 4875
rect 10199 4849 10409 4875
rect 10777 4849 10807 4875
rect 11027 4849 11237 4875
rect 11395 4849 11425 4875
rect 11483 4849 11513 4875
rect 11671 4849 11881 4875
rect 12679 4849 12709 4875
rect 12867 4849 13077 4875
rect 13235 4849 13265 4875
rect 13323 4849 13353 4875
rect 13511 4849 13905 4875
rect 14155 4849 15101 4875
rect 15469 4849 15499 4875
rect 15719 4849 15929 4875
rect 16087 4849 16117 4875
rect 16175 4849 16205 4875
rect 16363 4849 16573 4875
rect 16731 4849 16761 4875
rect 16819 4849 16849 4875
rect 17007 4849 17953 4875
rect 18111 4849 18505 4875
rect 18663 4849 18781 4875
rect 1183 4645 1301 4675
rect 1459 4649 2037 4675
rect 1183 4643 1221 4645
rect 1155 4627 1221 4643
rect 1155 4593 1171 4627
rect 1205 4593 1221 4627
rect 1459 4627 1723 4649
rect 2195 4645 2313 4675
rect 2195 4643 2233 4645
rect 1155 4577 1221 4593
rect 1263 4587 1329 4603
rect 1263 4553 1279 4587
rect 1313 4553 1329 4587
rect 1459 4593 1475 4627
rect 1509 4593 1574 4627
rect 1608 4593 1673 4627
rect 1707 4593 1723 4627
rect 2167 4627 2233 4643
rect 1459 4577 1723 4593
rect 1765 4591 2037 4607
rect 1263 4537 1329 4553
rect 1765 4557 1781 4591
rect 1815 4557 1884 4591
rect 1918 4557 1987 4591
rect 2021 4557 2037 4591
rect 2167 4593 2183 4627
rect 2217 4593 2233 4627
rect 2490 4617 2520 4649
rect 2585 4617 2685 4765
rect 2167 4577 2233 4593
rect 2275 4587 2341 4603
rect 1263 4535 1301 4537
rect 1765 4535 2037 4557
rect 2275 4553 2291 4587
rect 2325 4553 2341 4587
rect 2275 4537 2341 4553
rect 2489 4601 2543 4617
rect 2489 4567 2499 4601
rect 2533 4567 2543 4601
rect 2489 4551 2543 4567
rect 2585 4601 2739 4617
rect 2585 4567 2695 4601
rect 2729 4567 2739 4601
rect 2585 4551 2739 4567
rect 2843 4601 2943 4765
rect 2843 4567 2899 4601
rect 2933 4567 2943 4601
rect 2275 4535 2313 4537
rect 1183 4509 1301 4535
rect 1459 4509 2037 4535
rect 2195 4509 2313 4535
rect 2490 4529 2520 4551
rect 2585 4483 2685 4551
rect 2843 4483 2943 4567
rect 2997 4617 3027 4765
rect 3207 4649 3601 4675
rect 4587 4649 4797 4675
rect 5139 4649 5717 4675
rect 6218 4733 6248 4759
rect 6290 4733 6320 4759
rect 6928 4733 6958 4759
rect 7000 4733 7030 4759
rect 6519 4649 6729 4675
rect 7347 4649 7741 4675
rect 8008 4810 8038 4836
rect 8111 4810 8141 4836
rect 8325 4810 8355 4836
rect 8397 4810 8427 4836
rect 8493 4810 8523 4836
rect 3207 4627 3383 4649
rect 2997 4601 3057 4617
rect 2997 4567 3013 4601
rect 3047 4567 3057 4601
rect 3207 4593 3223 4627
rect 3257 4593 3333 4627
rect 3367 4593 3383 4627
rect 4044 4611 4074 4649
rect 4130 4611 4160 4649
rect 4216 4611 4246 4649
rect 4302 4611 4332 4649
rect 4398 4617 4428 4649
rect 4587 4643 4671 4649
rect 4529 4627 4671 4643
rect 3207 4577 3383 4593
rect 3425 4591 3601 4607
rect 2997 4551 3057 4567
rect 3425 4557 3441 4591
rect 3475 4557 3551 4591
rect 3585 4557 3601 4591
rect 4044 4601 4332 4611
rect 4044 4589 4107 4601
rect 2997 4483 3027 4551
rect 3425 4535 3601 4557
rect 3207 4509 3601 4535
rect 4043 4567 4107 4589
rect 4141 4567 4175 4601
rect 4209 4567 4243 4601
rect 4277 4567 4332 4601
rect 4043 4562 4332 4567
rect 4379 4601 4439 4617
rect 4379 4567 4389 4601
rect 4423 4567 4439 4601
rect 4529 4593 4545 4627
rect 4579 4593 4671 4627
rect 5139 4627 5403 4649
rect 4529 4577 4671 4593
rect 4713 4591 4855 4607
rect 4043 4556 4331 4562
rect 4043 4483 4073 4556
rect 4129 4483 4159 4556
rect 4215 4483 4245 4556
rect 4301 4483 4331 4556
rect 4379 4551 4439 4567
rect 4713 4557 4805 4591
rect 4839 4557 4855 4591
rect 5139 4593 5155 4627
rect 5189 4593 5254 4627
rect 5288 4593 5353 4627
rect 5387 4593 5403 4627
rect 6121 4617 6151 4649
rect 6218 4617 6248 4649
rect 5139 4577 5403 4593
rect 5445 4591 5717 4607
rect 4398 4483 4428 4551
rect 4713 4541 4855 4557
rect 5445 4557 5461 4591
rect 5495 4557 5564 4591
rect 5598 4557 5667 4591
rect 5701 4557 5717 4591
rect 4713 4535 4797 4541
rect 5445 4535 5717 4557
rect 6085 4601 6151 4617
rect 6085 4567 6101 4601
rect 6135 4567 6151 4601
rect 6085 4551 6151 4567
rect 6194 4601 6248 4617
rect 6194 4567 6204 4601
rect 6238 4567 6248 4601
rect 6194 4551 6248 4567
rect 6290 4617 6320 4649
rect 6519 4643 6603 4649
rect 6461 4627 6603 4643
rect 6290 4601 6390 4617
rect 6290 4567 6340 4601
rect 6374 4567 6390 4601
rect 6461 4593 6477 4627
rect 6511 4593 6603 4627
rect 6928 4617 6958 4649
rect 6461 4577 6603 4593
rect 6645 4591 6787 4607
rect 6290 4551 6390 4567
rect 6645 4557 6737 4591
rect 6771 4557 6787 4591
rect 4587 4509 4797 4535
rect 5139 4509 5717 4535
rect 6121 4529 6151 4551
rect 1183 4373 1301 4399
rect 1459 4373 2037 4399
rect 2195 4373 2313 4399
rect 2490 4373 2520 4399
rect 2585 4373 2685 4399
rect 2843 4373 2943 4399
rect 2997 4373 3027 4399
rect 3207 4373 3601 4399
rect 4043 4373 4073 4399
rect 4129 4373 4159 4399
rect 4215 4373 4245 4399
rect 4301 4373 4331 4399
rect 4398 4373 4428 4399
rect 4587 4373 4797 4399
rect 6218 4483 6248 4551
rect 6302 4483 6332 4551
rect 6645 4541 6787 4557
rect 6858 4601 6958 4617
rect 6858 4567 6874 4601
rect 6908 4567 6958 4601
rect 6858 4551 6958 4567
rect 7000 4617 7030 4649
rect 7097 4617 7127 4649
rect 7347 4627 7523 4649
rect 7000 4601 7054 4617
rect 7000 4567 7010 4601
rect 7044 4567 7054 4601
rect 7000 4551 7054 4567
rect 7097 4601 7163 4617
rect 7097 4567 7113 4601
rect 7147 4567 7163 4601
rect 7347 4593 7363 4627
rect 7397 4593 7473 4627
rect 7507 4593 7523 4627
rect 7899 4617 7929 4649
rect 8008 4617 8038 4726
rect 8111 4711 8141 4726
rect 8111 4681 8259 4711
rect 8325 4694 8355 4726
rect 7347 4577 7523 4593
rect 7565 4591 7741 4607
rect 7097 4551 7163 4567
rect 7565 4557 7581 4591
rect 7615 4557 7691 4591
rect 7725 4557 7741 4591
rect 6645 4535 6729 4541
rect 6519 4509 6729 4535
rect 6916 4483 6946 4551
rect 7000 4483 7030 4551
rect 7097 4529 7127 4551
rect 7565 4535 7741 4557
rect 7896 4601 7950 4617
rect 7896 4567 7906 4601
rect 7940 4567 7950 4601
rect 7896 4551 7950 4567
rect 7992 4601 8046 4617
rect 7992 4567 8002 4601
rect 8036 4567 8046 4601
rect 8229 4581 8259 4681
rect 8301 4678 8355 4694
rect 8301 4644 8311 4678
rect 8345 4644 8355 4678
rect 8301 4628 8355 4644
rect 7992 4551 8046 4567
rect 8104 4565 8187 4581
rect 7347 4509 7741 4535
rect 7899 4529 7929 4551
rect 8008 4483 8038 4551
rect 8104 4531 8143 4565
rect 8177 4531 8187 4565
rect 8104 4515 8187 4531
rect 8229 4565 8283 4581
rect 8397 4575 8427 4726
rect 8493 4694 8523 4726
rect 8469 4678 8523 4694
rect 8469 4644 8479 4678
rect 8513 4644 8523 4678
rect 9228 4733 9258 4759
rect 9300 4733 9330 4759
rect 10608 4733 10638 4759
rect 10680 4733 10710 4759
rect 9647 4649 9857 4675
rect 10199 4649 10409 4675
rect 11395 4676 11425 4691
rect 11027 4649 11237 4675
rect 11389 4652 11425 4676
rect 8469 4628 8523 4644
rect 8229 4531 8239 4565
rect 8273 4531 8283 4565
rect 8385 4565 8451 4575
rect 8385 4551 8401 4565
rect 8229 4515 8283 4531
rect 8325 4531 8401 4551
rect 8435 4531 8451 4565
rect 8325 4521 8451 4531
rect 8104 4483 8134 4515
rect 8229 4483 8259 4515
rect 8325 4483 8355 4521
rect 8493 4483 8523 4628
rect 9228 4617 9258 4649
rect 9158 4601 9258 4617
rect 9158 4567 9174 4601
rect 9208 4567 9258 4601
rect 9158 4551 9258 4567
rect 9300 4617 9330 4649
rect 9397 4617 9427 4649
rect 9647 4643 9731 4649
rect 10199 4643 10283 4649
rect 9589 4627 9731 4643
rect 9300 4601 9354 4617
rect 9300 4567 9310 4601
rect 9344 4567 9354 4601
rect 9300 4551 9354 4567
rect 9397 4601 9463 4617
rect 9397 4567 9413 4601
rect 9447 4567 9463 4601
rect 9589 4593 9605 4627
rect 9639 4593 9731 4627
rect 10141 4627 10283 4643
rect 9589 4577 9731 4593
rect 9773 4591 9915 4607
rect 9397 4551 9463 4567
rect 9773 4557 9865 4591
rect 9899 4557 9915 4591
rect 10141 4593 10157 4627
rect 10191 4593 10283 4627
rect 10608 4617 10638 4649
rect 10141 4577 10283 4593
rect 10325 4591 10467 4607
rect 9216 4483 9246 4551
rect 9300 4483 9330 4551
rect 9397 4529 9427 4551
rect 9773 4541 9915 4557
rect 10325 4557 10417 4591
rect 10451 4557 10467 4591
rect 10325 4541 10467 4557
rect 10538 4601 10638 4617
rect 10538 4567 10554 4601
rect 10588 4567 10638 4601
rect 10538 4551 10638 4567
rect 10680 4617 10710 4649
rect 10777 4617 10807 4649
rect 11027 4643 11111 4649
rect 10969 4627 11111 4643
rect 10680 4601 10734 4617
rect 10680 4567 10690 4601
rect 10724 4567 10734 4601
rect 10680 4551 10734 4567
rect 10777 4601 10843 4617
rect 10777 4567 10793 4601
rect 10827 4567 10843 4601
rect 10969 4593 10985 4627
rect 11019 4593 11111 4627
rect 11389 4617 11419 4652
rect 11483 4630 11513 4691
rect 12085 4810 12115 4836
rect 12181 4810 12211 4836
rect 12253 4810 12283 4836
rect 12467 4810 12497 4836
rect 12570 4810 12600 4836
rect 12085 4694 12115 4726
rect 12085 4678 12139 4694
rect 11671 4649 11881 4675
rect 11671 4643 11755 4649
rect 10969 4577 11111 4593
rect 11153 4591 11295 4607
rect 10777 4551 10843 4567
rect 11153 4557 11245 4591
rect 11279 4557 11295 4591
rect 9773 4535 9857 4541
rect 10325 4535 10409 4541
rect 9647 4509 9857 4535
rect 10199 4509 10409 4535
rect 5139 4373 5717 4399
rect 6121 4373 6151 4399
rect 6218 4373 6248 4399
rect 6302 4373 6332 4399
rect 6519 4373 6729 4399
rect 6916 4373 6946 4399
rect 7000 4373 7030 4399
rect 7097 4373 7127 4399
rect 7347 4373 7741 4399
rect 7899 4373 7929 4399
rect 8008 4373 8038 4399
rect 8104 4373 8134 4399
rect 8229 4373 8259 4399
rect 8325 4373 8355 4399
rect 8493 4373 8523 4399
rect 9216 4373 9246 4399
rect 9300 4373 9330 4399
rect 9397 4373 9427 4399
rect 9647 4373 9857 4399
rect 10596 4483 10626 4551
rect 10680 4483 10710 4551
rect 10777 4529 10807 4551
rect 11153 4541 11295 4557
rect 11343 4601 11419 4617
rect 11343 4567 11353 4601
rect 11387 4567 11419 4601
rect 11343 4551 11419 4567
rect 11463 4614 11517 4630
rect 11463 4580 11473 4614
rect 11507 4580 11517 4614
rect 11463 4564 11517 4580
rect 11613 4627 11755 4643
rect 11613 4593 11629 4627
rect 11663 4593 11755 4627
rect 12085 4644 12095 4678
rect 12129 4644 12139 4678
rect 12085 4628 12139 4644
rect 11613 4577 11755 4593
rect 11797 4591 11939 4607
rect 11389 4542 11419 4551
rect 11153 4535 11237 4541
rect 11027 4509 11237 4535
rect 11389 4518 11425 4542
rect 11395 4503 11425 4518
rect 11483 4503 11513 4564
rect 11797 4557 11889 4591
rect 11923 4557 11939 4591
rect 11797 4541 11939 4557
rect 11797 4535 11881 4541
rect 11671 4509 11881 4535
rect 12085 4483 12115 4628
rect 12181 4575 12211 4726
rect 12253 4694 12283 4726
rect 12467 4711 12497 4726
rect 12253 4678 12307 4694
rect 12253 4644 12263 4678
rect 12297 4644 12307 4678
rect 12253 4628 12307 4644
rect 12349 4681 12497 4711
rect 12349 4581 12379 4681
rect 12570 4617 12600 4726
rect 12867 4649 13077 4675
rect 12679 4617 12709 4649
rect 12867 4643 12951 4649
rect 12809 4627 12951 4643
rect 13235 4630 13265 4691
rect 13323 4676 13353 4691
rect 13323 4652 13359 4676
rect 12562 4601 12616 4617
rect 12157 4565 12223 4575
rect 12157 4531 12173 4565
rect 12207 4551 12223 4565
rect 12325 4565 12379 4581
rect 12207 4531 12283 4551
rect 12157 4521 12283 4531
rect 12253 4483 12283 4521
rect 12325 4531 12335 4565
rect 12369 4531 12379 4565
rect 12325 4515 12379 4531
rect 12421 4565 12504 4581
rect 12421 4531 12431 4565
rect 12465 4531 12504 4565
rect 12562 4567 12572 4601
rect 12606 4567 12616 4601
rect 12562 4551 12616 4567
rect 12658 4601 12712 4617
rect 12658 4567 12668 4601
rect 12702 4567 12712 4601
rect 12809 4593 12825 4627
rect 12859 4593 12951 4627
rect 13231 4614 13285 4630
rect 12809 4577 12951 4593
rect 12993 4591 13135 4607
rect 12658 4551 12712 4567
rect 12993 4557 13085 4591
rect 13119 4557 13135 4591
rect 13231 4580 13241 4614
rect 13275 4580 13285 4614
rect 13231 4564 13285 4580
rect 13329 4617 13359 4652
rect 13511 4649 13905 4675
rect 15300 4733 15330 4759
rect 15372 4733 15402 4759
rect 14155 4649 15101 4675
rect 15719 4649 15929 4675
rect 13511 4627 13687 4649
rect 13329 4601 13405 4617
rect 13329 4567 13361 4601
rect 13395 4567 13405 4601
rect 13511 4593 13527 4627
rect 13561 4593 13637 4627
rect 13671 4593 13687 4627
rect 14155 4627 14605 4649
rect 13511 4577 13687 4593
rect 13729 4591 13905 4607
rect 12421 4515 12504 4531
rect 12349 4483 12379 4515
rect 12474 4483 12504 4515
rect 12570 4483 12600 4551
rect 12679 4529 12709 4551
rect 12993 4541 13135 4557
rect 12993 4535 13077 4541
rect 12867 4509 13077 4535
rect 13235 4503 13265 4564
rect 13329 4551 13405 4567
rect 13729 4557 13745 4591
rect 13779 4557 13855 4591
rect 13889 4557 13905 4591
rect 14155 4593 14427 4627
rect 14461 4593 14605 4627
rect 15300 4617 15330 4649
rect 14155 4577 14605 4593
rect 14647 4591 15101 4607
rect 13329 4542 13359 4551
rect 13323 4518 13359 4542
rect 13729 4535 13905 4557
rect 14647 4557 14791 4591
rect 14825 4557 15101 4591
rect 14647 4535 15101 4557
rect 15230 4601 15330 4617
rect 15230 4567 15246 4601
rect 15280 4567 15330 4601
rect 15230 4551 15330 4567
rect 15372 4617 15402 4649
rect 15469 4617 15499 4649
rect 15719 4643 15803 4649
rect 15661 4627 15803 4643
rect 16087 4630 16117 4691
rect 16175 4676 16205 4691
rect 16175 4652 16211 4676
rect 15372 4601 15426 4617
rect 15372 4567 15382 4601
rect 15416 4567 15426 4601
rect 15372 4551 15426 4567
rect 15469 4601 15535 4617
rect 15469 4567 15485 4601
rect 15519 4567 15535 4601
rect 15661 4593 15677 4627
rect 15711 4593 15803 4627
rect 16083 4614 16137 4630
rect 15661 4577 15803 4593
rect 15845 4591 15987 4607
rect 15469 4551 15535 4567
rect 15845 4557 15937 4591
rect 15971 4557 15987 4591
rect 16083 4580 16093 4614
rect 16127 4580 16137 4614
rect 16083 4564 16137 4580
rect 16181 4617 16211 4652
rect 16363 4649 16573 4675
rect 16363 4643 16447 4649
rect 16305 4627 16447 4643
rect 16731 4630 16761 4691
rect 16819 4676 16849 4691
rect 16819 4652 16855 4676
rect 16181 4601 16257 4617
rect 16181 4567 16213 4601
rect 16247 4567 16257 4601
rect 16305 4593 16321 4627
rect 16355 4593 16447 4627
rect 16727 4614 16781 4630
rect 16305 4577 16447 4593
rect 16489 4591 16631 4607
rect 13323 4503 13353 4518
rect 13511 4509 13905 4535
rect 14155 4509 15101 4535
rect 15288 4483 15318 4551
rect 15372 4483 15402 4551
rect 15469 4529 15499 4551
rect 15845 4541 15987 4557
rect 15845 4535 15929 4541
rect 15719 4509 15929 4535
rect 16087 4503 16117 4564
rect 16181 4551 16257 4567
rect 16489 4557 16581 4591
rect 16615 4557 16631 4591
rect 16727 4580 16737 4614
rect 16771 4580 16781 4614
rect 16727 4564 16781 4580
rect 16825 4617 16855 4652
rect 17007 4649 17953 4675
rect 18111 4649 18505 4675
rect 17007 4627 17457 4649
rect 16825 4601 16901 4617
rect 16825 4567 16857 4601
rect 16891 4567 16901 4601
rect 17007 4593 17279 4627
rect 17313 4593 17457 4627
rect 18111 4627 18287 4649
rect 18663 4645 18781 4675
rect 17007 4577 17457 4593
rect 17499 4591 17953 4607
rect 16181 4542 16211 4551
rect 16175 4518 16211 4542
rect 16489 4541 16631 4557
rect 16489 4535 16573 4541
rect 16175 4503 16205 4518
rect 16363 4509 16573 4535
rect 16731 4503 16761 4564
rect 16825 4551 16901 4567
rect 17499 4557 17643 4591
rect 17677 4557 17953 4591
rect 18111 4593 18127 4627
rect 18161 4593 18237 4627
rect 18271 4593 18287 4627
rect 18743 4643 18781 4645
rect 18743 4627 18809 4643
rect 18111 4577 18287 4593
rect 18329 4591 18505 4607
rect 16825 4542 16855 4551
rect 16819 4518 16855 4542
rect 17499 4535 17953 4557
rect 18329 4557 18345 4591
rect 18379 4557 18455 4591
rect 18489 4557 18505 4591
rect 18329 4535 18505 4557
rect 18635 4587 18701 4603
rect 18635 4553 18651 4587
rect 18685 4553 18701 4587
rect 18743 4593 18759 4627
rect 18793 4593 18809 4627
rect 18743 4577 18809 4593
rect 18635 4537 18701 4553
rect 16819 4503 16849 4518
rect 17007 4509 17953 4535
rect 18111 4509 18505 4535
rect 18663 4535 18701 4537
rect 18663 4509 18781 4535
rect 10199 4373 10409 4399
rect 10596 4373 10626 4399
rect 10680 4373 10710 4399
rect 10777 4373 10807 4399
rect 11027 4373 11237 4399
rect 11395 4373 11425 4399
rect 11483 4373 11513 4399
rect 11671 4373 11881 4399
rect 12085 4373 12115 4399
rect 12253 4373 12283 4399
rect 12349 4373 12379 4399
rect 12474 4373 12504 4399
rect 12570 4373 12600 4399
rect 12679 4373 12709 4399
rect 12867 4373 13077 4399
rect 13235 4373 13265 4399
rect 13323 4373 13353 4399
rect 13511 4373 13905 4399
rect 14155 4373 15101 4399
rect 15288 4373 15318 4399
rect 15372 4373 15402 4399
rect 15469 4373 15499 4399
rect 15719 4373 15929 4399
rect 16087 4373 16117 4399
rect 16175 4373 16205 4399
rect 16363 4373 16573 4399
rect 16731 4373 16761 4399
rect 16819 4373 16849 4399
rect 17007 4373 17953 4399
rect 18111 4373 18505 4399
rect 18663 4373 18781 4399
rect 1183 4305 1301 4331
rect 1459 4305 2037 4331
rect 2287 4305 2317 4331
rect 2375 4305 2405 4331
rect 2563 4305 2773 4331
rect 2931 4305 2961 4331
rect 3015 4305 3045 4331
rect 3270 4305 3300 4331
rect 3365 4305 3395 4331
rect 3461 4305 3491 4331
rect 3627 4305 3657 4331
rect 3699 4305 3729 4331
rect 3831 4305 3861 4331
rect 3930 4305 3960 4331
rect 4039 4305 4069 4331
rect 4135 4305 4165 4331
rect 4284 4305 4314 4331
rect 4375 4305 4405 4331
rect 4583 4305 4613 4331
rect 4771 4305 4981 4331
rect 5081 4305 5177 4331
rect 1183 4169 1301 4195
rect 1459 4169 2037 4195
rect 2287 4186 2317 4201
rect 1263 4167 1301 4169
rect 1263 4151 1329 4167
rect 1155 4111 1221 4127
rect 1155 4077 1171 4111
rect 1205 4077 1221 4111
rect 1263 4117 1279 4151
rect 1313 4117 1329 4151
rect 1765 4147 2037 4169
rect 2281 4162 2317 4186
rect 2281 4153 2311 4162
rect 1263 4101 1329 4117
rect 1459 4111 1723 4127
rect 1155 4061 1221 4077
rect 1183 4059 1221 4061
rect 1459 4077 1475 4111
rect 1509 4077 1574 4111
rect 1608 4077 1673 4111
rect 1707 4077 1723 4111
rect 1765 4113 1781 4147
rect 1815 4113 1884 4147
rect 1918 4113 1987 4147
rect 2021 4113 2037 4147
rect 1765 4097 2037 4113
rect 2235 4137 2311 4153
rect 2375 4140 2405 4201
rect 2931 4206 2961 4221
rect 2563 4169 2773 4195
rect 2689 4163 2773 4169
rect 2898 4176 2961 4206
rect 2689 4147 2831 4163
rect 2898 4153 2928 4176
rect 2235 4103 2245 4137
rect 2279 4103 2311 4137
rect 2235 4087 2311 4103
rect 1183 4029 1301 4059
rect 1459 4055 1723 4077
rect 1459 4029 2037 4055
rect 2281 4052 2311 4087
rect 2355 4124 2409 4140
rect 2355 4090 2365 4124
rect 2399 4090 2409 4124
rect 2355 4074 2409 4090
rect 2505 4111 2647 4127
rect 2505 4077 2521 4111
rect 2555 4077 2647 4111
rect 2689 4113 2781 4147
rect 2815 4113 2831 4147
rect 2689 4097 2831 4113
rect 2874 4137 2928 4153
rect 2874 4103 2884 4137
rect 2918 4103 2928 4137
rect 3015 4132 3045 4221
rect 2874 4087 2928 4103
rect 2281 4028 2317 4052
rect 2287 4013 2317 4028
rect 2375 4013 2405 4074
rect 2505 4061 2647 4077
rect 2563 4055 2647 4061
rect 2563 4029 2773 4055
rect 2898 4034 2928 4087
rect 2970 4122 3045 4132
rect 2970 4088 2986 4122
rect 3020 4088 3045 4122
rect 3270 4092 3300 4221
rect 3365 4199 3395 4233
rect 3461 4199 3491 4233
rect 3342 4183 3396 4199
rect 3342 4149 3352 4183
rect 3386 4149 3396 4183
rect 3342 4133 3396 4149
rect 3438 4189 3504 4199
rect 3438 4155 3454 4189
rect 3488 4155 3504 4189
rect 3438 4145 3504 4155
rect 2970 4078 3045 4088
rect 2898 4004 2961 4034
rect 2931 3989 2961 4004
rect 3015 3989 3045 4078
rect 3183 4076 3300 4092
rect 3183 4042 3193 4076
rect 3227 4056 3300 4076
rect 3365 4103 3396 4133
rect 3365 4073 3503 4103
rect 3227 4042 3312 4056
rect 3183 4026 3312 4042
rect 3282 3939 3312 4026
rect 3358 4021 3424 4031
rect 3358 3987 3374 4021
rect 3408 3987 3424 4021
rect 3358 3977 3424 3987
rect 3374 3939 3404 3977
rect 3473 3939 3503 4073
rect 3627 4063 3657 4221
rect 3699 4199 3729 4221
rect 3699 4183 3753 4199
rect 3699 4149 3709 4183
rect 3743 4149 3753 4183
rect 3930 4211 3960 4233
rect 3930 4195 3997 4211
rect 3831 4151 3861 4177
rect 3699 4133 3753 4149
rect 3795 4135 3861 4151
rect 3930 4161 3953 4195
rect 3987 4161 3997 4195
rect 3930 4145 3997 4161
rect 4039 4163 4069 4233
rect 4135 4189 4165 4221
rect 4135 4173 4237 4189
rect 4039 4147 4093 4163
rect 4135 4159 4193 4173
rect 3613 4047 3668 4063
rect 3613 4013 3623 4047
rect 3657 4013 3668 4047
rect 3613 3997 3668 4013
rect 3613 3939 3643 3997
rect 3710 3939 3740 4133
rect 3795 4101 3805 4135
rect 3839 4101 3861 4135
rect 4039 4115 4049 4147
rect 4027 4113 4049 4115
rect 4083 4113 4093 4147
rect 4027 4103 4093 4113
rect 3795 4085 3861 4101
rect 3831 4068 3861 4085
rect 4006 4097 4093 4103
rect 4176 4139 4193 4159
rect 4227 4139 4237 4173
rect 4284 4161 4314 4221
rect 4176 4123 4237 4139
rect 4279 4145 4333 4161
rect 4006 4085 4069 4097
rect 4006 4073 4056 4085
rect 3831 4038 3937 4068
rect 3907 4023 3937 4038
rect 1183 3829 1301 3855
rect 1459 3829 2037 3855
rect 2287 3829 2317 3855
rect 2375 3829 2405 3855
rect 2563 3829 2773 3855
rect 2931 3835 2961 3861
rect 3015 3835 3045 3861
rect 4006 3939 4036 4073
rect 4078 4021 4132 4037
rect 4078 3987 4088 4021
rect 4122 3987 4132 4021
rect 4078 3971 4132 3987
rect 4092 3939 4122 3971
rect 4176 3939 4206 4123
rect 4279 4111 4289 4145
rect 4323 4111 4333 4145
rect 4279 4095 4333 4111
rect 4284 3939 4314 4095
rect 4375 4053 4405 4221
rect 5081 4271 5131 4305
rect 5165 4271 5177 4305
rect 5081 4237 5177 4271
rect 5081 4203 5131 4237
rect 5165 4203 5177 4237
rect 4583 4153 4613 4175
rect 4771 4169 4981 4195
rect 4554 4137 4613 4153
rect 4554 4103 4564 4137
rect 4598 4103 4613 4137
rect 4897 4163 4981 4169
rect 4897 4147 5039 4163
rect 4554 4087 4613 4103
rect 4583 4055 4613 4087
rect 4713 4111 4855 4127
rect 4713 4077 4729 4111
rect 4763 4077 4855 4111
rect 4897 4113 4989 4147
rect 5023 4113 5039 4147
rect 4897 4097 5039 4113
rect 5081 4120 5177 4203
rect 4713 4061 4855 4077
rect 4771 4055 4855 4061
rect 4356 4037 4410 4053
rect 4356 4003 4366 4037
rect 4400 4003 4410 4037
rect 4356 3987 4410 4003
rect 4368 3939 4398 3987
rect 4771 4029 4981 4055
rect 5081 3970 5177 4111
rect 5081 3936 5131 3970
rect 5165 3936 5177 3970
rect 5081 3902 5177 3936
rect 5081 3868 5131 3902
rect 5165 3868 5177 3902
rect 3282 3829 3312 3855
rect 3374 3829 3404 3855
rect 3473 3829 3503 3855
rect 3613 3829 3643 3855
rect 3710 3829 3740 3855
rect 3907 3829 3937 3855
rect 4006 3829 4036 3855
rect 4092 3829 4122 3855
rect 4176 3829 4206 3855
rect 4284 3829 4314 3855
rect 4368 3829 4398 3855
rect 4583 3829 4613 3855
rect 4771 3829 4981 3855
rect 5081 3829 5177 3868
rect 5219 4301 5315 4331
rect 5415 4305 5993 4331
rect 6427 4305 6545 4331
rect 6703 4305 6733 4331
rect 6791 4305 6821 4331
rect 6979 4305 7557 4331
rect 7761 4305 7791 4331
rect 7929 4305 7959 4331
rect 8025 4305 8055 4331
rect 8150 4305 8180 4331
rect 8246 4305 8276 4331
rect 8355 4305 8385 4331
rect 8543 4305 8753 4331
rect 9004 4305 9034 4331
rect 9090 4305 9120 4331
rect 9176 4305 9206 4331
rect 9262 4305 9292 4331
rect 9348 4305 9378 4331
rect 9434 4305 9464 4331
rect 9520 4305 9550 4331
rect 9606 4305 9636 4331
rect 9692 4305 9722 4331
rect 9778 4305 9808 4331
rect 9864 4305 9894 4331
rect 9950 4305 9980 4331
rect 10035 4305 10065 4331
rect 10121 4305 10151 4331
rect 10207 4305 10237 4331
rect 10293 4305 10323 4331
rect 10379 4305 10409 4331
rect 10465 4305 10495 4331
rect 10551 4305 10581 4331
rect 10637 4305 10667 4331
rect 10843 4305 11237 4331
rect 11763 4305 11793 4331
rect 11971 4305 12001 4331
rect 12062 4305 12092 4331
rect 12211 4305 12241 4331
rect 12307 4305 12337 4331
rect 12416 4305 12446 4331
rect 12515 4305 12545 4331
rect 12647 4305 12677 4331
rect 12719 4305 12749 4331
rect 12885 4305 12915 4331
rect 12981 4305 13011 4331
rect 13076 4305 13106 4331
rect 13331 4305 13361 4331
rect 13415 4305 13445 4331
rect 13603 4305 13813 4331
rect 13971 4305 14001 4331
rect 14055 4305 14085 4331
rect 14310 4305 14340 4331
rect 14405 4305 14435 4331
rect 14501 4305 14531 4331
rect 14667 4305 14697 4331
rect 14739 4305 14769 4331
rect 14871 4305 14901 4331
rect 14970 4305 15000 4331
rect 15079 4305 15109 4331
rect 15175 4305 15205 4331
rect 15324 4305 15354 4331
rect 15415 4305 15445 4331
rect 15623 4305 15653 4331
rect 15811 4305 16389 4331
rect 16731 4305 17677 4331
rect 17835 4305 18413 4331
rect 18663 4305 18781 4331
rect 5219 4267 5231 4301
rect 5265 4267 5315 4301
rect 5219 4233 5315 4267
rect 5219 4199 5231 4233
rect 5265 4199 5315 4233
rect 5219 4120 5315 4199
rect 5415 4169 5993 4195
rect 6427 4169 6545 4195
rect 5721 4147 5993 4169
rect 5219 3970 5315 4111
rect 5415 4111 5679 4127
rect 5415 4077 5431 4111
rect 5465 4077 5530 4111
rect 5564 4077 5629 4111
rect 5663 4077 5679 4111
rect 5721 4113 5737 4147
rect 5771 4113 5840 4147
rect 5874 4113 5943 4147
rect 5977 4113 5993 4147
rect 6507 4167 6545 4169
rect 6507 4151 6573 4167
rect 5721 4097 5993 4113
rect 6399 4111 6465 4127
rect 5415 4055 5679 4077
rect 6399 4077 6415 4111
rect 6449 4077 6465 4111
rect 6507 4117 6523 4151
rect 6557 4117 6573 4151
rect 6703 4140 6733 4201
rect 6791 4186 6821 4201
rect 6791 4162 6827 4186
rect 6979 4169 7557 4195
rect 6797 4153 6827 4162
rect 6507 4101 6573 4117
rect 6699 4124 6753 4140
rect 6399 4061 6465 4077
rect 6699 4090 6709 4124
rect 6743 4090 6753 4124
rect 6699 4074 6753 4090
rect 6797 4137 6873 4153
rect 6797 4103 6829 4137
rect 6863 4103 6873 4137
rect 7285 4147 7557 4169
rect 6797 4087 6873 4103
rect 6979 4111 7243 4127
rect 6427 4059 6465 4061
rect 5415 4029 5993 4055
rect 5219 3936 5231 3970
rect 5265 3936 5315 3970
rect 5219 3902 5315 3936
rect 5219 3868 5231 3902
rect 5265 3868 5315 3902
rect 5219 3829 5315 3868
rect 6427 4029 6545 4059
rect 6703 4013 6733 4074
rect 6797 4052 6827 4087
rect 6791 4028 6827 4052
rect 6979 4077 6995 4111
rect 7029 4077 7094 4111
rect 7128 4077 7193 4111
rect 7227 4077 7243 4111
rect 7285 4113 7301 4147
rect 7335 4113 7404 4147
rect 7438 4113 7507 4147
rect 7541 4113 7557 4147
rect 7285 4097 7557 4113
rect 6979 4055 7243 4077
rect 7761 4076 7791 4221
rect 7929 4183 7959 4221
rect 8025 4189 8055 4221
rect 8150 4189 8180 4221
rect 7833 4173 7959 4183
rect 7833 4139 7849 4173
rect 7883 4153 7959 4173
rect 8001 4173 8055 4189
rect 7883 4139 7899 4153
rect 7833 4129 7899 4139
rect 8001 4139 8011 4173
rect 8045 4139 8055 4173
rect 7761 4060 7815 4076
rect 6979 4029 7557 4055
rect 6791 4013 6821 4028
rect 7761 4026 7771 4060
rect 7805 4026 7815 4060
rect 7761 4010 7815 4026
rect 7761 3978 7791 4010
rect 7857 3978 7887 4129
rect 8001 4123 8055 4139
rect 8097 4173 8180 4189
rect 8097 4139 8107 4173
rect 8141 4139 8180 4173
rect 8246 4153 8276 4221
rect 8355 4153 8385 4175
rect 8543 4169 8753 4195
rect 9004 4172 9034 4221
rect 9090 4172 9120 4221
rect 9176 4172 9206 4221
rect 9262 4172 9292 4221
rect 8669 4163 8753 4169
rect 8097 4123 8180 4139
rect 8238 4137 8292 4153
rect 7929 4060 7983 4076
rect 7929 4026 7939 4060
rect 7973 4026 7983 4060
rect 7929 4010 7983 4026
rect 8025 4023 8055 4123
rect 8238 4103 8248 4137
rect 8282 4103 8292 4137
rect 8238 4087 8292 4103
rect 8334 4137 8388 4153
rect 8334 4103 8344 4137
rect 8378 4103 8388 4137
rect 8669 4147 8811 4163
rect 8334 4087 8388 4103
rect 8485 4111 8627 4127
rect 7929 3978 7959 4010
rect 8025 3993 8173 4023
rect 8143 3978 8173 3993
rect 8246 3978 8276 4087
rect 8355 4055 8385 4087
rect 8485 4077 8501 4111
rect 8535 4077 8627 4111
rect 8669 4113 8761 4147
rect 8795 4113 8811 4147
rect 8669 4097 8811 4113
rect 8945 4137 9292 4172
rect 8945 4103 8961 4137
rect 8995 4103 9292 4137
rect 8485 4061 8627 4077
rect 8945 4070 9292 4103
rect 8543 4055 8627 4061
rect 9004 4055 9034 4070
rect 9090 4055 9120 4070
rect 9176 4055 9206 4070
rect 9262 4055 9292 4070
rect 9348 4162 9378 4221
rect 9434 4162 9464 4221
rect 9520 4162 9550 4221
rect 9606 4162 9636 4221
rect 9692 4162 9722 4221
rect 9778 4162 9808 4221
rect 9864 4162 9894 4221
rect 9950 4162 9980 4221
rect 10035 4162 10065 4221
rect 10121 4162 10151 4221
rect 10207 4162 10237 4221
rect 10293 4162 10323 4221
rect 10379 4162 10409 4221
rect 10465 4162 10495 4221
rect 10551 4162 10581 4221
rect 10637 4162 10667 4221
rect 10843 4169 11237 4195
rect 9348 4137 10667 4162
rect 9348 4103 9388 4137
rect 9422 4103 9456 4137
rect 9490 4103 9524 4137
rect 9558 4103 9592 4137
rect 9626 4103 9660 4137
rect 9694 4103 9728 4137
rect 9762 4103 9796 4137
rect 9830 4103 9864 4137
rect 9898 4103 9932 4137
rect 9966 4103 10000 4137
rect 10034 4103 10068 4137
rect 10102 4103 10136 4137
rect 10170 4103 10204 4137
rect 10238 4103 10272 4137
rect 10306 4103 10340 4137
rect 10374 4103 10408 4137
rect 10442 4103 10667 4137
rect 11061 4147 11237 4169
rect 9348 4087 10667 4103
rect 9348 4055 9378 4087
rect 9434 4055 9464 4087
rect 9520 4055 9550 4087
rect 9606 4055 9636 4087
rect 9692 4055 9722 4087
rect 9778 4055 9808 4087
rect 9864 4055 9894 4087
rect 9950 4055 9980 4087
rect 10035 4055 10065 4087
rect 10121 4055 10151 4087
rect 10207 4055 10237 4087
rect 10293 4055 10323 4087
rect 10379 4055 10409 4087
rect 10465 4055 10495 4087
rect 10551 4055 10581 4087
rect 10637 4055 10667 4087
rect 10843 4111 11019 4127
rect 10843 4077 10859 4111
rect 10893 4077 10969 4111
rect 11003 4077 11019 4111
rect 11061 4113 11077 4147
rect 11111 4113 11187 4147
rect 11221 4113 11237 4147
rect 11061 4097 11237 4113
rect 11763 4153 11793 4175
rect 11763 4137 11822 4153
rect 11763 4103 11778 4137
rect 11812 4103 11822 4137
rect 10843 4055 11019 4077
rect 11763 4087 11822 4103
rect 11763 4055 11793 4087
rect 7761 3868 7791 3894
rect 7857 3868 7887 3894
rect 7929 3868 7959 3894
rect 8143 3868 8173 3894
rect 8246 3868 8276 3894
rect 8543 4029 8753 4055
rect 10843 4029 11237 4055
rect 11971 4053 12001 4221
rect 12062 4161 12092 4221
rect 12211 4189 12241 4221
rect 12139 4173 12241 4189
rect 12043 4145 12097 4161
rect 12043 4111 12053 4145
rect 12087 4111 12097 4145
rect 12139 4139 12149 4173
rect 12183 4159 12241 4173
rect 12307 4163 12337 4233
rect 12416 4211 12446 4233
rect 12183 4139 12200 4159
rect 12139 4123 12200 4139
rect 12043 4095 12097 4111
rect 11966 4037 12020 4053
rect 11966 4003 11976 4037
rect 12010 4003 12020 4037
rect 11966 3987 12020 4003
rect 11978 3939 12008 3987
rect 12062 3939 12092 4095
rect 12170 3939 12200 4123
rect 12283 4147 12337 4163
rect 12283 4113 12293 4147
rect 12327 4115 12337 4147
rect 12379 4195 12446 4211
rect 12379 4161 12389 4195
rect 12423 4161 12446 4195
rect 12647 4199 12677 4221
rect 12623 4183 12677 4199
rect 12379 4145 12446 4161
rect 12515 4151 12545 4177
rect 12515 4135 12581 4151
rect 12327 4113 12349 4115
rect 12283 4103 12349 4113
rect 12283 4097 12370 4103
rect 12307 4085 12370 4097
rect 12320 4073 12370 4085
rect 12244 4021 12298 4037
rect 12244 3987 12254 4021
rect 12288 3987 12298 4021
rect 12244 3971 12298 3987
rect 12254 3939 12284 3971
rect 12340 3939 12370 4073
rect 12515 4101 12537 4135
rect 12571 4101 12581 4135
rect 12623 4149 12633 4183
rect 12667 4149 12677 4183
rect 12623 4133 12677 4149
rect 12515 4085 12581 4101
rect 12515 4068 12545 4085
rect 12439 4038 12545 4068
rect 12439 4023 12469 4038
rect 12636 3939 12666 4133
rect 12719 4063 12749 4221
rect 12885 4199 12915 4233
rect 12981 4199 13011 4233
rect 12872 4189 12938 4199
rect 12872 4155 12888 4189
rect 12922 4155 12938 4189
rect 12872 4145 12938 4155
rect 12980 4183 13034 4199
rect 12980 4149 12990 4183
rect 13024 4149 13034 4183
rect 12980 4133 13034 4149
rect 12980 4103 13011 4133
rect 12873 4073 13011 4103
rect 13076 4092 13106 4221
rect 13331 4132 13361 4221
rect 13415 4206 13445 4221
rect 13415 4176 13478 4206
rect 13971 4206 14001 4221
rect 13448 4153 13478 4176
rect 13603 4169 13813 4195
rect 13729 4163 13813 4169
rect 13938 4176 14001 4206
rect 13448 4137 13502 4153
rect 13331 4122 13406 4132
rect 13076 4076 13193 4092
rect 12708 4047 12763 4063
rect 12708 4013 12719 4047
rect 12753 4013 12763 4047
rect 12708 3997 12763 4013
rect 12733 3939 12763 3997
rect 12873 3939 12903 4073
rect 13076 4056 13149 4076
rect 13064 4042 13149 4056
rect 13183 4042 13193 4076
rect 12952 4021 13018 4031
rect 12952 3987 12968 4021
rect 13002 3987 13018 4021
rect 12952 3977 13018 3987
rect 13064 4026 13193 4042
rect 13331 4088 13356 4122
rect 13390 4088 13406 4122
rect 13331 4078 13406 4088
rect 13448 4103 13458 4137
rect 13492 4103 13502 4137
rect 13729 4147 13871 4163
rect 13938 4153 13968 4176
rect 13448 4087 13502 4103
rect 13545 4111 13687 4127
rect 12972 3939 13002 3977
rect 13064 3939 13094 4026
rect 13331 3989 13361 4078
rect 13448 4034 13478 4087
rect 13545 4077 13561 4111
rect 13595 4077 13687 4111
rect 13729 4113 13821 4147
rect 13855 4113 13871 4147
rect 13729 4097 13871 4113
rect 13914 4137 13968 4153
rect 13914 4103 13924 4137
rect 13958 4103 13968 4137
rect 14055 4132 14085 4221
rect 13914 4087 13968 4103
rect 13545 4061 13687 4077
rect 13415 4004 13478 4034
rect 13603 4055 13687 4061
rect 13603 4029 13813 4055
rect 13938 4034 13968 4087
rect 14010 4122 14085 4132
rect 14010 4088 14026 4122
rect 14060 4088 14085 4122
rect 14310 4092 14340 4221
rect 14405 4199 14435 4233
rect 14501 4199 14531 4233
rect 14382 4183 14436 4199
rect 14382 4149 14392 4183
rect 14426 4149 14436 4183
rect 14382 4133 14436 4149
rect 14478 4189 14544 4199
rect 14478 4155 14494 4189
rect 14528 4155 14544 4189
rect 14478 4145 14544 4155
rect 14010 4078 14085 4088
rect 13415 3989 13445 4004
rect 5415 3829 5993 3855
rect 6427 3829 6545 3855
rect 6703 3829 6733 3855
rect 6791 3829 6821 3855
rect 6979 3829 7557 3855
rect 8355 3829 8385 3855
rect 8543 3829 8753 3855
rect 9004 3829 9034 3855
rect 9090 3829 9120 3855
rect 9176 3829 9206 3855
rect 9262 3829 9292 3855
rect 9348 3829 9378 3855
rect 9434 3829 9464 3855
rect 9520 3829 9550 3855
rect 9606 3829 9636 3855
rect 9692 3829 9722 3855
rect 9778 3829 9808 3855
rect 9864 3829 9894 3855
rect 9950 3829 9980 3855
rect 10035 3829 10065 3855
rect 10121 3829 10151 3855
rect 10207 3829 10237 3855
rect 10293 3829 10323 3855
rect 10379 3829 10409 3855
rect 10465 3829 10495 3855
rect 10551 3829 10581 3855
rect 10637 3829 10667 3855
rect 10843 3829 11237 3855
rect 11763 3829 11793 3855
rect 11978 3829 12008 3855
rect 12062 3829 12092 3855
rect 12170 3829 12200 3855
rect 12254 3829 12284 3855
rect 12340 3829 12370 3855
rect 12439 3829 12469 3855
rect 12636 3829 12666 3855
rect 12733 3829 12763 3855
rect 12873 3829 12903 3855
rect 12972 3829 13002 3855
rect 13064 3829 13094 3855
rect 13331 3835 13361 3861
rect 13415 3835 13445 3861
rect 13938 4004 14001 4034
rect 13971 3989 14001 4004
rect 14055 3989 14085 4078
rect 14223 4076 14340 4092
rect 14223 4042 14233 4076
rect 14267 4056 14340 4076
rect 14405 4103 14436 4133
rect 14405 4073 14543 4103
rect 14267 4042 14352 4056
rect 14223 4026 14352 4042
rect 14322 3939 14352 4026
rect 14398 4021 14464 4031
rect 14398 3987 14414 4021
rect 14448 3987 14464 4021
rect 14398 3977 14464 3987
rect 14414 3939 14444 3977
rect 14513 3939 14543 4073
rect 14667 4063 14697 4221
rect 14739 4199 14769 4221
rect 14739 4183 14793 4199
rect 14739 4149 14749 4183
rect 14783 4149 14793 4183
rect 14970 4211 15000 4233
rect 14970 4195 15037 4211
rect 14871 4151 14901 4177
rect 14739 4133 14793 4149
rect 14835 4135 14901 4151
rect 14970 4161 14993 4195
rect 15027 4161 15037 4195
rect 14970 4145 15037 4161
rect 15079 4163 15109 4233
rect 15175 4189 15205 4221
rect 15175 4173 15277 4189
rect 15079 4147 15133 4163
rect 15175 4159 15233 4173
rect 14653 4047 14708 4063
rect 14653 4013 14663 4047
rect 14697 4013 14708 4047
rect 14653 3997 14708 4013
rect 14653 3939 14683 3997
rect 14750 3939 14780 4133
rect 14835 4101 14845 4135
rect 14879 4101 14901 4135
rect 15079 4115 15089 4147
rect 15067 4113 15089 4115
rect 15123 4113 15133 4147
rect 15067 4103 15133 4113
rect 14835 4085 14901 4101
rect 14871 4068 14901 4085
rect 15046 4097 15133 4103
rect 15216 4139 15233 4159
rect 15267 4139 15277 4173
rect 15324 4161 15354 4221
rect 15216 4123 15277 4139
rect 15319 4145 15373 4161
rect 15046 4085 15109 4097
rect 15046 4073 15096 4085
rect 14871 4038 14977 4068
rect 14947 4023 14977 4038
rect 13603 3829 13813 3855
rect 13971 3835 14001 3861
rect 14055 3835 14085 3861
rect 15046 3939 15076 4073
rect 15118 4021 15172 4037
rect 15118 3987 15128 4021
rect 15162 3987 15172 4021
rect 15118 3971 15172 3987
rect 15132 3939 15162 3971
rect 15216 3939 15246 4123
rect 15319 4111 15329 4145
rect 15363 4111 15373 4145
rect 15319 4095 15373 4111
rect 15324 3939 15354 4095
rect 15415 4053 15445 4221
rect 15623 4153 15653 4175
rect 15811 4169 16389 4195
rect 16731 4169 17677 4195
rect 17835 4169 18413 4195
rect 15594 4137 15653 4153
rect 15594 4103 15604 4137
rect 15638 4103 15653 4137
rect 16117 4147 16389 4169
rect 15594 4087 15653 4103
rect 15623 4055 15653 4087
rect 15811 4111 16075 4127
rect 15811 4077 15827 4111
rect 15861 4077 15926 4111
rect 15960 4077 16025 4111
rect 16059 4077 16075 4111
rect 16117 4113 16133 4147
rect 16167 4113 16236 4147
rect 16270 4113 16339 4147
rect 16373 4113 16389 4147
rect 17223 4147 17677 4169
rect 16117 4097 16389 4113
rect 16731 4111 17181 4127
rect 15811 4055 16075 4077
rect 16731 4077 17003 4111
rect 17037 4077 17181 4111
rect 17223 4113 17367 4147
rect 17401 4113 17677 4147
rect 18141 4147 18413 4169
rect 18663 4169 18781 4195
rect 18663 4167 18701 4169
rect 17223 4097 17677 4113
rect 17835 4111 18099 4127
rect 16731 4055 17181 4077
rect 17835 4077 17851 4111
rect 17885 4077 17950 4111
rect 17984 4077 18049 4111
rect 18083 4077 18099 4111
rect 18141 4113 18157 4147
rect 18191 4113 18260 4147
rect 18294 4113 18363 4147
rect 18397 4113 18413 4147
rect 18141 4097 18413 4113
rect 18635 4151 18701 4167
rect 18635 4117 18651 4151
rect 18685 4117 18701 4151
rect 18635 4101 18701 4117
rect 18743 4111 18809 4127
rect 17835 4055 18099 4077
rect 18743 4077 18759 4111
rect 18793 4077 18809 4111
rect 18743 4061 18809 4077
rect 18743 4059 18781 4061
rect 15396 4037 15450 4053
rect 15396 4003 15406 4037
rect 15440 4003 15450 4037
rect 15396 3987 15450 4003
rect 15408 3939 15438 3987
rect 15811 4029 16389 4055
rect 16731 4029 17677 4055
rect 17835 4029 18413 4055
rect 18663 4029 18781 4059
rect 14322 3829 14352 3855
rect 14414 3829 14444 3855
rect 14513 3829 14543 3855
rect 14653 3829 14683 3855
rect 14750 3829 14780 3855
rect 14947 3829 14977 3855
rect 15046 3829 15076 3855
rect 15132 3829 15162 3855
rect 15216 3829 15246 3855
rect 15324 3829 15354 3855
rect 15408 3829 15438 3855
rect 15623 3829 15653 3855
rect 15811 3829 16389 3855
rect 16731 3829 17677 3855
rect 17835 3829 18413 3855
rect 18663 3829 18781 3855
rect 1183 3761 1301 3787
rect 1459 3761 1577 3787
rect 1735 3755 1765 3781
rect 1819 3755 1849 3781
rect 2086 3761 2116 3787
rect 2178 3761 2208 3787
rect 2277 3761 2307 3787
rect 2417 3761 2447 3787
rect 2514 3761 2544 3787
rect 2711 3761 2741 3787
rect 2810 3761 2840 3787
rect 2896 3761 2926 3787
rect 2980 3761 3010 3787
rect 3088 3761 3118 3787
rect 3172 3761 3202 3787
rect 3387 3761 3417 3787
rect 3851 3761 4429 3787
rect 4605 3761 4635 3787
rect 4691 3761 4721 3787
rect 4777 3761 4807 3787
rect 4863 3761 4893 3787
rect 4949 3761 4979 3787
rect 5035 3761 5065 3787
rect 5121 3761 5151 3787
rect 5207 3761 5237 3787
rect 5292 3761 5322 3787
rect 5378 3761 5408 3787
rect 5464 3761 5494 3787
rect 5550 3761 5580 3787
rect 5636 3761 5666 3787
rect 5722 3761 5752 3787
rect 5808 3761 5838 3787
rect 5894 3761 5924 3787
rect 5980 3761 6010 3787
rect 6066 3761 6096 3787
rect 6152 3761 6182 3787
rect 6238 3761 6268 3787
rect 6427 3761 6637 3787
rect 1735 3612 1765 3627
rect 1183 3557 1301 3587
rect 1459 3557 1577 3587
rect 1702 3582 1765 3612
rect 1183 3555 1221 3557
rect 1459 3555 1497 3557
rect 1155 3539 1221 3555
rect 1155 3505 1171 3539
rect 1205 3505 1221 3539
rect 1431 3539 1497 3555
rect 1155 3489 1221 3505
rect 1263 3499 1329 3515
rect 1263 3465 1279 3499
rect 1313 3465 1329 3499
rect 1431 3505 1447 3539
rect 1481 3505 1497 3539
rect 1702 3529 1732 3582
rect 1819 3538 1849 3627
rect 2086 3590 2116 3677
rect 2178 3639 2208 3677
rect 1431 3489 1497 3505
rect 1539 3499 1605 3515
rect 1263 3449 1329 3465
rect 1539 3465 1555 3499
rect 1589 3465 1605 3499
rect 1539 3449 1605 3465
rect 1678 3513 1732 3529
rect 1678 3479 1688 3513
rect 1722 3479 1732 3513
rect 1774 3528 1849 3538
rect 1774 3494 1790 3528
rect 1824 3494 1849 3528
rect 1987 3574 2116 3590
rect 2162 3629 2228 3639
rect 2162 3595 2178 3629
rect 2212 3595 2228 3629
rect 2162 3585 2228 3595
rect 1987 3540 1997 3574
rect 2031 3560 2116 3574
rect 2031 3540 2104 3560
rect 2277 3543 2307 3677
rect 2417 3619 2447 3677
rect 2417 3603 2472 3619
rect 2417 3569 2427 3603
rect 2461 3569 2472 3603
rect 2417 3553 2472 3569
rect 1987 3524 2104 3540
rect 1774 3484 1849 3494
rect 1678 3463 1732 3479
rect 1263 3447 1301 3449
rect 1539 3447 1577 3449
rect 1183 3421 1301 3447
rect 1459 3421 1577 3447
rect 1702 3440 1732 3463
rect 1702 3410 1765 3440
rect 1735 3395 1765 3410
rect 1819 3395 1849 3484
rect 2074 3395 2104 3524
rect 2169 3513 2307 3543
rect 2169 3483 2200 3513
rect 2146 3467 2200 3483
rect 2146 3433 2156 3467
rect 2190 3433 2200 3467
rect 2146 3417 2200 3433
rect 2242 3461 2308 3471
rect 2242 3427 2258 3461
rect 2292 3427 2308 3461
rect 2242 3417 2308 3427
rect 2169 3383 2199 3417
rect 2265 3383 2295 3417
rect 2431 3395 2461 3553
rect 2514 3483 2544 3677
rect 2711 3578 2741 3593
rect 2635 3548 2741 3578
rect 2635 3531 2665 3548
rect 2599 3515 2665 3531
rect 2503 3467 2557 3483
rect 2503 3433 2513 3467
rect 2547 3433 2557 3467
rect 2599 3481 2609 3515
rect 2643 3481 2665 3515
rect 2810 3543 2840 3677
rect 2896 3645 2926 3677
rect 2882 3629 2936 3645
rect 2882 3595 2892 3629
rect 2926 3595 2936 3629
rect 2882 3579 2936 3595
rect 2810 3531 2860 3543
rect 2810 3519 2873 3531
rect 2810 3513 2897 3519
rect 2831 3503 2897 3513
rect 2831 3501 2853 3503
rect 2599 3465 2665 3481
rect 2635 3439 2665 3465
rect 2734 3455 2801 3471
rect 2503 3417 2557 3433
rect 2503 3395 2533 3417
rect 2734 3421 2757 3455
rect 2791 3421 2801 3455
rect 2734 3405 2801 3421
rect 2843 3469 2853 3501
rect 2887 3469 2897 3503
rect 2843 3453 2897 3469
rect 2980 3493 3010 3677
rect 3088 3521 3118 3677
rect 3172 3629 3202 3677
rect 3160 3613 3214 3629
rect 3160 3579 3170 3613
rect 3204 3579 3214 3613
rect 3160 3563 3214 3579
rect 3083 3505 3137 3521
rect 2980 3477 3041 3493
rect 2980 3457 2997 3477
rect 2734 3383 2764 3405
rect 2843 3383 2873 3453
rect 2939 3443 2997 3457
rect 3031 3443 3041 3477
rect 3083 3471 3093 3505
rect 3127 3471 3137 3505
rect 3083 3455 3137 3471
rect 2939 3427 3041 3443
rect 2939 3395 2969 3427
rect 3088 3395 3118 3455
rect 3179 3395 3209 3563
rect 3851 3561 4429 3587
rect 6795 3755 6825 3781
rect 6879 3755 6909 3781
rect 7146 3761 7176 3787
rect 7238 3761 7268 3787
rect 7337 3761 7367 3787
rect 7477 3761 7507 3787
rect 7574 3761 7604 3787
rect 7771 3761 7801 3787
rect 7870 3761 7900 3787
rect 7956 3761 7986 3787
rect 8040 3761 8070 3787
rect 8148 3761 8178 3787
rect 8232 3761 8262 3787
rect 8447 3761 8477 3787
rect 8635 3761 8753 3787
rect 6795 3612 6825 3627
rect 6427 3561 6637 3587
rect 6762 3582 6825 3612
rect 3387 3529 3417 3561
rect 3358 3513 3417 3529
rect 3358 3479 3368 3513
rect 3402 3479 3417 3513
rect 3851 3539 4115 3561
rect 3851 3505 3867 3539
rect 3901 3505 3966 3539
rect 4000 3505 4065 3539
rect 4099 3505 4115 3539
rect 4605 3529 4635 3561
rect 4691 3529 4721 3561
rect 4777 3529 4807 3561
rect 4863 3529 4893 3561
rect 4949 3529 4979 3561
rect 5035 3529 5065 3561
rect 5121 3529 5151 3561
rect 5207 3529 5237 3561
rect 5292 3529 5322 3561
rect 5378 3529 5408 3561
rect 5464 3529 5494 3561
rect 5550 3529 5580 3561
rect 5636 3529 5666 3561
rect 5722 3529 5752 3561
rect 5808 3529 5838 3561
rect 5894 3529 5924 3561
rect 3851 3489 4115 3505
rect 4157 3503 4429 3519
rect 3358 3463 3417 3479
rect 3387 3441 3417 3463
rect 4157 3469 4173 3503
rect 4207 3469 4276 3503
rect 4310 3469 4379 3503
rect 4413 3469 4429 3503
rect 4157 3447 4429 3469
rect 3851 3421 4429 3447
rect 4605 3513 5924 3529
rect 4605 3479 4830 3513
rect 4864 3479 4898 3513
rect 4932 3479 4966 3513
rect 5000 3479 5034 3513
rect 5068 3479 5102 3513
rect 5136 3479 5170 3513
rect 5204 3479 5238 3513
rect 5272 3479 5306 3513
rect 5340 3479 5374 3513
rect 5408 3479 5442 3513
rect 5476 3479 5510 3513
rect 5544 3479 5578 3513
rect 5612 3479 5646 3513
rect 5680 3479 5714 3513
rect 5748 3479 5782 3513
rect 5816 3479 5850 3513
rect 5884 3479 5924 3513
rect 4605 3454 5924 3479
rect 4605 3395 4635 3454
rect 4691 3395 4721 3454
rect 4777 3395 4807 3454
rect 4863 3395 4893 3454
rect 4949 3395 4979 3454
rect 5035 3395 5065 3454
rect 5121 3395 5151 3454
rect 5207 3395 5237 3454
rect 5292 3395 5322 3454
rect 5378 3395 5408 3454
rect 5464 3395 5494 3454
rect 5550 3395 5580 3454
rect 5636 3395 5666 3454
rect 5722 3395 5752 3454
rect 5808 3395 5838 3454
rect 5894 3395 5924 3454
rect 5980 3546 6010 3561
rect 6066 3546 6096 3561
rect 6152 3546 6182 3561
rect 6238 3546 6268 3561
rect 6427 3555 6511 3561
rect 5980 3513 6327 3546
rect 5980 3479 6277 3513
rect 6311 3479 6327 3513
rect 6369 3539 6511 3555
rect 6369 3505 6385 3539
rect 6419 3505 6511 3539
rect 6762 3529 6792 3582
rect 6879 3538 6909 3627
rect 7146 3590 7176 3677
rect 7238 3639 7268 3677
rect 6369 3489 6511 3505
rect 6553 3503 6695 3519
rect 5980 3444 6327 3479
rect 6553 3469 6645 3503
rect 6679 3469 6695 3503
rect 6553 3453 6695 3469
rect 6738 3513 6792 3529
rect 6738 3479 6748 3513
rect 6782 3479 6792 3513
rect 6834 3528 6909 3538
rect 6834 3494 6850 3528
rect 6884 3494 6909 3528
rect 7047 3574 7176 3590
rect 7222 3629 7288 3639
rect 7222 3595 7238 3629
rect 7272 3595 7288 3629
rect 7222 3585 7288 3595
rect 7047 3540 7057 3574
rect 7091 3560 7176 3574
rect 7091 3540 7164 3560
rect 7337 3543 7367 3677
rect 7477 3619 7507 3677
rect 7477 3603 7532 3619
rect 7477 3569 7487 3603
rect 7521 3569 7532 3603
rect 7477 3553 7532 3569
rect 7047 3524 7164 3540
rect 6834 3484 6909 3494
rect 6738 3463 6792 3479
rect 6553 3447 6637 3453
rect 5980 3395 6010 3444
rect 6066 3395 6096 3444
rect 6152 3395 6182 3444
rect 6238 3395 6268 3444
rect 6427 3421 6637 3447
rect 6762 3440 6792 3463
rect 6762 3410 6825 3440
rect 6795 3395 6825 3410
rect 6879 3395 6909 3484
rect 7134 3395 7164 3524
rect 7229 3513 7367 3543
rect 7229 3483 7260 3513
rect 7206 3467 7260 3483
rect 7206 3433 7216 3467
rect 7250 3433 7260 3467
rect 7206 3417 7260 3433
rect 7302 3461 7368 3471
rect 7302 3427 7318 3461
rect 7352 3427 7368 3461
rect 7302 3417 7368 3427
rect 7229 3383 7259 3417
rect 7325 3383 7355 3417
rect 7491 3395 7521 3553
rect 7574 3483 7604 3677
rect 7771 3578 7801 3593
rect 7695 3548 7801 3578
rect 7695 3531 7725 3548
rect 7659 3515 7725 3531
rect 7563 3467 7617 3483
rect 7563 3433 7573 3467
rect 7607 3433 7617 3467
rect 7659 3481 7669 3515
rect 7703 3481 7725 3515
rect 7870 3543 7900 3677
rect 7956 3645 7986 3677
rect 7942 3629 7996 3645
rect 7942 3595 7952 3629
rect 7986 3595 7996 3629
rect 7942 3579 7996 3595
rect 7870 3531 7920 3543
rect 7870 3519 7933 3531
rect 7870 3513 7957 3519
rect 7891 3503 7957 3513
rect 7891 3501 7913 3503
rect 7659 3465 7725 3481
rect 7695 3439 7725 3465
rect 7794 3455 7861 3471
rect 7563 3417 7617 3433
rect 7563 3395 7593 3417
rect 7794 3421 7817 3455
rect 7851 3421 7861 3455
rect 7794 3405 7861 3421
rect 7903 3469 7913 3501
rect 7947 3469 7957 3503
rect 7903 3453 7957 3469
rect 8040 3493 8070 3677
rect 8148 3521 8178 3677
rect 8232 3629 8262 3677
rect 8220 3613 8274 3629
rect 8220 3579 8230 3613
rect 8264 3579 8274 3613
rect 8220 3563 8274 3579
rect 8143 3505 8197 3521
rect 8040 3477 8101 3493
rect 8040 3457 8057 3477
rect 7794 3383 7824 3405
rect 7903 3383 7933 3453
rect 7999 3443 8057 3457
rect 8091 3443 8101 3477
rect 8143 3471 8153 3505
rect 8187 3471 8197 3505
rect 8143 3455 8197 3471
rect 7999 3427 8101 3443
rect 7999 3395 8029 3427
rect 8148 3395 8178 3455
rect 8239 3395 8269 3563
rect 9187 3753 9217 3779
rect 9282 3761 9312 3787
rect 9366 3761 9396 3787
rect 9555 3761 9949 3787
rect 10107 3761 10137 3787
rect 10195 3761 10225 3787
rect 10383 3761 10777 3787
rect 11027 3761 11057 3787
rect 11115 3761 11145 3787
rect 11303 3761 11881 3787
rect 12039 3761 12069 3787
rect 12254 3761 12284 3787
rect 12338 3761 12368 3787
rect 12446 3761 12476 3787
rect 12530 3761 12560 3787
rect 12616 3761 12646 3787
rect 12715 3761 12745 3787
rect 12912 3761 12942 3787
rect 13009 3761 13039 3787
rect 13149 3761 13179 3787
rect 13248 3761 13278 3787
rect 13340 3761 13370 3787
rect 8447 3529 8477 3561
rect 8635 3557 8753 3587
rect 8635 3555 8673 3557
rect 8418 3513 8477 3529
rect 8418 3479 8428 3513
rect 8462 3479 8477 3513
rect 8607 3539 8673 3555
rect 8607 3505 8623 3539
rect 8657 3505 8673 3539
rect 9187 3529 9217 3625
rect 9555 3561 9949 3587
rect 9282 3529 9312 3561
rect 9366 3529 9396 3561
rect 8607 3489 8673 3505
rect 8715 3499 8781 3515
rect 8418 3463 8477 3479
rect 8447 3441 8477 3463
rect 8715 3465 8731 3499
rect 8765 3465 8781 3499
rect 8715 3449 8781 3465
rect 9135 3513 9217 3529
rect 9135 3479 9145 3513
rect 9179 3479 9217 3513
rect 9135 3463 9217 3479
rect 9259 3513 9396 3529
rect 9259 3479 9269 3513
rect 9303 3479 9396 3513
rect 9555 3539 9731 3561
rect 10107 3542 10137 3603
rect 10195 3588 10225 3603
rect 10195 3564 10231 3588
rect 11027 3588 11057 3603
rect 9555 3505 9571 3539
rect 9605 3505 9681 3539
rect 9715 3505 9731 3539
rect 10103 3526 10157 3542
rect 9555 3489 9731 3505
rect 9773 3503 9949 3519
rect 9259 3463 9396 3479
rect 8715 3447 8753 3449
rect 8635 3421 8753 3447
rect 9187 3395 9217 3463
rect 9282 3441 9312 3463
rect 9366 3441 9396 3463
rect 9773 3469 9789 3503
rect 9823 3469 9899 3503
rect 9933 3469 9949 3503
rect 10103 3492 10113 3526
rect 10147 3492 10157 3526
rect 10103 3476 10157 3492
rect 10201 3529 10231 3564
rect 10383 3561 10777 3587
rect 11021 3564 11057 3588
rect 10383 3539 10559 3561
rect 10201 3513 10277 3529
rect 10201 3479 10233 3513
rect 10267 3479 10277 3513
rect 10383 3505 10399 3539
rect 10433 3505 10509 3539
rect 10543 3505 10559 3539
rect 11021 3529 11051 3564
rect 11115 3542 11145 3603
rect 11303 3561 11881 3587
rect 12254 3629 12284 3677
rect 12242 3613 12296 3629
rect 12242 3579 12252 3613
rect 12286 3579 12296 3613
rect 12242 3563 12296 3579
rect 10383 3489 10559 3505
rect 10601 3503 10777 3519
rect 9773 3447 9949 3469
rect 9555 3421 9949 3447
rect 10107 3415 10137 3476
rect 10201 3463 10277 3479
rect 10601 3469 10617 3503
rect 10651 3469 10727 3503
rect 10761 3469 10777 3503
rect 10201 3454 10231 3463
rect 10195 3430 10231 3454
rect 10601 3447 10777 3469
rect 10975 3513 11051 3529
rect 10975 3479 10985 3513
rect 11019 3479 11051 3513
rect 10975 3463 11051 3479
rect 11095 3526 11149 3542
rect 11095 3492 11105 3526
rect 11139 3492 11149 3526
rect 11095 3476 11149 3492
rect 11303 3539 11567 3561
rect 11303 3505 11319 3539
rect 11353 3505 11418 3539
rect 11452 3505 11517 3539
rect 11551 3505 11567 3539
rect 12039 3529 12069 3561
rect 11303 3489 11567 3505
rect 11609 3503 11881 3519
rect 10195 3415 10225 3430
rect 10383 3421 10777 3447
rect 11021 3454 11051 3463
rect 11021 3430 11057 3454
rect 11027 3415 11057 3430
rect 11115 3415 11145 3476
rect 11609 3469 11625 3503
rect 11659 3469 11728 3503
rect 11762 3469 11831 3503
rect 11865 3469 11881 3503
rect 11609 3447 11881 3469
rect 11303 3421 11881 3447
rect 12039 3513 12098 3529
rect 12039 3479 12054 3513
rect 12088 3479 12098 3513
rect 12039 3463 12098 3479
rect 12039 3441 12069 3463
rect 12247 3395 12277 3563
rect 12338 3521 12368 3677
rect 12319 3505 12373 3521
rect 12319 3471 12329 3505
rect 12363 3471 12373 3505
rect 12446 3493 12476 3677
rect 12530 3645 12560 3677
rect 12520 3629 12574 3645
rect 12520 3595 12530 3629
rect 12564 3595 12574 3629
rect 12520 3579 12574 3595
rect 12616 3543 12646 3677
rect 13607 3755 13637 3781
rect 13691 3755 13721 3781
rect 14155 3761 15101 3787
rect 15259 3761 16205 3787
rect 16363 3761 17309 3787
rect 17467 3761 18413 3787
rect 18663 3761 18781 3787
rect 12715 3578 12745 3593
rect 12715 3548 12821 3578
rect 12596 3531 12646 3543
rect 12583 3519 12646 3531
rect 12319 3455 12373 3471
rect 12415 3477 12476 3493
rect 12338 3395 12368 3455
rect 12415 3443 12425 3477
rect 12459 3457 12476 3477
rect 12559 3513 12646 3519
rect 12791 3531 12821 3548
rect 12791 3515 12857 3531
rect 12559 3503 12625 3513
rect 12559 3469 12569 3503
rect 12603 3501 12625 3503
rect 12603 3469 12613 3501
rect 12791 3481 12813 3515
rect 12847 3481 12857 3515
rect 12912 3483 12942 3677
rect 13009 3619 13039 3677
rect 12984 3603 13039 3619
rect 12984 3569 12995 3603
rect 13029 3569 13039 3603
rect 12984 3553 13039 3569
rect 12459 3443 12517 3457
rect 12559 3453 12613 3469
rect 12415 3427 12517 3443
rect 12487 3395 12517 3427
rect 12583 3383 12613 3453
rect 12655 3455 12722 3471
rect 12655 3421 12665 3455
rect 12699 3421 12722 3455
rect 12791 3465 12857 3481
rect 12899 3467 12953 3483
rect 12791 3439 12821 3465
rect 12655 3405 12722 3421
rect 12692 3383 12722 3405
rect 12899 3433 12909 3467
rect 12943 3433 12953 3467
rect 12899 3417 12953 3433
rect 12923 3395 12953 3417
rect 12995 3395 13025 3553
rect 13149 3543 13179 3677
rect 13248 3639 13278 3677
rect 13228 3629 13294 3639
rect 13228 3595 13244 3629
rect 13278 3595 13294 3629
rect 13228 3585 13294 3595
rect 13340 3590 13370 3677
rect 13340 3574 13469 3590
rect 13340 3560 13425 3574
rect 13149 3513 13287 3543
rect 13256 3483 13287 3513
rect 13352 3540 13425 3560
rect 13459 3540 13469 3574
rect 13352 3524 13469 3540
rect 13607 3538 13637 3627
rect 13691 3612 13721 3627
rect 13691 3582 13754 3612
rect 13607 3528 13682 3538
rect 13148 3461 13214 3471
rect 13148 3427 13164 3461
rect 13198 3427 13214 3461
rect 13148 3417 13214 3427
rect 13256 3467 13310 3483
rect 13256 3433 13266 3467
rect 13300 3433 13310 3467
rect 13256 3417 13310 3433
rect 13161 3383 13191 3417
rect 13257 3383 13287 3417
rect 13352 3395 13382 3524
rect 13607 3494 13632 3528
rect 13666 3494 13682 3528
rect 13607 3484 13682 3494
rect 13724 3529 13754 3582
rect 14155 3561 15101 3587
rect 15259 3561 16205 3587
rect 16363 3561 17309 3587
rect 17467 3561 18413 3587
rect 14155 3539 14605 3561
rect 13724 3513 13778 3529
rect 13607 3395 13637 3484
rect 13724 3479 13734 3513
rect 13768 3479 13778 3513
rect 14155 3505 14427 3539
rect 14461 3505 14605 3539
rect 15259 3539 15709 3561
rect 14155 3489 14605 3505
rect 14647 3503 15101 3519
rect 13724 3463 13778 3479
rect 14647 3469 14791 3503
rect 14825 3469 15101 3503
rect 15259 3505 15531 3539
rect 15565 3505 15709 3539
rect 16363 3539 16813 3561
rect 15259 3489 15709 3505
rect 15751 3503 16205 3519
rect 13724 3440 13754 3463
rect 14647 3447 15101 3469
rect 15751 3469 15895 3503
rect 15929 3469 16205 3503
rect 16363 3505 16635 3539
rect 16669 3505 16813 3539
rect 17467 3539 17917 3561
rect 18663 3557 18781 3587
rect 16363 3489 16813 3505
rect 16855 3503 17309 3519
rect 15751 3447 16205 3469
rect 16855 3469 16999 3503
rect 17033 3469 17309 3503
rect 17467 3505 17739 3539
rect 17773 3505 17917 3539
rect 18743 3555 18781 3557
rect 18743 3539 18809 3555
rect 17467 3489 17917 3505
rect 17959 3503 18413 3519
rect 16855 3447 17309 3469
rect 17959 3469 18103 3503
rect 18137 3469 18413 3503
rect 17959 3447 18413 3469
rect 18635 3499 18701 3515
rect 18635 3465 18651 3499
rect 18685 3465 18701 3499
rect 18743 3505 18759 3539
rect 18793 3505 18809 3539
rect 18743 3489 18809 3505
rect 18635 3449 18701 3465
rect 13691 3410 13754 3440
rect 13691 3395 13721 3410
rect 14155 3421 15101 3447
rect 15259 3421 16205 3447
rect 16363 3421 17309 3447
rect 17467 3421 18413 3447
rect 18663 3447 18701 3449
rect 18663 3421 18781 3447
rect 1183 3285 1301 3311
rect 1459 3285 1577 3311
rect 1735 3285 1765 3311
rect 1819 3285 1849 3311
rect 2074 3285 2104 3311
rect 2169 3285 2199 3311
rect 2265 3285 2295 3311
rect 2431 3285 2461 3311
rect 2503 3285 2533 3311
rect 2635 3285 2665 3311
rect 2734 3285 2764 3311
rect 2843 3285 2873 3311
rect 2939 3285 2969 3311
rect 3088 3285 3118 3311
rect 3179 3285 3209 3311
rect 3387 3285 3417 3311
rect 3851 3285 4429 3311
rect 4605 3285 4635 3311
rect 4691 3285 4721 3311
rect 4777 3285 4807 3311
rect 4863 3285 4893 3311
rect 4949 3285 4979 3311
rect 5035 3285 5065 3311
rect 5121 3285 5151 3311
rect 5207 3285 5237 3311
rect 5292 3285 5322 3311
rect 5378 3285 5408 3311
rect 5464 3285 5494 3311
rect 5550 3285 5580 3311
rect 5636 3285 5666 3311
rect 5722 3285 5752 3311
rect 5808 3285 5838 3311
rect 5894 3285 5924 3311
rect 5980 3285 6010 3311
rect 6066 3285 6096 3311
rect 6152 3285 6182 3311
rect 6238 3285 6268 3311
rect 6427 3285 6637 3311
rect 6795 3285 6825 3311
rect 6879 3285 6909 3311
rect 7134 3285 7164 3311
rect 7229 3285 7259 3311
rect 7325 3285 7355 3311
rect 7491 3285 7521 3311
rect 7563 3285 7593 3311
rect 7695 3285 7725 3311
rect 7794 3285 7824 3311
rect 7903 3285 7933 3311
rect 7999 3285 8029 3311
rect 8148 3285 8178 3311
rect 8239 3285 8269 3311
rect 8447 3285 8477 3311
rect 8635 3285 8753 3311
rect 9187 3285 9217 3311
rect 9282 3285 9312 3311
rect 9366 3285 9396 3311
rect 9555 3285 9949 3311
rect 10107 3285 10137 3311
rect 10195 3285 10225 3311
rect 10383 3285 10777 3311
rect 11027 3285 11057 3311
rect 11115 3285 11145 3311
rect 11303 3285 11881 3311
rect 12039 3285 12069 3311
rect 12247 3285 12277 3311
rect 12338 3285 12368 3311
rect 12487 3285 12517 3311
rect 12583 3285 12613 3311
rect 12692 3285 12722 3311
rect 12791 3285 12821 3311
rect 12923 3285 12953 3311
rect 12995 3285 13025 3311
rect 13161 3285 13191 3311
rect 13257 3285 13287 3311
rect 13352 3285 13382 3311
rect 13607 3285 13637 3311
rect 13691 3285 13721 3311
rect 14155 3285 15101 3311
rect 15259 3285 16205 3311
rect 16363 3285 17309 3311
rect 17467 3285 18413 3311
rect 18663 3285 18781 3311
rect 1183 3217 1301 3243
rect 1459 3217 1853 3243
rect 2011 3217 2041 3243
rect 2219 3217 2249 3243
rect 2310 3217 2340 3243
rect 2459 3217 2489 3243
rect 2555 3217 2585 3243
rect 2664 3217 2694 3243
rect 2763 3217 2793 3243
rect 2895 3217 2925 3243
rect 2967 3217 2997 3243
rect 3133 3217 3163 3243
rect 3229 3217 3259 3243
rect 3324 3217 3354 3243
rect 3579 3217 3609 3243
rect 3663 3217 3693 3243
rect 3851 3217 4061 3243
rect 4219 3217 4249 3243
rect 4303 3217 4333 3243
rect 4491 3217 4521 3243
rect 4586 3217 4616 3243
rect 4696 3217 4726 3243
rect 4792 3217 4822 3243
rect 4906 3217 4936 3243
rect 4978 3217 5008 3243
rect 5166 3217 5196 3243
rect 5238 3217 5268 3243
rect 5334 3217 5364 3243
rect 5406 3217 5436 3243
rect 5482 3217 5512 3243
rect 5606 3217 5636 3243
rect 5794 3217 5824 3243
rect 5889 3217 5919 3243
rect 6427 3217 7005 3243
rect 7255 3217 7285 3243
rect 7463 3217 7493 3243
rect 7554 3217 7584 3243
rect 7703 3217 7733 3243
rect 7799 3217 7829 3243
rect 7908 3217 7938 3243
rect 8007 3217 8037 3243
rect 8139 3217 8169 3243
rect 8211 3217 8241 3243
rect 8377 3217 8407 3243
rect 8473 3217 8503 3243
rect 8568 3217 8598 3243
rect 8823 3217 8853 3243
rect 8907 3217 8937 3243
rect 9095 3217 9305 3243
rect 9464 3217 9494 3243
rect 9550 3217 9580 3243
rect 9636 3217 9666 3243
rect 9722 3217 9752 3243
rect 9808 3217 9838 3243
rect 9894 3217 9924 3243
rect 9980 3217 10010 3243
rect 10066 3217 10096 3243
rect 10152 3217 10182 3243
rect 10238 3217 10268 3243
rect 10324 3217 10354 3243
rect 10410 3217 10440 3243
rect 10495 3217 10525 3243
rect 10581 3217 10611 3243
rect 10667 3217 10697 3243
rect 10753 3217 10783 3243
rect 10839 3217 10869 3243
rect 10925 3217 10955 3243
rect 11011 3217 11041 3243
rect 11097 3217 11127 3243
rect 11763 3217 11793 3243
rect 11971 3217 12001 3243
rect 12062 3217 12092 3243
rect 12211 3217 12241 3243
rect 12307 3217 12337 3243
rect 12416 3217 12446 3243
rect 12515 3217 12545 3243
rect 12647 3217 12677 3243
rect 12719 3217 12749 3243
rect 12885 3217 12915 3243
rect 12981 3217 13011 3243
rect 13076 3217 13106 3243
rect 13331 3217 13361 3243
rect 13415 3217 13445 3243
rect 13603 3217 13813 3243
rect 13971 3217 14001 3243
rect 14066 3217 14096 3243
rect 14150 3217 14180 3243
rect 14339 3217 15285 3243
rect 15443 3217 16389 3243
rect 16731 3217 17677 3243
rect 17835 3217 18413 3243
rect 18663 3217 18781 3243
rect 1183 3081 1301 3107
rect 1459 3081 1853 3107
rect 1263 3079 1301 3081
rect 1263 3063 1329 3079
rect 1155 3023 1221 3039
rect 1155 2989 1171 3023
rect 1205 2989 1221 3023
rect 1263 3029 1279 3063
rect 1313 3029 1329 3063
rect 1677 3059 1853 3081
rect 1263 3013 1329 3029
rect 1459 3023 1635 3039
rect 1155 2973 1221 2989
rect 1183 2971 1221 2973
rect 1459 2989 1475 3023
rect 1509 2989 1585 3023
rect 1619 2989 1635 3023
rect 1677 3025 1693 3059
rect 1727 3025 1803 3059
rect 1837 3025 1853 3059
rect 1677 3009 1853 3025
rect 2011 3065 2041 3087
rect 2011 3049 2070 3065
rect 2011 3015 2026 3049
rect 2060 3015 2070 3049
rect 1183 2941 1301 2971
rect 1459 2967 1635 2989
rect 2011 2999 2070 3015
rect 2011 2967 2041 2999
rect 1459 2941 1853 2967
rect 2219 2965 2249 3133
rect 2310 3073 2340 3133
rect 2459 3101 2489 3133
rect 2387 3085 2489 3101
rect 2291 3057 2345 3073
rect 2291 3023 2301 3057
rect 2335 3023 2345 3057
rect 2387 3051 2397 3085
rect 2431 3071 2489 3085
rect 2555 3075 2585 3145
rect 2664 3123 2694 3145
rect 2431 3051 2448 3071
rect 2387 3035 2448 3051
rect 2291 3007 2345 3023
rect 2214 2949 2268 2965
rect 2214 2915 2224 2949
rect 2258 2915 2268 2949
rect 2214 2899 2268 2915
rect 2226 2851 2256 2899
rect 2310 2851 2340 3007
rect 2418 2851 2448 3035
rect 2531 3059 2585 3075
rect 2531 3025 2541 3059
rect 2575 3027 2585 3059
rect 2627 3107 2694 3123
rect 2627 3073 2637 3107
rect 2671 3073 2694 3107
rect 2895 3111 2925 3133
rect 2871 3095 2925 3111
rect 2627 3057 2694 3073
rect 2763 3063 2793 3089
rect 2763 3047 2829 3063
rect 2575 3025 2597 3027
rect 2531 3015 2597 3025
rect 2531 3009 2618 3015
rect 2555 2997 2618 3009
rect 2568 2985 2618 2997
rect 2492 2933 2546 2949
rect 2492 2899 2502 2933
rect 2536 2899 2546 2933
rect 2492 2883 2546 2899
rect 2502 2851 2532 2883
rect 2588 2851 2618 2985
rect 2763 3013 2785 3047
rect 2819 3013 2829 3047
rect 2871 3061 2881 3095
rect 2915 3061 2925 3095
rect 2871 3045 2925 3061
rect 2763 2997 2829 3013
rect 2763 2980 2793 2997
rect 2687 2950 2793 2980
rect 2687 2935 2717 2950
rect 2884 2851 2914 3045
rect 2967 2975 2997 3133
rect 3133 3111 3163 3145
rect 3229 3111 3259 3145
rect 3120 3101 3186 3111
rect 3120 3067 3136 3101
rect 3170 3067 3186 3101
rect 3120 3057 3186 3067
rect 3228 3095 3282 3111
rect 3228 3061 3238 3095
rect 3272 3061 3282 3095
rect 3228 3045 3282 3061
rect 3228 3015 3259 3045
rect 3121 2985 3259 3015
rect 3324 3004 3354 3133
rect 3579 3044 3609 3133
rect 3663 3118 3693 3133
rect 3663 3088 3726 3118
rect 4219 3118 4249 3133
rect 3696 3065 3726 3088
rect 3851 3081 4061 3107
rect 3977 3075 4061 3081
rect 4186 3088 4249 3118
rect 3696 3049 3750 3065
rect 3579 3034 3654 3044
rect 3324 2988 3441 3004
rect 2956 2959 3011 2975
rect 2956 2925 2967 2959
rect 3001 2925 3011 2959
rect 2956 2909 3011 2925
rect 2981 2851 3011 2909
rect 3121 2851 3151 2985
rect 3324 2968 3397 2988
rect 3312 2954 3397 2968
rect 3431 2954 3441 2988
rect 3200 2933 3266 2943
rect 3200 2899 3216 2933
rect 3250 2899 3266 2933
rect 3200 2889 3266 2899
rect 3312 2938 3441 2954
rect 3579 3000 3604 3034
rect 3638 3000 3654 3034
rect 3579 2990 3654 3000
rect 3696 3015 3706 3049
rect 3740 3015 3750 3049
rect 3977 3059 4119 3075
rect 3696 2999 3750 3015
rect 3793 3023 3935 3039
rect 3220 2851 3250 2889
rect 3312 2851 3342 2938
rect 3579 2901 3609 2990
rect 3696 2946 3726 2999
rect 3793 2989 3809 3023
rect 3843 2989 3935 3023
rect 3977 3025 4069 3059
rect 4103 3025 4119 3059
rect 4186 3050 4216 3088
rect 3977 3009 4119 3025
rect 4162 3034 4216 3050
rect 4303 3044 4333 3133
rect 4586 3123 4616 3145
rect 4586 3107 4654 3123
rect 4491 3063 4521 3089
rect 4586 3073 4610 3107
rect 4644 3073 4654 3107
rect 3793 2973 3935 2989
rect 4162 3000 4172 3034
rect 4206 3000 4216 3034
rect 4162 2984 4216 3000
rect 4258 3034 4333 3044
rect 4258 3000 4274 3034
rect 4308 3000 4333 3034
rect 4258 2990 4333 3000
rect 4484 3047 4538 3063
rect 4586 3057 4654 3073
rect 4696 3111 4726 3145
rect 4696 3095 4750 3111
rect 4696 3061 4706 3095
rect 4740 3061 4750 3095
rect 4484 3013 4494 3047
rect 4528 3013 4538 3047
rect 4696 3045 4750 3061
rect 4696 3015 4726 3045
rect 4484 2997 4538 3013
rect 3663 2916 3726 2946
rect 3851 2967 3935 2973
rect 3851 2941 4061 2967
rect 4186 2946 4216 2984
rect 3663 2901 3693 2916
rect 1183 2741 1301 2767
rect 1459 2741 1853 2767
rect 2011 2741 2041 2767
rect 2226 2741 2256 2767
rect 2310 2741 2340 2767
rect 2418 2741 2448 2767
rect 2502 2741 2532 2767
rect 2588 2741 2618 2767
rect 2687 2741 2717 2767
rect 2884 2741 2914 2767
rect 2981 2741 3011 2767
rect 3121 2741 3151 2767
rect 3220 2741 3250 2767
rect 3312 2741 3342 2767
rect 3579 2747 3609 2773
rect 3663 2747 3693 2773
rect 4186 2916 4249 2946
rect 4219 2901 4249 2916
rect 4303 2901 4333 2990
rect 4491 2935 4521 2997
rect 4588 2985 4726 3015
rect 3851 2741 4061 2767
rect 4219 2747 4249 2773
rect 4303 2747 4333 2773
rect 4588 2851 4618 2985
rect 4792 2949 4822 3133
rect 4906 3101 4936 3133
rect 4868 3085 4936 3101
rect 4868 3051 4878 3085
rect 4912 3071 4936 3085
rect 4978 3117 5008 3133
rect 5166 3117 5196 3133
rect 4978 3081 5196 3117
rect 4912 3051 4928 3071
rect 4868 3035 4928 3051
rect 4660 2933 4726 2943
rect 4660 2899 4676 2933
rect 4710 2899 4726 2933
rect 4660 2889 4726 2899
rect 4792 2933 4856 2949
rect 4792 2899 4812 2933
rect 4846 2899 4856 2933
rect 4672 2851 4702 2889
rect 4792 2883 4856 2899
rect 4792 2851 4822 2883
rect 4898 2851 4928 3035
rect 4978 3017 5008 3081
rect 5238 3039 5268 3133
rect 5334 3111 5364 3133
rect 5310 3095 5364 3111
rect 5310 3061 5320 3095
rect 5354 3061 5364 3095
rect 5310 3045 5364 3061
rect 5174 3029 5268 3039
rect 4970 3001 5096 3017
rect 4970 2967 4980 3001
rect 5014 2967 5096 3001
rect 5174 2995 5190 3029
rect 5224 3003 5268 3029
rect 5406 3003 5436 3133
rect 5482 3101 5512 3133
rect 5482 3085 5536 3101
rect 5482 3051 5492 3085
rect 5526 3051 5536 3085
rect 5482 3035 5536 3051
rect 5606 3045 5636 3109
rect 5794 3045 5824 3133
rect 5889 3065 5919 3087
rect 6427 3081 7005 3107
rect 5224 2995 5280 3003
rect 5174 2985 5280 2995
rect 5238 2973 5280 2985
rect 4970 2951 5096 2967
rect 4982 2851 5012 2951
rect 5066 2851 5096 2951
rect 5142 2933 5208 2943
rect 5142 2899 5158 2933
rect 5192 2899 5208 2933
rect 5142 2889 5208 2899
rect 5142 2851 5172 2889
rect 5250 2851 5280 2973
rect 5322 2973 5436 3003
rect 5322 2949 5386 2973
rect 5322 2915 5342 2949
rect 5376 2915 5386 2949
rect 5506 2957 5536 3035
rect 5578 3029 5824 3045
rect 5578 2995 5588 3029
rect 5622 2995 5824 3029
rect 5866 3049 5920 3065
rect 5866 3015 5876 3049
rect 5910 3015 5920 3049
rect 6733 3059 7005 3081
rect 5866 2999 5920 3015
rect 6427 3023 6691 3039
rect 5578 2979 5824 2995
rect 5506 2927 5540 2957
rect 5606 2935 5636 2979
rect 5322 2899 5386 2915
rect 5322 2851 5352 2899
rect 5510 2851 5540 2927
rect 5794 2895 5824 2979
rect 5889 2967 5919 2999
rect 6427 2989 6443 3023
rect 6477 2989 6542 3023
rect 6576 2989 6641 3023
rect 6675 2989 6691 3023
rect 6733 3025 6749 3059
rect 6783 3025 6852 3059
rect 6886 3025 6955 3059
rect 6989 3025 7005 3059
rect 6733 3009 7005 3025
rect 7255 3065 7285 3087
rect 7255 3049 7314 3065
rect 7255 3015 7270 3049
rect 7304 3015 7314 3049
rect 6427 2967 6691 2989
rect 7255 2999 7314 3015
rect 7255 2967 7285 2999
rect 6427 2941 7005 2967
rect 7463 2965 7493 3133
rect 7554 3073 7584 3133
rect 7703 3101 7733 3133
rect 7631 3085 7733 3101
rect 7535 3057 7589 3073
rect 7535 3023 7545 3057
rect 7579 3023 7589 3057
rect 7631 3051 7641 3085
rect 7675 3071 7733 3085
rect 7799 3075 7829 3145
rect 7908 3123 7938 3145
rect 7675 3051 7692 3071
rect 7631 3035 7692 3051
rect 7535 3007 7589 3023
rect 7458 2949 7512 2965
rect 7458 2915 7468 2949
rect 7502 2915 7512 2949
rect 7458 2899 7512 2915
rect 7470 2851 7500 2899
rect 7554 2851 7584 3007
rect 7662 2851 7692 3035
rect 7775 3059 7829 3075
rect 7775 3025 7785 3059
rect 7819 3027 7829 3059
rect 7871 3107 7938 3123
rect 7871 3073 7881 3107
rect 7915 3073 7938 3107
rect 8139 3111 8169 3133
rect 8115 3095 8169 3111
rect 7871 3057 7938 3073
rect 8007 3063 8037 3089
rect 8007 3047 8073 3063
rect 7819 3025 7841 3027
rect 7775 3015 7841 3025
rect 7775 3009 7862 3015
rect 7799 2997 7862 3009
rect 7812 2985 7862 2997
rect 7736 2933 7790 2949
rect 7736 2899 7746 2933
rect 7780 2899 7790 2933
rect 7736 2883 7790 2899
rect 7746 2851 7776 2883
rect 7832 2851 7862 2985
rect 8007 3013 8029 3047
rect 8063 3013 8073 3047
rect 8115 3061 8125 3095
rect 8159 3061 8169 3095
rect 8115 3045 8169 3061
rect 8007 2997 8073 3013
rect 8007 2980 8037 2997
rect 7931 2950 8037 2980
rect 7931 2935 7961 2950
rect 8128 2851 8158 3045
rect 8211 2975 8241 3133
rect 8377 3111 8407 3145
rect 8473 3111 8503 3145
rect 8364 3101 8430 3111
rect 8364 3067 8380 3101
rect 8414 3067 8430 3101
rect 8364 3057 8430 3067
rect 8472 3095 8526 3111
rect 8472 3061 8482 3095
rect 8516 3061 8526 3095
rect 8472 3045 8526 3061
rect 8472 3015 8503 3045
rect 8365 2985 8503 3015
rect 8568 3004 8598 3133
rect 8823 3044 8853 3133
rect 8907 3118 8937 3133
rect 8907 3088 8970 3118
rect 8940 3065 8970 3088
rect 9095 3081 9305 3107
rect 9464 3084 9494 3133
rect 9550 3084 9580 3133
rect 9636 3084 9666 3133
rect 9722 3084 9752 3133
rect 9221 3075 9305 3081
rect 8940 3049 8994 3065
rect 8823 3034 8898 3044
rect 8568 2988 8685 3004
rect 8200 2959 8255 2975
rect 8200 2925 8211 2959
rect 8245 2925 8255 2959
rect 8200 2909 8255 2925
rect 8225 2851 8255 2909
rect 8365 2851 8395 2985
rect 8568 2968 8641 2988
rect 8556 2954 8641 2968
rect 8675 2954 8685 2988
rect 8444 2933 8510 2943
rect 8444 2899 8460 2933
rect 8494 2899 8510 2933
rect 8444 2889 8510 2899
rect 8556 2938 8685 2954
rect 8823 3000 8848 3034
rect 8882 3000 8898 3034
rect 8823 2990 8898 3000
rect 8940 3015 8950 3049
rect 8984 3015 8994 3049
rect 9221 3059 9363 3075
rect 8940 2999 8994 3015
rect 9037 3023 9179 3039
rect 8464 2851 8494 2889
rect 8556 2851 8586 2938
rect 8823 2901 8853 2990
rect 8940 2946 8970 2999
rect 9037 2989 9053 3023
rect 9087 2989 9179 3023
rect 9221 3025 9313 3059
rect 9347 3025 9363 3059
rect 9221 3009 9363 3025
rect 9405 3049 9752 3084
rect 9405 3015 9421 3049
rect 9455 3015 9752 3049
rect 9037 2973 9179 2989
rect 9405 2982 9752 3015
rect 8907 2916 8970 2946
rect 9095 2967 9179 2973
rect 9464 2967 9494 2982
rect 9550 2967 9580 2982
rect 9636 2967 9666 2982
rect 9722 2967 9752 2982
rect 9808 3074 9838 3133
rect 9894 3074 9924 3133
rect 9980 3074 10010 3133
rect 10066 3074 10096 3133
rect 10152 3074 10182 3133
rect 10238 3074 10268 3133
rect 10324 3074 10354 3133
rect 10410 3074 10440 3133
rect 10495 3074 10525 3133
rect 10581 3074 10611 3133
rect 10667 3074 10697 3133
rect 10753 3074 10783 3133
rect 10839 3074 10869 3133
rect 10925 3074 10955 3133
rect 11011 3074 11041 3133
rect 11097 3074 11127 3133
rect 9808 3049 11127 3074
rect 9808 3015 9848 3049
rect 9882 3015 9916 3049
rect 9950 3015 9984 3049
rect 10018 3015 10052 3049
rect 10086 3015 10120 3049
rect 10154 3015 10188 3049
rect 10222 3015 10256 3049
rect 10290 3015 10324 3049
rect 10358 3015 10392 3049
rect 10426 3015 10460 3049
rect 10494 3015 10528 3049
rect 10562 3015 10596 3049
rect 10630 3015 10664 3049
rect 10698 3015 10732 3049
rect 10766 3015 10800 3049
rect 10834 3015 10868 3049
rect 10902 3015 11127 3049
rect 9808 2999 11127 3015
rect 9808 2967 9838 2999
rect 9894 2967 9924 2999
rect 9980 2967 10010 2999
rect 10066 2967 10096 2999
rect 10152 2967 10182 2999
rect 10238 2967 10268 2999
rect 10324 2967 10354 2999
rect 10410 2967 10440 2999
rect 10495 2967 10525 2999
rect 10581 2967 10611 2999
rect 10667 2967 10697 2999
rect 10753 2967 10783 2999
rect 10839 2967 10869 2999
rect 10925 2967 10955 2999
rect 11011 2967 11041 2999
rect 11097 2967 11127 2999
rect 11763 3065 11793 3087
rect 11763 3049 11822 3065
rect 11763 3015 11778 3049
rect 11812 3015 11822 3049
rect 11763 2999 11822 3015
rect 11763 2967 11793 2999
rect 9095 2941 9305 2967
rect 8907 2901 8937 2916
rect 4491 2741 4521 2767
rect 4588 2741 4618 2767
rect 4672 2741 4702 2767
rect 4792 2741 4822 2767
rect 4898 2741 4928 2767
rect 4982 2741 5012 2767
rect 5066 2741 5096 2767
rect 5142 2741 5172 2767
rect 5250 2741 5280 2767
rect 5322 2741 5352 2767
rect 5510 2741 5540 2767
rect 5606 2741 5636 2767
rect 5794 2741 5824 2767
rect 5889 2741 5919 2767
rect 6427 2741 7005 2767
rect 7255 2741 7285 2767
rect 7470 2741 7500 2767
rect 7554 2741 7584 2767
rect 7662 2741 7692 2767
rect 7746 2741 7776 2767
rect 7832 2741 7862 2767
rect 7931 2741 7961 2767
rect 8128 2741 8158 2767
rect 8225 2741 8255 2767
rect 8365 2741 8395 2767
rect 8464 2741 8494 2767
rect 8556 2741 8586 2767
rect 8823 2747 8853 2773
rect 8907 2747 8937 2773
rect 11971 2965 12001 3133
rect 12062 3073 12092 3133
rect 12211 3101 12241 3133
rect 12139 3085 12241 3101
rect 12043 3057 12097 3073
rect 12043 3023 12053 3057
rect 12087 3023 12097 3057
rect 12139 3051 12149 3085
rect 12183 3071 12241 3085
rect 12307 3075 12337 3145
rect 12416 3123 12446 3145
rect 12183 3051 12200 3071
rect 12139 3035 12200 3051
rect 12043 3007 12097 3023
rect 11966 2949 12020 2965
rect 11966 2915 11976 2949
rect 12010 2915 12020 2949
rect 11966 2899 12020 2915
rect 11978 2851 12008 2899
rect 12062 2851 12092 3007
rect 12170 2851 12200 3035
rect 12283 3059 12337 3075
rect 12283 3025 12293 3059
rect 12327 3027 12337 3059
rect 12379 3107 12446 3123
rect 12379 3073 12389 3107
rect 12423 3073 12446 3107
rect 12647 3111 12677 3133
rect 12623 3095 12677 3111
rect 12379 3057 12446 3073
rect 12515 3063 12545 3089
rect 12515 3047 12581 3063
rect 12327 3025 12349 3027
rect 12283 3015 12349 3025
rect 12283 3009 12370 3015
rect 12307 2997 12370 3009
rect 12320 2985 12370 2997
rect 12244 2933 12298 2949
rect 12244 2899 12254 2933
rect 12288 2899 12298 2933
rect 12244 2883 12298 2899
rect 12254 2851 12284 2883
rect 12340 2851 12370 2985
rect 12515 3013 12537 3047
rect 12571 3013 12581 3047
rect 12623 3061 12633 3095
rect 12667 3061 12677 3095
rect 12623 3045 12677 3061
rect 12515 2997 12581 3013
rect 12515 2980 12545 2997
rect 12439 2950 12545 2980
rect 12439 2935 12469 2950
rect 12636 2851 12666 3045
rect 12719 2975 12749 3133
rect 12885 3111 12915 3145
rect 12981 3111 13011 3145
rect 12872 3101 12938 3111
rect 12872 3067 12888 3101
rect 12922 3067 12938 3101
rect 12872 3057 12938 3067
rect 12980 3095 13034 3111
rect 12980 3061 12990 3095
rect 13024 3061 13034 3095
rect 12980 3045 13034 3061
rect 12980 3015 13011 3045
rect 12873 2985 13011 3015
rect 13076 3004 13106 3133
rect 13331 3044 13361 3133
rect 13415 3118 13445 3133
rect 13415 3088 13478 3118
rect 13448 3065 13478 3088
rect 13603 3081 13813 3107
rect 13729 3075 13813 3081
rect 13448 3049 13502 3065
rect 13331 3034 13406 3044
rect 13076 2988 13193 3004
rect 12708 2959 12763 2975
rect 12708 2925 12719 2959
rect 12753 2925 12763 2959
rect 12708 2909 12763 2925
rect 12733 2851 12763 2909
rect 12873 2851 12903 2985
rect 13076 2968 13149 2988
rect 13064 2954 13149 2968
rect 13183 2954 13193 2988
rect 12952 2933 13018 2943
rect 12952 2899 12968 2933
rect 13002 2899 13018 2933
rect 12952 2889 13018 2899
rect 13064 2938 13193 2954
rect 13331 3000 13356 3034
rect 13390 3000 13406 3034
rect 13331 2990 13406 3000
rect 13448 3015 13458 3049
rect 13492 3015 13502 3049
rect 13729 3059 13871 3075
rect 13971 3065 14001 3133
rect 14066 3065 14096 3087
rect 14150 3065 14180 3087
rect 14339 3081 15285 3107
rect 15443 3081 16389 3107
rect 16731 3081 17677 3107
rect 17835 3081 18413 3107
rect 13448 2999 13502 3015
rect 13545 3023 13687 3039
rect 12972 2851 13002 2889
rect 13064 2851 13094 2938
rect 13331 2901 13361 2990
rect 13448 2946 13478 2999
rect 13545 2989 13561 3023
rect 13595 2989 13687 3023
rect 13729 3025 13821 3059
rect 13855 3025 13871 3059
rect 13729 3009 13871 3025
rect 13919 3049 14001 3065
rect 13919 3015 13929 3049
rect 13963 3015 14001 3049
rect 13919 2999 14001 3015
rect 14043 3049 14180 3065
rect 14043 3015 14053 3049
rect 14087 3015 14180 3049
rect 14831 3059 15285 3081
rect 14043 2999 14180 3015
rect 13545 2973 13687 2989
rect 13415 2916 13478 2946
rect 13603 2967 13687 2973
rect 13603 2941 13813 2967
rect 13415 2901 13445 2916
rect 9095 2741 9305 2767
rect 9464 2741 9494 2767
rect 9550 2741 9580 2767
rect 9636 2741 9666 2767
rect 9722 2741 9752 2767
rect 9808 2741 9838 2767
rect 9894 2741 9924 2767
rect 9980 2741 10010 2767
rect 10066 2741 10096 2767
rect 10152 2741 10182 2767
rect 10238 2741 10268 2767
rect 10324 2741 10354 2767
rect 10410 2741 10440 2767
rect 10495 2741 10525 2767
rect 10581 2741 10611 2767
rect 10667 2741 10697 2767
rect 10753 2741 10783 2767
rect 10839 2741 10869 2767
rect 10925 2741 10955 2767
rect 11011 2741 11041 2767
rect 11097 2741 11127 2767
rect 11763 2741 11793 2767
rect 11978 2741 12008 2767
rect 12062 2741 12092 2767
rect 12170 2741 12200 2767
rect 12254 2741 12284 2767
rect 12340 2741 12370 2767
rect 12439 2741 12469 2767
rect 12636 2741 12666 2767
rect 12733 2741 12763 2767
rect 12873 2741 12903 2767
rect 12972 2741 13002 2767
rect 13064 2741 13094 2767
rect 13331 2747 13361 2773
rect 13415 2747 13445 2773
rect 13971 2903 14001 2999
rect 14066 2967 14096 2999
rect 14150 2967 14180 2999
rect 14339 3023 14789 3039
rect 14339 2989 14611 3023
rect 14645 2989 14789 3023
rect 14831 3025 14975 3059
rect 15009 3025 15285 3059
rect 15935 3059 16389 3081
rect 14831 3009 15285 3025
rect 15443 3023 15893 3039
rect 14339 2967 14789 2989
rect 15443 2989 15715 3023
rect 15749 2989 15893 3023
rect 15935 3025 16079 3059
rect 16113 3025 16389 3059
rect 17223 3059 17677 3081
rect 15935 3009 16389 3025
rect 16731 3023 17181 3039
rect 15443 2967 15893 2989
rect 16731 2989 17003 3023
rect 17037 2989 17181 3023
rect 17223 3025 17367 3059
rect 17401 3025 17677 3059
rect 18141 3059 18413 3081
rect 18663 3081 18781 3107
rect 18663 3079 18701 3081
rect 17223 3009 17677 3025
rect 17835 3023 18099 3039
rect 16731 2967 17181 2989
rect 17835 2989 17851 3023
rect 17885 2989 17950 3023
rect 17984 2989 18049 3023
rect 18083 2989 18099 3023
rect 18141 3025 18157 3059
rect 18191 3025 18260 3059
rect 18294 3025 18363 3059
rect 18397 3025 18413 3059
rect 18141 3009 18413 3025
rect 18635 3063 18701 3079
rect 18635 3029 18651 3063
rect 18685 3029 18701 3063
rect 18635 3013 18701 3029
rect 18743 3023 18809 3039
rect 17835 2967 18099 2989
rect 18743 2989 18759 3023
rect 18793 2989 18809 3023
rect 18743 2973 18809 2989
rect 18743 2971 18781 2973
rect 13603 2741 13813 2767
rect 13971 2749 14001 2775
rect 14339 2941 15285 2967
rect 15443 2941 16389 2967
rect 16731 2941 17677 2967
rect 17835 2941 18413 2967
rect 18663 2941 18781 2971
rect 14066 2741 14096 2767
rect 14150 2741 14180 2767
rect 14339 2741 15285 2767
rect 15443 2741 16389 2767
rect 16731 2741 17677 2767
rect 17835 2741 18413 2767
rect 18663 2741 18781 2767
rect 1183 2673 1301 2699
rect 1459 2673 1577 2699
rect 1735 2667 1765 2693
rect 1819 2667 1849 2693
rect 2086 2673 2116 2699
rect 2178 2673 2208 2699
rect 2277 2673 2307 2699
rect 2417 2673 2447 2699
rect 2514 2673 2544 2699
rect 2711 2673 2741 2699
rect 2810 2673 2840 2699
rect 2896 2673 2926 2699
rect 2980 2673 3010 2699
rect 3088 2673 3118 2699
rect 3172 2673 3202 2699
rect 3387 2673 3417 2699
rect 3851 2673 4061 2699
rect 1735 2524 1765 2539
rect 1183 2469 1301 2499
rect 1459 2469 1577 2499
rect 1702 2494 1765 2524
rect 1183 2467 1221 2469
rect 1459 2467 1497 2469
rect 1155 2451 1221 2467
rect 1155 2417 1171 2451
rect 1205 2417 1221 2451
rect 1431 2451 1497 2467
rect 1155 2401 1221 2417
rect 1263 2411 1329 2427
rect 1263 2377 1279 2411
rect 1313 2377 1329 2411
rect 1431 2417 1447 2451
rect 1481 2417 1497 2451
rect 1702 2441 1732 2494
rect 1819 2450 1849 2539
rect 2086 2502 2116 2589
rect 2178 2551 2208 2589
rect 1431 2401 1497 2417
rect 1539 2411 1605 2427
rect 1263 2361 1329 2377
rect 1539 2377 1555 2411
rect 1589 2377 1605 2411
rect 1539 2361 1605 2377
rect 1678 2425 1732 2441
rect 1678 2391 1688 2425
rect 1722 2391 1732 2425
rect 1774 2440 1849 2450
rect 1774 2406 1790 2440
rect 1824 2406 1849 2440
rect 1987 2486 2116 2502
rect 2162 2541 2228 2551
rect 2162 2507 2178 2541
rect 2212 2507 2228 2541
rect 2162 2497 2228 2507
rect 1987 2452 1997 2486
rect 2031 2472 2116 2486
rect 2031 2452 2104 2472
rect 2277 2455 2307 2589
rect 2417 2531 2447 2589
rect 2417 2515 2472 2531
rect 2417 2481 2427 2515
rect 2461 2481 2472 2515
rect 2417 2465 2472 2481
rect 1987 2436 2104 2452
rect 1774 2396 1849 2406
rect 1678 2375 1732 2391
rect 1263 2359 1301 2361
rect 1539 2359 1577 2361
rect 1183 2333 1301 2359
rect 1459 2333 1577 2359
rect 1702 2352 1732 2375
rect 1702 2322 1765 2352
rect 1735 2307 1765 2322
rect 1819 2307 1849 2396
rect 2074 2307 2104 2436
rect 2169 2425 2307 2455
rect 2169 2395 2200 2425
rect 2146 2379 2200 2395
rect 2146 2345 2156 2379
rect 2190 2345 2200 2379
rect 2146 2329 2200 2345
rect 2242 2373 2308 2383
rect 2242 2339 2258 2373
rect 2292 2339 2308 2373
rect 2242 2329 2308 2339
rect 2169 2295 2199 2329
rect 2265 2295 2295 2329
rect 2431 2307 2461 2465
rect 2514 2395 2544 2589
rect 2711 2490 2741 2505
rect 2635 2460 2741 2490
rect 2635 2443 2665 2460
rect 2599 2427 2665 2443
rect 2503 2379 2557 2395
rect 2503 2345 2513 2379
rect 2547 2345 2557 2379
rect 2599 2393 2609 2427
rect 2643 2393 2665 2427
rect 2810 2455 2840 2589
rect 2896 2557 2926 2589
rect 2882 2541 2936 2557
rect 2882 2507 2892 2541
rect 2926 2507 2936 2541
rect 2882 2491 2936 2507
rect 2810 2443 2860 2455
rect 2810 2431 2873 2443
rect 2810 2425 2897 2431
rect 2831 2415 2897 2425
rect 2831 2413 2853 2415
rect 2599 2377 2665 2393
rect 2635 2351 2665 2377
rect 2734 2367 2801 2383
rect 2503 2329 2557 2345
rect 2503 2307 2533 2329
rect 2734 2333 2757 2367
rect 2791 2333 2801 2367
rect 2734 2317 2801 2333
rect 2843 2381 2853 2413
rect 2887 2381 2897 2415
rect 2843 2365 2897 2381
rect 2980 2405 3010 2589
rect 3088 2433 3118 2589
rect 3172 2541 3202 2589
rect 3160 2525 3214 2541
rect 3160 2491 3170 2525
rect 3204 2491 3214 2525
rect 3160 2475 3214 2491
rect 3083 2417 3137 2433
rect 2980 2389 3041 2405
rect 2980 2369 2997 2389
rect 2734 2295 2764 2317
rect 2843 2295 2873 2365
rect 2939 2355 2997 2369
rect 3031 2355 3041 2389
rect 3083 2383 3093 2417
rect 3127 2383 3137 2417
rect 3083 2367 3137 2383
rect 2939 2339 3041 2355
rect 2939 2307 2969 2339
rect 3088 2307 3118 2367
rect 3179 2307 3209 2475
rect 4311 2667 4341 2693
rect 4395 2667 4425 2693
rect 4662 2673 4692 2699
rect 4754 2673 4784 2699
rect 4853 2673 4883 2699
rect 4993 2673 5023 2699
rect 5090 2673 5120 2699
rect 5287 2673 5317 2699
rect 5386 2673 5416 2699
rect 5472 2673 5502 2699
rect 5556 2673 5586 2699
rect 5664 2673 5694 2699
rect 5748 2673 5778 2699
rect 5963 2673 5993 2699
rect 6427 2673 7373 2699
rect 7531 2673 8477 2699
rect 8635 2673 8753 2699
rect 9187 2673 9217 2699
rect 9402 2673 9432 2699
rect 9486 2673 9516 2699
rect 9594 2673 9624 2699
rect 9678 2673 9708 2699
rect 9764 2673 9794 2699
rect 9863 2673 9893 2699
rect 10060 2673 10090 2699
rect 10157 2673 10187 2699
rect 10297 2673 10327 2699
rect 10396 2673 10426 2699
rect 10488 2673 10518 2699
rect 4311 2524 4341 2539
rect 3851 2473 4061 2499
rect 4278 2494 4341 2524
rect 3387 2441 3417 2473
rect 3851 2467 3935 2473
rect 3358 2425 3417 2441
rect 3358 2391 3368 2425
rect 3402 2391 3417 2425
rect 3793 2451 3935 2467
rect 3793 2417 3809 2451
rect 3843 2417 3935 2451
rect 4278 2441 4308 2494
rect 4395 2450 4425 2539
rect 4662 2502 4692 2589
rect 4754 2551 4784 2589
rect 3793 2401 3935 2417
rect 3977 2415 4119 2431
rect 3358 2375 3417 2391
rect 3387 2353 3417 2375
rect 3977 2381 4069 2415
rect 4103 2381 4119 2415
rect 3977 2365 4119 2381
rect 4254 2425 4308 2441
rect 4254 2391 4264 2425
rect 4298 2391 4308 2425
rect 4350 2440 4425 2450
rect 4350 2406 4366 2440
rect 4400 2406 4425 2440
rect 4563 2486 4692 2502
rect 4738 2541 4804 2551
rect 4738 2507 4754 2541
rect 4788 2507 4804 2541
rect 4738 2497 4804 2507
rect 4563 2452 4573 2486
rect 4607 2472 4692 2486
rect 4607 2452 4680 2472
rect 4853 2455 4883 2589
rect 4993 2531 5023 2589
rect 4993 2515 5048 2531
rect 4993 2481 5003 2515
rect 5037 2481 5048 2515
rect 4993 2465 5048 2481
rect 4563 2436 4680 2452
rect 4350 2396 4425 2406
rect 4254 2375 4308 2391
rect 3977 2359 4061 2365
rect 3851 2333 4061 2359
rect 4278 2352 4308 2375
rect 4278 2322 4341 2352
rect 4311 2307 4341 2322
rect 4395 2307 4425 2396
rect 4650 2307 4680 2436
rect 4745 2425 4883 2455
rect 4745 2395 4776 2425
rect 4722 2379 4776 2395
rect 4722 2345 4732 2379
rect 4766 2345 4776 2379
rect 4722 2329 4776 2345
rect 4818 2373 4884 2383
rect 4818 2339 4834 2373
rect 4868 2339 4884 2373
rect 4818 2329 4884 2339
rect 4745 2295 4775 2329
rect 4841 2295 4871 2329
rect 5007 2307 5037 2465
rect 5090 2395 5120 2589
rect 5287 2490 5317 2505
rect 5211 2460 5317 2490
rect 5211 2443 5241 2460
rect 5175 2427 5241 2443
rect 5079 2379 5133 2395
rect 5079 2345 5089 2379
rect 5123 2345 5133 2379
rect 5175 2393 5185 2427
rect 5219 2393 5241 2427
rect 5386 2455 5416 2589
rect 5472 2557 5502 2589
rect 5458 2541 5512 2557
rect 5458 2507 5468 2541
rect 5502 2507 5512 2541
rect 5458 2491 5512 2507
rect 5386 2443 5436 2455
rect 5386 2431 5449 2443
rect 5386 2425 5473 2431
rect 5407 2415 5473 2425
rect 5407 2413 5429 2415
rect 5175 2377 5241 2393
rect 5211 2351 5241 2377
rect 5310 2367 5377 2383
rect 5079 2329 5133 2345
rect 5079 2307 5109 2329
rect 5310 2333 5333 2367
rect 5367 2333 5377 2367
rect 5310 2317 5377 2333
rect 5419 2381 5429 2413
rect 5463 2381 5473 2415
rect 5419 2365 5473 2381
rect 5556 2405 5586 2589
rect 5664 2433 5694 2589
rect 5748 2541 5778 2589
rect 5736 2525 5790 2541
rect 5736 2491 5746 2525
rect 5780 2491 5790 2525
rect 5736 2475 5790 2491
rect 5659 2417 5713 2433
rect 5556 2389 5617 2405
rect 5556 2369 5573 2389
rect 5310 2295 5340 2317
rect 5419 2295 5449 2365
rect 5515 2355 5573 2369
rect 5607 2355 5617 2389
rect 5659 2383 5669 2417
rect 5703 2383 5713 2417
rect 5659 2367 5713 2383
rect 5515 2339 5617 2355
rect 5515 2307 5545 2339
rect 5664 2307 5694 2367
rect 5755 2307 5785 2475
rect 6427 2473 7373 2499
rect 7531 2473 8477 2499
rect 5963 2441 5993 2473
rect 5934 2425 5993 2441
rect 5934 2391 5944 2425
rect 5978 2391 5993 2425
rect 6427 2451 6877 2473
rect 6427 2417 6699 2451
rect 6733 2417 6877 2451
rect 7531 2451 7981 2473
rect 8635 2469 8753 2499
rect 9402 2541 9432 2589
rect 9390 2525 9444 2541
rect 9390 2491 9400 2525
rect 9434 2491 9444 2525
rect 9390 2475 9444 2491
rect 8635 2467 8673 2469
rect 6427 2401 6877 2417
rect 6919 2415 7373 2431
rect 5934 2375 5993 2391
rect 5963 2353 5993 2375
rect 6919 2381 7063 2415
rect 7097 2381 7373 2415
rect 7531 2417 7803 2451
rect 7837 2417 7981 2451
rect 8607 2451 8673 2467
rect 7531 2401 7981 2417
rect 8023 2415 8477 2431
rect 6919 2359 7373 2381
rect 8023 2381 8167 2415
rect 8201 2381 8477 2415
rect 8607 2417 8623 2451
rect 8657 2417 8673 2451
rect 9187 2441 9217 2473
rect 8607 2401 8673 2417
rect 8715 2411 8781 2427
rect 8023 2359 8477 2381
rect 8715 2377 8731 2411
rect 8765 2377 8781 2411
rect 8715 2361 8781 2377
rect 9187 2425 9246 2441
rect 9187 2391 9202 2425
rect 9236 2391 9246 2425
rect 9187 2375 9246 2391
rect 8715 2359 8753 2361
rect 6427 2333 7373 2359
rect 7531 2333 8477 2359
rect 8635 2333 8753 2359
rect 9187 2353 9217 2375
rect 9395 2307 9425 2475
rect 9486 2433 9516 2589
rect 9467 2417 9521 2433
rect 9467 2383 9477 2417
rect 9511 2383 9521 2417
rect 9594 2405 9624 2589
rect 9678 2557 9708 2589
rect 9668 2541 9722 2557
rect 9668 2507 9678 2541
rect 9712 2507 9722 2541
rect 9668 2491 9722 2507
rect 9764 2455 9794 2589
rect 10755 2667 10785 2693
rect 10839 2667 10869 2693
rect 11027 2673 11237 2699
rect 11579 2673 11789 2699
rect 12039 2673 12069 2699
rect 12254 2673 12284 2699
rect 12338 2673 12368 2699
rect 12446 2673 12476 2699
rect 12530 2673 12560 2699
rect 12616 2673 12646 2699
rect 12715 2673 12745 2699
rect 12912 2673 12942 2699
rect 13009 2673 13039 2699
rect 13149 2673 13179 2699
rect 13248 2673 13278 2699
rect 13340 2673 13370 2699
rect 9863 2490 9893 2505
rect 9863 2460 9969 2490
rect 9744 2443 9794 2455
rect 9731 2431 9794 2443
rect 9467 2367 9521 2383
rect 9563 2389 9624 2405
rect 9486 2307 9516 2367
rect 9563 2355 9573 2389
rect 9607 2369 9624 2389
rect 9707 2425 9794 2431
rect 9939 2443 9969 2460
rect 9939 2427 10005 2443
rect 9707 2415 9773 2425
rect 9707 2381 9717 2415
rect 9751 2413 9773 2415
rect 9751 2381 9761 2413
rect 9939 2393 9961 2427
rect 9995 2393 10005 2427
rect 10060 2395 10090 2589
rect 10157 2531 10187 2589
rect 10132 2515 10187 2531
rect 10132 2481 10143 2515
rect 10177 2481 10187 2515
rect 10132 2465 10187 2481
rect 9607 2355 9665 2369
rect 9707 2365 9761 2381
rect 9563 2339 9665 2355
rect 9635 2307 9665 2339
rect 9731 2295 9761 2365
rect 9803 2367 9870 2383
rect 9803 2333 9813 2367
rect 9847 2333 9870 2367
rect 9939 2377 10005 2393
rect 10047 2379 10101 2395
rect 9939 2351 9969 2377
rect 9803 2317 9870 2333
rect 9840 2295 9870 2317
rect 10047 2345 10057 2379
rect 10091 2345 10101 2379
rect 10047 2329 10101 2345
rect 10071 2307 10101 2329
rect 10143 2307 10173 2465
rect 10297 2455 10327 2589
rect 10396 2551 10426 2589
rect 10376 2541 10442 2551
rect 10376 2507 10392 2541
rect 10426 2507 10442 2541
rect 10376 2497 10442 2507
rect 10488 2502 10518 2589
rect 10488 2486 10617 2502
rect 10488 2472 10573 2486
rect 10297 2425 10435 2455
rect 10404 2395 10435 2425
rect 10500 2452 10573 2472
rect 10607 2452 10617 2486
rect 10500 2436 10617 2452
rect 10755 2450 10785 2539
rect 10839 2524 10869 2539
rect 10839 2494 10902 2524
rect 10755 2440 10830 2450
rect 10296 2373 10362 2383
rect 10296 2339 10312 2373
rect 10346 2339 10362 2373
rect 10296 2329 10362 2339
rect 10404 2379 10458 2395
rect 10404 2345 10414 2379
rect 10448 2345 10458 2379
rect 10404 2329 10458 2345
rect 10309 2295 10339 2329
rect 10405 2295 10435 2329
rect 10500 2307 10530 2436
rect 10755 2406 10780 2440
rect 10814 2406 10830 2440
rect 10755 2396 10830 2406
rect 10872 2441 10902 2494
rect 11027 2473 11237 2499
rect 11579 2473 11789 2499
rect 12254 2541 12284 2589
rect 12242 2525 12296 2541
rect 12242 2491 12252 2525
rect 12286 2491 12296 2525
rect 12242 2475 12296 2491
rect 11027 2467 11111 2473
rect 11579 2467 11663 2473
rect 10969 2451 11111 2467
rect 10872 2425 10926 2441
rect 10755 2307 10785 2396
rect 10872 2391 10882 2425
rect 10916 2391 10926 2425
rect 10969 2417 10985 2451
rect 11019 2417 11111 2451
rect 11521 2451 11663 2467
rect 10969 2401 11111 2417
rect 11153 2415 11295 2431
rect 10872 2375 10926 2391
rect 11153 2381 11245 2415
rect 11279 2381 11295 2415
rect 11521 2417 11537 2451
rect 11571 2417 11663 2451
rect 12039 2441 12069 2473
rect 11521 2401 11663 2417
rect 11705 2415 11847 2431
rect 10872 2352 10902 2375
rect 11153 2365 11295 2381
rect 11705 2381 11797 2415
rect 11831 2381 11847 2415
rect 11705 2365 11847 2381
rect 12039 2425 12098 2441
rect 12039 2391 12054 2425
rect 12088 2391 12098 2425
rect 12039 2375 12098 2391
rect 11153 2359 11237 2365
rect 11705 2359 11789 2365
rect 10839 2322 10902 2352
rect 11027 2333 11237 2359
rect 10839 2307 10869 2322
rect 11579 2333 11789 2359
rect 12039 2353 12069 2375
rect 12247 2307 12277 2475
rect 12338 2433 12368 2589
rect 12319 2417 12373 2433
rect 12319 2383 12329 2417
rect 12363 2383 12373 2417
rect 12446 2405 12476 2589
rect 12530 2557 12560 2589
rect 12520 2541 12574 2557
rect 12520 2507 12530 2541
rect 12564 2507 12574 2541
rect 12520 2491 12574 2507
rect 12616 2455 12646 2589
rect 13607 2667 13637 2693
rect 13691 2667 13721 2693
rect 14339 2673 14369 2699
rect 14554 2673 14584 2699
rect 14638 2673 14668 2699
rect 14746 2673 14776 2699
rect 14830 2673 14860 2699
rect 14916 2673 14946 2699
rect 15015 2673 15045 2699
rect 15212 2673 15242 2699
rect 15309 2673 15339 2699
rect 15449 2673 15479 2699
rect 15548 2673 15578 2699
rect 15640 2673 15670 2699
rect 12715 2490 12745 2505
rect 12715 2460 12821 2490
rect 12596 2443 12646 2455
rect 12583 2431 12646 2443
rect 12319 2367 12373 2383
rect 12415 2389 12476 2405
rect 12338 2307 12368 2367
rect 12415 2355 12425 2389
rect 12459 2369 12476 2389
rect 12559 2425 12646 2431
rect 12791 2443 12821 2460
rect 12791 2427 12857 2443
rect 12559 2415 12625 2425
rect 12559 2381 12569 2415
rect 12603 2413 12625 2415
rect 12603 2381 12613 2413
rect 12791 2393 12813 2427
rect 12847 2393 12857 2427
rect 12912 2395 12942 2589
rect 13009 2531 13039 2589
rect 12984 2515 13039 2531
rect 12984 2481 12995 2515
rect 13029 2481 13039 2515
rect 12984 2465 13039 2481
rect 12459 2355 12517 2369
rect 12559 2365 12613 2381
rect 12415 2339 12517 2355
rect 12487 2307 12517 2339
rect 12583 2295 12613 2365
rect 12655 2367 12722 2383
rect 12655 2333 12665 2367
rect 12699 2333 12722 2367
rect 12791 2377 12857 2393
rect 12899 2379 12953 2395
rect 12791 2351 12821 2377
rect 12655 2317 12722 2333
rect 12692 2295 12722 2317
rect 12899 2345 12909 2379
rect 12943 2345 12953 2379
rect 12899 2329 12953 2345
rect 12923 2307 12953 2329
rect 12995 2307 13025 2465
rect 13149 2455 13179 2589
rect 13248 2551 13278 2589
rect 13228 2541 13294 2551
rect 13228 2507 13244 2541
rect 13278 2507 13294 2541
rect 13228 2497 13294 2507
rect 13340 2502 13370 2589
rect 13340 2486 13469 2502
rect 13340 2472 13425 2486
rect 13149 2425 13287 2455
rect 13256 2395 13287 2425
rect 13352 2452 13425 2472
rect 13459 2452 13469 2486
rect 13352 2436 13469 2452
rect 13607 2450 13637 2539
rect 13691 2524 13721 2539
rect 13691 2494 13754 2524
rect 13607 2440 13682 2450
rect 13148 2373 13214 2383
rect 13148 2339 13164 2373
rect 13198 2339 13214 2373
rect 13148 2329 13214 2339
rect 13256 2379 13310 2395
rect 13256 2345 13266 2379
rect 13300 2345 13310 2379
rect 13256 2329 13310 2345
rect 13161 2295 13191 2329
rect 13257 2295 13287 2329
rect 13352 2307 13382 2436
rect 13607 2406 13632 2440
rect 13666 2406 13682 2440
rect 13607 2396 13682 2406
rect 13724 2441 13754 2494
rect 14554 2541 14584 2589
rect 14542 2525 14596 2541
rect 14542 2491 14552 2525
rect 14586 2491 14596 2525
rect 14542 2475 14596 2491
rect 14339 2441 14369 2473
rect 13724 2425 13778 2441
rect 13607 2307 13637 2396
rect 13724 2391 13734 2425
rect 13768 2391 13778 2425
rect 13724 2375 13778 2391
rect 14339 2425 14398 2441
rect 14339 2391 14354 2425
rect 14388 2391 14398 2425
rect 14339 2375 14398 2391
rect 13724 2352 13754 2375
rect 14339 2353 14369 2375
rect 13691 2322 13754 2352
rect 13691 2307 13721 2322
rect 14547 2307 14577 2475
rect 14638 2433 14668 2589
rect 14619 2417 14673 2433
rect 14619 2383 14629 2417
rect 14663 2383 14673 2417
rect 14746 2405 14776 2589
rect 14830 2557 14860 2589
rect 14820 2541 14874 2557
rect 14820 2507 14830 2541
rect 14864 2507 14874 2541
rect 14820 2491 14874 2507
rect 14916 2455 14946 2589
rect 15907 2667 15937 2693
rect 15991 2667 16021 2693
rect 16179 2673 16389 2699
rect 16731 2673 17309 2699
rect 15015 2490 15045 2505
rect 15015 2460 15121 2490
rect 14896 2443 14946 2455
rect 14883 2431 14946 2443
rect 14619 2367 14673 2383
rect 14715 2389 14776 2405
rect 14638 2307 14668 2367
rect 14715 2355 14725 2389
rect 14759 2369 14776 2389
rect 14859 2425 14946 2431
rect 15091 2443 15121 2460
rect 15091 2427 15157 2443
rect 14859 2415 14925 2425
rect 14859 2381 14869 2415
rect 14903 2413 14925 2415
rect 14903 2381 14913 2413
rect 15091 2393 15113 2427
rect 15147 2393 15157 2427
rect 15212 2395 15242 2589
rect 15309 2531 15339 2589
rect 15284 2515 15339 2531
rect 15284 2481 15295 2515
rect 15329 2481 15339 2515
rect 15284 2465 15339 2481
rect 14759 2355 14817 2369
rect 14859 2365 14913 2381
rect 14715 2339 14817 2355
rect 14787 2307 14817 2339
rect 14883 2295 14913 2365
rect 14955 2367 15022 2383
rect 14955 2333 14965 2367
rect 14999 2333 15022 2367
rect 15091 2377 15157 2393
rect 15199 2379 15253 2395
rect 15091 2351 15121 2377
rect 14955 2317 15022 2333
rect 14992 2295 15022 2317
rect 15199 2345 15209 2379
rect 15243 2345 15253 2379
rect 15199 2329 15253 2345
rect 15223 2307 15253 2329
rect 15295 2307 15325 2465
rect 15449 2455 15479 2589
rect 15548 2551 15578 2589
rect 15528 2541 15594 2551
rect 15528 2507 15544 2541
rect 15578 2507 15594 2541
rect 15528 2497 15594 2507
rect 15640 2502 15670 2589
rect 15640 2486 15769 2502
rect 15640 2472 15725 2486
rect 15449 2425 15587 2455
rect 15556 2395 15587 2425
rect 15652 2452 15725 2472
rect 15759 2452 15769 2486
rect 15652 2436 15769 2452
rect 15907 2450 15937 2539
rect 15991 2524 16021 2539
rect 15991 2494 16054 2524
rect 15907 2440 15982 2450
rect 15448 2373 15514 2383
rect 15448 2339 15464 2373
rect 15498 2339 15514 2373
rect 15448 2329 15514 2339
rect 15556 2379 15610 2395
rect 15556 2345 15566 2379
rect 15600 2345 15610 2379
rect 15556 2329 15610 2345
rect 15461 2295 15491 2329
rect 15557 2295 15587 2329
rect 15652 2307 15682 2436
rect 15907 2406 15932 2440
rect 15966 2406 15982 2440
rect 15907 2396 15982 2406
rect 16024 2441 16054 2494
rect 16179 2473 16389 2499
rect 17559 2665 17589 2691
rect 17654 2673 17684 2699
rect 17738 2673 17768 2699
rect 17927 2673 18505 2699
rect 18663 2673 18781 2699
rect 16731 2473 17309 2499
rect 16179 2467 16263 2473
rect 16121 2451 16263 2467
rect 16024 2425 16078 2441
rect 15907 2307 15937 2396
rect 16024 2391 16034 2425
rect 16068 2391 16078 2425
rect 16121 2417 16137 2451
rect 16171 2417 16263 2451
rect 16731 2451 16995 2473
rect 16121 2401 16263 2417
rect 16305 2415 16447 2431
rect 16024 2375 16078 2391
rect 16305 2381 16397 2415
rect 16431 2381 16447 2415
rect 16731 2417 16747 2451
rect 16781 2417 16846 2451
rect 16880 2417 16945 2451
rect 16979 2417 16995 2451
rect 17559 2441 17589 2537
rect 17927 2473 18505 2499
rect 17654 2441 17684 2473
rect 17738 2441 17768 2473
rect 16731 2401 16995 2417
rect 17037 2415 17309 2431
rect 16024 2352 16054 2375
rect 16305 2365 16447 2381
rect 17037 2381 17053 2415
rect 17087 2381 17156 2415
rect 17190 2381 17259 2415
rect 17293 2381 17309 2415
rect 16305 2359 16389 2365
rect 17037 2359 17309 2381
rect 17507 2425 17589 2441
rect 17507 2391 17517 2425
rect 17551 2391 17589 2425
rect 17507 2375 17589 2391
rect 17631 2425 17768 2441
rect 17631 2391 17641 2425
rect 17675 2391 17768 2425
rect 17927 2451 18191 2473
rect 18663 2469 18781 2499
rect 17927 2417 17943 2451
rect 17977 2417 18042 2451
rect 18076 2417 18141 2451
rect 18175 2417 18191 2451
rect 18743 2467 18781 2469
rect 18743 2451 18809 2467
rect 17927 2401 18191 2417
rect 18233 2415 18505 2431
rect 17631 2375 17768 2391
rect 15991 2322 16054 2352
rect 16179 2333 16389 2359
rect 15991 2307 16021 2322
rect 16731 2333 17309 2359
rect 17559 2307 17589 2375
rect 17654 2353 17684 2375
rect 17738 2353 17768 2375
rect 18233 2381 18249 2415
rect 18283 2381 18352 2415
rect 18386 2381 18455 2415
rect 18489 2381 18505 2415
rect 18233 2359 18505 2381
rect 18635 2411 18701 2427
rect 18635 2377 18651 2411
rect 18685 2377 18701 2411
rect 18743 2417 18759 2451
rect 18793 2417 18809 2451
rect 18743 2401 18809 2417
rect 18635 2361 18701 2377
rect 17927 2333 18505 2359
rect 18663 2359 18701 2361
rect 18663 2333 18781 2359
rect 1183 2197 1301 2223
rect 1459 2197 1577 2223
rect 1735 2197 1765 2223
rect 1819 2197 1849 2223
rect 2074 2197 2104 2223
rect 2169 2197 2199 2223
rect 2265 2197 2295 2223
rect 2431 2197 2461 2223
rect 2503 2197 2533 2223
rect 2635 2197 2665 2223
rect 2734 2197 2764 2223
rect 2843 2197 2873 2223
rect 2939 2197 2969 2223
rect 3088 2197 3118 2223
rect 3179 2197 3209 2223
rect 3387 2197 3417 2223
rect 3851 2197 4061 2223
rect 4311 2197 4341 2223
rect 4395 2197 4425 2223
rect 4650 2197 4680 2223
rect 4745 2197 4775 2223
rect 4841 2197 4871 2223
rect 5007 2197 5037 2223
rect 5079 2197 5109 2223
rect 5211 2197 5241 2223
rect 5310 2197 5340 2223
rect 5419 2197 5449 2223
rect 5515 2197 5545 2223
rect 5664 2197 5694 2223
rect 5755 2197 5785 2223
rect 5963 2197 5993 2223
rect 6427 2197 7373 2223
rect 7531 2197 8477 2223
rect 8635 2197 8753 2223
rect 9187 2197 9217 2223
rect 9395 2197 9425 2223
rect 9486 2197 9516 2223
rect 9635 2197 9665 2223
rect 9731 2197 9761 2223
rect 9840 2197 9870 2223
rect 9939 2197 9969 2223
rect 10071 2197 10101 2223
rect 10143 2197 10173 2223
rect 10309 2197 10339 2223
rect 10405 2197 10435 2223
rect 10500 2197 10530 2223
rect 10755 2197 10785 2223
rect 10839 2197 10869 2223
rect 11027 2197 11237 2223
rect 11579 2197 11789 2223
rect 12039 2197 12069 2223
rect 12247 2197 12277 2223
rect 12338 2197 12368 2223
rect 12487 2197 12517 2223
rect 12583 2197 12613 2223
rect 12692 2197 12722 2223
rect 12791 2197 12821 2223
rect 12923 2197 12953 2223
rect 12995 2197 13025 2223
rect 13161 2197 13191 2223
rect 13257 2197 13287 2223
rect 13352 2197 13382 2223
rect 13607 2197 13637 2223
rect 13691 2197 13721 2223
rect 14339 2197 14369 2223
rect 14547 2197 14577 2223
rect 14638 2197 14668 2223
rect 14787 2197 14817 2223
rect 14883 2197 14913 2223
rect 14992 2197 15022 2223
rect 15091 2197 15121 2223
rect 15223 2197 15253 2223
rect 15295 2197 15325 2223
rect 15461 2197 15491 2223
rect 15557 2197 15587 2223
rect 15652 2197 15682 2223
rect 15907 2197 15937 2223
rect 15991 2197 16021 2223
rect 16179 2197 16389 2223
rect 16731 2197 17309 2223
rect 17559 2197 17589 2223
rect 17654 2197 17684 2223
rect 17738 2197 17768 2223
rect 17927 2197 18505 2223
rect 18663 2197 18781 2223
<< polycont >>
rect 1171 7341 1205 7375
rect 1279 7381 1313 7415
rect 1737 7367 1771 7401
rect 1861 7367 1895 7401
rect 2283 7341 2317 7375
rect 2647 7377 2681 7411
rect 3131 7341 3165 7375
rect 3241 7341 3275 7375
rect 3349 7377 3383 7411
rect 3459 7377 3493 7411
rect 4129 7367 4163 7401
rect 4253 7367 4287 7401
rect 4675 7341 4709 7375
rect 5039 7377 5073 7411
rect 5785 7367 5819 7401
rect 5909 7367 5943 7401
rect 6047 7341 6081 7375
rect 6155 7381 6189 7415
rect 6699 7341 6733 7375
rect 7063 7377 7097 7411
rect 7489 7341 7523 7375
rect 7749 7377 7783 7411
rect 7993 7367 8027 7401
rect 8117 7367 8151 7401
rect 8283 7341 8317 7375
rect 8393 7341 8427 7375
rect 8501 7377 8535 7411
rect 8611 7377 8645 7411
rect 9019 7341 9053 7375
rect 9129 7341 9163 7375
rect 9237 7377 9271 7411
rect 9347 7377 9381 7411
rect 9697 7341 9731 7375
rect 9957 7377 9991 7411
rect 10117 7367 10151 7401
rect 10221 7367 10255 7401
rect 10491 7341 10525 7375
rect 10590 7341 10624 7375
rect 10689 7341 10723 7375
rect 10797 7377 10831 7411
rect 10900 7377 10934 7411
rect 11003 7377 11037 7411
rect 11199 7341 11233 7375
rect 11307 7381 11341 7415
rect 11595 7341 11629 7375
rect 11694 7341 11728 7375
rect 11793 7341 11827 7375
rect 11901 7377 11935 7411
rect 12004 7377 12038 7411
rect 12107 7377 12141 7411
rect 12273 7367 12307 7401
rect 12397 7367 12431 7401
rect 12955 7341 12989 7375
rect 13319 7377 13353 7411
rect 13775 7341 13809 7375
rect 13883 7381 13917 7415
rect 14113 7341 14147 7375
rect 14373 7377 14407 7411
rect 14481 7367 14515 7401
rect 14605 7367 14639 7401
rect 15163 7341 15197 7375
rect 15527 7377 15561 7411
rect 16011 7341 16045 7375
rect 16121 7341 16155 7375
rect 16229 7377 16263 7411
rect 16339 7377 16373 7411
rect 16873 7367 16907 7401
rect 16997 7367 17031 7401
rect 17299 7341 17333 7375
rect 17398 7341 17432 7375
rect 17497 7341 17531 7375
rect 17605 7377 17639 7411
rect 17708 7377 17742 7411
rect 17811 7377 17845 7411
rect 18069 7367 18103 7401
rect 18193 7367 18227 7401
rect 18651 7381 18685 7415
rect 18759 7341 18793 7375
rect 1171 6769 1205 6803
rect 1279 6729 1313 6763
rect 1731 6769 1765 6803
rect 2095 6733 2129 6767
rect 2835 6769 2869 6803
rect 3199 6733 3233 6767
rect 4123 6769 4157 6803
rect 4487 6733 4521 6767
rect 5227 6769 5261 6803
rect 5591 6733 5625 6767
rect 6331 6769 6365 6803
rect 6695 6733 6729 6767
rect 7435 6769 7469 6803
rect 7799 6733 7833 6767
rect 8283 6769 8317 6803
rect 8393 6769 8427 6803
rect 8501 6733 8535 6767
rect 8611 6733 8645 6767
rect 9275 6769 9309 6803
rect 9639 6733 9673 6767
rect 10379 6769 10413 6803
rect 10743 6733 10777 6767
rect 11483 6769 11517 6803
rect 11847 6733 11881 6767
rect 12587 6769 12621 6803
rect 12951 6733 12985 6767
rect 13435 6769 13469 6803
rect 13545 6769 13579 6803
rect 13653 6733 13687 6767
rect 13763 6733 13797 6767
rect 14427 6769 14461 6803
rect 14791 6733 14825 6767
rect 15531 6769 15565 6803
rect 15895 6733 15929 6767
rect 16635 6769 16669 6803
rect 16999 6733 17033 6767
rect 17739 6769 17773 6803
rect 18103 6733 18137 6767
rect 18651 6729 18685 6763
rect 18759 6769 18793 6803
rect 1171 6253 1205 6287
rect 1279 6293 1313 6327
rect 1731 6253 1765 6287
rect 2095 6289 2129 6323
rect 2835 6253 2869 6287
rect 3199 6289 3233 6323
rect 3939 6253 3973 6287
rect 4303 6289 4337 6323
rect 5043 6253 5077 6287
rect 5407 6289 5441 6323
rect 5833 6253 5867 6287
rect 6093 6289 6127 6323
rect 6699 6253 6733 6287
rect 7063 6289 7097 6323
rect 7547 6253 7581 6287
rect 7657 6253 7691 6287
rect 7765 6289 7799 6323
rect 7875 6289 7909 6323
rect 8070 6279 8104 6313
rect 8206 6279 8240 6313
rect 8309 6279 8343 6313
rect 8815 6253 8849 6287
rect 9179 6289 9213 6323
rect 9919 6253 9953 6287
rect 10283 6289 10317 6323
rect 10767 6253 10801 6287
rect 10866 6253 10900 6287
rect 10965 6253 10999 6287
rect 11073 6289 11107 6323
rect 11176 6289 11210 6323
rect 11279 6289 11313 6323
rect 11851 6253 11885 6287
rect 12215 6289 12249 6323
rect 12955 6253 12989 6287
rect 13319 6289 13353 6323
rect 14059 6253 14093 6287
rect 14423 6289 14457 6323
rect 15163 6253 15197 6287
rect 15527 6289 15561 6323
rect 16011 6253 16045 6287
rect 16121 6253 16155 6287
rect 16229 6289 16263 6323
rect 16339 6289 16373 6323
rect 17003 6253 17037 6287
rect 17367 6289 17401 6323
rect 17851 6253 17885 6287
rect 17950 6253 17984 6287
rect 18049 6253 18083 6287
rect 18157 6289 18191 6323
rect 18260 6289 18294 6323
rect 18363 6289 18397 6323
rect 18651 6293 18685 6327
rect 18759 6253 18793 6287
rect 1171 5681 1205 5715
rect 1279 5641 1313 5675
rect 1731 5681 1765 5715
rect 2095 5645 2129 5679
rect 2835 5681 2869 5715
rect 3199 5645 3233 5679
rect 4123 5681 4157 5715
rect 4487 5645 4521 5679
rect 5227 5681 5261 5715
rect 5591 5645 5625 5679
rect 6075 5681 6109 5715
rect 6174 5681 6208 5715
rect 6273 5681 6307 5715
rect 6381 5645 6415 5679
rect 6484 5645 6518 5679
rect 6587 5645 6621 5679
rect 6801 5668 6835 5702
rect 6921 5655 6955 5689
rect 7087 5681 7121 5715
rect 7197 5681 7231 5715
rect 7679 5732 7713 5766
rect 7305 5645 7339 5679
rect 7415 5645 7449 5679
rect 7847 5732 7881 5766
rect 7757 5619 7791 5653
rect 7919 5619 7953 5653
rect 8015 5619 8049 5653
rect 8156 5655 8190 5689
rect 8252 5655 8286 5689
rect 8409 5681 8443 5715
rect 8669 5645 8703 5679
rect 9275 5681 9309 5715
rect 9639 5645 9673 5679
rect 10379 5681 10413 5715
rect 10743 5645 10777 5679
rect 11169 5681 11203 5715
rect 11429 5645 11463 5679
rect 11566 5655 11600 5689
rect 11702 5655 11736 5689
rect 11805 5655 11839 5689
rect 12055 5681 12089 5715
rect 12154 5681 12188 5715
rect 12253 5681 12287 5715
rect 12361 5645 12395 5679
rect 12464 5645 12498 5679
rect 12567 5645 12601 5679
rect 12854 5655 12888 5689
rect 12990 5655 13024 5689
rect 13093 5655 13127 5689
rect 13343 5681 13377 5715
rect 13442 5681 13476 5715
rect 13541 5681 13575 5715
rect 13649 5645 13683 5679
rect 13752 5645 13786 5679
rect 13855 5645 13889 5679
rect 14427 5681 14461 5715
rect 14791 5645 14825 5679
rect 15531 5681 15565 5715
rect 15895 5645 15929 5679
rect 16635 5681 16669 5715
rect 16999 5645 17033 5679
rect 17739 5681 17773 5715
rect 18103 5645 18137 5679
rect 18651 5641 18685 5675
rect 18759 5681 18793 5715
rect 1171 5165 1205 5199
rect 1279 5205 1313 5239
rect 1731 5165 1765 5199
rect 2095 5201 2129 5235
rect 2551 5165 2585 5199
rect 2659 5205 2693 5239
rect 2792 5191 2826 5225
rect 2894 5176 2928 5210
rect 3260 5237 3294 5271
rect 3362 5243 3396 5277
rect 3101 5130 3135 5164
rect 3282 5075 3316 5109
rect 3617 5237 3651 5271
rect 3861 5249 3895 5283
rect 3531 5101 3565 5135
rect 3713 5189 3747 5223
rect 3957 5201 3991 5235
rect 4101 5227 4135 5261
rect 3996 5075 4030 5109
rect 4197 5199 4231 5233
rect 4472 5191 4506 5225
rect 4951 5165 4985 5199
rect 5315 5201 5349 5235
rect 5799 5165 5833 5199
rect 5909 5165 5943 5199
rect 6017 5201 6051 5235
rect 6127 5201 6161 5235
rect 6415 5165 6449 5199
rect 6523 5205 6557 5239
rect 6710 5191 6744 5225
rect 6806 5191 6840 5225
rect 6947 5227 6981 5261
rect 7043 5227 7077 5261
rect 7205 5227 7239 5261
rect 4274 5091 4308 5125
rect 7115 5114 7149 5148
rect 7489 5165 7523 5199
rect 7749 5201 7783 5235
rect 7852 5191 7886 5225
rect 7283 5114 7317 5148
rect 7954 5176 7988 5210
rect 8320 5237 8354 5271
rect 8422 5243 8456 5277
rect 8161 5130 8195 5164
rect 8342 5075 8376 5109
rect 8677 5237 8711 5271
rect 8921 5249 8955 5283
rect 8591 5101 8625 5135
rect 8773 5189 8807 5223
rect 9017 5201 9051 5235
rect 9161 5227 9195 5261
rect 9056 5075 9090 5109
rect 9257 5199 9291 5233
rect 9532 5191 9566 5225
rect 9697 5165 9731 5199
rect 9957 5201 9991 5235
rect 10241 5227 10275 5261
rect 10403 5227 10437 5261
rect 9334 5091 9368 5125
rect 10163 5114 10197 5148
rect 10499 5227 10533 5261
rect 10331 5114 10365 5148
rect 10640 5191 10674 5225
rect 10736 5191 10770 5225
rect 10951 5165 10985 5199
rect 11061 5165 11095 5199
rect 11169 5201 11203 5235
rect 11279 5201 11313 5235
rect 11770 5191 11804 5225
rect 11866 5191 11900 5225
rect 12007 5227 12041 5261
rect 12103 5227 12137 5261
rect 12265 5227 12299 5261
rect 12175 5114 12209 5148
rect 12549 5165 12583 5199
rect 12809 5201 12843 5235
rect 12343 5114 12377 5148
rect 13093 5227 13127 5261
rect 13255 5227 13289 5261
rect 13015 5114 13049 5148
rect 13351 5227 13385 5261
rect 13183 5114 13217 5148
rect 13492 5191 13526 5225
rect 13588 5191 13622 5225
rect 14059 5165 14093 5199
rect 14423 5201 14457 5235
rect 15163 5165 15197 5199
rect 15527 5201 15561 5235
rect 16011 5165 16045 5199
rect 16121 5165 16155 5199
rect 16229 5201 16263 5235
rect 16339 5201 16373 5235
rect 17003 5165 17037 5199
rect 17367 5201 17401 5235
rect 17851 5165 17885 5199
rect 17950 5165 17984 5199
rect 18049 5165 18083 5199
rect 18157 5201 18191 5235
rect 18260 5201 18294 5235
rect 18363 5201 18397 5235
rect 18651 5205 18685 5239
rect 18759 5165 18793 5199
rect 1171 4593 1205 4627
rect 1279 4553 1313 4587
rect 1475 4593 1509 4627
rect 1574 4593 1608 4627
rect 1673 4593 1707 4627
rect 1781 4557 1815 4591
rect 1884 4557 1918 4591
rect 1987 4557 2021 4591
rect 2183 4593 2217 4627
rect 2291 4553 2325 4587
rect 2499 4567 2533 4601
rect 2695 4567 2729 4601
rect 2899 4567 2933 4601
rect 3013 4567 3047 4601
rect 3223 4593 3257 4627
rect 3333 4593 3367 4627
rect 3441 4557 3475 4591
rect 3551 4557 3585 4591
rect 4107 4567 4141 4601
rect 4175 4567 4209 4601
rect 4243 4567 4277 4601
rect 4389 4567 4423 4601
rect 4545 4593 4579 4627
rect 4805 4557 4839 4591
rect 5155 4593 5189 4627
rect 5254 4593 5288 4627
rect 5353 4593 5387 4627
rect 5461 4557 5495 4591
rect 5564 4557 5598 4591
rect 5667 4557 5701 4591
rect 6101 4567 6135 4601
rect 6204 4567 6238 4601
rect 6340 4567 6374 4601
rect 6477 4593 6511 4627
rect 6737 4557 6771 4591
rect 6874 4567 6908 4601
rect 7010 4567 7044 4601
rect 7113 4567 7147 4601
rect 7363 4593 7397 4627
rect 7473 4593 7507 4627
rect 7581 4557 7615 4591
rect 7691 4557 7725 4591
rect 7906 4567 7940 4601
rect 8002 4567 8036 4601
rect 8311 4644 8345 4678
rect 8143 4531 8177 4565
rect 8479 4644 8513 4678
rect 8239 4531 8273 4565
rect 8401 4531 8435 4565
rect 9174 4567 9208 4601
rect 9310 4567 9344 4601
rect 9413 4567 9447 4601
rect 9605 4593 9639 4627
rect 9865 4557 9899 4591
rect 10157 4593 10191 4627
rect 10417 4557 10451 4591
rect 10554 4567 10588 4601
rect 10690 4567 10724 4601
rect 10793 4567 10827 4601
rect 10985 4593 11019 4627
rect 11245 4557 11279 4591
rect 11353 4567 11387 4601
rect 11473 4580 11507 4614
rect 11629 4593 11663 4627
rect 12095 4644 12129 4678
rect 11889 4557 11923 4591
rect 12263 4644 12297 4678
rect 12173 4531 12207 4565
rect 12335 4531 12369 4565
rect 12431 4531 12465 4565
rect 12572 4567 12606 4601
rect 12668 4567 12702 4601
rect 12825 4593 12859 4627
rect 13085 4557 13119 4591
rect 13241 4580 13275 4614
rect 13361 4567 13395 4601
rect 13527 4593 13561 4627
rect 13637 4593 13671 4627
rect 13745 4557 13779 4591
rect 13855 4557 13889 4591
rect 14427 4593 14461 4627
rect 14791 4557 14825 4591
rect 15246 4567 15280 4601
rect 15382 4567 15416 4601
rect 15485 4567 15519 4601
rect 15677 4593 15711 4627
rect 15937 4557 15971 4591
rect 16093 4580 16127 4614
rect 16213 4567 16247 4601
rect 16321 4593 16355 4627
rect 16581 4557 16615 4591
rect 16737 4580 16771 4614
rect 16857 4567 16891 4601
rect 17279 4593 17313 4627
rect 17643 4557 17677 4591
rect 18127 4593 18161 4627
rect 18237 4593 18271 4627
rect 18345 4557 18379 4591
rect 18455 4557 18489 4591
rect 18651 4553 18685 4587
rect 18759 4593 18793 4627
rect 1171 4077 1205 4111
rect 1279 4117 1313 4151
rect 1475 4077 1509 4111
rect 1574 4077 1608 4111
rect 1673 4077 1707 4111
rect 1781 4113 1815 4147
rect 1884 4113 1918 4147
rect 1987 4113 2021 4147
rect 2245 4103 2279 4137
rect 2365 4090 2399 4124
rect 2521 4077 2555 4111
rect 2781 4113 2815 4147
rect 2884 4103 2918 4137
rect 2986 4088 3020 4122
rect 3352 4149 3386 4183
rect 3454 4155 3488 4189
rect 3193 4042 3227 4076
rect 3374 3987 3408 4021
rect 3709 4149 3743 4183
rect 3953 4161 3987 4195
rect 3623 4013 3657 4047
rect 3805 4101 3839 4135
rect 4049 4113 4083 4147
rect 4193 4139 4227 4173
rect 4088 3987 4122 4021
rect 4289 4111 4323 4145
rect 5131 4271 5165 4305
rect 5131 4203 5165 4237
rect 4564 4103 4598 4137
rect 4729 4077 4763 4111
rect 4989 4113 5023 4147
rect 4366 4003 4400 4037
rect 5131 3936 5165 3970
rect 5131 3868 5165 3902
rect 5231 4267 5265 4301
rect 5231 4199 5265 4233
rect 5431 4077 5465 4111
rect 5530 4077 5564 4111
rect 5629 4077 5663 4111
rect 5737 4113 5771 4147
rect 5840 4113 5874 4147
rect 5943 4113 5977 4147
rect 6415 4077 6449 4111
rect 6523 4117 6557 4151
rect 6709 4090 6743 4124
rect 6829 4103 6863 4137
rect 5231 3936 5265 3970
rect 5231 3868 5265 3902
rect 6995 4077 7029 4111
rect 7094 4077 7128 4111
rect 7193 4077 7227 4111
rect 7301 4113 7335 4147
rect 7404 4113 7438 4147
rect 7507 4113 7541 4147
rect 7849 4139 7883 4173
rect 8011 4139 8045 4173
rect 7771 4026 7805 4060
rect 8107 4139 8141 4173
rect 7939 4026 7973 4060
rect 8248 4103 8282 4137
rect 8344 4103 8378 4137
rect 8501 4077 8535 4111
rect 8761 4113 8795 4147
rect 8961 4103 8995 4137
rect 9388 4103 9422 4137
rect 9456 4103 9490 4137
rect 9524 4103 9558 4137
rect 9592 4103 9626 4137
rect 9660 4103 9694 4137
rect 9728 4103 9762 4137
rect 9796 4103 9830 4137
rect 9864 4103 9898 4137
rect 9932 4103 9966 4137
rect 10000 4103 10034 4137
rect 10068 4103 10102 4137
rect 10136 4103 10170 4137
rect 10204 4103 10238 4137
rect 10272 4103 10306 4137
rect 10340 4103 10374 4137
rect 10408 4103 10442 4137
rect 10859 4077 10893 4111
rect 10969 4077 11003 4111
rect 11077 4113 11111 4147
rect 11187 4113 11221 4147
rect 11778 4103 11812 4137
rect 12053 4111 12087 4145
rect 12149 4139 12183 4173
rect 11976 4003 12010 4037
rect 12293 4113 12327 4147
rect 12389 4161 12423 4195
rect 12254 3987 12288 4021
rect 12537 4101 12571 4135
rect 12633 4149 12667 4183
rect 12888 4155 12922 4189
rect 12990 4149 13024 4183
rect 12719 4013 12753 4047
rect 13149 4042 13183 4076
rect 12968 3987 13002 4021
rect 13356 4088 13390 4122
rect 13458 4103 13492 4137
rect 13561 4077 13595 4111
rect 13821 4113 13855 4147
rect 13924 4103 13958 4137
rect 14026 4088 14060 4122
rect 14392 4149 14426 4183
rect 14494 4155 14528 4189
rect 14233 4042 14267 4076
rect 14414 3987 14448 4021
rect 14749 4149 14783 4183
rect 14993 4161 15027 4195
rect 14663 4013 14697 4047
rect 14845 4101 14879 4135
rect 15089 4113 15123 4147
rect 15233 4139 15267 4173
rect 15128 3987 15162 4021
rect 15329 4111 15363 4145
rect 15604 4103 15638 4137
rect 15827 4077 15861 4111
rect 15926 4077 15960 4111
rect 16025 4077 16059 4111
rect 16133 4113 16167 4147
rect 16236 4113 16270 4147
rect 16339 4113 16373 4147
rect 17003 4077 17037 4111
rect 17367 4113 17401 4147
rect 17851 4077 17885 4111
rect 17950 4077 17984 4111
rect 18049 4077 18083 4111
rect 18157 4113 18191 4147
rect 18260 4113 18294 4147
rect 18363 4113 18397 4147
rect 18651 4117 18685 4151
rect 18759 4077 18793 4111
rect 15406 4003 15440 4037
rect 1171 3505 1205 3539
rect 1279 3465 1313 3499
rect 1447 3505 1481 3539
rect 1555 3465 1589 3499
rect 1688 3479 1722 3513
rect 1790 3494 1824 3528
rect 2178 3595 2212 3629
rect 1997 3540 2031 3574
rect 2427 3569 2461 3603
rect 2156 3433 2190 3467
rect 2258 3427 2292 3461
rect 2513 3433 2547 3467
rect 2609 3481 2643 3515
rect 2892 3595 2926 3629
rect 2757 3421 2791 3455
rect 2853 3469 2887 3503
rect 3170 3579 3204 3613
rect 2997 3443 3031 3477
rect 3093 3471 3127 3505
rect 3368 3479 3402 3513
rect 3867 3505 3901 3539
rect 3966 3505 4000 3539
rect 4065 3505 4099 3539
rect 4173 3469 4207 3503
rect 4276 3469 4310 3503
rect 4379 3469 4413 3503
rect 4830 3479 4864 3513
rect 4898 3479 4932 3513
rect 4966 3479 5000 3513
rect 5034 3479 5068 3513
rect 5102 3479 5136 3513
rect 5170 3479 5204 3513
rect 5238 3479 5272 3513
rect 5306 3479 5340 3513
rect 5374 3479 5408 3513
rect 5442 3479 5476 3513
rect 5510 3479 5544 3513
rect 5578 3479 5612 3513
rect 5646 3479 5680 3513
rect 5714 3479 5748 3513
rect 5782 3479 5816 3513
rect 5850 3479 5884 3513
rect 6277 3479 6311 3513
rect 6385 3505 6419 3539
rect 6645 3469 6679 3503
rect 6748 3479 6782 3513
rect 6850 3494 6884 3528
rect 7238 3595 7272 3629
rect 7057 3540 7091 3574
rect 7487 3569 7521 3603
rect 7216 3433 7250 3467
rect 7318 3427 7352 3461
rect 7573 3433 7607 3467
rect 7669 3481 7703 3515
rect 7952 3595 7986 3629
rect 7817 3421 7851 3455
rect 7913 3469 7947 3503
rect 8230 3579 8264 3613
rect 8057 3443 8091 3477
rect 8153 3471 8187 3505
rect 8428 3479 8462 3513
rect 8623 3505 8657 3539
rect 8731 3465 8765 3499
rect 9145 3479 9179 3513
rect 9269 3479 9303 3513
rect 9571 3505 9605 3539
rect 9681 3505 9715 3539
rect 9789 3469 9823 3503
rect 9899 3469 9933 3503
rect 10113 3492 10147 3526
rect 10233 3479 10267 3513
rect 10399 3505 10433 3539
rect 10509 3505 10543 3539
rect 12252 3579 12286 3613
rect 10617 3469 10651 3503
rect 10727 3469 10761 3503
rect 10985 3479 11019 3513
rect 11105 3492 11139 3526
rect 11319 3505 11353 3539
rect 11418 3505 11452 3539
rect 11517 3505 11551 3539
rect 11625 3469 11659 3503
rect 11728 3469 11762 3503
rect 11831 3469 11865 3503
rect 12054 3479 12088 3513
rect 12329 3471 12363 3505
rect 12530 3595 12564 3629
rect 12425 3443 12459 3477
rect 12569 3469 12603 3503
rect 12813 3481 12847 3515
rect 12995 3569 13029 3603
rect 12665 3421 12699 3455
rect 12909 3433 12943 3467
rect 13244 3595 13278 3629
rect 13425 3540 13459 3574
rect 13164 3427 13198 3461
rect 13266 3433 13300 3467
rect 13632 3494 13666 3528
rect 13734 3479 13768 3513
rect 14427 3505 14461 3539
rect 14791 3469 14825 3503
rect 15531 3505 15565 3539
rect 15895 3469 15929 3503
rect 16635 3505 16669 3539
rect 16999 3469 17033 3503
rect 17739 3505 17773 3539
rect 18103 3469 18137 3503
rect 18651 3465 18685 3499
rect 18759 3505 18793 3539
rect 1171 2989 1205 3023
rect 1279 3029 1313 3063
rect 1475 2989 1509 3023
rect 1585 2989 1619 3023
rect 1693 3025 1727 3059
rect 1803 3025 1837 3059
rect 2026 3015 2060 3049
rect 2301 3023 2335 3057
rect 2397 3051 2431 3085
rect 2224 2915 2258 2949
rect 2541 3025 2575 3059
rect 2637 3073 2671 3107
rect 2502 2899 2536 2933
rect 2785 3013 2819 3047
rect 2881 3061 2915 3095
rect 3136 3067 3170 3101
rect 3238 3061 3272 3095
rect 2967 2925 3001 2959
rect 3397 2954 3431 2988
rect 3216 2899 3250 2933
rect 3604 3000 3638 3034
rect 3706 3015 3740 3049
rect 3809 2989 3843 3023
rect 4069 3025 4103 3059
rect 4610 3073 4644 3107
rect 4172 3000 4206 3034
rect 4274 3000 4308 3034
rect 4706 3061 4740 3095
rect 4494 3013 4528 3047
rect 4878 3051 4912 3085
rect 4676 2899 4710 2933
rect 4812 2899 4846 2933
rect 5320 3061 5354 3095
rect 4980 2967 5014 3001
rect 5190 2995 5224 3029
rect 5492 3051 5526 3085
rect 5158 2899 5192 2933
rect 5342 2915 5376 2949
rect 5588 2995 5622 3029
rect 5876 3015 5910 3049
rect 6443 2989 6477 3023
rect 6542 2989 6576 3023
rect 6641 2989 6675 3023
rect 6749 3025 6783 3059
rect 6852 3025 6886 3059
rect 6955 3025 6989 3059
rect 7270 3015 7304 3049
rect 7545 3023 7579 3057
rect 7641 3051 7675 3085
rect 7468 2915 7502 2949
rect 7785 3025 7819 3059
rect 7881 3073 7915 3107
rect 7746 2899 7780 2933
rect 8029 3013 8063 3047
rect 8125 3061 8159 3095
rect 8380 3067 8414 3101
rect 8482 3061 8516 3095
rect 8211 2925 8245 2959
rect 8641 2954 8675 2988
rect 8460 2899 8494 2933
rect 8848 3000 8882 3034
rect 8950 3015 8984 3049
rect 9053 2989 9087 3023
rect 9313 3025 9347 3059
rect 9421 3015 9455 3049
rect 9848 3015 9882 3049
rect 9916 3015 9950 3049
rect 9984 3015 10018 3049
rect 10052 3015 10086 3049
rect 10120 3015 10154 3049
rect 10188 3015 10222 3049
rect 10256 3015 10290 3049
rect 10324 3015 10358 3049
rect 10392 3015 10426 3049
rect 10460 3015 10494 3049
rect 10528 3015 10562 3049
rect 10596 3015 10630 3049
rect 10664 3015 10698 3049
rect 10732 3015 10766 3049
rect 10800 3015 10834 3049
rect 10868 3015 10902 3049
rect 11778 3015 11812 3049
rect 12053 3023 12087 3057
rect 12149 3051 12183 3085
rect 11976 2915 12010 2949
rect 12293 3025 12327 3059
rect 12389 3073 12423 3107
rect 12254 2899 12288 2933
rect 12537 3013 12571 3047
rect 12633 3061 12667 3095
rect 12888 3067 12922 3101
rect 12990 3061 13024 3095
rect 12719 2925 12753 2959
rect 13149 2954 13183 2988
rect 12968 2899 13002 2933
rect 13356 3000 13390 3034
rect 13458 3015 13492 3049
rect 13561 2989 13595 3023
rect 13821 3025 13855 3059
rect 13929 3015 13963 3049
rect 14053 3015 14087 3049
rect 14611 2989 14645 3023
rect 14975 3025 15009 3059
rect 15715 2989 15749 3023
rect 16079 3025 16113 3059
rect 17003 2989 17037 3023
rect 17367 3025 17401 3059
rect 17851 2989 17885 3023
rect 17950 2989 17984 3023
rect 18049 2989 18083 3023
rect 18157 3025 18191 3059
rect 18260 3025 18294 3059
rect 18363 3025 18397 3059
rect 18651 3029 18685 3063
rect 18759 2989 18793 3023
rect 1171 2417 1205 2451
rect 1279 2377 1313 2411
rect 1447 2417 1481 2451
rect 1555 2377 1589 2411
rect 1688 2391 1722 2425
rect 1790 2406 1824 2440
rect 2178 2507 2212 2541
rect 1997 2452 2031 2486
rect 2427 2481 2461 2515
rect 2156 2345 2190 2379
rect 2258 2339 2292 2373
rect 2513 2345 2547 2379
rect 2609 2393 2643 2427
rect 2892 2507 2926 2541
rect 2757 2333 2791 2367
rect 2853 2381 2887 2415
rect 3170 2491 3204 2525
rect 2997 2355 3031 2389
rect 3093 2383 3127 2417
rect 3368 2391 3402 2425
rect 3809 2417 3843 2451
rect 4069 2381 4103 2415
rect 4264 2391 4298 2425
rect 4366 2406 4400 2440
rect 4754 2507 4788 2541
rect 4573 2452 4607 2486
rect 5003 2481 5037 2515
rect 4732 2345 4766 2379
rect 4834 2339 4868 2373
rect 5089 2345 5123 2379
rect 5185 2393 5219 2427
rect 5468 2507 5502 2541
rect 5333 2333 5367 2367
rect 5429 2381 5463 2415
rect 5746 2491 5780 2525
rect 5573 2355 5607 2389
rect 5669 2383 5703 2417
rect 5944 2391 5978 2425
rect 6699 2417 6733 2451
rect 9400 2491 9434 2525
rect 7063 2381 7097 2415
rect 7803 2417 7837 2451
rect 8167 2381 8201 2415
rect 8623 2417 8657 2451
rect 8731 2377 8765 2411
rect 9202 2391 9236 2425
rect 9477 2383 9511 2417
rect 9678 2507 9712 2541
rect 9573 2355 9607 2389
rect 9717 2381 9751 2415
rect 9961 2393 9995 2427
rect 10143 2481 10177 2515
rect 9813 2333 9847 2367
rect 10057 2345 10091 2379
rect 10392 2507 10426 2541
rect 10573 2452 10607 2486
rect 10312 2339 10346 2373
rect 10414 2345 10448 2379
rect 10780 2406 10814 2440
rect 12252 2491 12286 2525
rect 10882 2391 10916 2425
rect 10985 2417 11019 2451
rect 11245 2381 11279 2415
rect 11537 2417 11571 2451
rect 11797 2381 11831 2415
rect 12054 2391 12088 2425
rect 12329 2383 12363 2417
rect 12530 2507 12564 2541
rect 12425 2355 12459 2389
rect 12569 2381 12603 2415
rect 12813 2393 12847 2427
rect 12995 2481 13029 2515
rect 12665 2333 12699 2367
rect 12909 2345 12943 2379
rect 13244 2507 13278 2541
rect 13425 2452 13459 2486
rect 13164 2339 13198 2373
rect 13266 2345 13300 2379
rect 13632 2406 13666 2440
rect 14552 2491 14586 2525
rect 13734 2391 13768 2425
rect 14354 2391 14388 2425
rect 14629 2383 14663 2417
rect 14830 2507 14864 2541
rect 14725 2355 14759 2389
rect 14869 2381 14903 2415
rect 15113 2393 15147 2427
rect 15295 2481 15329 2515
rect 14965 2333 14999 2367
rect 15209 2345 15243 2379
rect 15544 2507 15578 2541
rect 15725 2452 15759 2486
rect 15464 2339 15498 2373
rect 15566 2345 15600 2379
rect 15932 2406 15966 2440
rect 16034 2391 16068 2425
rect 16137 2417 16171 2451
rect 16397 2381 16431 2415
rect 16747 2417 16781 2451
rect 16846 2417 16880 2451
rect 16945 2417 16979 2451
rect 17053 2381 17087 2415
rect 17156 2381 17190 2415
rect 17259 2381 17293 2415
rect 17517 2391 17551 2425
rect 17641 2391 17675 2425
rect 17943 2417 17977 2451
rect 18042 2417 18076 2451
rect 18141 2417 18175 2451
rect 18249 2381 18283 2415
rect 18352 2381 18386 2415
rect 18455 2381 18489 2415
rect 18651 2377 18685 2411
rect 18759 2417 18793 2451
<< rmp >>
rect 5081 4111 5177 4120
rect 5219 4111 5315 4120
<< ndiode >>
rect 9503 7559 9629 7577
rect 9503 7525 9511 7559
rect 9545 7525 9586 7559
rect 9620 7525 9629 7559
rect 9503 7491 9629 7525
rect 9503 7457 9511 7491
rect 9545 7457 9586 7491
rect 9620 7457 9629 7491
rect 9503 7439 9629 7457
rect 4903 4511 5029 4529
rect 4903 4477 4911 4511
rect 4945 4477 4986 4511
rect 5020 4477 5029 4511
rect 4903 4443 5029 4477
rect 4903 4409 4911 4443
rect 4945 4409 4986 4443
rect 5020 4409 5029 4443
rect 4903 4391 5029 4409
rect 9963 4511 10089 4529
rect 9963 4477 9971 4511
rect 10005 4477 10046 4511
rect 10080 4477 10089 4511
rect 9963 4443 10089 4477
rect 9963 4409 9971 4443
rect 10005 4409 10046 4443
rect 10080 4409 10089 4443
rect 9963 4391 10089 4409
<< ndiodec >>
rect 9511 7525 9545 7559
rect 9586 7525 9620 7559
rect 9511 7457 9545 7491
rect 9586 7457 9620 7491
rect 4911 4477 4945 4511
rect 4986 4477 5020 4511
rect 4911 4409 4945 4443
rect 4986 4409 5020 4443
rect 9971 4477 10005 4511
rect 10046 4477 10080 4511
rect 9971 4409 10005 4443
rect 10046 4409 10080 4443
<< locali >>
rect 1104 7599 1133 7633
rect 1167 7599 1225 7633
rect 1259 7599 1317 7633
rect 1351 7599 1409 7633
rect 1443 7599 1501 7633
rect 1535 7599 1593 7633
rect 1627 7599 1685 7633
rect 1719 7599 1777 7633
rect 1811 7599 1869 7633
rect 1903 7599 1961 7633
rect 1995 7599 2053 7633
rect 2087 7599 2145 7633
rect 2179 7599 2237 7633
rect 2271 7599 2329 7633
rect 2363 7599 2421 7633
rect 2455 7599 2513 7633
rect 2547 7599 2605 7633
rect 2639 7599 2697 7633
rect 2731 7599 2789 7633
rect 2823 7599 2881 7633
rect 2915 7599 2973 7633
rect 3007 7599 3065 7633
rect 3099 7599 3157 7633
rect 3191 7599 3249 7633
rect 3283 7599 3341 7633
rect 3375 7599 3433 7633
rect 3467 7599 3525 7633
rect 3559 7599 3617 7633
rect 3651 7599 3709 7633
rect 3743 7599 3801 7633
rect 3835 7599 3893 7633
rect 3927 7599 3985 7633
rect 4019 7599 4077 7633
rect 4111 7599 4169 7633
rect 4203 7599 4261 7633
rect 4295 7599 4353 7633
rect 4387 7599 4445 7633
rect 4479 7599 4537 7633
rect 4571 7599 4629 7633
rect 4663 7599 4721 7633
rect 4755 7599 4813 7633
rect 4847 7599 4905 7633
rect 4939 7599 4997 7633
rect 5031 7599 5089 7633
rect 5123 7599 5181 7633
rect 5215 7599 5273 7633
rect 5307 7599 5365 7633
rect 5399 7599 5457 7633
rect 5491 7599 5549 7633
rect 5583 7599 5641 7633
rect 5675 7599 5733 7633
rect 5767 7599 5825 7633
rect 5859 7599 5917 7633
rect 5951 7599 6009 7633
rect 6043 7599 6101 7633
rect 6135 7599 6193 7633
rect 6227 7599 6285 7633
rect 6319 7599 6377 7633
rect 6411 7599 6469 7633
rect 6503 7599 6561 7633
rect 6595 7599 6653 7633
rect 6687 7599 6745 7633
rect 6779 7599 6837 7633
rect 6871 7599 6929 7633
rect 6963 7599 7021 7633
rect 7055 7599 7113 7633
rect 7147 7599 7205 7633
rect 7239 7599 7297 7633
rect 7331 7599 7389 7633
rect 7423 7599 7481 7633
rect 7515 7599 7573 7633
rect 7607 7599 7665 7633
rect 7699 7599 7757 7633
rect 7791 7599 7849 7633
rect 7883 7599 7941 7633
rect 7975 7599 8033 7633
rect 8067 7599 8125 7633
rect 8159 7599 8217 7633
rect 8251 7599 8309 7633
rect 8343 7599 8401 7633
rect 8435 7599 8493 7633
rect 8527 7599 8585 7633
rect 8619 7599 8677 7633
rect 8711 7599 8769 7633
rect 8803 7599 8861 7633
rect 8895 7599 8953 7633
rect 8987 7599 9045 7633
rect 9079 7599 9137 7633
rect 9171 7599 9229 7633
rect 9263 7599 9321 7633
rect 9355 7599 9413 7633
rect 9447 7599 9505 7633
rect 9539 7599 9597 7633
rect 9631 7599 9689 7633
rect 9723 7599 9781 7633
rect 9815 7599 9873 7633
rect 9907 7599 9965 7633
rect 9999 7599 10057 7633
rect 10091 7599 10149 7633
rect 10183 7599 10241 7633
rect 10275 7599 10333 7633
rect 10367 7599 10425 7633
rect 10459 7599 10517 7633
rect 10551 7599 10609 7633
rect 10643 7599 10701 7633
rect 10735 7599 10793 7633
rect 10827 7599 10885 7633
rect 10919 7599 10977 7633
rect 11011 7599 11069 7633
rect 11103 7599 11161 7633
rect 11195 7599 11253 7633
rect 11287 7599 11345 7633
rect 11379 7599 11437 7633
rect 11471 7599 11529 7633
rect 11563 7599 11621 7633
rect 11655 7599 11713 7633
rect 11747 7599 11805 7633
rect 11839 7599 11897 7633
rect 11931 7599 11989 7633
rect 12023 7599 12081 7633
rect 12115 7599 12173 7633
rect 12207 7599 12265 7633
rect 12299 7599 12357 7633
rect 12391 7599 12449 7633
rect 12483 7599 12541 7633
rect 12575 7599 12633 7633
rect 12667 7599 12725 7633
rect 12759 7599 12817 7633
rect 12851 7599 12909 7633
rect 12943 7599 13001 7633
rect 13035 7599 13093 7633
rect 13127 7599 13185 7633
rect 13219 7599 13277 7633
rect 13311 7599 13369 7633
rect 13403 7599 13461 7633
rect 13495 7599 13553 7633
rect 13587 7599 13645 7633
rect 13679 7599 13737 7633
rect 13771 7599 13829 7633
rect 13863 7599 13921 7633
rect 13955 7599 14013 7633
rect 14047 7599 14105 7633
rect 14139 7599 14197 7633
rect 14231 7599 14289 7633
rect 14323 7599 14381 7633
rect 14415 7599 14473 7633
rect 14507 7599 14565 7633
rect 14599 7599 14657 7633
rect 14691 7599 14749 7633
rect 14783 7599 14841 7633
rect 14875 7599 14933 7633
rect 14967 7599 15025 7633
rect 15059 7599 15117 7633
rect 15151 7599 15209 7633
rect 15243 7599 15301 7633
rect 15335 7599 15393 7633
rect 15427 7599 15485 7633
rect 15519 7599 15577 7633
rect 15611 7599 15669 7633
rect 15703 7599 15761 7633
rect 15795 7599 15853 7633
rect 15887 7599 15945 7633
rect 15979 7599 16037 7633
rect 16071 7599 16129 7633
rect 16163 7599 16221 7633
rect 16255 7599 16313 7633
rect 16347 7599 16405 7633
rect 16439 7599 16497 7633
rect 16531 7599 16589 7633
rect 16623 7599 16681 7633
rect 16715 7599 16773 7633
rect 16807 7599 16865 7633
rect 16899 7599 16957 7633
rect 16991 7599 17049 7633
rect 17083 7599 17141 7633
rect 17175 7599 17233 7633
rect 17267 7599 17325 7633
rect 17359 7599 17417 7633
rect 17451 7599 17509 7633
rect 17543 7599 17601 7633
rect 17635 7599 17693 7633
rect 17727 7599 17785 7633
rect 17819 7599 17877 7633
rect 17911 7599 17969 7633
rect 18003 7599 18061 7633
rect 18095 7599 18153 7633
rect 18187 7599 18245 7633
rect 18279 7599 18337 7633
rect 18371 7599 18429 7633
rect 18463 7599 18521 7633
rect 18555 7599 18613 7633
rect 18647 7599 18705 7633
rect 18739 7599 18797 7633
rect 18831 7599 18860 7633
rect 1121 7536 1363 7599
rect 1121 7502 1139 7536
rect 1173 7502 1311 7536
rect 1345 7502 1363 7536
rect 1121 7449 1363 7502
rect 1582 7553 1634 7599
rect 1582 7519 1600 7553
rect 1582 7485 1634 7519
rect 1582 7451 1600 7485
rect 1121 7375 1225 7449
rect 1582 7431 1634 7451
rect 1669 7531 1720 7565
rect 1669 7527 1685 7531
rect 1669 7493 1684 7527
rect 1719 7497 1720 7531
rect 1754 7557 1820 7599
rect 1754 7523 1770 7557
rect 1804 7523 1820 7557
rect 1863 7544 1897 7565
rect 1718 7493 1720 7497
rect 1669 7450 1720 7493
rect 1863 7489 1897 7510
rect 1949 7538 3018 7599
rect 1949 7504 1967 7538
rect 2001 7504 2967 7538
rect 3001 7504 3018 7538
rect 1949 7490 3018 7504
rect 3053 7538 3571 7599
rect 3053 7504 3071 7538
rect 3105 7504 3519 7538
rect 3553 7504 3571 7538
rect 1754 7455 1897 7489
rect 1121 7341 1171 7375
rect 1205 7341 1225 7375
rect 1259 7381 1279 7415
rect 1313 7381 1363 7415
rect 1259 7307 1363 7381
rect 1121 7260 1363 7307
rect 1121 7226 1139 7260
rect 1173 7226 1311 7260
rect 1345 7226 1363 7260
rect 1121 7165 1363 7226
rect 1121 7131 1139 7165
rect 1173 7131 1311 7165
rect 1345 7131 1363 7165
rect 1121 7089 1363 7131
rect 1582 7301 1634 7319
rect 1582 7267 1600 7301
rect 1582 7233 1634 7267
rect 1582 7199 1600 7233
rect 1582 7165 1634 7199
rect 1582 7131 1600 7165
rect 1582 7089 1634 7131
rect 1669 7304 1703 7450
rect 1754 7417 1788 7455
rect 1737 7401 1788 7417
rect 1771 7367 1788 7401
rect 1737 7351 1788 7367
rect 1754 7309 1788 7351
rect 1844 7401 1915 7419
rect 1844 7367 1861 7401
rect 1895 7395 1915 7401
rect 1844 7361 1869 7367
rect 1903 7361 1915 7395
rect 1844 7345 1915 7361
rect 2266 7375 2334 7490
rect 3053 7445 3571 7504
rect 3697 7505 3755 7599
rect 3697 7471 3709 7505
rect 3743 7471 3755 7505
rect 3697 7454 3755 7471
rect 3974 7553 4026 7599
rect 3974 7519 3992 7553
rect 3974 7485 4026 7519
rect 3974 7451 3992 7485
rect 2266 7341 2283 7375
rect 2317 7341 2334 7375
rect 2266 7324 2334 7341
rect 2630 7411 2700 7426
rect 2630 7377 2647 7411
rect 2681 7377 2700 7411
rect 1669 7270 1720 7304
rect 1754 7275 1897 7309
rect 1669 7236 1684 7270
rect 1718 7236 1720 7270
rect 1863 7241 1897 7275
rect 1669 7189 1720 7236
rect 1669 7155 1684 7189
rect 1718 7155 1720 7189
rect 1669 7123 1720 7155
rect 1754 7207 1770 7241
rect 1804 7207 1820 7241
rect 1754 7173 1820 7207
rect 1754 7139 1770 7173
rect 1804 7139 1820 7173
rect 1754 7089 1820 7139
rect 1863 7173 1897 7207
rect 2630 7176 2700 7377
rect 3053 7375 3295 7445
rect 3974 7431 4026 7451
rect 4061 7531 4112 7565
rect 4061 7527 4077 7531
rect 4061 7493 4076 7527
rect 4111 7497 4112 7531
rect 4146 7557 4212 7599
rect 4146 7523 4162 7557
rect 4196 7523 4212 7557
rect 4255 7544 4289 7565
rect 4110 7493 4112 7497
rect 4061 7450 4112 7493
rect 4255 7489 4289 7510
rect 4341 7538 5410 7599
rect 4341 7504 4359 7538
rect 4393 7504 5359 7538
rect 5393 7504 5410 7538
rect 4341 7490 5410 7504
rect 5630 7553 5682 7599
rect 5630 7519 5648 7553
rect 4146 7455 4289 7489
rect 3053 7341 3131 7375
rect 3165 7341 3241 7375
rect 3275 7341 3295 7375
rect 3329 7377 3349 7411
rect 3383 7377 3459 7411
rect 3493 7377 3571 7411
rect 3329 7307 3571 7377
rect 3053 7267 3571 7307
rect 3053 7233 3071 7267
rect 3105 7233 3519 7267
rect 3553 7233 3571 7267
rect 1863 7123 1897 7139
rect 1949 7165 3018 7176
rect 1949 7131 1967 7165
rect 2001 7131 2967 7165
rect 3001 7131 3018 7165
rect 1949 7089 3018 7131
rect 3053 7165 3571 7233
rect 3053 7131 3071 7165
rect 3105 7131 3519 7165
rect 3553 7131 3571 7165
rect 3053 7089 3571 7131
rect 3697 7287 3755 7322
rect 3697 7253 3709 7287
rect 3743 7253 3755 7287
rect 3697 7194 3755 7253
rect 3697 7160 3709 7194
rect 3743 7160 3755 7194
rect 3697 7089 3755 7160
rect 3974 7301 4026 7319
rect 3974 7267 3992 7301
rect 3974 7233 4026 7267
rect 3974 7199 3992 7233
rect 3974 7165 4026 7199
rect 3974 7131 3992 7165
rect 3974 7089 4026 7131
rect 4061 7304 4095 7450
rect 4146 7417 4180 7455
rect 4129 7401 4180 7417
rect 4163 7367 4180 7401
rect 4129 7351 4180 7367
rect 4146 7309 4180 7351
rect 4236 7401 4307 7419
rect 4236 7367 4253 7401
rect 4287 7395 4307 7401
rect 4236 7361 4261 7367
rect 4295 7361 4307 7395
rect 4236 7345 4307 7361
rect 4658 7375 4726 7490
rect 5630 7485 5682 7519
rect 5630 7451 5648 7485
rect 5630 7431 5682 7451
rect 5717 7531 5768 7565
rect 5717 7527 5733 7531
rect 5717 7493 5732 7527
rect 5767 7497 5768 7531
rect 5802 7557 5868 7599
rect 5802 7523 5818 7557
rect 5852 7523 5868 7557
rect 5911 7544 5945 7565
rect 5766 7493 5768 7497
rect 5717 7450 5768 7493
rect 5911 7489 5945 7510
rect 5802 7455 5945 7489
rect 5997 7536 6239 7599
rect 5997 7502 6015 7536
rect 6049 7502 6187 7536
rect 6221 7502 6239 7536
rect 4658 7341 4675 7375
rect 4709 7341 4726 7375
rect 4658 7324 4726 7341
rect 5022 7411 5092 7426
rect 5022 7377 5039 7411
rect 5073 7377 5092 7411
rect 4061 7270 4112 7304
rect 4146 7275 4289 7309
rect 4061 7236 4076 7270
rect 4110 7236 4112 7270
rect 4255 7241 4289 7275
rect 4061 7189 4112 7236
rect 4061 7155 4076 7189
rect 4110 7155 4112 7189
rect 4061 7123 4112 7155
rect 4146 7207 4162 7241
rect 4196 7207 4212 7241
rect 4146 7173 4212 7207
rect 4146 7139 4162 7173
rect 4196 7139 4212 7173
rect 4146 7089 4212 7139
rect 4255 7173 4289 7207
rect 5022 7176 5092 7377
rect 5630 7301 5682 7319
rect 5630 7267 5648 7301
rect 5630 7233 5682 7267
rect 5630 7199 5648 7233
rect 4255 7123 4289 7139
rect 4341 7165 5410 7176
rect 4341 7131 4359 7165
rect 4393 7131 5359 7165
rect 5393 7131 5410 7165
rect 4341 7089 5410 7131
rect 5630 7165 5682 7199
rect 5630 7131 5648 7165
rect 5630 7089 5682 7131
rect 5717 7304 5751 7450
rect 5802 7417 5836 7455
rect 5997 7449 6239 7502
rect 6273 7505 6331 7599
rect 6273 7471 6285 7505
rect 6319 7471 6331 7505
rect 6365 7538 7434 7599
rect 6365 7504 6383 7538
rect 6417 7504 7383 7538
rect 7417 7504 7434 7538
rect 6365 7490 7434 7504
rect 7469 7531 7803 7599
rect 7469 7497 7487 7531
rect 7521 7497 7751 7531
rect 7785 7497 7803 7531
rect 6273 7454 6331 7471
rect 5785 7401 5836 7417
rect 5819 7367 5836 7401
rect 5785 7351 5836 7367
rect 5802 7309 5836 7351
rect 5892 7401 5963 7419
rect 5892 7367 5909 7401
rect 5943 7395 5963 7401
rect 5892 7361 5917 7367
rect 5951 7361 5963 7395
rect 5892 7345 5963 7361
rect 5997 7375 6101 7449
rect 5997 7341 6047 7375
rect 6081 7341 6101 7375
rect 6135 7381 6155 7415
rect 6189 7381 6239 7415
rect 5717 7270 5768 7304
rect 5802 7275 5945 7309
rect 6135 7307 6239 7381
rect 6682 7375 6750 7490
rect 7469 7445 7803 7497
rect 7838 7553 7890 7599
rect 7838 7519 7856 7553
rect 7838 7485 7890 7519
rect 7838 7451 7856 7485
rect 6682 7341 6699 7375
rect 6733 7341 6750 7375
rect 6682 7324 6750 7341
rect 7046 7411 7116 7426
rect 7046 7377 7063 7411
rect 7097 7377 7116 7411
rect 5717 7236 5732 7270
rect 5766 7236 5768 7270
rect 5911 7241 5945 7275
rect 5717 7189 5768 7236
rect 5717 7155 5732 7189
rect 5766 7155 5768 7189
rect 5717 7123 5768 7155
rect 5802 7207 5818 7241
rect 5852 7207 5868 7241
rect 5802 7173 5868 7207
rect 5802 7139 5818 7173
rect 5852 7139 5868 7173
rect 5802 7089 5868 7139
rect 5911 7173 5945 7207
rect 5911 7123 5945 7139
rect 5997 7260 6239 7307
rect 5997 7226 6015 7260
rect 6049 7226 6187 7260
rect 6221 7226 6239 7260
rect 5997 7165 6239 7226
rect 5997 7131 6015 7165
rect 6049 7131 6187 7165
rect 6221 7131 6239 7165
rect 5997 7089 6239 7131
rect 6273 7287 6331 7322
rect 6273 7253 6285 7287
rect 6319 7253 6331 7287
rect 6273 7194 6331 7253
rect 6273 7160 6285 7194
rect 6319 7160 6331 7194
rect 7046 7176 7116 7377
rect 7469 7375 7619 7445
rect 7838 7431 7890 7451
rect 7925 7531 7976 7565
rect 7925 7527 7941 7531
rect 7925 7493 7940 7527
rect 7975 7497 7976 7531
rect 8010 7557 8076 7599
rect 8010 7523 8026 7557
rect 8060 7523 8076 7557
rect 8119 7544 8153 7565
rect 7974 7493 7976 7497
rect 7925 7450 7976 7493
rect 8119 7489 8153 7510
rect 8010 7455 8153 7489
rect 8205 7538 8723 7599
rect 8205 7504 8223 7538
rect 8257 7504 8671 7538
rect 8705 7504 8723 7538
rect 7469 7341 7489 7375
rect 7523 7341 7619 7375
rect 7653 7377 7749 7411
rect 7783 7377 7803 7411
rect 7653 7307 7803 7377
rect 7469 7267 7803 7307
rect 7469 7233 7487 7267
rect 7521 7233 7751 7267
rect 7785 7233 7803 7267
rect 6273 7089 6331 7160
rect 6365 7165 7434 7176
rect 6365 7131 6383 7165
rect 6417 7131 7383 7165
rect 7417 7131 7434 7165
rect 6365 7089 7434 7131
rect 7469 7165 7803 7233
rect 7469 7131 7487 7165
rect 7521 7131 7751 7165
rect 7785 7131 7803 7165
rect 7469 7089 7803 7131
rect 7838 7301 7890 7319
rect 7838 7267 7856 7301
rect 7838 7233 7890 7267
rect 7838 7199 7856 7233
rect 7838 7165 7890 7199
rect 7838 7131 7856 7165
rect 7838 7089 7890 7131
rect 7925 7304 7959 7450
rect 8010 7417 8044 7455
rect 8205 7445 8723 7504
rect 8849 7505 8907 7599
rect 8849 7471 8861 7505
rect 8895 7471 8907 7505
rect 8849 7454 8907 7471
rect 8941 7538 9459 7599
rect 8941 7504 8959 7538
rect 8993 7504 9407 7538
rect 9441 7504 9459 7538
rect 8941 7445 9459 7504
rect 9493 7559 9643 7565
rect 9493 7525 9511 7559
rect 9545 7525 9586 7559
rect 9620 7525 9643 7559
rect 9493 7491 9643 7525
rect 9493 7457 9511 7491
rect 9545 7457 9586 7491
rect 9620 7463 9643 7491
rect 7993 7401 8044 7417
rect 8027 7367 8044 7401
rect 7993 7351 8044 7367
rect 8010 7309 8044 7351
rect 8100 7401 8171 7419
rect 8100 7367 8117 7401
rect 8151 7395 8171 7401
rect 8100 7361 8125 7367
rect 8159 7361 8171 7395
rect 8100 7345 8171 7361
rect 8205 7375 8447 7445
rect 8205 7341 8283 7375
rect 8317 7341 8393 7375
rect 8427 7341 8447 7375
rect 8481 7377 8501 7411
rect 8535 7377 8611 7411
rect 8645 7377 8723 7411
rect 7925 7270 7976 7304
rect 8010 7275 8153 7309
rect 8481 7307 8723 7377
rect 8941 7375 9183 7445
rect 9493 7429 9597 7457
rect 9631 7429 9643 7463
rect 8941 7341 9019 7375
rect 9053 7341 9129 7375
rect 9163 7341 9183 7375
rect 9217 7377 9237 7411
rect 9271 7377 9347 7411
rect 9381 7377 9459 7411
rect 7925 7236 7940 7270
rect 7974 7236 7976 7270
rect 8119 7241 8153 7275
rect 7925 7189 7976 7236
rect 7925 7155 7940 7189
rect 7974 7155 7976 7189
rect 7925 7123 7976 7155
rect 8010 7207 8026 7241
rect 8060 7207 8076 7241
rect 8010 7173 8076 7207
rect 8010 7139 8026 7173
rect 8060 7139 8076 7173
rect 8010 7089 8076 7139
rect 8119 7173 8153 7207
rect 8119 7123 8153 7139
rect 8205 7267 8723 7307
rect 8205 7233 8223 7267
rect 8257 7233 8671 7267
rect 8705 7233 8723 7267
rect 8205 7165 8723 7233
rect 8205 7131 8223 7165
rect 8257 7131 8671 7165
rect 8705 7131 8723 7165
rect 8205 7089 8723 7131
rect 8849 7287 8907 7322
rect 9217 7307 9459 7377
rect 8849 7253 8861 7287
rect 8895 7253 8907 7287
rect 8849 7194 8907 7253
rect 8849 7160 8861 7194
rect 8895 7160 8907 7194
rect 8849 7089 8907 7160
rect 8941 7267 9459 7307
rect 8941 7233 8959 7267
rect 8993 7233 9407 7267
rect 9441 7233 9459 7267
rect 8941 7165 9459 7233
rect 8941 7131 8959 7165
rect 8993 7131 9407 7165
rect 9441 7131 9459 7165
rect 8941 7089 9459 7131
rect 9493 7123 9643 7429
rect 9677 7531 10011 7599
rect 9677 7497 9695 7531
rect 9729 7497 9959 7531
rect 9993 7497 10011 7531
rect 9677 7445 10011 7497
rect 10045 7549 10097 7565
rect 10045 7515 10063 7549
rect 10045 7499 10097 7515
rect 10139 7553 10194 7599
rect 10139 7519 10149 7553
rect 10183 7519 10194 7553
rect 10139 7503 10194 7519
rect 10236 7549 10277 7565
rect 10236 7515 10243 7549
rect 10311 7553 10378 7599
rect 10311 7519 10327 7553
rect 10361 7519 10378 7553
rect 10413 7538 11115 7599
rect 9677 7375 9827 7445
rect 9677 7341 9697 7375
rect 9731 7341 9827 7375
rect 9861 7377 9957 7411
rect 9991 7377 10011 7411
rect 9861 7307 10011 7377
rect 9677 7267 10011 7307
rect 9677 7233 9695 7267
rect 9729 7233 9959 7267
rect 9993 7233 10011 7267
rect 9677 7165 10011 7233
rect 9677 7131 9695 7165
rect 9729 7131 9959 7165
rect 9993 7131 10011 7165
rect 9677 7089 10011 7131
rect 10045 7317 10079 7499
rect 10236 7485 10277 7515
rect 10413 7504 10431 7538
rect 10465 7504 11063 7538
rect 11097 7504 11115 7538
rect 10113 7463 10185 7467
rect 10113 7429 10149 7463
rect 10183 7429 10185 7463
rect 10236 7451 10373 7485
rect 10113 7401 10185 7429
rect 10113 7367 10117 7401
rect 10151 7367 10185 7401
rect 10113 7351 10185 7367
rect 10221 7401 10271 7417
rect 10255 7367 10271 7401
rect 10221 7317 10271 7367
rect 10045 7284 10271 7317
rect 10045 7250 10063 7284
rect 10097 7283 10271 7284
rect 10097 7250 10099 7283
rect 10045 7179 10099 7250
rect 10305 7259 10373 7451
rect 10413 7445 11115 7504
rect 11149 7536 11391 7599
rect 11149 7502 11167 7536
rect 11201 7502 11339 7536
rect 11373 7502 11391 7536
rect 11149 7449 11391 7502
rect 11425 7505 11483 7599
rect 11425 7471 11437 7505
rect 11471 7471 11483 7505
rect 11425 7454 11483 7471
rect 11517 7538 12219 7599
rect 11517 7504 11535 7538
rect 11569 7504 12167 7538
rect 12201 7504 12219 7538
rect 10413 7375 10743 7445
rect 10413 7341 10491 7375
rect 10525 7341 10590 7375
rect 10624 7341 10689 7375
rect 10723 7341 10743 7375
rect 10777 7377 10797 7411
rect 10831 7377 10900 7411
rect 10934 7377 11003 7411
rect 11037 7377 11115 7411
rect 10777 7307 11115 7377
rect 11149 7375 11253 7449
rect 11517 7445 12219 7504
rect 12271 7544 12305 7565
rect 12348 7557 12414 7599
rect 12348 7523 12364 7557
rect 12398 7523 12414 7557
rect 12448 7531 12499 7565
rect 12271 7489 12305 7510
rect 12448 7497 12449 7531
rect 12483 7527 12499 7531
rect 12448 7493 12450 7497
rect 12484 7493 12499 7527
rect 12271 7455 12414 7489
rect 11149 7341 11199 7375
rect 11233 7341 11253 7375
rect 11287 7381 11307 7415
rect 11341 7381 11391 7415
rect 11287 7307 11391 7381
rect 11517 7375 11847 7445
rect 11517 7341 11595 7375
rect 11629 7341 11694 7375
rect 11728 7341 11793 7375
rect 11827 7341 11847 7375
rect 11881 7377 11901 7411
rect 11935 7377 12004 7411
rect 12038 7377 12107 7411
rect 12141 7377 12219 7411
rect 10305 7245 10333 7259
rect 10045 7145 10063 7179
rect 10097 7145 10099 7179
rect 10045 7129 10099 7145
rect 10133 7211 10149 7245
rect 10183 7211 10199 7245
rect 10133 7177 10199 7211
rect 10133 7143 10149 7177
rect 10183 7143 10199 7177
rect 10133 7089 10199 7143
rect 10240 7225 10333 7245
rect 10367 7225 10373 7259
rect 10240 7210 10373 7225
rect 10413 7267 11115 7307
rect 10413 7233 10431 7267
rect 10465 7233 11063 7267
rect 11097 7233 11115 7267
rect 10240 7179 10277 7210
rect 10240 7145 10243 7179
rect 10240 7129 10277 7145
rect 10311 7140 10327 7174
rect 10361 7140 10378 7174
rect 10311 7089 10378 7140
rect 10413 7165 11115 7233
rect 10413 7131 10431 7165
rect 10465 7131 11063 7165
rect 11097 7131 11115 7165
rect 10413 7089 11115 7131
rect 11149 7260 11391 7307
rect 11149 7226 11167 7260
rect 11201 7226 11339 7260
rect 11373 7226 11391 7260
rect 11149 7165 11391 7226
rect 11149 7131 11167 7165
rect 11201 7131 11339 7165
rect 11373 7131 11391 7165
rect 11149 7089 11391 7131
rect 11425 7287 11483 7322
rect 11881 7307 12219 7377
rect 12253 7401 12324 7419
rect 12253 7395 12273 7401
rect 12253 7361 12265 7395
rect 12307 7367 12324 7401
rect 12299 7361 12324 7367
rect 12253 7345 12324 7361
rect 12380 7417 12414 7455
rect 12448 7450 12499 7493
rect 12380 7401 12431 7417
rect 12380 7367 12397 7401
rect 12380 7351 12431 7367
rect 12380 7309 12414 7351
rect 11425 7253 11437 7287
rect 11471 7253 11483 7287
rect 11425 7194 11483 7253
rect 11425 7160 11437 7194
rect 11471 7160 11483 7194
rect 11425 7089 11483 7160
rect 11517 7267 12219 7307
rect 11517 7233 11535 7267
rect 11569 7233 12167 7267
rect 12201 7233 12219 7267
rect 11517 7165 12219 7233
rect 11517 7131 11535 7165
rect 11569 7131 12167 7165
rect 12201 7131 12219 7165
rect 11517 7089 12219 7131
rect 12271 7275 12414 7309
rect 12465 7304 12499 7450
rect 12534 7553 12586 7599
rect 12568 7519 12586 7553
rect 12534 7485 12586 7519
rect 12621 7538 13690 7599
rect 12621 7504 12639 7538
rect 12673 7504 13639 7538
rect 13673 7504 13690 7538
rect 12621 7490 13690 7504
rect 13725 7536 13967 7599
rect 13725 7502 13743 7536
rect 13777 7502 13915 7536
rect 13949 7502 13967 7536
rect 12568 7451 12586 7485
rect 12534 7431 12586 7451
rect 12938 7375 13006 7490
rect 13725 7449 13967 7502
rect 14001 7505 14059 7599
rect 14001 7471 14013 7505
rect 14047 7471 14059 7505
rect 14001 7454 14059 7471
rect 14093 7531 14427 7599
rect 14093 7497 14111 7531
rect 14145 7497 14375 7531
rect 14409 7497 14427 7531
rect 12938 7341 12955 7375
rect 12989 7341 13006 7375
rect 12938 7324 13006 7341
rect 13302 7411 13372 7426
rect 13302 7377 13319 7411
rect 13353 7377 13372 7411
rect 12271 7241 12305 7275
rect 12448 7270 12499 7304
rect 12271 7173 12305 7207
rect 12271 7123 12305 7139
rect 12348 7207 12364 7241
rect 12398 7207 12414 7241
rect 12348 7173 12414 7207
rect 12348 7139 12364 7173
rect 12398 7139 12414 7173
rect 12348 7089 12414 7139
rect 12448 7236 12450 7270
rect 12484 7236 12499 7270
rect 12448 7189 12499 7236
rect 12448 7155 12450 7189
rect 12484 7155 12499 7189
rect 12448 7123 12499 7155
rect 12534 7301 12586 7319
rect 12568 7267 12586 7301
rect 12534 7233 12586 7267
rect 12568 7199 12586 7233
rect 12534 7165 12586 7199
rect 13302 7176 13372 7377
rect 13725 7375 13829 7449
rect 14093 7445 14427 7497
rect 14479 7544 14513 7565
rect 14556 7557 14622 7599
rect 14556 7523 14572 7557
rect 14606 7523 14622 7557
rect 14656 7531 14707 7565
rect 14479 7489 14513 7510
rect 14656 7497 14657 7531
rect 14691 7527 14707 7531
rect 14656 7493 14658 7497
rect 14692 7493 14707 7527
rect 14479 7455 14622 7489
rect 13725 7341 13775 7375
rect 13809 7341 13829 7375
rect 13863 7381 13883 7415
rect 13917 7381 13967 7415
rect 13863 7307 13967 7381
rect 14093 7375 14243 7445
rect 14093 7341 14113 7375
rect 14147 7341 14243 7375
rect 14277 7377 14373 7411
rect 14407 7377 14427 7411
rect 13725 7260 13967 7307
rect 13725 7226 13743 7260
rect 13777 7226 13915 7260
rect 13949 7226 13967 7260
rect 12568 7131 12586 7165
rect 12534 7089 12586 7131
rect 12621 7165 13690 7176
rect 12621 7131 12639 7165
rect 12673 7131 13639 7165
rect 13673 7131 13690 7165
rect 12621 7089 13690 7131
rect 13725 7165 13967 7226
rect 13725 7131 13743 7165
rect 13777 7131 13915 7165
rect 13949 7131 13967 7165
rect 13725 7089 13967 7131
rect 14001 7287 14059 7322
rect 14277 7307 14427 7377
rect 14461 7401 14532 7419
rect 14461 7395 14481 7401
rect 14461 7361 14473 7395
rect 14515 7367 14532 7401
rect 14507 7361 14532 7367
rect 14461 7345 14532 7361
rect 14588 7417 14622 7455
rect 14656 7450 14707 7493
rect 14588 7401 14639 7417
rect 14588 7367 14605 7401
rect 14588 7351 14639 7367
rect 14588 7309 14622 7351
rect 14001 7253 14013 7287
rect 14047 7253 14059 7287
rect 14001 7194 14059 7253
rect 14001 7160 14013 7194
rect 14047 7160 14059 7194
rect 14001 7089 14059 7160
rect 14093 7267 14427 7307
rect 14093 7233 14111 7267
rect 14145 7233 14375 7267
rect 14409 7233 14427 7267
rect 14093 7165 14427 7233
rect 14093 7131 14111 7165
rect 14145 7131 14375 7165
rect 14409 7131 14427 7165
rect 14093 7089 14427 7131
rect 14479 7275 14622 7309
rect 14673 7304 14707 7450
rect 14742 7553 14794 7599
rect 14776 7519 14794 7553
rect 14742 7485 14794 7519
rect 14829 7538 15898 7599
rect 14829 7504 14847 7538
rect 14881 7504 15847 7538
rect 15881 7504 15898 7538
rect 14829 7490 15898 7504
rect 15933 7538 16451 7599
rect 15933 7504 15951 7538
rect 15985 7504 16399 7538
rect 16433 7504 16451 7538
rect 14776 7451 14794 7485
rect 14742 7431 14794 7451
rect 15146 7375 15214 7490
rect 15933 7445 16451 7504
rect 16577 7505 16635 7599
rect 16577 7471 16589 7505
rect 16623 7471 16635 7505
rect 16577 7454 16635 7471
rect 16871 7544 16905 7565
rect 16948 7557 17014 7599
rect 16948 7523 16964 7557
rect 16998 7523 17014 7557
rect 17048 7531 17099 7565
rect 16871 7489 16905 7510
rect 17048 7497 17049 7531
rect 17083 7527 17099 7531
rect 17048 7493 17050 7497
rect 17084 7493 17099 7527
rect 16871 7455 17014 7489
rect 15146 7341 15163 7375
rect 15197 7341 15214 7375
rect 15146 7324 15214 7341
rect 15510 7411 15580 7426
rect 15510 7377 15527 7411
rect 15561 7377 15580 7411
rect 14479 7241 14513 7275
rect 14656 7270 14707 7304
rect 14479 7173 14513 7207
rect 14479 7123 14513 7139
rect 14556 7207 14572 7241
rect 14606 7207 14622 7241
rect 14556 7173 14622 7207
rect 14556 7139 14572 7173
rect 14606 7139 14622 7173
rect 14556 7089 14622 7139
rect 14656 7236 14658 7270
rect 14692 7236 14707 7270
rect 14656 7189 14707 7236
rect 14656 7155 14658 7189
rect 14692 7155 14707 7189
rect 14656 7123 14707 7155
rect 14742 7301 14794 7319
rect 14776 7267 14794 7301
rect 14742 7233 14794 7267
rect 14776 7199 14794 7233
rect 14742 7165 14794 7199
rect 15510 7176 15580 7377
rect 15933 7375 16175 7445
rect 15933 7341 16011 7375
rect 16045 7341 16121 7375
rect 16155 7341 16175 7375
rect 16209 7377 16229 7411
rect 16263 7377 16339 7411
rect 16373 7377 16451 7411
rect 16209 7307 16451 7377
rect 16853 7401 16924 7419
rect 16853 7395 16873 7401
rect 16853 7361 16865 7395
rect 16907 7367 16924 7401
rect 16899 7361 16924 7367
rect 16853 7345 16924 7361
rect 16980 7417 17014 7455
rect 17048 7450 17099 7493
rect 16980 7401 17031 7417
rect 16980 7367 16997 7401
rect 16980 7351 17031 7367
rect 15933 7267 16451 7307
rect 15933 7233 15951 7267
rect 15985 7233 16399 7267
rect 16433 7233 16451 7267
rect 14776 7131 14794 7165
rect 14742 7089 14794 7131
rect 14829 7165 15898 7176
rect 14829 7131 14847 7165
rect 14881 7131 15847 7165
rect 15881 7131 15898 7165
rect 14829 7089 15898 7131
rect 15933 7165 16451 7233
rect 15933 7131 15951 7165
rect 15985 7131 16399 7165
rect 16433 7131 16451 7165
rect 15933 7089 16451 7131
rect 16577 7287 16635 7322
rect 16980 7309 17014 7351
rect 16577 7253 16589 7287
rect 16623 7253 16635 7287
rect 16577 7194 16635 7253
rect 16577 7160 16589 7194
rect 16623 7160 16635 7194
rect 16577 7089 16635 7160
rect 16871 7275 17014 7309
rect 17065 7304 17099 7450
rect 17134 7553 17186 7599
rect 17168 7519 17186 7553
rect 17134 7485 17186 7519
rect 17168 7451 17186 7485
rect 17134 7431 17186 7451
rect 17221 7538 17923 7599
rect 17221 7504 17239 7538
rect 17273 7504 17871 7538
rect 17905 7504 17923 7538
rect 17221 7445 17923 7504
rect 18067 7544 18101 7565
rect 18144 7557 18210 7599
rect 18144 7523 18160 7557
rect 18194 7523 18210 7557
rect 18244 7531 18295 7565
rect 18067 7489 18101 7510
rect 18244 7497 18245 7531
rect 18279 7527 18295 7531
rect 18244 7493 18246 7497
rect 18280 7493 18295 7527
rect 18067 7455 18210 7489
rect 17221 7375 17551 7445
rect 17221 7341 17299 7375
rect 17333 7341 17398 7375
rect 17432 7341 17497 7375
rect 17531 7341 17551 7375
rect 17585 7377 17605 7411
rect 17639 7377 17708 7411
rect 17742 7377 17811 7411
rect 17845 7377 17923 7411
rect 16871 7241 16905 7275
rect 17048 7270 17099 7304
rect 16871 7173 16905 7207
rect 16871 7123 16905 7139
rect 16948 7207 16964 7241
rect 16998 7207 17014 7241
rect 16948 7173 17014 7207
rect 16948 7139 16964 7173
rect 16998 7139 17014 7173
rect 16948 7089 17014 7139
rect 17048 7236 17050 7270
rect 17084 7236 17099 7270
rect 17048 7189 17099 7236
rect 17048 7155 17050 7189
rect 17084 7155 17099 7189
rect 17048 7123 17099 7155
rect 17134 7301 17186 7319
rect 17585 7307 17923 7377
rect 18049 7401 18120 7419
rect 18049 7395 18069 7401
rect 18049 7361 18061 7395
rect 18103 7367 18120 7401
rect 18095 7361 18120 7367
rect 18049 7345 18120 7361
rect 18176 7417 18210 7455
rect 18244 7450 18295 7493
rect 18176 7401 18227 7417
rect 18176 7367 18193 7401
rect 18176 7351 18227 7367
rect 18176 7309 18210 7351
rect 17168 7267 17186 7301
rect 17134 7233 17186 7267
rect 17168 7199 17186 7233
rect 17134 7165 17186 7199
rect 17168 7131 17186 7165
rect 17134 7089 17186 7131
rect 17221 7267 17923 7307
rect 17221 7233 17239 7267
rect 17273 7233 17871 7267
rect 17905 7233 17923 7267
rect 17221 7165 17923 7233
rect 17221 7131 17239 7165
rect 17273 7131 17871 7165
rect 17905 7131 17923 7165
rect 17221 7089 17923 7131
rect 18067 7275 18210 7309
rect 18261 7304 18295 7450
rect 18330 7553 18382 7599
rect 18364 7519 18382 7553
rect 18330 7485 18382 7519
rect 18364 7451 18382 7485
rect 18330 7431 18382 7451
rect 18601 7536 18843 7599
rect 18601 7502 18619 7536
rect 18653 7502 18791 7536
rect 18825 7502 18843 7536
rect 18601 7449 18843 7502
rect 18601 7381 18651 7415
rect 18685 7381 18705 7415
rect 18067 7241 18101 7275
rect 18244 7270 18295 7304
rect 18067 7173 18101 7207
rect 18067 7123 18101 7139
rect 18144 7207 18160 7241
rect 18194 7207 18210 7241
rect 18144 7173 18210 7207
rect 18144 7139 18160 7173
rect 18194 7139 18210 7173
rect 18144 7089 18210 7139
rect 18244 7236 18246 7270
rect 18280 7236 18295 7270
rect 18244 7189 18295 7236
rect 18244 7155 18246 7189
rect 18280 7155 18295 7189
rect 18244 7123 18295 7155
rect 18330 7301 18382 7319
rect 18364 7267 18382 7301
rect 18330 7233 18382 7267
rect 18364 7199 18382 7233
rect 18330 7165 18382 7199
rect 18364 7131 18382 7165
rect 18330 7089 18382 7131
rect 18601 7307 18705 7381
rect 18739 7375 18843 7449
rect 18739 7341 18759 7375
rect 18793 7341 18843 7375
rect 18601 7260 18843 7307
rect 18601 7226 18619 7260
rect 18653 7226 18791 7260
rect 18825 7226 18843 7260
rect 18601 7165 18843 7226
rect 18601 7131 18619 7165
rect 18653 7131 18791 7165
rect 18825 7131 18843 7165
rect 18601 7089 18843 7131
rect 1104 7055 1133 7089
rect 1167 7055 1225 7089
rect 1259 7055 1317 7089
rect 1351 7055 1409 7089
rect 1443 7055 1501 7089
rect 1535 7055 1593 7089
rect 1627 7055 1685 7089
rect 1719 7055 1777 7089
rect 1811 7055 1869 7089
rect 1903 7055 1961 7089
rect 1995 7055 2053 7089
rect 2087 7055 2145 7089
rect 2179 7055 2237 7089
rect 2271 7055 2329 7089
rect 2363 7055 2421 7089
rect 2455 7055 2513 7089
rect 2547 7055 2605 7089
rect 2639 7055 2697 7089
rect 2731 7055 2789 7089
rect 2823 7055 2881 7089
rect 2915 7055 2973 7089
rect 3007 7055 3065 7089
rect 3099 7055 3157 7089
rect 3191 7055 3249 7089
rect 3283 7055 3341 7089
rect 3375 7055 3433 7089
rect 3467 7055 3525 7089
rect 3559 7055 3617 7089
rect 3651 7055 3709 7089
rect 3743 7055 3801 7089
rect 3835 7055 3893 7089
rect 3927 7055 3985 7089
rect 4019 7055 4077 7089
rect 4111 7055 4169 7089
rect 4203 7055 4261 7089
rect 4295 7055 4353 7089
rect 4387 7055 4445 7089
rect 4479 7055 4537 7089
rect 4571 7055 4629 7089
rect 4663 7055 4721 7089
rect 4755 7055 4813 7089
rect 4847 7055 4905 7089
rect 4939 7055 4997 7089
rect 5031 7055 5089 7089
rect 5123 7055 5181 7089
rect 5215 7055 5273 7089
rect 5307 7055 5365 7089
rect 5399 7055 5457 7089
rect 5491 7055 5549 7089
rect 5583 7055 5641 7089
rect 5675 7055 5733 7089
rect 5767 7055 5825 7089
rect 5859 7055 5917 7089
rect 5951 7055 6009 7089
rect 6043 7055 6101 7089
rect 6135 7055 6193 7089
rect 6227 7055 6285 7089
rect 6319 7055 6377 7089
rect 6411 7055 6469 7089
rect 6503 7055 6561 7089
rect 6595 7055 6653 7089
rect 6687 7055 6745 7089
rect 6779 7055 6837 7089
rect 6871 7055 6929 7089
rect 6963 7055 7021 7089
rect 7055 7055 7113 7089
rect 7147 7055 7205 7089
rect 7239 7055 7297 7089
rect 7331 7055 7389 7089
rect 7423 7055 7481 7089
rect 7515 7055 7573 7089
rect 7607 7055 7665 7089
rect 7699 7055 7757 7089
rect 7791 7055 7849 7089
rect 7883 7055 7941 7089
rect 7975 7055 8033 7089
rect 8067 7055 8125 7089
rect 8159 7055 8217 7089
rect 8251 7055 8309 7089
rect 8343 7055 8401 7089
rect 8435 7055 8493 7089
rect 8527 7055 8585 7089
rect 8619 7055 8677 7089
rect 8711 7055 8769 7089
rect 8803 7055 8861 7089
rect 8895 7055 8953 7089
rect 8987 7055 9045 7089
rect 9079 7055 9137 7089
rect 9171 7055 9229 7089
rect 9263 7055 9321 7089
rect 9355 7055 9413 7089
rect 9447 7055 9505 7089
rect 9539 7055 9597 7089
rect 9631 7055 9689 7089
rect 9723 7055 9781 7089
rect 9815 7055 9873 7089
rect 9907 7055 9965 7089
rect 9999 7055 10057 7089
rect 10091 7055 10149 7089
rect 10183 7055 10241 7089
rect 10275 7055 10333 7089
rect 10367 7055 10425 7089
rect 10459 7055 10517 7089
rect 10551 7055 10609 7089
rect 10643 7055 10701 7089
rect 10735 7055 10793 7089
rect 10827 7055 10885 7089
rect 10919 7055 10977 7089
rect 11011 7055 11069 7089
rect 11103 7055 11161 7089
rect 11195 7055 11253 7089
rect 11287 7055 11345 7089
rect 11379 7055 11437 7089
rect 11471 7055 11529 7089
rect 11563 7055 11621 7089
rect 11655 7055 11713 7089
rect 11747 7055 11805 7089
rect 11839 7055 11897 7089
rect 11931 7055 11989 7089
rect 12023 7055 12081 7089
rect 12115 7055 12173 7089
rect 12207 7055 12265 7089
rect 12299 7055 12357 7089
rect 12391 7055 12449 7089
rect 12483 7055 12541 7089
rect 12575 7055 12633 7089
rect 12667 7055 12725 7089
rect 12759 7055 12817 7089
rect 12851 7055 12909 7089
rect 12943 7055 13001 7089
rect 13035 7055 13093 7089
rect 13127 7055 13185 7089
rect 13219 7055 13277 7089
rect 13311 7055 13369 7089
rect 13403 7055 13461 7089
rect 13495 7055 13553 7089
rect 13587 7055 13645 7089
rect 13679 7055 13737 7089
rect 13771 7055 13829 7089
rect 13863 7055 13921 7089
rect 13955 7055 14013 7089
rect 14047 7055 14105 7089
rect 14139 7055 14197 7089
rect 14231 7055 14289 7089
rect 14323 7055 14381 7089
rect 14415 7055 14473 7089
rect 14507 7055 14565 7089
rect 14599 7055 14657 7089
rect 14691 7055 14749 7089
rect 14783 7055 14841 7089
rect 14875 7055 14933 7089
rect 14967 7055 15025 7089
rect 15059 7055 15117 7089
rect 15151 7055 15209 7089
rect 15243 7055 15301 7089
rect 15335 7055 15393 7089
rect 15427 7055 15485 7089
rect 15519 7055 15577 7089
rect 15611 7055 15669 7089
rect 15703 7055 15761 7089
rect 15795 7055 15853 7089
rect 15887 7055 15945 7089
rect 15979 7055 16037 7089
rect 16071 7055 16129 7089
rect 16163 7055 16221 7089
rect 16255 7055 16313 7089
rect 16347 7055 16405 7089
rect 16439 7055 16497 7089
rect 16531 7055 16589 7089
rect 16623 7055 16681 7089
rect 16715 7055 16773 7089
rect 16807 7055 16865 7089
rect 16899 7055 16957 7089
rect 16991 7055 17049 7089
rect 17083 7055 17141 7089
rect 17175 7055 17233 7089
rect 17267 7055 17325 7089
rect 17359 7055 17417 7089
rect 17451 7055 17509 7089
rect 17543 7055 17601 7089
rect 17635 7055 17693 7089
rect 17727 7055 17785 7089
rect 17819 7055 17877 7089
rect 17911 7055 17969 7089
rect 18003 7055 18061 7089
rect 18095 7055 18153 7089
rect 18187 7055 18245 7089
rect 18279 7055 18337 7089
rect 18371 7055 18429 7089
rect 18463 7055 18521 7089
rect 18555 7055 18613 7089
rect 18647 7055 18705 7089
rect 18739 7055 18797 7089
rect 18831 7055 18860 7089
rect 1121 7013 1363 7055
rect 1121 6979 1139 7013
rect 1173 6979 1311 7013
rect 1345 6979 1363 7013
rect 1121 6918 1363 6979
rect 1397 7013 2466 7055
rect 1397 6979 1415 7013
rect 1449 6979 2415 7013
rect 2449 6979 2466 7013
rect 1397 6968 2466 6979
rect 2501 7013 3570 7055
rect 2501 6979 2519 7013
rect 2553 6979 3519 7013
rect 3553 6979 3570 7013
rect 2501 6968 3570 6979
rect 3697 6984 3755 7055
rect 1121 6884 1139 6918
rect 1173 6884 1311 6918
rect 1345 6884 1363 6918
rect 1121 6837 1363 6884
rect 1121 6769 1171 6803
rect 1205 6769 1225 6803
rect 1121 6695 1225 6769
rect 1259 6763 1363 6837
rect 1259 6729 1279 6763
rect 1313 6729 1363 6763
rect 1714 6803 1782 6820
rect 1714 6769 1731 6803
rect 1765 6769 1782 6803
rect 1121 6642 1363 6695
rect 1714 6654 1782 6769
rect 2078 6767 2148 6968
rect 2078 6733 2095 6767
rect 2129 6733 2148 6767
rect 2078 6718 2148 6733
rect 2818 6803 2886 6820
rect 2818 6769 2835 6803
rect 2869 6769 2886 6803
rect 2818 6654 2886 6769
rect 3182 6767 3252 6968
rect 3697 6950 3709 6984
rect 3743 6950 3755 6984
rect 3789 7013 4858 7055
rect 3789 6979 3807 7013
rect 3841 6979 4807 7013
rect 4841 6979 4858 7013
rect 3789 6968 4858 6979
rect 4893 7013 5962 7055
rect 4893 6979 4911 7013
rect 4945 6979 5911 7013
rect 5945 6979 5962 7013
rect 4893 6968 5962 6979
rect 5997 7013 7066 7055
rect 5997 6979 6015 7013
rect 6049 6979 7015 7013
rect 7049 6979 7066 7013
rect 5997 6968 7066 6979
rect 7101 7013 8170 7055
rect 7101 6979 7119 7013
rect 7153 6979 8119 7013
rect 8153 6979 8170 7013
rect 7101 6968 8170 6979
rect 8205 7013 8723 7055
rect 8205 6979 8223 7013
rect 8257 6979 8671 7013
rect 8705 6979 8723 7013
rect 3697 6891 3755 6950
rect 3697 6857 3709 6891
rect 3743 6857 3755 6891
rect 3697 6822 3755 6857
rect 3182 6733 3199 6767
rect 3233 6733 3252 6767
rect 3182 6718 3252 6733
rect 4106 6803 4174 6820
rect 4106 6769 4123 6803
rect 4157 6769 4174 6803
rect 3697 6673 3755 6690
rect 1121 6608 1139 6642
rect 1173 6608 1311 6642
rect 1345 6608 1363 6642
rect 1121 6545 1363 6608
rect 1397 6640 2466 6654
rect 1397 6606 1415 6640
rect 1449 6606 2415 6640
rect 2449 6606 2466 6640
rect 1397 6545 2466 6606
rect 2501 6640 3570 6654
rect 2501 6606 2519 6640
rect 2553 6606 3519 6640
rect 3553 6606 3570 6640
rect 2501 6545 3570 6606
rect 3697 6639 3709 6673
rect 3743 6639 3755 6673
rect 4106 6654 4174 6769
rect 4470 6767 4540 6968
rect 4470 6733 4487 6767
rect 4521 6733 4540 6767
rect 4470 6718 4540 6733
rect 5210 6803 5278 6820
rect 5210 6769 5227 6803
rect 5261 6769 5278 6803
rect 5210 6654 5278 6769
rect 5574 6767 5644 6968
rect 5574 6733 5591 6767
rect 5625 6733 5644 6767
rect 5574 6718 5644 6733
rect 6314 6803 6382 6820
rect 6314 6769 6331 6803
rect 6365 6769 6382 6803
rect 6314 6654 6382 6769
rect 6678 6767 6748 6968
rect 6678 6733 6695 6767
rect 6729 6733 6748 6767
rect 6678 6718 6748 6733
rect 7418 6803 7486 6820
rect 7418 6769 7435 6803
rect 7469 6769 7486 6803
rect 7418 6654 7486 6769
rect 7782 6767 7852 6968
rect 8205 6911 8723 6979
rect 8205 6877 8223 6911
rect 8257 6877 8671 6911
rect 8705 6877 8723 6911
rect 8205 6837 8723 6877
rect 7782 6733 7799 6767
rect 7833 6733 7852 6767
rect 7782 6718 7852 6733
rect 8205 6769 8283 6803
rect 8317 6769 8393 6803
rect 8427 6769 8447 6803
rect 8205 6699 8447 6769
rect 8481 6767 8723 6837
rect 8849 6984 8907 7055
rect 8849 6950 8861 6984
rect 8895 6950 8907 6984
rect 8941 7013 10010 7055
rect 8941 6979 8959 7013
rect 8993 6979 9959 7013
rect 9993 6979 10010 7013
rect 8941 6968 10010 6979
rect 10045 7013 11114 7055
rect 10045 6979 10063 7013
rect 10097 6979 11063 7013
rect 11097 6979 11114 7013
rect 10045 6968 11114 6979
rect 11149 7013 12218 7055
rect 11149 6979 11167 7013
rect 11201 6979 12167 7013
rect 12201 6979 12218 7013
rect 11149 6968 12218 6979
rect 12253 7013 13322 7055
rect 12253 6979 12271 7013
rect 12305 6979 13271 7013
rect 13305 6979 13322 7013
rect 12253 6968 13322 6979
rect 13357 7013 13875 7055
rect 13357 6979 13375 7013
rect 13409 6979 13823 7013
rect 13857 6979 13875 7013
rect 8849 6891 8907 6950
rect 8849 6857 8861 6891
rect 8895 6857 8907 6891
rect 8849 6822 8907 6857
rect 8481 6733 8501 6767
rect 8535 6733 8611 6767
rect 8645 6733 8723 6767
rect 9258 6803 9326 6820
rect 9258 6769 9275 6803
rect 9309 6769 9326 6803
rect 3697 6545 3755 6639
rect 3789 6640 4858 6654
rect 3789 6606 3807 6640
rect 3841 6606 4807 6640
rect 4841 6606 4858 6640
rect 3789 6545 4858 6606
rect 4893 6640 5962 6654
rect 4893 6606 4911 6640
rect 4945 6606 5911 6640
rect 5945 6606 5962 6640
rect 4893 6545 5962 6606
rect 5997 6640 7066 6654
rect 5997 6606 6015 6640
rect 6049 6606 7015 6640
rect 7049 6606 7066 6640
rect 5997 6545 7066 6606
rect 7101 6640 8170 6654
rect 7101 6606 7119 6640
rect 7153 6606 8119 6640
rect 8153 6606 8170 6640
rect 7101 6545 8170 6606
rect 8205 6640 8723 6699
rect 8205 6606 8223 6640
rect 8257 6606 8671 6640
rect 8705 6606 8723 6640
rect 8205 6545 8723 6606
rect 8849 6673 8907 6690
rect 8849 6639 8861 6673
rect 8895 6639 8907 6673
rect 9258 6654 9326 6769
rect 9622 6767 9692 6968
rect 9622 6733 9639 6767
rect 9673 6733 9692 6767
rect 9622 6718 9692 6733
rect 10362 6803 10430 6820
rect 10362 6769 10379 6803
rect 10413 6769 10430 6803
rect 10362 6654 10430 6769
rect 10726 6767 10796 6968
rect 10726 6733 10743 6767
rect 10777 6733 10796 6767
rect 10726 6718 10796 6733
rect 11466 6803 11534 6820
rect 11466 6769 11483 6803
rect 11517 6769 11534 6803
rect 11466 6654 11534 6769
rect 11830 6767 11900 6968
rect 11830 6733 11847 6767
rect 11881 6733 11900 6767
rect 11830 6718 11900 6733
rect 12570 6803 12638 6820
rect 12570 6769 12587 6803
rect 12621 6769 12638 6803
rect 12570 6654 12638 6769
rect 12934 6767 13004 6968
rect 13357 6911 13875 6979
rect 13357 6877 13375 6911
rect 13409 6877 13823 6911
rect 13857 6877 13875 6911
rect 13357 6837 13875 6877
rect 12934 6733 12951 6767
rect 12985 6733 13004 6767
rect 12934 6718 13004 6733
rect 13357 6769 13435 6803
rect 13469 6769 13545 6803
rect 13579 6769 13599 6803
rect 13357 6699 13599 6769
rect 13633 6767 13875 6837
rect 14001 6984 14059 7055
rect 14001 6950 14013 6984
rect 14047 6950 14059 6984
rect 14093 7013 15162 7055
rect 14093 6979 14111 7013
rect 14145 6979 15111 7013
rect 15145 6979 15162 7013
rect 14093 6968 15162 6979
rect 15197 7013 16266 7055
rect 15197 6979 15215 7013
rect 15249 6979 16215 7013
rect 16249 6979 16266 7013
rect 15197 6968 16266 6979
rect 16301 7013 17370 7055
rect 16301 6979 16319 7013
rect 16353 6979 17319 7013
rect 17353 6979 17370 7013
rect 16301 6968 17370 6979
rect 17405 7013 18474 7055
rect 17405 6979 17423 7013
rect 17457 6979 18423 7013
rect 18457 6979 18474 7013
rect 17405 6968 18474 6979
rect 18601 7013 18843 7055
rect 18601 6979 18619 7013
rect 18653 6979 18791 7013
rect 18825 6979 18843 7013
rect 14001 6891 14059 6950
rect 14001 6857 14013 6891
rect 14047 6857 14059 6891
rect 14001 6822 14059 6857
rect 13633 6733 13653 6767
rect 13687 6733 13763 6767
rect 13797 6733 13875 6767
rect 14410 6803 14478 6820
rect 14410 6769 14427 6803
rect 14461 6769 14478 6803
rect 8849 6545 8907 6639
rect 8941 6640 10010 6654
rect 8941 6606 8959 6640
rect 8993 6606 9959 6640
rect 9993 6606 10010 6640
rect 8941 6545 10010 6606
rect 10045 6640 11114 6654
rect 10045 6606 10063 6640
rect 10097 6606 11063 6640
rect 11097 6606 11114 6640
rect 10045 6545 11114 6606
rect 11149 6640 12218 6654
rect 11149 6606 11167 6640
rect 11201 6606 12167 6640
rect 12201 6606 12218 6640
rect 11149 6545 12218 6606
rect 12253 6640 13322 6654
rect 12253 6606 12271 6640
rect 12305 6606 13271 6640
rect 13305 6606 13322 6640
rect 12253 6545 13322 6606
rect 13357 6640 13875 6699
rect 13357 6606 13375 6640
rect 13409 6606 13823 6640
rect 13857 6606 13875 6640
rect 13357 6545 13875 6606
rect 14001 6673 14059 6690
rect 14001 6639 14013 6673
rect 14047 6639 14059 6673
rect 14410 6654 14478 6769
rect 14774 6767 14844 6968
rect 14774 6733 14791 6767
rect 14825 6733 14844 6767
rect 14774 6718 14844 6733
rect 15514 6803 15582 6820
rect 15514 6769 15531 6803
rect 15565 6769 15582 6803
rect 15514 6654 15582 6769
rect 15878 6767 15948 6968
rect 15878 6733 15895 6767
rect 15929 6733 15948 6767
rect 15878 6718 15948 6733
rect 16618 6803 16686 6820
rect 16618 6769 16635 6803
rect 16669 6769 16686 6803
rect 16618 6654 16686 6769
rect 16982 6767 17052 6968
rect 16982 6733 16999 6767
rect 17033 6733 17052 6767
rect 16982 6718 17052 6733
rect 17722 6803 17790 6820
rect 17722 6769 17739 6803
rect 17773 6769 17790 6803
rect 17722 6654 17790 6769
rect 18086 6767 18156 6968
rect 18086 6733 18103 6767
rect 18137 6733 18156 6767
rect 18086 6718 18156 6733
rect 18601 6918 18843 6979
rect 18601 6884 18619 6918
rect 18653 6884 18791 6918
rect 18825 6884 18843 6918
rect 18601 6837 18843 6884
rect 18601 6763 18705 6837
rect 18601 6729 18651 6763
rect 18685 6729 18705 6763
rect 18739 6769 18759 6803
rect 18793 6769 18843 6803
rect 18739 6695 18843 6769
rect 14001 6545 14059 6639
rect 14093 6640 15162 6654
rect 14093 6606 14111 6640
rect 14145 6606 15111 6640
rect 15145 6606 15162 6640
rect 14093 6545 15162 6606
rect 15197 6640 16266 6654
rect 15197 6606 15215 6640
rect 15249 6606 16215 6640
rect 16249 6606 16266 6640
rect 15197 6545 16266 6606
rect 16301 6640 17370 6654
rect 16301 6606 16319 6640
rect 16353 6606 17319 6640
rect 17353 6606 17370 6640
rect 16301 6545 17370 6606
rect 17405 6640 18474 6654
rect 17405 6606 17423 6640
rect 17457 6606 18423 6640
rect 18457 6606 18474 6640
rect 17405 6545 18474 6606
rect 18601 6642 18843 6695
rect 18601 6608 18619 6642
rect 18653 6608 18791 6642
rect 18825 6608 18843 6642
rect 18601 6545 18843 6608
rect 1104 6511 1133 6545
rect 1167 6511 1225 6545
rect 1259 6511 1317 6545
rect 1351 6511 1409 6545
rect 1443 6511 1501 6545
rect 1535 6511 1593 6545
rect 1627 6511 1685 6545
rect 1719 6511 1777 6545
rect 1811 6511 1869 6545
rect 1903 6511 1961 6545
rect 1995 6511 2053 6545
rect 2087 6511 2145 6545
rect 2179 6511 2237 6545
rect 2271 6511 2329 6545
rect 2363 6511 2421 6545
rect 2455 6511 2513 6545
rect 2547 6511 2605 6545
rect 2639 6511 2697 6545
rect 2731 6511 2789 6545
rect 2823 6511 2881 6545
rect 2915 6511 2973 6545
rect 3007 6511 3065 6545
rect 3099 6511 3157 6545
rect 3191 6511 3249 6545
rect 3283 6511 3341 6545
rect 3375 6511 3433 6545
rect 3467 6511 3525 6545
rect 3559 6511 3617 6545
rect 3651 6511 3709 6545
rect 3743 6511 3801 6545
rect 3835 6511 3893 6545
rect 3927 6511 3985 6545
rect 4019 6511 4077 6545
rect 4111 6511 4169 6545
rect 4203 6511 4261 6545
rect 4295 6511 4353 6545
rect 4387 6511 4445 6545
rect 4479 6511 4537 6545
rect 4571 6511 4629 6545
rect 4663 6511 4721 6545
rect 4755 6511 4813 6545
rect 4847 6511 4905 6545
rect 4939 6511 4997 6545
rect 5031 6511 5089 6545
rect 5123 6511 5181 6545
rect 5215 6511 5273 6545
rect 5307 6511 5365 6545
rect 5399 6511 5457 6545
rect 5491 6511 5549 6545
rect 5583 6511 5641 6545
rect 5675 6511 5733 6545
rect 5767 6511 5825 6545
rect 5859 6511 5917 6545
rect 5951 6511 6009 6545
rect 6043 6511 6101 6545
rect 6135 6511 6193 6545
rect 6227 6511 6285 6545
rect 6319 6511 6377 6545
rect 6411 6511 6469 6545
rect 6503 6511 6561 6545
rect 6595 6511 6653 6545
rect 6687 6511 6745 6545
rect 6779 6511 6837 6545
rect 6871 6511 6929 6545
rect 6963 6511 7021 6545
rect 7055 6511 7113 6545
rect 7147 6511 7205 6545
rect 7239 6511 7297 6545
rect 7331 6511 7389 6545
rect 7423 6511 7481 6545
rect 7515 6511 7573 6545
rect 7607 6511 7665 6545
rect 7699 6511 7757 6545
rect 7791 6511 7849 6545
rect 7883 6511 7941 6545
rect 7975 6511 8033 6545
rect 8067 6511 8125 6545
rect 8159 6511 8217 6545
rect 8251 6511 8309 6545
rect 8343 6511 8401 6545
rect 8435 6511 8493 6545
rect 8527 6511 8585 6545
rect 8619 6511 8677 6545
rect 8711 6511 8769 6545
rect 8803 6511 8861 6545
rect 8895 6511 8953 6545
rect 8987 6511 9045 6545
rect 9079 6511 9137 6545
rect 9171 6511 9229 6545
rect 9263 6511 9321 6545
rect 9355 6511 9413 6545
rect 9447 6511 9505 6545
rect 9539 6511 9597 6545
rect 9631 6511 9689 6545
rect 9723 6511 9781 6545
rect 9815 6511 9873 6545
rect 9907 6511 9965 6545
rect 9999 6511 10057 6545
rect 10091 6511 10149 6545
rect 10183 6511 10241 6545
rect 10275 6511 10333 6545
rect 10367 6511 10425 6545
rect 10459 6511 10517 6545
rect 10551 6511 10609 6545
rect 10643 6511 10701 6545
rect 10735 6511 10793 6545
rect 10827 6511 10885 6545
rect 10919 6511 10977 6545
rect 11011 6511 11069 6545
rect 11103 6511 11161 6545
rect 11195 6511 11253 6545
rect 11287 6511 11345 6545
rect 11379 6511 11437 6545
rect 11471 6511 11529 6545
rect 11563 6511 11621 6545
rect 11655 6511 11713 6545
rect 11747 6511 11805 6545
rect 11839 6511 11897 6545
rect 11931 6511 11989 6545
rect 12023 6511 12081 6545
rect 12115 6511 12173 6545
rect 12207 6511 12265 6545
rect 12299 6511 12357 6545
rect 12391 6511 12449 6545
rect 12483 6511 12541 6545
rect 12575 6511 12633 6545
rect 12667 6511 12725 6545
rect 12759 6511 12817 6545
rect 12851 6511 12909 6545
rect 12943 6511 13001 6545
rect 13035 6511 13093 6545
rect 13127 6511 13185 6545
rect 13219 6511 13277 6545
rect 13311 6511 13369 6545
rect 13403 6511 13461 6545
rect 13495 6511 13553 6545
rect 13587 6511 13645 6545
rect 13679 6511 13737 6545
rect 13771 6511 13829 6545
rect 13863 6511 13921 6545
rect 13955 6511 14013 6545
rect 14047 6511 14105 6545
rect 14139 6511 14197 6545
rect 14231 6511 14289 6545
rect 14323 6511 14381 6545
rect 14415 6511 14473 6545
rect 14507 6511 14565 6545
rect 14599 6511 14657 6545
rect 14691 6511 14749 6545
rect 14783 6511 14841 6545
rect 14875 6511 14933 6545
rect 14967 6511 15025 6545
rect 15059 6511 15117 6545
rect 15151 6511 15209 6545
rect 15243 6511 15301 6545
rect 15335 6511 15393 6545
rect 15427 6511 15485 6545
rect 15519 6511 15577 6545
rect 15611 6511 15669 6545
rect 15703 6511 15761 6545
rect 15795 6511 15853 6545
rect 15887 6511 15945 6545
rect 15979 6511 16037 6545
rect 16071 6511 16129 6545
rect 16163 6511 16221 6545
rect 16255 6511 16313 6545
rect 16347 6511 16405 6545
rect 16439 6511 16497 6545
rect 16531 6511 16589 6545
rect 16623 6511 16681 6545
rect 16715 6511 16773 6545
rect 16807 6511 16865 6545
rect 16899 6511 16957 6545
rect 16991 6511 17049 6545
rect 17083 6511 17141 6545
rect 17175 6511 17233 6545
rect 17267 6511 17325 6545
rect 17359 6511 17417 6545
rect 17451 6511 17509 6545
rect 17543 6511 17601 6545
rect 17635 6511 17693 6545
rect 17727 6511 17785 6545
rect 17819 6511 17877 6545
rect 17911 6511 17969 6545
rect 18003 6511 18061 6545
rect 18095 6511 18153 6545
rect 18187 6511 18245 6545
rect 18279 6511 18337 6545
rect 18371 6511 18429 6545
rect 18463 6511 18521 6545
rect 18555 6511 18613 6545
rect 18647 6511 18705 6545
rect 18739 6511 18797 6545
rect 18831 6511 18860 6545
rect 1121 6448 1363 6511
rect 1121 6414 1139 6448
rect 1173 6414 1311 6448
rect 1345 6414 1363 6448
rect 1121 6361 1363 6414
rect 1397 6450 2466 6511
rect 1397 6416 1415 6450
rect 1449 6416 2415 6450
rect 2449 6416 2466 6450
rect 1397 6402 2466 6416
rect 2501 6450 3570 6511
rect 2501 6416 2519 6450
rect 2553 6416 3519 6450
rect 3553 6416 3570 6450
rect 2501 6402 3570 6416
rect 3605 6450 4674 6511
rect 3605 6416 3623 6450
rect 3657 6416 4623 6450
rect 4657 6416 4674 6450
rect 3605 6402 4674 6416
rect 4709 6450 5778 6511
rect 4709 6416 4727 6450
rect 4761 6416 5727 6450
rect 5761 6416 5778 6450
rect 4709 6402 5778 6416
rect 5813 6443 6147 6511
rect 5813 6409 5831 6443
rect 5865 6409 6095 6443
rect 6129 6409 6147 6443
rect 1121 6287 1225 6361
rect 1121 6253 1171 6287
rect 1205 6253 1225 6287
rect 1259 6293 1279 6327
rect 1313 6293 1363 6327
rect 1259 6219 1363 6293
rect 1714 6287 1782 6402
rect 1714 6253 1731 6287
rect 1765 6253 1782 6287
rect 1714 6236 1782 6253
rect 2078 6323 2148 6338
rect 2078 6289 2095 6323
rect 2129 6289 2148 6323
rect 1121 6172 1363 6219
rect 1121 6138 1139 6172
rect 1173 6138 1311 6172
rect 1345 6138 1363 6172
rect 1121 6077 1363 6138
rect 2078 6088 2148 6289
rect 2818 6287 2886 6402
rect 2818 6253 2835 6287
rect 2869 6253 2886 6287
rect 2818 6236 2886 6253
rect 3182 6323 3252 6338
rect 3182 6289 3199 6323
rect 3233 6289 3252 6323
rect 3182 6088 3252 6289
rect 3922 6287 3990 6402
rect 3922 6253 3939 6287
rect 3973 6253 3990 6287
rect 3922 6236 3990 6253
rect 4286 6323 4356 6338
rect 4286 6289 4303 6323
rect 4337 6289 4356 6323
rect 4286 6088 4356 6289
rect 5026 6287 5094 6402
rect 5813 6357 6147 6409
rect 6273 6417 6331 6511
rect 6273 6383 6285 6417
rect 6319 6383 6331 6417
rect 6365 6450 7434 6511
rect 6365 6416 6383 6450
rect 6417 6416 7383 6450
rect 7417 6416 7434 6450
rect 6365 6402 7434 6416
rect 7469 6450 7987 6511
rect 7469 6416 7487 6450
rect 7521 6416 7935 6450
rect 7969 6416 7987 6450
rect 6273 6366 6331 6383
rect 5026 6253 5043 6287
rect 5077 6253 5094 6287
rect 5026 6236 5094 6253
rect 5390 6323 5460 6338
rect 5390 6289 5407 6323
rect 5441 6289 5460 6323
rect 5390 6088 5460 6289
rect 5813 6287 5963 6357
rect 5813 6253 5833 6287
rect 5867 6253 5963 6287
rect 5997 6289 6093 6323
rect 6127 6289 6147 6323
rect 5997 6219 6147 6289
rect 6682 6287 6750 6402
rect 7469 6357 7987 6416
rect 8054 6459 8102 6511
rect 8054 6425 8068 6459
rect 8054 6409 8102 6425
rect 8138 6459 8194 6475
rect 8138 6425 8152 6459
rect 8186 6425 8194 6459
rect 8138 6409 8194 6425
rect 8240 6459 8283 6511
rect 8240 6425 8248 6459
rect 8282 6425 8283 6459
rect 8240 6409 8283 6425
rect 8317 6467 8440 6477
rect 8317 6433 8333 6467
rect 8367 6433 8440 6467
rect 6682 6253 6699 6287
rect 6733 6253 6750 6287
rect 6682 6236 6750 6253
rect 7046 6323 7116 6338
rect 7046 6289 7063 6323
rect 7097 6289 7116 6323
rect 5813 6179 6147 6219
rect 5813 6145 5831 6179
rect 5865 6145 6095 6179
rect 6129 6145 6147 6179
rect 1121 6043 1139 6077
rect 1173 6043 1311 6077
rect 1345 6043 1363 6077
rect 1121 6001 1363 6043
rect 1397 6077 2466 6088
rect 1397 6043 1415 6077
rect 1449 6043 2415 6077
rect 2449 6043 2466 6077
rect 1397 6001 2466 6043
rect 2501 6077 3570 6088
rect 2501 6043 2519 6077
rect 2553 6043 3519 6077
rect 3553 6043 3570 6077
rect 2501 6001 3570 6043
rect 3605 6077 4674 6088
rect 3605 6043 3623 6077
rect 3657 6043 4623 6077
rect 4657 6043 4674 6077
rect 3605 6001 4674 6043
rect 4709 6077 5778 6088
rect 4709 6043 4727 6077
rect 4761 6043 5727 6077
rect 5761 6043 5778 6077
rect 4709 6001 5778 6043
rect 5813 6077 6147 6145
rect 5813 6043 5831 6077
rect 5865 6043 6095 6077
rect 6129 6043 6147 6077
rect 5813 6001 6147 6043
rect 6273 6199 6331 6234
rect 6273 6165 6285 6199
rect 6319 6165 6331 6199
rect 6273 6106 6331 6165
rect 6273 6072 6285 6106
rect 6319 6072 6331 6106
rect 7046 6088 7116 6289
rect 7469 6287 7711 6357
rect 7469 6253 7547 6287
rect 7581 6253 7657 6287
rect 7691 6253 7711 6287
rect 7745 6289 7765 6323
rect 7799 6289 7875 6323
rect 7909 6289 7987 6323
rect 7745 6219 7987 6289
rect 8033 6313 8104 6375
rect 8033 6307 8070 6313
rect 8067 6279 8070 6307
rect 8067 6273 8104 6279
rect 8033 6263 8104 6273
rect 8138 6229 8172 6409
rect 8317 6399 8440 6433
rect 8481 6450 9550 6511
rect 8481 6416 8499 6450
rect 8533 6416 9499 6450
rect 9533 6416 9550 6450
rect 8481 6402 9550 6416
rect 9585 6450 10654 6511
rect 9585 6416 9603 6450
rect 9637 6416 10603 6450
rect 10637 6416 10654 6450
rect 9585 6402 10654 6416
rect 10689 6450 11391 6511
rect 10689 6416 10707 6450
rect 10741 6416 11339 6450
rect 11373 6416 11391 6450
rect 8206 6313 8259 6375
rect 8317 6365 8333 6399
rect 8367 6365 8440 6399
rect 8317 6363 8440 6365
rect 8240 6307 8259 6313
rect 8206 6273 8217 6279
rect 8251 6273 8259 6307
rect 8206 6263 8259 6273
rect 8309 6313 8343 6329
rect 8309 6229 8343 6279
rect 7469 6179 7987 6219
rect 7469 6145 7487 6179
rect 7521 6145 7935 6179
rect 7969 6145 7987 6179
rect 8058 6213 8343 6229
rect 8058 6179 8080 6213
rect 8114 6195 8343 6213
rect 8114 6179 8136 6195
rect 8058 6160 8136 6179
rect 6273 6001 6331 6072
rect 6365 6077 7434 6088
rect 6365 6043 6383 6077
rect 6417 6043 7383 6077
rect 7417 6043 7434 6077
rect 6365 6001 7434 6043
rect 7469 6077 7987 6145
rect 7469 6043 7487 6077
rect 7521 6043 7935 6077
rect 7969 6043 7987 6077
rect 7469 6001 7987 6043
rect 8233 6127 8249 6161
rect 8283 6127 8299 6161
rect 8377 6159 8440 6363
rect 8798 6287 8866 6402
rect 8798 6253 8815 6287
rect 8849 6253 8866 6287
rect 8798 6236 8866 6253
rect 9162 6323 9232 6338
rect 9162 6289 9179 6323
rect 9213 6289 9232 6323
rect 8233 6093 8299 6127
rect 8233 6059 8249 6093
rect 8283 6059 8299 6093
rect 8233 6001 8299 6059
rect 8333 6145 8440 6159
rect 8333 6111 8349 6145
rect 8383 6111 8440 6145
rect 8333 6103 8440 6111
rect 8333 6077 8401 6103
rect 8333 6043 8349 6077
rect 8383 6069 8401 6077
rect 8435 6069 8440 6103
rect 9162 6088 9232 6289
rect 9902 6287 9970 6402
rect 10689 6357 11391 6416
rect 11425 6417 11483 6511
rect 11425 6383 11437 6417
rect 11471 6383 11483 6417
rect 11517 6450 12586 6511
rect 11517 6416 11535 6450
rect 11569 6416 12535 6450
rect 12569 6416 12586 6450
rect 11517 6402 12586 6416
rect 12621 6450 13690 6511
rect 12621 6416 12639 6450
rect 12673 6416 13639 6450
rect 13673 6416 13690 6450
rect 12621 6402 13690 6416
rect 13725 6450 14794 6511
rect 13725 6416 13743 6450
rect 13777 6416 14743 6450
rect 14777 6416 14794 6450
rect 13725 6402 14794 6416
rect 14829 6450 15898 6511
rect 14829 6416 14847 6450
rect 14881 6416 15847 6450
rect 15881 6416 15898 6450
rect 14829 6402 15898 6416
rect 15933 6450 16451 6511
rect 15933 6416 15951 6450
rect 15985 6416 16399 6450
rect 16433 6416 16451 6450
rect 11425 6366 11483 6383
rect 9902 6253 9919 6287
rect 9953 6253 9970 6287
rect 9902 6236 9970 6253
rect 10266 6323 10336 6338
rect 10266 6289 10283 6323
rect 10317 6289 10336 6323
rect 10266 6088 10336 6289
rect 10689 6287 11019 6357
rect 10689 6253 10767 6287
rect 10801 6253 10866 6287
rect 10900 6253 10965 6287
rect 10999 6253 11019 6287
rect 11053 6289 11073 6323
rect 11107 6289 11176 6323
rect 11210 6289 11279 6323
rect 11313 6289 11391 6323
rect 11053 6219 11391 6289
rect 11834 6287 11902 6402
rect 11834 6253 11851 6287
rect 11885 6253 11902 6287
rect 11834 6236 11902 6253
rect 12198 6323 12268 6338
rect 12198 6289 12215 6323
rect 12249 6289 12268 6323
rect 10689 6179 11391 6219
rect 10689 6145 10707 6179
rect 10741 6145 11339 6179
rect 11373 6145 11391 6179
rect 8383 6043 8440 6069
rect 8333 6035 8440 6043
rect 8481 6077 9550 6088
rect 8481 6043 8499 6077
rect 8533 6043 9499 6077
rect 9533 6043 9550 6077
rect 8481 6001 9550 6043
rect 9585 6077 10654 6088
rect 9585 6043 9603 6077
rect 9637 6043 10603 6077
rect 10637 6043 10654 6077
rect 9585 6001 10654 6043
rect 10689 6077 11391 6145
rect 10689 6043 10707 6077
rect 10741 6043 11339 6077
rect 11373 6043 11391 6077
rect 10689 6001 11391 6043
rect 11425 6199 11483 6234
rect 11425 6165 11437 6199
rect 11471 6165 11483 6199
rect 11425 6106 11483 6165
rect 11425 6072 11437 6106
rect 11471 6072 11483 6106
rect 12198 6088 12268 6289
rect 12938 6287 13006 6402
rect 12938 6253 12955 6287
rect 12989 6253 13006 6287
rect 12938 6236 13006 6253
rect 13302 6323 13372 6338
rect 13302 6289 13319 6323
rect 13353 6289 13372 6323
rect 13302 6088 13372 6289
rect 14042 6287 14110 6402
rect 14042 6253 14059 6287
rect 14093 6253 14110 6287
rect 14042 6236 14110 6253
rect 14406 6323 14476 6338
rect 14406 6289 14423 6323
rect 14457 6289 14476 6323
rect 14406 6088 14476 6289
rect 15146 6287 15214 6402
rect 15933 6357 16451 6416
rect 16577 6417 16635 6511
rect 16577 6383 16589 6417
rect 16623 6383 16635 6417
rect 16669 6450 17738 6511
rect 16669 6416 16687 6450
rect 16721 6416 17687 6450
rect 17721 6416 17738 6450
rect 16669 6402 17738 6416
rect 17773 6450 18475 6511
rect 17773 6416 17791 6450
rect 17825 6416 18423 6450
rect 18457 6416 18475 6450
rect 16577 6366 16635 6383
rect 15146 6253 15163 6287
rect 15197 6253 15214 6287
rect 15146 6236 15214 6253
rect 15510 6323 15580 6338
rect 15510 6289 15527 6323
rect 15561 6289 15580 6323
rect 15510 6088 15580 6289
rect 15933 6287 16175 6357
rect 15933 6253 16011 6287
rect 16045 6253 16121 6287
rect 16155 6253 16175 6287
rect 16209 6289 16229 6323
rect 16263 6289 16339 6323
rect 16373 6289 16451 6323
rect 16209 6219 16451 6289
rect 16986 6287 17054 6402
rect 17773 6357 18475 6416
rect 18601 6448 18843 6511
rect 18601 6414 18619 6448
rect 18653 6414 18791 6448
rect 18825 6414 18843 6448
rect 18601 6361 18843 6414
rect 16986 6253 17003 6287
rect 17037 6253 17054 6287
rect 16986 6236 17054 6253
rect 17350 6323 17420 6338
rect 17350 6289 17367 6323
rect 17401 6289 17420 6323
rect 15933 6179 16451 6219
rect 15933 6145 15951 6179
rect 15985 6145 16399 6179
rect 16433 6145 16451 6179
rect 11425 6001 11483 6072
rect 11517 6077 12586 6088
rect 11517 6043 11535 6077
rect 11569 6043 12535 6077
rect 12569 6043 12586 6077
rect 11517 6001 12586 6043
rect 12621 6077 13690 6088
rect 12621 6043 12639 6077
rect 12673 6043 13639 6077
rect 13673 6043 13690 6077
rect 12621 6001 13690 6043
rect 13725 6077 14794 6088
rect 13725 6043 13743 6077
rect 13777 6043 14743 6077
rect 14777 6043 14794 6077
rect 13725 6001 14794 6043
rect 14829 6077 15898 6088
rect 14829 6043 14847 6077
rect 14881 6043 15847 6077
rect 15881 6043 15898 6077
rect 14829 6001 15898 6043
rect 15933 6077 16451 6145
rect 15933 6043 15951 6077
rect 15985 6043 16399 6077
rect 16433 6043 16451 6077
rect 15933 6001 16451 6043
rect 16577 6199 16635 6234
rect 16577 6165 16589 6199
rect 16623 6165 16635 6199
rect 16577 6106 16635 6165
rect 16577 6072 16589 6106
rect 16623 6072 16635 6106
rect 17350 6088 17420 6289
rect 17773 6287 18103 6357
rect 17773 6253 17851 6287
rect 17885 6253 17950 6287
rect 17984 6253 18049 6287
rect 18083 6253 18103 6287
rect 18137 6289 18157 6323
rect 18191 6289 18260 6323
rect 18294 6289 18363 6323
rect 18397 6289 18475 6323
rect 18137 6219 18475 6289
rect 17773 6179 18475 6219
rect 17773 6145 17791 6179
rect 17825 6145 18423 6179
rect 18457 6145 18475 6179
rect 16577 6001 16635 6072
rect 16669 6077 17738 6088
rect 16669 6043 16687 6077
rect 16721 6043 17687 6077
rect 17721 6043 17738 6077
rect 16669 6001 17738 6043
rect 17773 6077 18475 6145
rect 17773 6043 17791 6077
rect 17825 6043 18423 6077
rect 18457 6043 18475 6077
rect 17773 6001 18475 6043
rect 18601 6293 18651 6327
rect 18685 6293 18705 6327
rect 18601 6219 18705 6293
rect 18739 6287 18843 6361
rect 18739 6253 18759 6287
rect 18793 6253 18843 6287
rect 18601 6172 18843 6219
rect 18601 6138 18619 6172
rect 18653 6138 18791 6172
rect 18825 6138 18843 6172
rect 18601 6077 18843 6138
rect 18601 6043 18619 6077
rect 18653 6043 18791 6077
rect 18825 6043 18843 6077
rect 18601 6001 18843 6043
rect 1104 5967 1133 6001
rect 1167 5967 1225 6001
rect 1259 5967 1317 6001
rect 1351 5967 1409 6001
rect 1443 5967 1501 6001
rect 1535 5967 1593 6001
rect 1627 5967 1685 6001
rect 1719 5967 1777 6001
rect 1811 5967 1869 6001
rect 1903 5967 1961 6001
rect 1995 5967 2053 6001
rect 2087 5967 2145 6001
rect 2179 5967 2237 6001
rect 2271 5967 2329 6001
rect 2363 5967 2421 6001
rect 2455 5967 2513 6001
rect 2547 5967 2605 6001
rect 2639 5967 2697 6001
rect 2731 5967 2789 6001
rect 2823 5967 2881 6001
rect 2915 5967 2973 6001
rect 3007 5967 3065 6001
rect 3099 5967 3157 6001
rect 3191 5967 3249 6001
rect 3283 5967 3341 6001
rect 3375 5967 3433 6001
rect 3467 5967 3525 6001
rect 3559 5967 3617 6001
rect 3651 5967 3709 6001
rect 3743 5967 3801 6001
rect 3835 5967 3893 6001
rect 3927 5967 3985 6001
rect 4019 5967 4077 6001
rect 4111 5967 4169 6001
rect 4203 5967 4261 6001
rect 4295 5967 4353 6001
rect 4387 5967 4445 6001
rect 4479 5967 4537 6001
rect 4571 5967 4629 6001
rect 4663 5967 4721 6001
rect 4755 5967 4813 6001
rect 4847 5967 4905 6001
rect 4939 5967 4997 6001
rect 5031 5967 5089 6001
rect 5123 5967 5181 6001
rect 5215 5967 5273 6001
rect 5307 5967 5365 6001
rect 5399 5967 5457 6001
rect 5491 5967 5549 6001
rect 5583 5967 5641 6001
rect 5675 5967 5733 6001
rect 5767 5967 5825 6001
rect 5859 5967 5917 6001
rect 5951 5967 6009 6001
rect 6043 5967 6101 6001
rect 6135 5967 6193 6001
rect 6227 5967 6285 6001
rect 6319 5967 6377 6001
rect 6411 5967 6469 6001
rect 6503 5967 6561 6001
rect 6595 5967 6653 6001
rect 6687 5967 6745 6001
rect 6779 5967 6837 6001
rect 6871 5967 6929 6001
rect 6963 5967 7021 6001
rect 7055 5967 7113 6001
rect 7147 5967 7205 6001
rect 7239 5967 7297 6001
rect 7331 5967 7389 6001
rect 7423 5967 7481 6001
rect 7515 5967 7573 6001
rect 7607 5967 7665 6001
rect 7699 5967 7757 6001
rect 7791 5967 7849 6001
rect 7883 5967 7941 6001
rect 7975 5967 8033 6001
rect 8067 5967 8125 6001
rect 8159 5967 8217 6001
rect 8251 5967 8309 6001
rect 8343 5967 8401 6001
rect 8435 5967 8493 6001
rect 8527 5967 8585 6001
rect 8619 5967 8677 6001
rect 8711 5967 8769 6001
rect 8803 5967 8861 6001
rect 8895 5967 8953 6001
rect 8987 5967 9045 6001
rect 9079 5967 9137 6001
rect 9171 5967 9229 6001
rect 9263 5967 9321 6001
rect 9355 5967 9413 6001
rect 9447 5967 9505 6001
rect 9539 5967 9597 6001
rect 9631 5967 9689 6001
rect 9723 5967 9781 6001
rect 9815 5967 9873 6001
rect 9907 5967 9965 6001
rect 9999 5967 10057 6001
rect 10091 5967 10149 6001
rect 10183 5967 10241 6001
rect 10275 5967 10333 6001
rect 10367 5967 10425 6001
rect 10459 5967 10517 6001
rect 10551 5967 10609 6001
rect 10643 5967 10701 6001
rect 10735 5967 10793 6001
rect 10827 5967 10885 6001
rect 10919 5967 10977 6001
rect 11011 5967 11069 6001
rect 11103 5967 11161 6001
rect 11195 5967 11253 6001
rect 11287 5967 11345 6001
rect 11379 5967 11437 6001
rect 11471 5967 11529 6001
rect 11563 5967 11621 6001
rect 11655 5967 11713 6001
rect 11747 5967 11805 6001
rect 11839 5967 11897 6001
rect 11931 5967 11989 6001
rect 12023 5967 12081 6001
rect 12115 5967 12173 6001
rect 12207 5967 12265 6001
rect 12299 5967 12357 6001
rect 12391 5967 12449 6001
rect 12483 5967 12541 6001
rect 12575 5967 12633 6001
rect 12667 5967 12725 6001
rect 12759 5967 12817 6001
rect 12851 5967 12909 6001
rect 12943 5967 13001 6001
rect 13035 5967 13093 6001
rect 13127 5967 13185 6001
rect 13219 5967 13277 6001
rect 13311 5967 13369 6001
rect 13403 5967 13461 6001
rect 13495 5967 13553 6001
rect 13587 5967 13645 6001
rect 13679 5967 13737 6001
rect 13771 5967 13829 6001
rect 13863 5967 13921 6001
rect 13955 5967 14013 6001
rect 14047 5967 14105 6001
rect 14139 5967 14197 6001
rect 14231 5967 14289 6001
rect 14323 5967 14381 6001
rect 14415 5967 14473 6001
rect 14507 5967 14565 6001
rect 14599 5967 14657 6001
rect 14691 5967 14749 6001
rect 14783 5967 14841 6001
rect 14875 5967 14933 6001
rect 14967 5967 15025 6001
rect 15059 5967 15117 6001
rect 15151 5967 15209 6001
rect 15243 5967 15301 6001
rect 15335 5967 15393 6001
rect 15427 5967 15485 6001
rect 15519 5967 15577 6001
rect 15611 5967 15669 6001
rect 15703 5967 15761 6001
rect 15795 5967 15853 6001
rect 15887 5967 15945 6001
rect 15979 5967 16037 6001
rect 16071 5967 16129 6001
rect 16163 5967 16221 6001
rect 16255 5967 16313 6001
rect 16347 5967 16405 6001
rect 16439 5967 16497 6001
rect 16531 5967 16589 6001
rect 16623 5967 16681 6001
rect 16715 5967 16773 6001
rect 16807 5967 16865 6001
rect 16899 5967 16957 6001
rect 16991 5967 17049 6001
rect 17083 5967 17141 6001
rect 17175 5967 17233 6001
rect 17267 5967 17325 6001
rect 17359 5967 17417 6001
rect 17451 5967 17509 6001
rect 17543 5967 17601 6001
rect 17635 5967 17693 6001
rect 17727 5967 17785 6001
rect 17819 5967 17877 6001
rect 17911 5967 17969 6001
rect 18003 5967 18061 6001
rect 18095 5967 18153 6001
rect 18187 5967 18245 6001
rect 18279 5967 18337 6001
rect 18371 5967 18429 6001
rect 18463 5967 18521 6001
rect 18555 5967 18613 6001
rect 18647 5967 18705 6001
rect 18739 5967 18797 6001
rect 18831 5967 18860 6001
rect 1121 5925 1363 5967
rect 1121 5891 1139 5925
rect 1173 5891 1311 5925
rect 1345 5891 1363 5925
rect 1121 5830 1363 5891
rect 1397 5925 2466 5967
rect 1397 5891 1415 5925
rect 1449 5891 2415 5925
rect 2449 5891 2466 5925
rect 1397 5880 2466 5891
rect 2501 5925 3570 5967
rect 2501 5891 2519 5925
rect 2553 5891 3519 5925
rect 3553 5891 3570 5925
rect 2501 5880 3570 5891
rect 3697 5896 3755 5967
rect 1121 5796 1139 5830
rect 1173 5796 1311 5830
rect 1345 5796 1363 5830
rect 1121 5749 1363 5796
rect 1121 5681 1171 5715
rect 1205 5681 1225 5715
rect 1121 5607 1225 5681
rect 1259 5675 1363 5749
rect 1259 5641 1279 5675
rect 1313 5641 1363 5675
rect 1714 5715 1782 5732
rect 1714 5681 1731 5715
rect 1765 5681 1782 5715
rect 1121 5554 1363 5607
rect 1714 5566 1782 5681
rect 2078 5679 2148 5880
rect 2078 5645 2095 5679
rect 2129 5645 2148 5679
rect 2078 5630 2148 5645
rect 2818 5715 2886 5732
rect 2818 5681 2835 5715
rect 2869 5681 2886 5715
rect 2818 5566 2886 5681
rect 3182 5679 3252 5880
rect 3697 5862 3709 5896
rect 3743 5862 3755 5896
rect 3789 5925 4858 5967
rect 3789 5891 3807 5925
rect 3841 5891 4807 5925
rect 4841 5891 4858 5925
rect 3789 5880 4858 5891
rect 4893 5925 5962 5967
rect 4893 5891 4911 5925
rect 4945 5891 5911 5925
rect 5945 5891 5962 5925
rect 4893 5880 5962 5891
rect 5997 5925 6699 5967
rect 5997 5891 6015 5925
rect 6049 5891 6647 5925
rect 6681 5891 6699 5925
rect 3697 5803 3755 5862
rect 3697 5769 3709 5803
rect 3743 5769 3755 5803
rect 3697 5734 3755 5769
rect 3182 5645 3199 5679
rect 3233 5645 3252 5679
rect 3182 5630 3252 5645
rect 4106 5715 4174 5732
rect 4106 5681 4123 5715
rect 4157 5681 4174 5715
rect 3697 5585 3755 5602
rect 1121 5520 1139 5554
rect 1173 5520 1311 5554
rect 1345 5520 1363 5554
rect 1121 5457 1363 5520
rect 1397 5552 2466 5566
rect 1397 5518 1415 5552
rect 1449 5518 2415 5552
rect 2449 5518 2466 5552
rect 1397 5457 2466 5518
rect 2501 5552 3570 5566
rect 2501 5518 2519 5552
rect 2553 5518 3519 5552
rect 3553 5518 3570 5552
rect 2501 5457 3570 5518
rect 3697 5551 3709 5585
rect 3743 5551 3755 5585
rect 4106 5566 4174 5681
rect 4470 5679 4540 5880
rect 4470 5645 4487 5679
rect 4521 5645 4540 5679
rect 4470 5630 4540 5645
rect 5210 5715 5278 5732
rect 5210 5681 5227 5715
rect 5261 5681 5278 5715
rect 5210 5566 5278 5681
rect 5574 5679 5644 5880
rect 5997 5823 6699 5891
rect 5997 5789 6015 5823
rect 6049 5789 6647 5823
rect 6681 5789 6699 5823
rect 5997 5749 6699 5789
rect 5574 5645 5591 5679
rect 5625 5645 5644 5679
rect 5574 5630 5644 5645
rect 5997 5681 6075 5715
rect 6109 5681 6174 5715
rect 6208 5681 6273 5715
rect 6307 5681 6327 5715
rect 5997 5611 6327 5681
rect 6361 5679 6699 5749
rect 6361 5645 6381 5679
rect 6415 5645 6484 5679
rect 6518 5645 6587 5679
rect 6621 5645 6699 5679
rect 6733 5917 6787 5933
rect 6733 5883 6751 5917
rect 6785 5883 6787 5917
rect 6733 5836 6787 5883
rect 6733 5802 6751 5836
rect 6785 5802 6787 5836
rect 6821 5917 6887 5967
rect 6821 5883 6837 5917
rect 6871 5883 6887 5917
rect 6821 5849 6887 5883
rect 6821 5815 6837 5849
rect 6871 5815 6887 5849
rect 6923 5917 6957 5933
rect 6923 5849 6957 5883
rect 6733 5752 6787 5802
rect 6923 5781 6957 5815
rect 3697 5457 3755 5551
rect 3789 5552 4858 5566
rect 3789 5518 3807 5552
rect 3841 5518 4807 5552
rect 4841 5518 4858 5552
rect 3789 5457 4858 5518
rect 4893 5552 5962 5566
rect 4893 5518 4911 5552
rect 4945 5518 5911 5552
rect 5945 5518 5962 5552
rect 4893 5457 5962 5518
rect 5997 5552 6699 5611
rect 5997 5518 6015 5552
rect 6049 5518 6647 5552
rect 6681 5518 6699 5552
rect 5997 5457 6699 5518
rect 6733 5592 6767 5752
rect 6824 5747 6957 5781
rect 7009 5925 7527 5967
rect 7009 5891 7027 5925
rect 7061 5891 7475 5925
rect 7509 5891 7527 5925
rect 7009 5823 7527 5891
rect 7009 5789 7027 5823
rect 7061 5789 7475 5823
rect 7509 5789 7527 5823
rect 7009 5749 7527 5789
rect 6824 5718 6858 5747
rect 6801 5702 6858 5718
rect 6835 5668 6858 5702
rect 6801 5652 6858 5668
rect 6824 5601 6858 5652
rect 6905 5695 6971 5711
rect 6905 5689 6929 5695
rect 6905 5655 6921 5689
rect 6963 5661 6971 5695
rect 6955 5655 6971 5661
rect 6905 5637 6971 5655
rect 7009 5681 7087 5715
rect 7121 5681 7197 5715
rect 7231 5681 7251 5715
rect 7009 5611 7251 5681
rect 7285 5679 7527 5749
rect 7285 5645 7305 5679
rect 7339 5645 7415 5679
rect 7449 5645 7527 5679
rect 7561 5865 7664 5897
rect 7561 5831 7625 5865
rect 7659 5831 7664 5865
rect 7561 5815 7664 5831
rect 7711 5865 7745 5967
rect 7711 5815 7745 5831
rect 7779 5899 8185 5933
rect 7561 5653 7629 5815
rect 7779 5766 7813 5899
rect 7892 5831 7908 5865
rect 7942 5831 7983 5865
rect 8017 5831 8117 5865
rect 7663 5732 7679 5766
rect 7713 5763 7813 5766
rect 7713 5732 7757 5763
rect 7663 5729 7757 5732
rect 7791 5729 7813 5763
rect 7663 5728 7813 5729
rect 7847 5766 8049 5797
rect 7881 5763 8049 5766
rect 7881 5732 7885 5763
rect 7561 5619 7757 5653
rect 7791 5619 7807 5653
rect 6733 5563 6785 5592
rect 6824 5567 6957 5601
rect 6733 5559 6751 5563
rect 6733 5525 6745 5559
rect 6923 5546 6957 5567
rect 6779 5525 6785 5529
rect 6733 5491 6785 5525
rect 6821 5499 6837 5533
rect 6871 5499 6887 5533
rect 6821 5457 6887 5499
rect 6923 5491 6957 5512
rect 7009 5552 7527 5611
rect 7009 5518 7027 5552
rect 7061 5518 7475 5552
rect 7509 5518 7527 5552
rect 7009 5457 7527 5518
rect 7616 5548 7665 5619
rect 7616 5514 7625 5548
rect 7659 5514 7665 5548
rect 7616 5498 7665 5514
rect 7709 5548 7811 5564
rect 7743 5514 7777 5548
rect 7709 5457 7811 5514
rect 7847 5559 7885 5732
rect 7847 5525 7849 5559
rect 7883 5525 7885 5559
rect 7847 5491 7885 5525
rect 7919 5653 7974 5723
rect 7953 5627 7974 5653
rect 8015 5653 8049 5763
rect 7919 5593 7941 5619
rect 8015 5603 8049 5619
rect 8083 5605 8117 5831
rect 8151 5705 8185 5899
rect 8219 5925 8253 5967
rect 8219 5857 8253 5891
rect 8219 5789 8253 5823
rect 8219 5739 8253 5755
rect 8287 5925 8354 5933
rect 8287 5891 8303 5925
rect 8337 5899 8354 5925
rect 8287 5865 8309 5891
rect 8343 5865 8354 5899
rect 8287 5857 8354 5865
rect 8287 5823 8303 5857
rect 8337 5823 8354 5857
rect 8287 5789 8354 5823
rect 8287 5755 8303 5789
rect 8337 5755 8354 5789
rect 8287 5739 8354 5755
rect 8389 5925 8723 5967
rect 8389 5891 8407 5925
rect 8441 5891 8671 5925
rect 8705 5891 8723 5925
rect 8389 5823 8723 5891
rect 8389 5789 8407 5823
rect 8441 5789 8671 5823
rect 8705 5789 8723 5823
rect 8389 5749 8723 5789
rect 8151 5689 8190 5705
rect 8151 5655 8156 5689
rect 8151 5639 8190 5655
rect 8235 5689 8286 5705
rect 8235 5655 8252 5689
rect 8235 5639 8286 5655
rect 8235 5605 8269 5639
rect 8320 5605 8354 5739
rect 7919 5491 7974 5593
rect 8083 5571 8269 5605
rect 8083 5564 8118 5571
rect 8012 5548 8118 5564
rect 8046 5514 8118 5548
rect 8303 5552 8354 5605
rect 8012 5491 8118 5514
rect 8203 5533 8269 5537
rect 8203 5499 8219 5533
rect 8253 5499 8269 5533
rect 8203 5457 8269 5499
rect 8337 5518 8354 5552
rect 8303 5491 8354 5518
rect 8389 5681 8409 5715
rect 8443 5681 8539 5715
rect 8389 5611 8539 5681
rect 8573 5679 8723 5749
rect 8849 5896 8907 5967
rect 8849 5862 8861 5896
rect 8895 5862 8907 5896
rect 8941 5925 10010 5967
rect 8941 5891 8959 5925
rect 8993 5891 9959 5925
rect 9993 5891 10010 5925
rect 8941 5880 10010 5891
rect 10045 5925 11114 5967
rect 10045 5891 10063 5925
rect 10097 5891 11063 5925
rect 11097 5891 11114 5925
rect 10045 5880 11114 5891
rect 11149 5925 11483 5967
rect 11149 5891 11167 5925
rect 11201 5891 11431 5925
rect 11465 5891 11483 5925
rect 8849 5803 8907 5862
rect 8849 5769 8861 5803
rect 8895 5769 8907 5803
rect 8849 5734 8907 5769
rect 8573 5645 8669 5679
rect 8703 5645 8723 5679
rect 9258 5715 9326 5732
rect 9258 5681 9275 5715
rect 9309 5681 9326 5715
rect 8389 5559 8723 5611
rect 8389 5525 8407 5559
rect 8441 5525 8671 5559
rect 8705 5525 8723 5559
rect 8389 5457 8723 5525
rect 8849 5585 8907 5602
rect 8849 5551 8861 5585
rect 8895 5551 8907 5585
rect 9258 5566 9326 5681
rect 9622 5679 9692 5880
rect 9622 5645 9639 5679
rect 9673 5645 9692 5679
rect 9622 5630 9692 5645
rect 10362 5715 10430 5732
rect 10362 5681 10379 5715
rect 10413 5681 10430 5715
rect 10362 5566 10430 5681
rect 10726 5679 10796 5880
rect 11149 5823 11483 5891
rect 11149 5789 11167 5823
rect 11201 5789 11431 5823
rect 11465 5789 11483 5823
rect 11729 5909 11795 5967
rect 11729 5875 11745 5909
rect 11779 5875 11795 5909
rect 11729 5841 11795 5875
rect 11149 5749 11483 5789
rect 10726 5645 10743 5679
rect 10777 5645 10796 5679
rect 10726 5630 10796 5645
rect 11149 5681 11169 5715
rect 11203 5681 11299 5715
rect 11149 5611 11299 5681
rect 11333 5679 11483 5749
rect 11554 5789 11632 5808
rect 11729 5807 11745 5841
rect 11779 5807 11795 5841
rect 11829 5925 11936 5933
rect 11829 5891 11845 5925
rect 11879 5891 11936 5925
rect 11829 5857 11936 5891
rect 11829 5823 11845 5857
rect 11879 5823 11936 5857
rect 11829 5809 11936 5823
rect 11554 5755 11576 5789
rect 11610 5773 11632 5789
rect 11610 5755 11839 5773
rect 11554 5739 11839 5755
rect 11333 5645 11429 5679
rect 11463 5645 11483 5679
rect 11529 5689 11600 5705
rect 11529 5655 11566 5689
rect 11529 5627 11600 5655
rect 8849 5457 8907 5551
rect 8941 5552 10010 5566
rect 8941 5518 8959 5552
rect 8993 5518 9959 5552
rect 9993 5518 10010 5552
rect 8941 5457 10010 5518
rect 10045 5552 11114 5566
rect 10045 5518 10063 5552
rect 10097 5518 11063 5552
rect 11097 5518 11114 5552
rect 10045 5457 11114 5518
rect 11149 5559 11483 5611
rect 11563 5593 11600 5627
rect 11634 5559 11668 5739
rect 11702 5689 11755 5705
rect 11736 5655 11755 5689
rect 11702 5627 11755 5655
rect 11805 5689 11839 5739
rect 11805 5639 11839 5655
rect 11702 5593 11713 5627
rect 11747 5593 11755 5627
rect 11873 5605 11936 5809
rect 11977 5925 12679 5967
rect 11977 5891 11995 5925
rect 12029 5891 12627 5925
rect 12661 5891 12679 5925
rect 11977 5823 12679 5891
rect 11977 5789 11995 5823
rect 12029 5789 12627 5823
rect 12661 5789 12679 5823
rect 13017 5909 13083 5967
rect 13017 5875 13033 5909
rect 13067 5875 13083 5909
rect 13017 5841 13083 5875
rect 11977 5749 12679 5789
rect 11813 5603 11936 5605
rect 11813 5569 11829 5603
rect 11863 5569 11936 5603
rect 11813 5559 11936 5569
rect 11149 5525 11167 5559
rect 11201 5525 11431 5559
rect 11465 5525 11483 5559
rect 11149 5457 11483 5525
rect 11550 5543 11598 5559
rect 11550 5509 11564 5543
rect 11550 5457 11598 5509
rect 11634 5543 11690 5559
rect 11634 5509 11648 5543
rect 11682 5509 11690 5543
rect 11634 5493 11690 5509
rect 11736 5543 11779 5559
rect 11736 5509 11744 5543
rect 11778 5509 11779 5543
rect 11736 5457 11779 5509
rect 11813 5535 11897 5559
rect 11813 5501 11829 5535
rect 11863 5525 11897 5535
rect 11931 5525 11936 5559
rect 11863 5501 11936 5525
rect 11813 5491 11936 5501
rect 11977 5681 12055 5715
rect 12089 5681 12154 5715
rect 12188 5681 12253 5715
rect 12287 5681 12307 5715
rect 11977 5611 12307 5681
rect 12341 5679 12679 5749
rect 12842 5789 12920 5808
rect 13017 5807 13033 5841
rect 13067 5807 13083 5841
rect 13117 5925 13224 5933
rect 13117 5891 13133 5925
rect 13167 5891 13224 5925
rect 13117 5857 13224 5891
rect 13117 5823 13133 5857
rect 13167 5823 13224 5857
rect 13117 5809 13224 5823
rect 12842 5755 12864 5789
rect 12898 5773 12920 5789
rect 12898 5755 13127 5773
rect 12842 5739 13127 5755
rect 12341 5645 12361 5679
rect 12395 5645 12464 5679
rect 12498 5645 12567 5679
rect 12601 5645 12679 5679
rect 12817 5689 12888 5705
rect 12817 5655 12854 5689
rect 12817 5627 12888 5655
rect 11977 5552 12679 5611
rect 12851 5593 12888 5627
rect 12922 5559 12956 5739
rect 12990 5689 13043 5705
rect 13024 5655 13043 5689
rect 12990 5627 13043 5655
rect 13093 5689 13127 5739
rect 13093 5639 13127 5655
rect 12990 5593 13001 5627
rect 13035 5593 13043 5627
rect 13161 5605 13224 5809
rect 13265 5925 13967 5967
rect 13265 5891 13283 5925
rect 13317 5891 13915 5925
rect 13949 5891 13967 5925
rect 13265 5823 13967 5891
rect 13265 5789 13283 5823
rect 13317 5789 13915 5823
rect 13949 5789 13967 5823
rect 13265 5749 13967 5789
rect 13101 5603 13224 5605
rect 13101 5569 13117 5603
rect 13151 5569 13224 5603
rect 13101 5559 13224 5569
rect 11977 5518 11995 5552
rect 12029 5518 12627 5552
rect 12661 5518 12679 5552
rect 11977 5457 12679 5518
rect 12838 5543 12886 5559
rect 12838 5509 12852 5543
rect 12838 5457 12886 5509
rect 12922 5543 12978 5559
rect 12922 5509 12936 5543
rect 12970 5509 12978 5543
rect 12922 5493 12978 5509
rect 13024 5543 13067 5559
rect 13024 5509 13032 5543
rect 13066 5509 13067 5543
rect 13024 5457 13067 5509
rect 13101 5535 13185 5559
rect 13101 5501 13117 5535
rect 13151 5525 13185 5535
rect 13219 5525 13224 5559
rect 13151 5501 13224 5525
rect 13101 5491 13224 5501
rect 13265 5681 13343 5715
rect 13377 5681 13442 5715
rect 13476 5681 13541 5715
rect 13575 5681 13595 5715
rect 13265 5611 13595 5681
rect 13629 5679 13967 5749
rect 14001 5896 14059 5967
rect 14001 5862 14013 5896
rect 14047 5862 14059 5896
rect 14093 5925 15162 5967
rect 14093 5891 14111 5925
rect 14145 5891 15111 5925
rect 15145 5891 15162 5925
rect 14093 5880 15162 5891
rect 15197 5925 16266 5967
rect 15197 5891 15215 5925
rect 15249 5891 16215 5925
rect 16249 5891 16266 5925
rect 15197 5880 16266 5891
rect 16301 5925 17370 5967
rect 16301 5891 16319 5925
rect 16353 5891 17319 5925
rect 17353 5891 17370 5925
rect 16301 5880 17370 5891
rect 17405 5925 18474 5967
rect 17405 5891 17423 5925
rect 17457 5891 18423 5925
rect 18457 5891 18474 5925
rect 17405 5880 18474 5891
rect 18601 5925 18843 5967
rect 18601 5891 18619 5925
rect 18653 5891 18791 5925
rect 18825 5891 18843 5925
rect 14001 5803 14059 5862
rect 14001 5769 14013 5803
rect 14047 5769 14059 5803
rect 14001 5734 14059 5769
rect 13629 5645 13649 5679
rect 13683 5645 13752 5679
rect 13786 5645 13855 5679
rect 13889 5645 13967 5679
rect 14410 5715 14478 5732
rect 14410 5681 14427 5715
rect 14461 5681 14478 5715
rect 13265 5552 13967 5611
rect 13265 5518 13283 5552
rect 13317 5518 13915 5552
rect 13949 5518 13967 5552
rect 13265 5457 13967 5518
rect 14001 5585 14059 5602
rect 14001 5551 14013 5585
rect 14047 5551 14059 5585
rect 14410 5566 14478 5681
rect 14774 5679 14844 5880
rect 14774 5645 14791 5679
rect 14825 5645 14844 5679
rect 14774 5630 14844 5645
rect 15514 5715 15582 5732
rect 15514 5681 15531 5715
rect 15565 5681 15582 5715
rect 15514 5566 15582 5681
rect 15878 5679 15948 5880
rect 15878 5645 15895 5679
rect 15929 5645 15948 5679
rect 15878 5630 15948 5645
rect 16618 5715 16686 5732
rect 16618 5681 16635 5715
rect 16669 5681 16686 5715
rect 16618 5566 16686 5681
rect 16982 5679 17052 5880
rect 16982 5645 16999 5679
rect 17033 5645 17052 5679
rect 16982 5630 17052 5645
rect 17722 5715 17790 5732
rect 17722 5681 17739 5715
rect 17773 5681 17790 5715
rect 17722 5566 17790 5681
rect 18086 5679 18156 5880
rect 18086 5645 18103 5679
rect 18137 5645 18156 5679
rect 18086 5630 18156 5645
rect 18601 5830 18843 5891
rect 18601 5796 18619 5830
rect 18653 5796 18791 5830
rect 18825 5796 18843 5830
rect 18601 5749 18843 5796
rect 18601 5675 18705 5749
rect 18601 5641 18651 5675
rect 18685 5641 18705 5675
rect 18739 5681 18759 5715
rect 18793 5681 18843 5715
rect 18739 5607 18843 5681
rect 14001 5457 14059 5551
rect 14093 5552 15162 5566
rect 14093 5518 14111 5552
rect 14145 5518 15111 5552
rect 15145 5518 15162 5552
rect 14093 5457 15162 5518
rect 15197 5552 16266 5566
rect 15197 5518 15215 5552
rect 15249 5518 16215 5552
rect 16249 5518 16266 5552
rect 15197 5457 16266 5518
rect 16301 5552 17370 5566
rect 16301 5518 16319 5552
rect 16353 5518 17319 5552
rect 17353 5518 17370 5552
rect 16301 5457 17370 5518
rect 17405 5552 18474 5566
rect 17405 5518 17423 5552
rect 17457 5518 18423 5552
rect 18457 5518 18474 5552
rect 17405 5457 18474 5518
rect 18601 5554 18843 5607
rect 18601 5520 18619 5554
rect 18653 5520 18791 5554
rect 18825 5520 18843 5554
rect 18601 5457 18843 5520
rect 1104 5423 1133 5457
rect 1167 5423 1225 5457
rect 1259 5423 1317 5457
rect 1351 5423 1409 5457
rect 1443 5423 1501 5457
rect 1535 5423 1593 5457
rect 1627 5423 1685 5457
rect 1719 5423 1777 5457
rect 1811 5423 1869 5457
rect 1903 5423 1961 5457
rect 1995 5423 2053 5457
rect 2087 5423 2145 5457
rect 2179 5423 2237 5457
rect 2271 5423 2329 5457
rect 2363 5423 2421 5457
rect 2455 5423 2513 5457
rect 2547 5423 2605 5457
rect 2639 5423 2697 5457
rect 2731 5423 2789 5457
rect 2823 5423 2881 5457
rect 2915 5423 2973 5457
rect 3007 5423 3065 5457
rect 3099 5423 3157 5457
rect 3191 5423 3249 5457
rect 3283 5423 3341 5457
rect 3375 5423 3433 5457
rect 3467 5423 3525 5457
rect 3559 5423 3617 5457
rect 3651 5423 3709 5457
rect 3743 5423 3801 5457
rect 3835 5423 3893 5457
rect 3927 5423 3985 5457
rect 4019 5423 4077 5457
rect 4111 5423 4169 5457
rect 4203 5423 4261 5457
rect 4295 5423 4353 5457
rect 4387 5423 4445 5457
rect 4479 5423 4537 5457
rect 4571 5423 4629 5457
rect 4663 5423 4721 5457
rect 4755 5423 4813 5457
rect 4847 5423 4905 5457
rect 4939 5423 4997 5457
rect 5031 5423 5089 5457
rect 5123 5423 5181 5457
rect 5215 5423 5273 5457
rect 5307 5423 5365 5457
rect 5399 5423 5457 5457
rect 5491 5423 5549 5457
rect 5583 5423 5641 5457
rect 5675 5423 5733 5457
rect 5767 5423 5825 5457
rect 5859 5423 5917 5457
rect 5951 5423 6009 5457
rect 6043 5423 6101 5457
rect 6135 5423 6193 5457
rect 6227 5423 6285 5457
rect 6319 5423 6377 5457
rect 6411 5423 6469 5457
rect 6503 5423 6561 5457
rect 6595 5423 6653 5457
rect 6687 5423 6745 5457
rect 6779 5423 6837 5457
rect 6871 5423 6929 5457
rect 6963 5423 7021 5457
rect 7055 5423 7113 5457
rect 7147 5423 7205 5457
rect 7239 5423 7297 5457
rect 7331 5423 7389 5457
rect 7423 5423 7481 5457
rect 7515 5423 7573 5457
rect 7607 5423 7665 5457
rect 7699 5423 7757 5457
rect 7791 5423 7849 5457
rect 7883 5423 7941 5457
rect 7975 5423 8033 5457
rect 8067 5423 8125 5457
rect 8159 5423 8217 5457
rect 8251 5423 8309 5457
rect 8343 5423 8401 5457
rect 8435 5423 8493 5457
rect 8527 5423 8585 5457
rect 8619 5423 8677 5457
rect 8711 5423 8769 5457
rect 8803 5423 8861 5457
rect 8895 5423 8953 5457
rect 8987 5423 9045 5457
rect 9079 5423 9137 5457
rect 9171 5423 9229 5457
rect 9263 5423 9321 5457
rect 9355 5423 9413 5457
rect 9447 5423 9505 5457
rect 9539 5423 9597 5457
rect 9631 5423 9689 5457
rect 9723 5423 9781 5457
rect 9815 5423 9873 5457
rect 9907 5423 9965 5457
rect 9999 5423 10057 5457
rect 10091 5423 10149 5457
rect 10183 5423 10241 5457
rect 10275 5423 10333 5457
rect 10367 5423 10425 5457
rect 10459 5423 10517 5457
rect 10551 5423 10609 5457
rect 10643 5423 10701 5457
rect 10735 5423 10793 5457
rect 10827 5423 10885 5457
rect 10919 5423 10977 5457
rect 11011 5423 11069 5457
rect 11103 5423 11161 5457
rect 11195 5423 11253 5457
rect 11287 5423 11345 5457
rect 11379 5423 11437 5457
rect 11471 5423 11529 5457
rect 11563 5423 11621 5457
rect 11655 5423 11713 5457
rect 11747 5423 11805 5457
rect 11839 5423 11897 5457
rect 11931 5423 11989 5457
rect 12023 5423 12081 5457
rect 12115 5423 12173 5457
rect 12207 5423 12265 5457
rect 12299 5423 12357 5457
rect 12391 5423 12449 5457
rect 12483 5423 12541 5457
rect 12575 5423 12633 5457
rect 12667 5423 12725 5457
rect 12759 5423 12817 5457
rect 12851 5423 12909 5457
rect 12943 5423 13001 5457
rect 13035 5423 13093 5457
rect 13127 5423 13185 5457
rect 13219 5423 13277 5457
rect 13311 5423 13369 5457
rect 13403 5423 13461 5457
rect 13495 5423 13553 5457
rect 13587 5423 13645 5457
rect 13679 5423 13737 5457
rect 13771 5423 13829 5457
rect 13863 5423 13921 5457
rect 13955 5423 14013 5457
rect 14047 5423 14105 5457
rect 14139 5423 14197 5457
rect 14231 5423 14289 5457
rect 14323 5423 14381 5457
rect 14415 5423 14473 5457
rect 14507 5423 14565 5457
rect 14599 5423 14657 5457
rect 14691 5423 14749 5457
rect 14783 5423 14841 5457
rect 14875 5423 14933 5457
rect 14967 5423 15025 5457
rect 15059 5423 15117 5457
rect 15151 5423 15209 5457
rect 15243 5423 15301 5457
rect 15335 5423 15393 5457
rect 15427 5423 15485 5457
rect 15519 5423 15577 5457
rect 15611 5423 15669 5457
rect 15703 5423 15761 5457
rect 15795 5423 15853 5457
rect 15887 5423 15945 5457
rect 15979 5423 16037 5457
rect 16071 5423 16129 5457
rect 16163 5423 16221 5457
rect 16255 5423 16313 5457
rect 16347 5423 16405 5457
rect 16439 5423 16497 5457
rect 16531 5423 16589 5457
rect 16623 5423 16681 5457
rect 16715 5423 16773 5457
rect 16807 5423 16865 5457
rect 16899 5423 16957 5457
rect 16991 5423 17049 5457
rect 17083 5423 17141 5457
rect 17175 5423 17233 5457
rect 17267 5423 17325 5457
rect 17359 5423 17417 5457
rect 17451 5423 17509 5457
rect 17543 5423 17601 5457
rect 17635 5423 17693 5457
rect 17727 5423 17785 5457
rect 17819 5423 17877 5457
rect 17911 5423 17969 5457
rect 18003 5423 18061 5457
rect 18095 5423 18153 5457
rect 18187 5423 18245 5457
rect 18279 5423 18337 5457
rect 18371 5423 18429 5457
rect 18463 5423 18521 5457
rect 18555 5423 18613 5457
rect 18647 5423 18705 5457
rect 18739 5423 18797 5457
rect 18831 5423 18860 5457
rect 1121 5360 1363 5423
rect 1121 5326 1139 5360
rect 1173 5326 1311 5360
rect 1345 5326 1363 5360
rect 1121 5273 1363 5326
rect 1397 5362 2466 5423
rect 1397 5328 1415 5362
rect 1449 5328 2415 5362
rect 2449 5328 2466 5362
rect 1397 5314 2466 5328
rect 2501 5360 2743 5423
rect 2863 5381 2929 5423
rect 2501 5326 2519 5360
rect 2553 5326 2691 5360
rect 2725 5326 2743 5360
rect 1121 5199 1225 5273
rect 1121 5165 1171 5199
rect 1205 5165 1225 5199
rect 1259 5205 1279 5239
rect 1313 5205 1363 5239
rect 1259 5131 1363 5205
rect 1714 5199 1782 5314
rect 2501 5273 2743 5326
rect 2778 5355 2829 5371
rect 2778 5321 2795 5355
rect 2863 5347 2879 5381
rect 2913 5347 2929 5381
rect 3069 5385 3135 5423
rect 2963 5355 2997 5371
rect 2778 5313 2829 5321
rect 3069 5351 3085 5385
rect 3119 5351 3135 5385
rect 3655 5381 3721 5423
rect 2778 5279 2928 5313
rect 1714 5165 1731 5199
rect 1765 5165 1782 5199
rect 1714 5148 1782 5165
rect 2078 5235 2148 5250
rect 2078 5201 2095 5235
rect 2129 5201 2148 5235
rect 1121 5084 1363 5131
rect 1121 5050 1139 5084
rect 1173 5050 1311 5084
rect 1345 5050 1363 5084
rect 1121 4989 1363 5050
rect 2078 5000 2148 5201
rect 2501 5199 2605 5273
rect 2501 5165 2551 5199
rect 2585 5165 2605 5199
rect 2639 5205 2659 5239
rect 2693 5205 2743 5239
rect 2639 5131 2743 5205
rect 2501 5084 2743 5131
rect 2778 5225 2848 5245
rect 2778 5191 2792 5225
rect 2826 5191 2848 5225
rect 2778 5151 2848 5191
rect 2778 5117 2789 5151
rect 2823 5117 2848 5151
rect 2778 5115 2848 5117
rect 2882 5219 2928 5279
rect 2916 5210 2928 5219
rect 2882 5176 2894 5185
rect 2501 5050 2519 5084
rect 2553 5050 2691 5084
rect 2725 5050 2743 5084
rect 2882 5081 2928 5176
rect 1121 4955 1139 4989
rect 1173 4955 1311 4989
rect 1345 4955 1363 4989
rect 1121 4913 1363 4955
rect 1397 4989 2466 5000
rect 1397 4955 1415 4989
rect 1449 4955 2415 4989
rect 2449 4955 2466 4989
rect 1397 4913 2466 4955
rect 2501 4989 2743 5050
rect 2501 4955 2519 4989
rect 2553 4955 2691 4989
rect 2725 4955 2743 4989
rect 2501 4913 2743 4955
rect 2778 5065 2928 5081
rect 2778 5031 2795 5065
rect 2829 5047 2928 5065
rect 2963 5083 2997 5321
rect 3169 5345 3218 5379
rect 3252 5345 3268 5379
rect 3309 5345 3325 5379
rect 3359 5345 3480 5379
rect 3043 5164 3135 5317
rect 3043 5151 3101 5164
rect 3043 5117 3065 5151
rect 3099 5130 3101 5151
rect 3099 5117 3135 5130
rect 3043 5107 3135 5117
rect 2778 4997 2829 5031
rect 2778 4963 2795 4997
rect 2778 4947 2829 4963
rect 2863 4979 2879 5013
rect 2913 4979 2929 5013
rect 2863 4913 2929 4979
rect 2963 4997 2997 5031
rect 2963 4947 2997 4963
rect 3031 4950 3096 5107
rect 3169 5073 3203 5345
rect 3237 5271 3307 5287
rect 3237 5237 3260 5271
rect 3294 5237 3307 5271
rect 3237 5219 3307 5237
rect 3237 5185 3249 5219
rect 3283 5185 3307 5219
rect 3237 5163 3307 5185
rect 3341 5277 3412 5287
rect 3341 5243 3362 5277
rect 3396 5243 3412 5277
rect 3341 5125 3375 5243
rect 3446 5203 3480 5345
rect 3655 5347 3671 5381
rect 3705 5347 3721 5381
rect 3655 5331 3721 5347
rect 3763 5351 3783 5385
rect 3817 5351 3833 5385
rect 3877 5381 4067 5389
rect 3555 5253 3593 5287
rect 3627 5271 3679 5287
rect 3763 5273 3815 5351
rect 3877 5347 3893 5381
rect 3927 5347 4067 5381
rect 3877 5333 4067 5347
rect 4101 5385 4139 5423
rect 4101 5351 4105 5385
rect 4436 5381 4497 5423
rect 4101 5335 4139 5351
rect 4173 5365 4387 5381
rect 4173 5347 4323 5365
rect 3521 5237 3617 5253
rect 3651 5237 3679 5271
rect 3713 5223 3747 5239
rect 3282 5109 3375 5125
rect 3316 5083 3375 5109
rect 3316 5075 3341 5083
rect 3169 5039 3248 5073
rect 3282 5049 3341 5075
rect 3282 5047 3375 5049
rect 3409 5189 3713 5203
rect 3409 5169 3747 5189
rect 3214 5013 3248 5039
rect 3409 5013 3443 5169
rect 3781 5135 3815 5273
rect 3515 5101 3531 5135
rect 3565 5101 3815 5135
rect 3853 5283 3895 5299
rect 3853 5249 3861 5283
rect 3853 5141 3895 5249
rect 3929 5235 3999 5299
rect 3929 5201 3957 5235
rect 3991 5219 3999 5235
rect 3929 5185 3965 5201
rect 3929 5175 3999 5185
rect 4033 5177 4067 5333
rect 4173 5301 4207 5347
rect 4357 5331 4387 5365
rect 4436 5347 4447 5381
rect 4481 5347 4497 5381
rect 4436 5331 4497 5347
rect 4531 5355 4582 5387
rect 4531 5331 4537 5355
rect 4101 5267 4207 5301
rect 4241 5287 4289 5313
rect 4101 5261 4145 5267
rect 4135 5227 4145 5261
rect 4275 5253 4289 5287
rect 4241 5233 4289 5253
rect 4101 5211 4145 5227
rect 4181 5224 4197 5233
rect 4231 5199 4289 5233
rect 4215 5190 4289 5199
rect 4033 5143 4114 5177
rect 4181 5159 4289 5190
rect 4323 5276 4387 5331
rect 4571 5321 4582 5355
rect 4565 5297 4582 5321
rect 4617 5362 5686 5423
rect 4617 5328 4635 5362
rect 4669 5328 5635 5362
rect 5669 5328 5686 5362
rect 4617 5314 5686 5328
rect 5721 5362 6239 5423
rect 5721 5328 5739 5362
rect 5773 5328 6187 5362
rect 6221 5328 6239 5362
rect 4531 5281 4582 5297
rect 4323 5241 4388 5276
rect 4323 5225 4506 5241
rect 4323 5191 4472 5225
rect 4323 5181 4506 5191
rect 4358 5175 4506 5181
rect 3853 5109 3988 5141
rect 4080 5125 4114 5143
rect 3853 5107 3996 5109
rect 3781 5073 3815 5101
rect 3954 5083 3996 5107
rect 3130 4989 3180 5005
rect 3130 4955 3146 4989
rect 3130 4913 3180 4955
rect 3214 4997 3264 5013
rect 3214 4963 3230 4997
rect 3214 4947 3264 4963
rect 3307 4991 3443 5013
rect 3307 4957 3323 4991
rect 3357 4957 3443 4991
rect 3477 5033 3692 5067
rect 3781 5039 3893 5073
rect 3954 5049 3965 5083
rect 4030 5075 4046 5109
rect 3999 5049 4046 5075
rect 4080 5091 4274 5125
rect 4308 5091 4324 5125
rect 3477 5015 3511 5033
rect 3658 5015 3692 5033
rect 3477 4965 3511 4981
rect 3558 4965 3574 4999
rect 3608 4965 3624 4999
rect 3658 4965 3692 4981
rect 3751 4989 3825 5005
rect 3307 4947 3443 4957
rect 3558 4913 3624 4965
rect 3751 4955 3771 4989
rect 3805 4955 3825 4989
rect 3751 4913 3825 4955
rect 3859 4997 3893 5039
rect 4080 5015 4114 5091
rect 4358 5057 4392 5175
rect 4540 5151 4582 5281
rect 3859 4947 3893 4963
rect 3940 4990 4114 5015
rect 4232 5023 4392 5057
rect 4436 5057 4497 5141
rect 4436 5023 4447 5057
rect 4481 5023 4497 5057
rect 4232 5015 4266 5023
rect 3940 4956 3956 4990
rect 3990 4956 4114 4990
rect 3940 4947 4114 4956
rect 4148 4989 4198 5005
rect 4182 4955 4198 4989
rect 4436 4989 4497 5023
rect 4232 4965 4266 4981
rect 4148 4913 4198 4955
rect 4302 4955 4318 4989
rect 4352 4955 4368 4989
rect 4302 4913 4368 4955
rect 4436 4955 4447 4989
rect 4481 4955 4497 4989
rect 4531 5093 4582 5151
rect 4934 5199 5002 5314
rect 5721 5269 6239 5328
rect 6273 5329 6331 5423
rect 6273 5295 6285 5329
rect 6319 5295 6331 5329
rect 6273 5278 6331 5295
rect 6365 5360 6607 5423
rect 6365 5326 6383 5360
rect 6417 5326 6555 5360
rect 6589 5326 6607 5360
rect 6365 5273 6607 5326
rect 6642 5362 6693 5389
rect 6642 5328 6659 5362
rect 6727 5381 6793 5423
rect 6727 5347 6743 5381
rect 6777 5347 6793 5381
rect 6727 5343 6793 5347
rect 6878 5366 6984 5389
rect 6642 5275 6693 5328
rect 6878 5332 6950 5366
rect 7022 5355 7077 5389
rect 6878 5316 6984 5332
rect 7055 5321 7077 5355
rect 6878 5309 6913 5316
rect 6727 5275 6913 5309
rect 4934 5165 4951 5199
rect 4985 5165 5002 5199
rect 4934 5148 5002 5165
rect 5298 5235 5368 5250
rect 5298 5201 5315 5235
rect 5349 5201 5368 5235
rect 4565 5059 4582 5093
rect 4531 5025 4582 5059
rect 4565 4991 4582 5025
rect 5298 5000 5368 5201
rect 5721 5199 5963 5269
rect 5721 5165 5799 5199
rect 5833 5165 5909 5199
rect 5943 5165 5963 5199
rect 5997 5201 6017 5235
rect 6051 5201 6127 5235
rect 6161 5201 6239 5235
rect 5997 5131 6239 5201
rect 6365 5199 6469 5273
rect 6365 5165 6415 5199
rect 6449 5165 6469 5199
rect 6503 5205 6523 5239
rect 6557 5205 6607 5239
rect 5721 5091 6239 5131
rect 5721 5057 5739 5091
rect 5773 5057 6187 5091
rect 6221 5057 6239 5091
rect 4531 4975 4582 4991
rect 4617 4989 5686 5000
rect 4436 4913 4497 4955
rect 4617 4955 4635 4989
rect 4669 4955 5635 4989
rect 5669 4955 5686 4989
rect 4617 4913 5686 4955
rect 5721 4989 6239 5057
rect 5721 4955 5739 4989
rect 5773 4955 6187 4989
rect 6221 4955 6239 4989
rect 5721 4913 6239 4955
rect 6273 5111 6331 5146
rect 6503 5131 6607 5205
rect 6273 5077 6285 5111
rect 6319 5077 6331 5111
rect 6273 5018 6331 5077
rect 6273 4984 6285 5018
rect 6319 4984 6331 5018
rect 6273 4913 6331 4984
rect 6365 5084 6607 5131
rect 6365 5050 6383 5084
rect 6417 5050 6555 5084
rect 6589 5050 6607 5084
rect 6365 4989 6607 5050
rect 6365 4955 6383 4989
rect 6417 4955 6555 4989
rect 6589 4955 6607 4989
rect 6365 4913 6607 4955
rect 6642 5141 6676 5275
rect 6727 5241 6761 5275
rect 6710 5225 6761 5241
rect 6744 5191 6761 5225
rect 6710 5175 6761 5191
rect 6806 5225 6845 5241
rect 6840 5191 6845 5225
rect 6806 5175 6845 5191
rect 6642 5125 6709 5141
rect 6642 5091 6659 5125
rect 6693 5091 6709 5125
rect 6642 5057 6709 5091
rect 6642 5023 6659 5057
rect 6693 5023 6709 5057
rect 6642 5015 6709 5023
rect 6642 4981 6653 5015
rect 6687 4989 6709 5015
rect 6642 4955 6659 4981
rect 6693 4955 6709 4989
rect 6642 4947 6709 4955
rect 6743 5125 6777 5141
rect 6743 5057 6777 5091
rect 6743 4989 6777 5023
rect 6743 4913 6777 4955
rect 6811 4981 6845 5175
rect 6879 5049 6913 5275
rect 6947 5261 6981 5277
rect 6947 5117 6981 5227
rect 7022 5261 7077 5321
rect 7022 5227 7043 5261
rect 7022 5157 7077 5227
rect 7111 5355 7149 5389
rect 7111 5321 7113 5355
rect 7147 5321 7149 5355
rect 7111 5148 7149 5321
rect 7185 5366 7287 5423
rect 7219 5332 7253 5366
rect 7185 5316 7287 5332
rect 7331 5366 7380 5382
rect 7331 5332 7337 5366
rect 7371 5332 7380 5366
rect 7331 5261 7380 5332
rect 7469 5355 7803 5423
rect 7923 5381 7989 5423
rect 7469 5321 7487 5355
rect 7521 5321 7751 5355
rect 7785 5321 7803 5355
rect 7469 5269 7803 5321
rect 7838 5355 7889 5371
rect 7838 5321 7855 5355
rect 7923 5347 7939 5381
rect 7973 5347 7989 5381
rect 8129 5385 8195 5423
rect 8023 5355 8057 5371
rect 7838 5313 7889 5321
rect 8129 5351 8145 5385
rect 8179 5351 8195 5385
rect 8715 5381 8781 5423
rect 7838 5279 7988 5313
rect 7189 5227 7205 5261
rect 7239 5227 7435 5261
rect 7111 5117 7115 5148
rect 6947 5114 7115 5117
rect 6947 5083 7149 5114
rect 7183 5151 7333 5152
rect 7183 5117 7205 5151
rect 7239 5148 7333 5151
rect 7239 5117 7283 5148
rect 7183 5114 7283 5117
rect 7317 5114 7333 5148
rect 6879 5015 6979 5049
rect 7013 5015 7054 5049
rect 7088 5015 7104 5049
rect 7183 4981 7217 5114
rect 7367 5065 7435 5227
rect 7469 5199 7619 5269
rect 7469 5165 7489 5199
rect 7523 5165 7619 5199
rect 7653 5201 7749 5235
rect 7783 5201 7803 5235
rect 7653 5131 7803 5201
rect 6811 4947 7217 4981
rect 7251 5049 7285 5065
rect 7251 4913 7285 5015
rect 7332 5049 7435 5065
rect 7332 5015 7337 5049
rect 7371 5015 7435 5049
rect 7332 4983 7435 5015
rect 7469 5091 7803 5131
rect 7838 5225 7908 5245
rect 7838 5191 7852 5225
rect 7886 5191 7908 5225
rect 7838 5151 7908 5191
rect 7838 5117 7849 5151
rect 7883 5117 7908 5151
rect 7838 5115 7908 5117
rect 7942 5219 7988 5279
rect 7976 5210 7988 5219
rect 7942 5176 7954 5185
rect 7469 5057 7487 5091
rect 7521 5057 7751 5091
rect 7785 5057 7803 5091
rect 7942 5081 7988 5176
rect 7469 4989 7803 5057
rect 7469 4955 7487 4989
rect 7521 4955 7751 4989
rect 7785 4955 7803 4989
rect 7469 4913 7803 4955
rect 7838 5065 7988 5081
rect 7838 5031 7855 5065
rect 7889 5047 7988 5065
rect 8023 5083 8057 5321
rect 8229 5345 8278 5379
rect 8312 5345 8328 5379
rect 8369 5345 8385 5379
rect 8419 5345 8540 5379
rect 8103 5164 8195 5317
rect 8103 5151 8161 5164
rect 8103 5117 8125 5151
rect 8159 5130 8161 5151
rect 8159 5117 8195 5130
rect 8103 5107 8195 5117
rect 7838 4997 7889 5031
rect 7838 4963 7855 4997
rect 7838 4947 7889 4963
rect 7923 4979 7939 5013
rect 7973 4979 7989 5013
rect 7923 4913 7989 4979
rect 8023 4997 8057 5031
rect 8023 4947 8057 4963
rect 8091 4950 8156 5107
rect 8229 5073 8263 5345
rect 8297 5271 8367 5287
rect 8297 5237 8320 5271
rect 8354 5237 8367 5271
rect 8297 5219 8367 5237
rect 8297 5185 8309 5219
rect 8343 5185 8367 5219
rect 8297 5163 8367 5185
rect 8401 5277 8472 5287
rect 8401 5243 8422 5277
rect 8456 5243 8472 5277
rect 8401 5125 8435 5243
rect 8506 5203 8540 5345
rect 8715 5347 8731 5381
rect 8765 5347 8781 5381
rect 8715 5331 8781 5347
rect 8823 5351 8843 5385
rect 8877 5351 8893 5385
rect 8937 5381 9127 5389
rect 8615 5253 8653 5287
rect 8687 5271 8739 5287
rect 8823 5273 8875 5351
rect 8937 5347 8953 5381
rect 8987 5347 9127 5381
rect 8937 5333 9127 5347
rect 9161 5385 9199 5423
rect 9161 5351 9165 5385
rect 9496 5381 9557 5423
rect 9161 5335 9199 5351
rect 9233 5365 9447 5381
rect 9233 5347 9383 5365
rect 8581 5237 8677 5253
rect 8711 5237 8739 5271
rect 8773 5223 8807 5239
rect 8342 5109 8435 5125
rect 8376 5083 8435 5109
rect 8376 5075 8401 5083
rect 8229 5039 8308 5073
rect 8342 5049 8401 5075
rect 8342 5047 8435 5049
rect 8469 5189 8773 5203
rect 8469 5169 8807 5189
rect 8274 5013 8308 5039
rect 8469 5013 8503 5169
rect 8841 5135 8875 5273
rect 8575 5101 8591 5135
rect 8625 5101 8875 5135
rect 8913 5283 8955 5299
rect 8913 5249 8921 5283
rect 8913 5141 8955 5249
rect 8989 5235 9059 5299
rect 8989 5201 9017 5235
rect 9051 5219 9059 5235
rect 8989 5185 9025 5201
rect 8989 5175 9059 5185
rect 9093 5177 9127 5333
rect 9233 5301 9267 5347
rect 9417 5331 9447 5365
rect 9496 5347 9507 5381
rect 9541 5347 9557 5381
rect 9496 5331 9557 5347
rect 9591 5331 9642 5387
rect 9161 5267 9267 5301
rect 9301 5287 9349 5313
rect 9161 5261 9205 5267
rect 9195 5227 9205 5261
rect 9335 5253 9349 5287
rect 9301 5233 9349 5253
rect 9161 5211 9205 5227
rect 9241 5224 9257 5233
rect 9291 5199 9349 5233
rect 9275 5190 9349 5199
rect 9093 5143 9174 5177
rect 9241 5159 9349 5190
rect 9383 5276 9447 5331
rect 9625 5297 9642 5331
rect 9591 5281 9642 5297
rect 9383 5241 9448 5276
rect 9383 5225 9566 5241
rect 9383 5191 9532 5225
rect 9383 5181 9566 5191
rect 9418 5175 9566 5181
rect 8913 5109 9048 5141
rect 9140 5125 9174 5143
rect 8913 5107 9056 5109
rect 8841 5073 8875 5101
rect 9014 5083 9056 5107
rect 8190 4989 8240 5005
rect 8190 4955 8206 4989
rect 8190 4913 8240 4955
rect 8274 4997 8324 5013
rect 8274 4963 8290 4997
rect 8274 4947 8324 4963
rect 8367 4991 8503 5013
rect 8367 4957 8383 4991
rect 8417 4957 8503 4991
rect 8537 5033 8752 5067
rect 8841 5039 8953 5073
rect 9014 5049 9025 5083
rect 9090 5075 9106 5109
rect 9059 5049 9106 5075
rect 9140 5091 9334 5125
rect 9368 5091 9384 5125
rect 8537 5015 8571 5033
rect 8718 5015 8752 5033
rect 8537 4965 8571 4981
rect 8618 4965 8634 4999
rect 8668 4965 8684 4999
rect 8718 4965 8752 4981
rect 8811 4989 8885 5005
rect 8367 4947 8503 4957
rect 8618 4913 8684 4965
rect 8811 4955 8831 4989
rect 8865 4955 8885 4989
rect 8811 4913 8885 4955
rect 8919 4997 8953 5039
rect 9140 5015 9174 5091
rect 9418 5057 9452 5175
rect 9600 5151 9642 5281
rect 9677 5355 10011 5423
rect 9677 5321 9695 5355
rect 9729 5321 9959 5355
rect 9993 5321 10011 5355
rect 9677 5269 10011 5321
rect 10100 5366 10149 5382
rect 10100 5332 10109 5366
rect 10143 5332 10149 5366
rect 9677 5199 9827 5269
rect 10100 5261 10149 5332
rect 10193 5366 10295 5423
rect 10227 5332 10261 5366
rect 10193 5316 10295 5332
rect 10331 5287 10369 5389
rect 9677 5165 9697 5199
rect 9731 5165 9827 5199
rect 9861 5201 9957 5235
rect 9991 5201 10011 5235
rect 8919 4947 8953 4963
rect 9000 4990 9174 5015
rect 9292 5023 9452 5057
rect 9496 5057 9557 5141
rect 9496 5023 9507 5057
rect 9541 5023 9557 5057
rect 9292 5015 9326 5023
rect 9000 4956 9016 4990
rect 9050 4956 9174 4990
rect 9000 4947 9174 4956
rect 9208 4989 9258 5005
rect 9242 4955 9258 4989
rect 9496 4989 9557 5023
rect 9292 4965 9326 4981
rect 9208 4913 9258 4955
rect 9362 4955 9378 4989
rect 9412 4955 9428 4989
rect 9362 4913 9428 4955
rect 9496 4955 9507 4989
rect 9541 4955 9557 4989
rect 9591 5093 9642 5151
rect 9861 5131 10011 5201
rect 9625 5059 9642 5093
rect 9591 5025 9642 5059
rect 9625 5015 9642 5025
rect 9591 4981 9597 4991
rect 9631 4981 9642 5015
rect 9591 4975 9642 4981
rect 9677 5091 10011 5131
rect 9677 5057 9695 5091
rect 9729 5057 9959 5091
rect 9993 5057 10011 5091
rect 9677 4989 10011 5057
rect 9496 4913 9557 4955
rect 9677 4955 9695 4989
rect 9729 4955 9959 4989
rect 9993 4955 10011 4989
rect 10045 5227 10241 5261
rect 10275 5227 10291 5261
rect 10331 5253 10333 5287
rect 10367 5253 10369 5287
rect 10045 5065 10113 5227
rect 10147 5151 10297 5152
rect 10147 5117 10149 5151
rect 10183 5148 10297 5151
rect 10147 5114 10163 5117
rect 10197 5114 10297 5148
rect 10045 5049 10148 5065
rect 10045 5015 10109 5049
rect 10143 5015 10148 5049
rect 10045 4983 10148 5015
rect 10195 5049 10229 5065
rect 9677 4913 10011 4955
rect 10195 4913 10229 5015
rect 10263 4981 10297 5114
rect 10331 5148 10369 5253
rect 10403 5355 10458 5389
rect 10496 5366 10602 5389
rect 10403 5321 10425 5355
rect 10530 5332 10602 5366
rect 10687 5381 10753 5423
rect 10687 5347 10703 5381
rect 10737 5347 10753 5381
rect 10687 5343 10753 5347
rect 10787 5362 10838 5389
rect 10403 5261 10458 5321
rect 10496 5316 10602 5332
rect 10567 5309 10602 5316
rect 10821 5328 10838 5362
rect 10437 5227 10458 5261
rect 10403 5157 10458 5227
rect 10499 5261 10533 5277
rect 10365 5117 10369 5148
rect 10499 5117 10533 5227
rect 10365 5114 10533 5117
rect 10331 5083 10533 5114
rect 10567 5275 10753 5309
rect 10787 5275 10838 5328
rect 10567 5049 10601 5275
rect 10719 5241 10753 5275
rect 10376 5015 10392 5049
rect 10426 5015 10467 5049
rect 10501 5015 10601 5049
rect 10635 5225 10674 5241
rect 10635 5191 10640 5225
rect 10635 5175 10674 5191
rect 10719 5225 10770 5241
rect 10719 5191 10736 5225
rect 10719 5175 10770 5191
rect 10635 4981 10669 5175
rect 10804 5141 10838 5275
rect 10873 5362 11391 5423
rect 10873 5328 10891 5362
rect 10925 5328 11339 5362
rect 11373 5328 11391 5362
rect 10873 5269 11391 5328
rect 11425 5329 11483 5423
rect 11425 5295 11437 5329
rect 11471 5295 11483 5329
rect 11425 5278 11483 5295
rect 11702 5362 11753 5389
rect 11702 5355 11719 5362
rect 11702 5321 11713 5355
rect 11787 5381 11853 5423
rect 11787 5347 11803 5381
rect 11837 5347 11853 5381
rect 11787 5343 11853 5347
rect 11938 5366 12044 5389
rect 11747 5321 11753 5328
rect 11702 5275 11753 5321
rect 11938 5332 12010 5366
rect 11938 5316 12044 5332
rect 11938 5309 11973 5316
rect 11787 5275 11973 5309
rect 12082 5287 12137 5389
rect 10873 5199 11115 5269
rect 10873 5165 10951 5199
rect 10985 5165 11061 5199
rect 11095 5165 11115 5199
rect 11149 5201 11169 5235
rect 11203 5201 11279 5235
rect 11313 5201 11391 5235
rect 10263 4947 10669 4981
rect 10703 5125 10737 5141
rect 10703 5057 10737 5091
rect 10703 4989 10737 5023
rect 10703 4913 10737 4955
rect 10771 5125 10838 5141
rect 11149 5131 11391 5201
rect 10771 5091 10787 5125
rect 10821 5091 10838 5125
rect 10771 5057 10838 5091
rect 10771 5023 10787 5057
rect 10821 5023 10838 5057
rect 10771 5015 10838 5023
rect 10771 4989 10793 5015
rect 10771 4955 10787 4989
rect 10827 4981 10838 5015
rect 10821 4955 10838 4981
rect 10771 4947 10838 4955
rect 10873 5091 11391 5131
rect 10873 5057 10891 5091
rect 10925 5057 11339 5091
rect 11373 5057 11391 5091
rect 10873 4989 11391 5057
rect 10873 4955 10891 4989
rect 10925 4955 11339 4989
rect 11373 4955 11391 4989
rect 10873 4913 11391 4955
rect 11425 5111 11483 5146
rect 11425 5077 11437 5111
rect 11471 5077 11483 5111
rect 11425 5018 11483 5077
rect 11425 4984 11437 5018
rect 11471 4984 11483 5018
rect 11425 4913 11483 4984
rect 11702 5141 11736 5275
rect 11787 5241 11821 5275
rect 11770 5225 11821 5241
rect 11804 5191 11821 5225
rect 11770 5175 11821 5191
rect 11866 5225 11905 5241
rect 11900 5191 11905 5225
rect 11866 5175 11905 5191
rect 11702 5125 11769 5141
rect 11702 5091 11719 5125
rect 11753 5091 11769 5125
rect 11702 5057 11769 5091
rect 11702 5023 11719 5057
rect 11753 5023 11769 5057
rect 11702 4989 11769 5023
rect 11702 4955 11719 4989
rect 11753 4955 11769 4989
rect 11702 4947 11769 4955
rect 11803 5125 11837 5141
rect 11803 5057 11837 5091
rect 11803 4989 11837 5023
rect 11803 4913 11837 4955
rect 11871 4981 11905 5175
rect 11939 5049 11973 5275
rect 12007 5261 12041 5277
rect 12115 5261 12137 5287
rect 12007 5117 12041 5227
rect 12082 5227 12103 5253
rect 12082 5157 12137 5227
rect 12171 5355 12209 5389
rect 12171 5321 12173 5355
rect 12207 5321 12209 5355
rect 12171 5148 12209 5321
rect 12245 5366 12347 5423
rect 12279 5332 12313 5366
rect 12245 5316 12347 5332
rect 12391 5366 12440 5382
rect 12391 5332 12397 5366
rect 12431 5332 12440 5366
rect 12391 5261 12440 5332
rect 12529 5355 12863 5423
rect 12529 5321 12547 5355
rect 12581 5321 12811 5355
rect 12845 5321 12863 5355
rect 12529 5269 12863 5321
rect 12952 5366 13001 5382
rect 12952 5332 12961 5366
rect 12995 5332 13001 5366
rect 12249 5227 12265 5261
rect 12299 5227 12495 5261
rect 12171 5117 12175 5148
rect 12007 5114 12175 5117
rect 12007 5083 12209 5114
rect 12243 5151 12393 5152
rect 12243 5117 12265 5151
rect 12299 5148 12393 5151
rect 12299 5117 12343 5148
rect 12243 5114 12343 5117
rect 12377 5114 12393 5148
rect 11939 5015 12039 5049
rect 12073 5015 12114 5049
rect 12148 5015 12164 5049
rect 12243 4981 12277 5114
rect 12427 5065 12495 5227
rect 12529 5199 12679 5269
rect 12952 5261 13001 5332
rect 13045 5366 13147 5423
rect 13079 5332 13113 5366
rect 13045 5316 13147 5332
rect 13183 5355 13221 5389
rect 13183 5321 13185 5355
rect 13219 5321 13221 5355
rect 12529 5165 12549 5199
rect 12583 5165 12679 5199
rect 12713 5201 12809 5235
rect 12843 5201 12863 5235
rect 12713 5131 12863 5201
rect 11871 4947 12277 4981
rect 12311 5049 12345 5065
rect 12311 4913 12345 5015
rect 12392 5049 12495 5065
rect 12392 5015 12397 5049
rect 12431 5015 12495 5049
rect 12392 4983 12495 5015
rect 12529 5091 12863 5131
rect 12529 5057 12547 5091
rect 12581 5057 12811 5091
rect 12845 5057 12863 5091
rect 12529 4989 12863 5057
rect 12529 4955 12547 4989
rect 12581 4955 12811 4989
rect 12845 4955 12863 4989
rect 12897 5227 13093 5261
rect 13127 5227 13143 5261
rect 12897 5065 12965 5227
rect 12999 5151 13149 5152
rect 12999 5148 13093 5151
rect 12999 5114 13015 5148
rect 13049 5117 13093 5148
rect 13127 5117 13149 5151
rect 13049 5114 13149 5117
rect 12897 5049 13000 5065
rect 12897 5015 12961 5049
rect 12995 5015 13000 5049
rect 12897 4983 13000 5015
rect 13047 5049 13081 5065
rect 12529 4913 12863 4955
rect 13047 4913 13081 5015
rect 13115 4981 13149 5114
rect 13183 5148 13221 5321
rect 13255 5261 13310 5389
rect 13348 5366 13454 5389
rect 13382 5332 13454 5366
rect 13539 5381 13605 5423
rect 13539 5347 13555 5381
rect 13589 5347 13605 5381
rect 13539 5343 13605 5347
rect 13639 5362 13690 5389
rect 13348 5316 13454 5332
rect 13419 5309 13454 5316
rect 13673 5328 13690 5362
rect 13289 5227 13310 5261
rect 13255 5219 13310 5227
rect 13351 5261 13385 5277
rect 13255 5185 13277 5219
rect 13255 5157 13310 5185
rect 13217 5117 13221 5148
rect 13351 5117 13385 5227
rect 13217 5114 13385 5117
rect 13183 5083 13385 5114
rect 13419 5275 13605 5309
rect 13639 5275 13690 5328
rect 13725 5362 14794 5423
rect 13725 5328 13743 5362
rect 13777 5328 14743 5362
rect 14777 5328 14794 5362
rect 13725 5314 14794 5328
rect 14829 5362 15898 5423
rect 14829 5328 14847 5362
rect 14881 5328 15847 5362
rect 15881 5328 15898 5362
rect 14829 5314 15898 5328
rect 15933 5362 16451 5423
rect 15933 5328 15951 5362
rect 15985 5328 16399 5362
rect 16433 5328 16451 5362
rect 13419 5049 13453 5275
rect 13571 5241 13605 5275
rect 13228 5015 13244 5049
rect 13278 5015 13319 5049
rect 13353 5015 13453 5049
rect 13487 5225 13526 5241
rect 13487 5191 13492 5225
rect 13487 5175 13526 5191
rect 13571 5225 13622 5241
rect 13571 5191 13588 5225
rect 13571 5175 13622 5191
rect 13487 4981 13521 5175
rect 13656 5141 13690 5275
rect 14042 5199 14110 5314
rect 14042 5165 14059 5199
rect 14093 5165 14110 5199
rect 14042 5148 14110 5165
rect 14406 5235 14476 5250
rect 14406 5201 14423 5235
rect 14457 5201 14476 5235
rect 13115 4947 13521 4981
rect 13555 5125 13589 5141
rect 13555 5057 13589 5091
rect 13555 4989 13589 5023
rect 13555 4913 13589 4955
rect 13623 5125 13690 5141
rect 13623 5091 13639 5125
rect 13673 5091 13690 5125
rect 13623 5057 13690 5091
rect 13623 5023 13639 5057
rect 13673 5023 13690 5057
rect 13623 5015 13690 5023
rect 13623 4989 13645 5015
rect 13623 4955 13639 4989
rect 13679 4981 13690 5015
rect 14406 5000 14476 5201
rect 15146 5199 15214 5314
rect 15933 5269 16451 5328
rect 16577 5329 16635 5423
rect 16577 5295 16589 5329
rect 16623 5295 16635 5329
rect 16669 5362 17738 5423
rect 16669 5328 16687 5362
rect 16721 5328 17687 5362
rect 17721 5328 17738 5362
rect 16669 5314 17738 5328
rect 17773 5362 18475 5423
rect 17773 5328 17791 5362
rect 17825 5328 18423 5362
rect 18457 5328 18475 5362
rect 16577 5278 16635 5295
rect 15146 5165 15163 5199
rect 15197 5165 15214 5199
rect 15146 5148 15214 5165
rect 15510 5235 15580 5250
rect 15510 5201 15527 5235
rect 15561 5201 15580 5235
rect 15510 5000 15580 5201
rect 15933 5199 16175 5269
rect 15933 5165 16011 5199
rect 16045 5165 16121 5199
rect 16155 5165 16175 5199
rect 16209 5201 16229 5235
rect 16263 5201 16339 5235
rect 16373 5201 16451 5235
rect 16209 5131 16451 5201
rect 16986 5199 17054 5314
rect 17773 5269 18475 5328
rect 18601 5360 18843 5423
rect 18601 5326 18619 5360
rect 18653 5326 18791 5360
rect 18825 5326 18843 5360
rect 18601 5273 18843 5326
rect 16986 5165 17003 5199
rect 17037 5165 17054 5199
rect 16986 5148 17054 5165
rect 17350 5235 17420 5250
rect 17350 5201 17367 5235
rect 17401 5201 17420 5235
rect 15933 5091 16451 5131
rect 15933 5057 15951 5091
rect 15985 5057 16399 5091
rect 16433 5057 16451 5091
rect 13673 4955 13690 4981
rect 13623 4947 13690 4955
rect 13725 4989 14794 5000
rect 13725 4955 13743 4989
rect 13777 4955 14743 4989
rect 14777 4955 14794 4989
rect 13725 4913 14794 4955
rect 14829 4989 15898 5000
rect 14829 4955 14847 4989
rect 14881 4955 15847 4989
rect 15881 4955 15898 4989
rect 14829 4913 15898 4955
rect 15933 4989 16451 5057
rect 15933 4955 15951 4989
rect 15985 4955 16399 4989
rect 16433 4955 16451 4989
rect 15933 4913 16451 4955
rect 16577 5111 16635 5146
rect 16577 5077 16589 5111
rect 16623 5077 16635 5111
rect 16577 5018 16635 5077
rect 16577 4984 16589 5018
rect 16623 4984 16635 5018
rect 17350 5000 17420 5201
rect 17773 5199 18103 5269
rect 17773 5165 17851 5199
rect 17885 5165 17950 5199
rect 17984 5165 18049 5199
rect 18083 5165 18103 5199
rect 18137 5201 18157 5235
rect 18191 5201 18260 5235
rect 18294 5201 18363 5235
rect 18397 5201 18475 5235
rect 18137 5131 18475 5201
rect 17773 5091 18475 5131
rect 17773 5057 17791 5091
rect 17825 5057 18423 5091
rect 18457 5057 18475 5091
rect 16577 4913 16635 4984
rect 16669 4989 17738 5000
rect 16669 4955 16687 4989
rect 16721 4955 17687 4989
rect 17721 4955 17738 4989
rect 16669 4913 17738 4955
rect 17773 4989 18475 5057
rect 17773 4955 17791 4989
rect 17825 4955 18423 4989
rect 18457 4955 18475 4989
rect 17773 4913 18475 4955
rect 18601 5205 18651 5239
rect 18685 5205 18705 5239
rect 18601 5131 18705 5205
rect 18739 5199 18843 5273
rect 18739 5165 18759 5199
rect 18793 5165 18843 5199
rect 18601 5084 18843 5131
rect 18601 5050 18619 5084
rect 18653 5050 18791 5084
rect 18825 5050 18843 5084
rect 18601 4989 18843 5050
rect 18601 4955 18619 4989
rect 18653 4955 18791 4989
rect 18825 4955 18843 4989
rect 18601 4913 18843 4955
rect 1104 4879 1133 4913
rect 1167 4879 1225 4913
rect 1259 4879 1317 4913
rect 1351 4879 1409 4913
rect 1443 4879 1501 4913
rect 1535 4879 1593 4913
rect 1627 4879 1685 4913
rect 1719 4879 1777 4913
rect 1811 4879 1869 4913
rect 1903 4879 1961 4913
rect 1995 4879 2053 4913
rect 2087 4879 2145 4913
rect 2179 4879 2237 4913
rect 2271 4879 2329 4913
rect 2363 4879 2421 4913
rect 2455 4879 2513 4913
rect 2547 4879 2605 4913
rect 2639 4879 2697 4913
rect 2731 4879 2789 4913
rect 2823 4879 2881 4913
rect 2915 4879 2973 4913
rect 3007 4879 3065 4913
rect 3099 4879 3157 4913
rect 3191 4879 3249 4913
rect 3283 4879 3341 4913
rect 3375 4879 3433 4913
rect 3467 4879 3525 4913
rect 3559 4879 3617 4913
rect 3651 4879 3709 4913
rect 3743 4879 3801 4913
rect 3835 4879 3893 4913
rect 3927 4879 3985 4913
rect 4019 4879 4077 4913
rect 4111 4879 4169 4913
rect 4203 4879 4261 4913
rect 4295 4879 4353 4913
rect 4387 4879 4445 4913
rect 4479 4879 4537 4913
rect 4571 4879 4629 4913
rect 4663 4879 4721 4913
rect 4755 4879 4813 4913
rect 4847 4879 4905 4913
rect 4939 4879 4997 4913
rect 5031 4879 5089 4913
rect 5123 4879 5181 4913
rect 5215 4879 5273 4913
rect 5307 4879 5365 4913
rect 5399 4879 5457 4913
rect 5491 4879 5549 4913
rect 5583 4879 5641 4913
rect 5675 4879 5733 4913
rect 5767 4879 5825 4913
rect 5859 4879 5917 4913
rect 5951 4879 6009 4913
rect 6043 4879 6101 4913
rect 6135 4879 6193 4913
rect 6227 4879 6285 4913
rect 6319 4879 6377 4913
rect 6411 4879 6469 4913
rect 6503 4879 6561 4913
rect 6595 4879 6653 4913
rect 6687 4879 6745 4913
rect 6779 4879 6837 4913
rect 6871 4879 6929 4913
rect 6963 4879 7021 4913
rect 7055 4879 7113 4913
rect 7147 4879 7205 4913
rect 7239 4879 7297 4913
rect 7331 4879 7389 4913
rect 7423 4879 7481 4913
rect 7515 4879 7573 4913
rect 7607 4879 7665 4913
rect 7699 4879 7757 4913
rect 7791 4879 7849 4913
rect 7883 4879 7941 4913
rect 7975 4879 8033 4913
rect 8067 4879 8125 4913
rect 8159 4879 8217 4913
rect 8251 4879 8309 4913
rect 8343 4879 8401 4913
rect 8435 4879 8493 4913
rect 8527 4879 8585 4913
rect 8619 4879 8677 4913
rect 8711 4879 8769 4913
rect 8803 4879 8861 4913
rect 8895 4879 8953 4913
rect 8987 4879 9045 4913
rect 9079 4879 9137 4913
rect 9171 4879 9229 4913
rect 9263 4879 9321 4913
rect 9355 4879 9413 4913
rect 9447 4879 9505 4913
rect 9539 4879 9597 4913
rect 9631 4879 9689 4913
rect 9723 4879 9781 4913
rect 9815 4879 9873 4913
rect 9907 4879 9965 4913
rect 9999 4879 10057 4913
rect 10091 4879 10149 4913
rect 10183 4879 10241 4913
rect 10275 4879 10333 4913
rect 10367 4879 10425 4913
rect 10459 4879 10517 4913
rect 10551 4879 10609 4913
rect 10643 4879 10701 4913
rect 10735 4879 10793 4913
rect 10827 4879 10885 4913
rect 10919 4879 10977 4913
rect 11011 4879 11069 4913
rect 11103 4879 11161 4913
rect 11195 4879 11253 4913
rect 11287 4879 11345 4913
rect 11379 4879 11437 4913
rect 11471 4879 11529 4913
rect 11563 4879 11621 4913
rect 11655 4879 11713 4913
rect 11747 4879 11805 4913
rect 11839 4879 11897 4913
rect 11931 4879 11989 4913
rect 12023 4879 12081 4913
rect 12115 4879 12173 4913
rect 12207 4879 12265 4913
rect 12299 4879 12357 4913
rect 12391 4879 12449 4913
rect 12483 4879 12541 4913
rect 12575 4879 12633 4913
rect 12667 4879 12725 4913
rect 12759 4879 12817 4913
rect 12851 4879 12909 4913
rect 12943 4879 13001 4913
rect 13035 4879 13093 4913
rect 13127 4879 13185 4913
rect 13219 4879 13277 4913
rect 13311 4879 13369 4913
rect 13403 4879 13461 4913
rect 13495 4879 13553 4913
rect 13587 4879 13645 4913
rect 13679 4879 13737 4913
rect 13771 4879 13829 4913
rect 13863 4879 13921 4913
rect 13955 4879 14013 4913
rect 14047 4879 14105 4913
rect 14139 4879 14197 4913
rect 14231 4879 14289 4913
rect 14323 4879 14381 4913
rect 14415 4879 14473 4913
rect 14507 4879 14565 4913
rect 14599 4879 14657 4913
rect 14691 4879 14749 4913
rect 14783 4879 14841 4913
rect 14875 4879 14933 4913
rect 14967 4879 15025 4913
rect 15059 4879 15117 4913
rect 15151 4879 15209 4913
rect 15243 4879 15301 4913
rect 15335 4879 15393 4913
rect 15427 4879 15485 4913
rect 15519 4879 15577 4913
rect 15611 4879 15669 4913
rect 15703 4879 15761 4913
rect 15795 4879 15853 4913
rect 15887 4879 15945 4913
rect 15979 4879 16037 4913
rect 16071 4879 16129 4913
rect 16163 4879 16221 4913
rect 16255 4879 16313 4913
rect 16347 4879 16405 4913
rect 16439 4879 16497 4913
rect 16531 4879 16589 4913
rect 16623 4879 16681 4913
rect 16715 4879 16773 4913
rect 16807 4879 16865 4913
rect 16899 4879 16957 4913
rect 16991 4879 17049 4913
rect 17083 4879 17141 4913
rect 17175 4879 17233 4913
rect 17267 4879 17325 4913
rect 17359 4879 17417 4913
rect 17451 4879 17509 4913
rect 17543 4879 17601 4913
rect 17635 4879 17693 4913
rect 17727 4879 17785 4913
rect 17819 4879 17877 4913
rect 17911 4879 17969 4913
rect 18003 4879 18061 4913
rect 18095 4879 18153 4913
rect 18187 4879 18245 4913
rect 18279 4879 18337 4913
rect 18371 4879 18429 4913
rect 18463 4879 18521 4913
rect 18555 4879 18613 4913
rect 18647 4879 18705 4913
rect 18739 4879 18797 4913
rect 18831 4879 18860 4913
rect 1121 4837 1363 4879
rect 1121 4803 1139 4837
rect 1173 4803 1311 4837
rect 1345 4803 1363 4837
rect 1121 4742 1363 4803
rect 1121 4708 1139 4742
rect 1173 4708 1311 4742
rect 1345 4708 1363 4742
rect 1121 4661 1363 4708
rect 1397 4837 2099 4879
rect 1397 4803 1415 4837
rect 1449 4803 2047 4837
rect 2081 4803 2099 4837
rect 1397 4735 2099 4803
rect 1397 4701 1415 4735
rect 1449 4701 2047 4735
rect 2081 4701 2099 4735
rect 1397 4661 2099 4701
rect 2133 4837 2375 4879
rect 2133 4803 2151 4837
rect 2185 4803 2323 4837
rect 2357 4803 2375 4837
rect 2133 4742 2375 4803
rect 2133 4708 2151 4742
rect 2185 4708 2323 4742
rect 2357 4708 2375 4742
rect 2133 4661 2375 4708
rect 1121 4593 1171 4627
rect 1205 4593 1225 4627
rect 1121 4519 1225 4593
rect 1259 4587 1363 4661
rect 1259 4553 1279 4587
rect 1313 4553 1363 4587
rect 1397 4593 1475 4627
rect 1509 4593 1574 4627
rect 1608 4593 1673 4627
rect 1707 4593 1727 4627
rect 1397 4523 1727 4593
rect 1761 4591 2099 4661
rect 1761 4557 1781 4591
rect 1815 4557 1884 4591
rect 1918 4557 1987 4591
rect 2021 4557 2099 4591
rect 2133 4593 2183 4627
rect 2217 4593 2237 4627
rect 1121 4466 1363 4519
rect 1121 4432 1139 4466
rect 1173 4432 1311 4466
rect 1345 4432 1363 4466
rect 1121 4369 1363 4432
rect 1397 4464 2099 4523
rect 1397 4430 1415 4464
rect 1449 4430 2047 4464
rect 2081 4430 2099 4464
rect 1397 4369 2099 4430
rect 2133 4519 2237 4593
rect 2271 4587 2375 4661
rect 2271 4553 2291 4587
rect 2325 4553 2375 4587
rect 2409 4811 2486 4845
rect 2409 4777 2446 4811
rect 2480 4777 2486 4811
rect 2520 4837 2585 4879
rect 2520 4803 2536 4837
rect 2570 4803 2585 4837
rect 2520 4787 2585 4803
rect 2689 4811 2745 4845
rect 2409 4651 2486 4777
rect 2689 4777 2695 4811
rect 2729 4777 2745 4811
rect 2689 4753 2745 4777
rect 2520 4709 2745 4753
rect 2783 4811 2863 4845
rect 2783 4777 2799 4811
rect 2833 4777 2863 4811
rect 2943 4837 2997 4879
rect 2943 4803 2953 4837
rect 2987 4803 2997 4837
rect 2943 4787 2997 4803
rect 3031 4811 3088 4845
rect 2133 4466 2375 4519
rect 2133 4432 2151 4466
rect 2185 4432 2323 4466
rect 2357 4432 2375 4466
rect 2133 4369 2375 4432
rect 2409 4517 2465 4651
rect 2520 4617 2610 4709
rect 2783 4675 2863 4777
rect 3031 4777 3037 4811
rect 3071 4777 3088 4811
rect 3031 4753 3088 4777
rect 2499 4601 2610 4617
rect 2533 4567 2610 4601
rect 2499 4551 2610 4567
rect 2644 4601 2863 4675
rect 2644 4567 2695 4601
rect 2729 4567 2863 4601
rect 2644 4563 2863 4567
rect 2520 4529 2610 4551
rect 2409 4471 2486 4517
rect 2520 4495 2745 4529
rect 2409 4437 2421 4471
rect 2480 4437 2486 4471
rect 2689 4471 2745 4495
rect 2409 4403 2486 4437
rect 2520 4445 2585 4461
rect 2520 4411 2536 4445
rect 2570 4411 2585 4445
rect 2520 4369 2585 4411
rect 2689 4437 2695 4471
rect 2729 4437 2745 4471
rect 2689 4403 2745 4437
rect 2783 4471 2863 4563
rect 2897 4709 3088 4753
rect 3145 4837 3663 4879
rect 3145 4803 3163 4837
rect 3197 4803 3611 4837
rect 3645 4803 3663 4837
rect 3145 4735 3663 4803
rect 2897 4601 2939 4709
rect 3145 4701 3163 4735
rect 3197 4701 3611 4735
rect 3645 4701 3663 4735
rect 2897 4567 2899 4601
rect 2933 4567 2939 4601
rect 2897 4529 2939 4567
rect 2973 4607 3111 4675
rect 3145 4661 3663 4701
rect 2973 4601 3065 4607
rect 2973 4567 3013 4601
rect 3047 4573 3065 4601
rect 3099 4573 3111 4607
rect 3047 4567 3111 4573
rect 2973 4563 3111 4567
rect 3145 4593 3223 4627
rect 3257 4593 3333 4627
rect 3367 4593 3387 4627
rect 2897 4495 3088 4529
rect 2783 4437 2799 4471
rect 2833 4437 2863 4471
rect 3031 4471 3088 4495
rect 2783 4403 2863 4437
rect 2943 4445 2997 4461
rect 2943 4411 2953 4445
rect 2987 4411 2997 4445
rect 2943 4369 2997 4411
rect 3031 4437 3037 4471
rect 3071 4437 3088 4471
rect 3031 4403 3088 4437
rect 3145 4523 3387 4593
rect 3421 4591 3663 4661
rect 3697 4808 3755 4879
rect 3697 4774 3709 4808
rect 3743 4774 3755 4808
rect 3697 4715 3755 4774
rect 3697 4681 3709 4715
rect 3743 4681 3755 4715
rect 3984 4823 4041 4879
rect 3984 4789 3999 4823
rect 4033 4789 4041 4823
rect 3984 4755 4041 4789
rect 3984 4721 3999 4755
rect 4033 4721 4041 4755
rect 3984 4705 4041 4721
rect 4075 4829 4127 4845
rect 4075 4795 4085 4829
rect 4119 4795 4127 4829
rect 4075 4761 4127 4795
rect 4162 4837 4213 4879
rect 4162 4803 4171 4837
rect 4205 4803 4213 4837
rect 4162 4787 4213 4803
rect 4247 4802 4299 4845
rect 4075 4727 4085 4761
rect 4119 4753 4127 4761
rect 4247 4768 4257 4802
rect 4291 4768 4299 4802
rect 4247 4753 4299 4768
rect 4119 4727 4299 4753
rect 4075 4719 4299 4727
rect 4333 4837 4395 4879
rect 4333 4803 4353 4837
rect 4387 4803 4395 4837
rect 4333 4769 4395 4803
rect 4333 4735 4353 4769
rect 4387 4735 4395 4769
rect 4333 4719 4395 4735
rect 4429 4829 4491 4845
rect 4429 4795 4439 4829
rect 4473 4795 4491 4829
rect 3697 4646 3755 4681
rect 4075 4693 4127 4719
rect 4075 4669 4085 4693
rect 3976 4659 4085 4669
rect 4119 4659 4127 4693
rect 4429 4707 4491 4795
rect 4429 4685 4439 4707
rect 3421 4557 3441 4591
rect 3475 4557 3551 4591
rect 3585 4557 3663 4591
rect 3976 4635 4127 4659
rect 4285 4673 4439 4685
rect 4473 4673 4491 4707
rect 4285 4651 4491 4673
rect 4525 4837 4859 4879
rect 4525 4803 4543 4837
rect 4577 4803 4807 4837
rect 4841 4803 4859 4837
rect 4525 4735 4859 4803
rect 4525 4701 4543 4735
rect 4577 4701 4807 4735
rect 4841 4701 4859 4735
rect 4525 4661 4859 4701
rect 3976 4533 4057 4635
rect 4285 4601 4319 4651
rect 4091 4567 4107 4601
rect 4141 4567 4175 4601
rect 4209 4567 4243 4601
rect 4277 4567 4319 4601
rect 4353 4601 4423 4617
rect 4353 4567 4389 4601
rect 4353 4539 4423 4567
rect 3145 4464 3663 4523
rect 3145 4430 3163 4464
rect 3197 4430 3611 4464
rect 3645 4430 3663 4464
rect 3145 4369 3663 4430
rect 3697 4497 3755 4514
rect 3976 4499 4306 4533
rect 4387 4505 4423 4539
rect 4353 4503 4423 4505
rect 3697 4463 3709 4497
rect 3743 4463 3755 4497
rect 4075 4471 4127 4499
rect 3697 4369 3755 4463
rect 3985 4449 4041 4465
rect 3985 4415 3998 4449
rect 4032 4415 4041 4449
rect 4075 4437 4077 4471
rect 4118 4437 4127 4471
rect 4247 4471 4306 4499
rect 4075 4421 4127 4437
rect 4162 4449 4213 4465
rect 3985 4369 4041 4415
rect 4162 4415 4170 4449
rect 4204 4415 4213 4449
rect 4247 4437 4256 4471
rect 4290 4437 4306 4471
rect 4457 4469 4491 4651
rect 4247 4421 4306 4437
rect 4342 4449 4397 4465
rect 4162 4369 4213 4415
rect 4342 4415 4353 4449
rect 4387 4415 4397 4449
rect 4342 4369 4397 4415
rect 4431 4453 4491 4469
rect 4431 4419 4439 4453
rect 4473 4419 4491 4453
rect 4431 4403 4491 4419
rect 4525 4593 4545 4627
rect 4579 4593 4675 4627
rect 4525 4523 4675 4593
rect 4709 4591 4859 4661
rect 4709 4557 4805 4591
rect 4839 4557 4859 4591
rect 4893 4607 5043 4845
rect 5077 4837 5779 4879
rect 5077 4803 5095 4837
rect 5129 4803 5727 4837
rect 5761 4803 5779 4837
rect 5077 4735 5779 4803
rect 5077 4701 5095 4735
rect 5129 4701 5727 4735
rect 5761 4701 5779 4735
rect 5077 4661 5779 4701
rect 4893 4573 4905 4607
rect 4939 4573 5043 4607
rect 4525 4471 4859 4523
rect 4525 4437 4543 4471
rect 4577 4437 4807 4471
rect 4841 4437 4859 4471
rect 4525 4369 4859 4437
rect 4893 4511 5043 4573
rect 4893 4477 4911 4511
rect 4945 4477 4986 4511
rect 5020 4477 5043 4511
rect 4893 4443 5043 4477
rect 4893 4409 4911 4443
rect 4945 4409 4986 4443
rect 5020 4409 5043 4443
rect 4893 4403 5043 4409
rect 5077 4593 5155 4627
rect 5189 4593 5254 4627
rect 5288 4593 5353 4627
rect 5387 4593 5407 4627
rect 5077 4523 5407 4593
rect 5441 4591 5779 4661
rect 5441 4557 5461 4591
rect 5495 4557 5564 4591
rect 5598 4557 5667 4591
rect 5701 4557 5779 4591
rect 6004 4837 6111 4845
rect 6004 4803 6061 4837
rect 6095 4803 6111 4837
rect 6004 4769 6111 4803
rect 6004 4735 6061 4769
rect 6095 4735 6111 4769
rect 6004 4721 6111 4735
rect 6145 4821 6211 4879
rect 6145 4787 6161 4821
rect 6195 4787 6211 4821
rect 6145 4753 6211 4787
rect 5077 4464 5779 4523
rect 5077 4430 5095 4464
rect 5129 4430 5727 4464
rect 5761 4430 5779 4464
rect 5077 4369 5779 4430
rect 6004 4517 6067 4721
rect 6145 4719 6161 4753
rect 6195 4719 6211 4753
rect 6457 4837 6791 4879
rect 6457 4803 6475 4837
rect 6509 4803 6739 4837
rect 6773 4803 6791 4837
rect 6457 4735 6791 4803
rect 6308 4701 6386 4720
rect 6308 4685 6330 4701
rect 6101 4667 6330 4685
rect 6364 4667 6386 4701
rect 6101 4651 6386 4667
rect 6457 4701 6475 4735
rect 6509 4701 6739 4735
rect 6773 4701 6791 4735
rect 7037 4821 7103 4879
rect 7037 4787 7053 4821
rect 7087 4787 7103 4821
rect 7037 4753 7103 4787
rect 6457 4661 6791 4701
rect 6101 4601 6135 4651
rect 6101 4551 6135 4567
rect 6185 4601 6238 4617
rect 6185 4567 6204 4601
rect 6185 4539 6238 4567
rect 6004 4515 6127 4517
rect 6004 4481 6077 4515
rect 6111 4481 6127 4515
rect 6185 4505 6193 4539
rect 6227 4505 6238 4539
rect 6004 4471 6127 4481
rect 6272 4471 6306 4651
rect 6340 4607 6411 4617
rect 6340 4601 6377 4607
rect 6374 4573 6377 4601
rect 6374 4567 6411 4573
rect 6340 4505 6411 4567
rect 6457 4593 6477 4627
rect 6511 4593 6607 4627
rect 6457 4523 6607 4593
rect 6641 4591 6791 4661
rect 6862 4701 6940 4720
rect 7037 4719 7053 4753
rect 7087 4719 7103 4753
rect 7137 4837 7244 4845
rect 7137 4803 7153 4837
rect 7187 4811 7244 4837
rect 7187 4803 7205 4811
rect 7137 4777 7205 4803
rect 7239 4777 7244 4811
rect 7137 4769 7244 4777
rect 7137 4735 7153 4769
rect 7187 4735 7244 4769
rect 7137 4721 7244 4735
rect 6862 4667 6884 4701
rect 6918 4685 6940 4701
rect 6918 4667 7147 4685
rect 6862 4651 7147 4667
rect 6641 4557 6737 4591
rect 6771 4557 6791 4591
rect 6837 4607 6908 4617
rect 6871 4601 6908 4607
rect 6871 4573 6874 4601
rect 6837 4567 6874 4573
rect 6457 4471 6791 4523
rect 6837 4505 6908 4567
rect 6942 4471 6976 4651
rect 7010 4601 7063 4617
rect 7044 4567 7063 4601
rect 7010 4539 7063 4567
rect 7113 4601 7147 4651
rect 7113 4551 7147 4567
rect 7010 4505 7021 4539
rect 7055 4505 7063 4539
rect 7181 4517 7244 4721
rect 7285 4837 7803 4879
rect 7285 4803 7303 4837
rect 7337 4803 7751 4837
rect 7785 4803 7803 4837
rect 7285 4735 7803 4803
rect 7285 4701 7303 4735
rect 7337 4701 7751 4735
rect 7785 4701 7803 4735
rect 7285 4661 7803 4701
rect 7121 4515 7244 4517
rect 7121 4481 7137 4515
rect 7171 4481 7244 4515
rect 6004 4437 6009 4471
rect 6043 4447 6127 4471
rect 6043 4437 6077 4447
rect 6004 4413 6077 4437
rect 6111 4413 6127 4447
rect 6004 4403 6127 4413
rect 6161 4455 6204 4471
rect 6161 4421 6162 4455
rect 6196 4421 6204 4455
rect 6161 4369 6204 4421
rect 6250 4455 6306 4471
rect 6250 4421 6258 4455
rect 6292 4421 6306 4455
rect 6250 4405 6306 4421
rect 6342 4455 6390 4471
rect 6376 4421 6390 4455
rect 6342 4369 6390 4421
rect 6457 4437 6475 4471
rect 6509 4437 6739 4471
rect 6773 4437 6791 4471
rect 6457 4369 6791 4437
rect 6858 4455 6906 4471
rect 6858 4421 6872 4455
rect 6858 4369 6906 4421
rect 6942 4455 6998 4471
rect 6942 4421 6956 4455
rect 6990 4421 6998 4455
rect 6942 4405 6998 4421
rect 7044 4455 7087 4471
rect 7044 4421 7052 4455
rect 7086 4421 7087 4455
rect 7044 4369 7087 4421
rect 7121 4447 7244 4481
rect 7121 4413 7137 4447
rect 7171 4413 7244 4447
rect 7121 4403 7244 4413
rect 7285 4593 7363 4627
rect 7397 4593 7473 4627
rect 7507 4593 7527 4627
rect 7285 4523 7527 4593
rect 7561 4591 7803 4661
rect 7561 4557 7581 4591
rect 7615 4557 7691 4591
rect 7725 4557 7803 4591
rect 7838 4837 7905 4845
rect 7838 4803 7855 4837
rect 7889 4803 7905 4837
rect 7838 4769 7905 4803
rect 7838 4743 7855 4769
rect 7838 4709 7849 4743
rect 7889 4735 7905 4769
rect 7883 4709 7905 4735
rect 7838 4701 7905 4709
rect 7838 4667 7855 4701
rect 7889 4667 7905 4701
rect 7838 4651 7905 4667
rect 7939 4837 7973 4879
rect 7939 4769 7973 4803
rect 7939 4701 7973 4735
rect 7939 4651 7973 4667
rect 8007 4811 8413 4845
rect 7285 4464 7803 4523
rect 7285 4430 7303 4464
rect 7337 4430 7751 4464
rect 7785 4430 7803 4464
rect 7285 4369 7803 4430
rect 7838 4517 7872 4651
rect 8007 4617 8041 4811
rect 7906 4601 7957 4617
rect 7940 4567 7957 4601
rect 7906 4551 7957 4567
rect 8002 4601 8041 4617
rect 8036 4567 8041 4601
rect 8002 4551 8041 4567
rect 8075 4743 8175 4777
rect 8209 4743 8250 4777
rect 8284 4743 8300 4777
rect 7923 4517 7957 4551
rect 8075 4517 8109 4743
rect 7838 4464 7889 4517
rect 7923 4483 8109 4517
rect 8143 4678 8345 4709
rect 8143 4675 8311 4678
rect 8143 4565 8177 4675
rect 8307 4644 8311 4675
rect 8143 4515 8177 4531
rect 8218 4565 8273 4635
rect 8218 4531 8239 4565
rect 7838 4430 7855 4464
rect 8074 4476 8109 4483
rect 8074 4460 8180 4476
rect 8218 4471 8273 4531
rect 7838 4403 7889 4430
rect 7923 4445 7989 4449
rect 7923 4411 7939 4445
rect 7973 4411 7989 4445
rect 7923 4369 7989 4411
rect 8074 4426 8146 4460
rect 8251 4437 8273 4471
rect 8074 4403 8180 4426
rect 8218 4403 8273 4437
rect 8307 4607 8345 4644
rect 8379 4678 8413 4811
rect 8447 4777 8481 4879
rect 8447 4727 8481 4743
rect 8528 4777 8631 4809
rect 8528 4743 8533 4777
rect 8567 4743 8631 4777
rect 8528 4727 8631 4743
rect 8379 4675 8479 4678
rect 8379 4641 8401 4675
rect 8435 4644 8479 4675
rect 8513 4644 8529 4678
rect 8435 4641 8529 4644
rect 8379 4640 8529 4641
rect 8307 4573 8309 4607
rect 8343 4573 8345 4607
rect 8307 4403 8345 4573
rect 8563 4565 8631 4727
rect 8849 4808 8907 4879
rect 8849 4774 8861 4808
rect 8895 4774 8907 4808
rect 8849 4715 8907 4774
rect 9337 4821 9403 4879
rect 9337 4787 9353 4821
rect 9387 4787 9403 4821
rect 9337 4753 9403 4787
rect 8849 4681 8861 4715
rect 8895 4681 8907 4715
rect 8849 4646 8907 4681
rect 9162 4701 9240 4720
rect 9337 4719 9353 4753
rect 9387 4719 9403 4753
rect 9437 4837 9544 4845
rect 9437 4803 9453 4837
rect 9487 4803 9544 4837
rect 9437 4769 9544 4803
rect 9437 4735 9453 4769
rect 9487 4735 9544 4769
rect 9437 4721 9544 4735
rect 9162 4667 9184 4701
rect 9218 4685 9240 4701
rect 9218 4667 9447 4685
rect 9162 4651 9447 4667
rect 8385 4531 8401 4565
rect 8435 4531 8631 4565
rect 9137 4601 9208 4617
rect 9137 4567 9174 4601
rect 9137 4539 9208 4567
rect 8381 4460 8483 4476
rect 8415 4426 8449 4460
rect 8381 4369 8483 4426
rect 8527 4460 8576 4531
rect 8527 4426 8533 4460
rect 8567 4426 8576 4460
rect 8527 4410 8576 4426
rect 8849 4497 8907 4514
rect 9171 4505 9208 4539
rect 8849 4463 8861 4497
rect 8895 4463 8907 4497
rect 9242 4471 9276 4651
rect 9310 4601 9363 4617
rect 9344 4567 9363 4601
rect 9310 4539 9363 4567
rect 9413 4601 9447 4651
rect 9413 4551 9447 4567
rect 9310 4505 9321 4539
rect 9355 4505 9363 4539
rect 9481 4517 9544 4721
rect 9585 4837 9919 4879
rect 9585 4803 9603 4837
rect 9637 4803 9867 4837
rect 9901 4803 9919 4837
rect 9585 4735 9919 4803
rect 9585 4701 9603 4735
rect 9637 4701 9867 4735
rect 9901 4701 9919 4735
rect 9585 4661 9919 4701
rect 9421 4515 9544 4517
rect 9421 4481 9437 4515
rect 9471 4481 9544 4515
rect 9421 4471 9544 4481
rect 8849 4369 8907 4463
rect 9158 4455 9206 4471
rect 9158 4421 9172 4455
rect 9158 4369 9206 4421
rect 9242 4455 9298 4471
rect 9242 4421 9256 4455
rect 9290 4421 9298 4455
rect 9242 4405 9298 4421
rect 9344 4455 9387 4471
rect 9344 4421 9352 4455
rect 9386 4421 9387 4455
rect 9344 4369 9387 4421
rect 9421 4447 9505 4471
rect 9421 4413 9437 4447
rect 9471 4437 9505 4447
rect 9539 4437 9544 4471
rect 9471 4413 9544 4437
rect 9421 4403 9544 4413
rect 9585 4593 9605 4627
rect 9639 4593 9735 4627
rect 9585 4523 9735 4593
rect 9769 4591 9919 4661
rect 9769 4557 9865 4591
rect 9899 4557 9919 4591
rect 9953 4607 10103 4845
rect 10137 4837 10471 4879
rect 10137 4803 10155 4837
rect 10189 4803 10419 4837
rect 10453 4803 10471 4837
rect 10137 4735 10471 4803
rect 10137 4701 10155 4735
rect 10189 4701 10419 4735
rect 10453 4701 10471 4735
rect 10717 4821 10783 4879
rect 10717 4787 10733 4821
rect 10767 4787 10783 4821
rect 10717 4753 10783 4787
rect 10137 4661 10471 4701
rect 9953 4573 9965 4607
rect 9999 4573 10103 4607
rect 9585 4471 9919 4523
rect 9585 4437 9603 4471
rect 9637 4437 9867 4471
rect 9901 4437 9919 4471
rect 9585 4369 9919 4437
rect 9953 4511 10103 4573
rect 9953 4477 9971 4511
rect 10005 4477 10046 4511
rect 10080 4477 10103 4511
rect 9953 4443 10103 4477
rect 9953 4409 9971 4443
rect 10005 4409 10046 4443
rect 10080 4409 10103 4443
rect 9953 4403 10103 4409
rect 10137 4593 10157 4627
rect 10191 4593 10287 4627
rect 10137 4523 10287 4593
rect 10321 4591 10471 4661
rect 10542 4701 10620 4720
rect 10717 4719 10733 4753
rect 10767 4719 10783 4753
rect 10817 4837 10924 4845
rect 10817 4803 10833 4837
rect 10867 4803 10924 4837
rect 10817 4769 10924 4803
rect 10817 4735 10833 4769
rect 10867 4735 10924 4769
rect 10817 4721 10924 4735
rect 10542 4667 10564 4701
rect 10598 4685 10620 4701
rect 10598 4667 10827 4685
rect 10542 4651 10827 4667
rect 10321 4557 10417 4591
rect 10451 4557 10471 4591
rect 10517 4607 10588 4617
rect 10551 4601 10588 4607
rect 10551 4573 10554 4601
rect 10517 4567 10554 4573
rect 10137 4471 10471 4523
rect 10517 4505 10588 4567
rect 10622 4471 10656 4651
rect 10690 4601 10743 4617
rect 10724 4567 10743 4601
rect 10690 4539 10743 4567
rect 10793 4601 10827 4651
rect 10793 4551 10827 4567
rect 10690 4505 10701 4539
rect 10735 4505 10743 4539
rect 10861 4517 10924 4721
rect 10965 4837 11299 4879
rect 10965 4803 10983 4837
rect 11017 4803 11247 4837
rect 11281 4803 11299 4837
rect 10965 4735 11299 4803
rect 10965 4701 10983 4735
rect 11017 4701 11247 4735
rect 11281 4701 11299 4735
rect 10965 4661 11299 4701
rect 10801 4515 10924 4517
rect 10801 4481 10817 4515
rect 10851 4481 10924 4515
rect 10801 4471 10924 4481
rect 10137 4437 10155 4471
rect 10189 4437 10419 4471
rect 10453 4437 10471 4471
rect 10137 4369 10471 4437
rect 10538 4455 10586 4471
rect 10538 4421 10552 4455
rect 10538 4369 10586 4421
rect 10622 4455 10678 4471
rect 10622 4421 10636 4455
rect 10670 4421 10678 4455
rect 10622 4405 10678 4421
rect 10724 4455 10767 4471
rect 10724 4421 10732 4455
rect 10766 4421 10767 4455
rect 10724 4369 10767 4421
rect 10801 4447 10885 4471
rect 10801 4413 10817 4447
rect 10851 4437 10885 4447
rect 10919 4437 10924 4471
rect 10851 4413 10924 4437
rect 10801 4403 10924 4413
rect 10965 4593 10985 4627
rect 11019 4593 11115 4627
rect 10965 4523 11115 4593
rect 11149 4591 11299 4661
rect 11351 4829 11385 4845
rect 11351 4761 11385 4795
rect 11421 4829 11487 4879
rect 11421 4795 11437 4829
rect 11471 4795 11487 4829
rect 11421 4761 11487 4795
rect 11421 4727 11437 4761
rect 11471 4727 11487 4761
rect 11521 4829 11575 4845
rect 11521 4795 11523 4829
rect 11557 4795 11575 4829
rect 11521 4748 11575 4795
rect 11351 4693 11385 4727
rect 11521 4714 11523 4748
rect 11557 4743 11575 4748
rect 11521 4709 11529 4714
rect 11563 4709 11575 4743
rect 11351 4659 11484 4693
rect 11521 4664 11575 4709
rect 11450 4630 11484 4659
rect 11149 4557 11245 4591
rect 11279 4557 11299 4591
rect 11337 4607 11403 4623
rect 11337 4573 11345 4607
rect 11379 4601 11403 4607
rect 11337 4567 11353 4573
rect 11387 4567 11403 4601
rect 11337 4549 11403 4567
rect 11450 4614 11507 4630
rect 11450 4580 11473 4614
rect 11450 4564 11507 4580
rect 10965 4471 11299 4523
rect 11450 4513 11484 4564
rect 10965 4437 10983 4471
rect 11017 4437 11247 4471
rect 11281 4437 11299 4471
rect 10965 4369 11299 4437
rect 11351 4479 11484 4513
rect 11541 4504 11575 4664
rect 11609 4837 11943 4879
rect 11609 4803 11627 4837
rect 11661 4803 11891 4837
rect 11925 4803 11943 4837
rect 11609 4735 11943 4803
rect 11609 4701 11627 4735
rect 11661 4701 11891 4735
rect 11925 4701 11943 4735
rect 11609 4661 11943 4701
rect 11351 4458 11385 4479
rect 11523 4475 11575 4504
rect 11351 4403 11385 4424
rect 11421 4411 11437 4445
rect 11471 4411 11487 4445
rect 11421 4369 11487 4411
rect 11557 4441 11575 4475
rect 11523 4403 11575 4441
rect 11609 4593 11629 4627
rect 11663 4593 11759 4627
rect 11609 4523 11759 4593
rect 11793 4591 11943 4661
rect 11793 4557 11889 4591
rect 11923 4557 11943 4591
rect 11977 4777 12080 4809
rect 11977 4743 12041 4777
rect 12075 4743 12080 4777
rect 11977 4727 12080 4743
rect 12127 4777 12161 4879
rect 12127 4727 12161 4743
rect 12195 4811 12601 4845
rect 11977 4565 12045 4727
rect 12195 4678 12229 4811
rect 12308 4743 12324 4777
rect 12358 4743 12399 4777
rect 12433 4743 12533 4777
rect 12079 4675 12095 4678
rect 12079 4641 12081 4675
rect 12129 4644 12229 4678
rect 12115 4641 12229 4644
rect 12079 4640 12229 4641
rect 12263 4678 12465 4709
rect 12297 4675 12465 4678
rect 12263 4641 12265 4644
rect 12299 4641 12301 4675
rect 11977 4531 12173 4565
rect 12207 4531 12223 4565
rect 11609 4471 11943 4523
rect 11609 4437 11627 4471
rect 11661 4437 11891 4471
rect 11925 4437 11943 4471
rect 11609 4369 11943 4437
rect 12032 4460 12081 4531
rect 12032 4426 12041 4460
rect 12075 4426 12081 4460
rect 12032 4410 12081 4426
rect 12125 4460 12227 4476
rect 12159 4426 12193 4460
rect 12125 4369 12227 4426
rect 12263 4403 12301 4641
rect 12335 4565 12390 4635
rect 12369 4531 12390 4565
rect 12335 4471 12390 4531
rect 12431 4565 12465 4675
rect 12431 4515 12465 4531
rect 12499 4517 12533 4743
rect 12567 4617 12601 4811
rect 12635 4837 12669 4879
rect 12635 4769 12669 4803
rect 12635 4701 12669 4735
rect 12635 4651 12669 4667
rect 12703 4837 12770 4845
rect 12703 4803 12719 4837
rect 12753 4811 12770 4837
rect 12703 4777 12725 4803
rect 12759 4777 12770 4811
rect 12703 4769 12770 4777
rect 12703 4735 12719 4769
rect 12753 4735 12770 4769
rect 12703 4701 12770 4735
rect 12703 4667 12719 4701
rect 12753 4667 12770 4701
rect 12703 4651 12770 4667
rect 12805 4837 13139 4879
rect 12805 4803 12823 4837
rect 12857 4803 13087 4837
rect 13121 4803 13139 4837
rect 12805 4735 13139 4803
rect 12805 4701 12823 4735
rect 12857 4701 13087 4735
rect 13121 4701 13139 4735
rect 12805 4661 13139 4701
rect 12567 4601 12606 4617
rect 12567 4567 12572 4601
rect 12567 4551 12606 4567
rect 12651 4601 12702 4617
rect 12651 4567 12668 4601
rect 12651 4551 12702 4567
rect 12651 4517 12685 4551
rect 12736 4517 12770 4651
rect 12499 4483 12685 4517
rect 12499 4476 12534 4483
rect 12335 4437 12357 4471
rect 12428 4460 12534 4476
rect 12335 4403 12390 4437
rect 12462 4426 12534 4460
rect 12719 4464 12770 4517
rect 12428 4403 12534 4426
rect 12619 4445 12685 4449
rect 12619 4411 12635 4445
rect 12669 4411 12685 4445
rect 12619 4369 12685 4411
rect 12753 4430 12770 4464
rect 12719 4403 12770 4430
rect 12805 4593 12825 4627
rect 12859 4593 12955 4627
rect 12805 4523 12955 4593
rect 12989 4591 13139 4661
rect 12989 4557 13085 4591
rect 13119 4557 13139 4591
rect 13173 4829 13227 4845
rect 13173 4795 13191 4829
rect 13225 4795 13227 4829
rect 13173 4748 13227 4795
rect 13173 4714 13191 4748
rect 13225 4714 13227 4748
rect 13261 4829 13327 4879
rect 13261 4795 13277 4829
rect 13311 4795 13327 4829
rect 13261 4761 13327 4795
rect 13261 4727 13277 4761
rect 13311 4727 13327 4761
rect 13363 4829 13397 4845
rect 13363 4761 13397 4795
rect 13173 4664 13227 4714
rect 13363 4693 13397 4727
rect 12805 4471 13139 4523
rect 12805 4437 12823 4471
rect 12857 4437 13087 4471
rect 13121 4437 13139 4471
rect 12805 4369 13139 4437
rect 13173 4504 13207 4664
rect 13264 4659 13397 4693
rect 13449 4837 13967 4879
rect 13449 4803 13467 4837
rect 13501 4803 13915 4837
rect 13949 4803 13967 4837
rect 13449 4735 13967 4803
rect 13449 4701 13467 4735
rect 13501 4701 13915 4735
rect 13949 4701 13967 4735
rect 13449 4661 13967 4701
rect 13264 4630 13298 4659
rect 13241 4614 13298 4630
rect 13275 4580 13298 4614
rect 13241 4564 13298 4580
rect 13264 4513 13298 4564
rect 13345 4607 13411 4623
rect 13345 4601 13369 4607
rect 13345 4567 13361 4601
rect 13403 4573 13411 4607
rect 13395 4567 13411 4573
rect 13345 4549 13411 4567
rect 13449 4593 13527 4627
rect 13561 4593 13637 4627
rect 13671 4593 13691 4627
rect 13449 4523 13691 4593
rect 13725 4591 13967 4661
rect 14001 4808 14059 4879
rect 14001 4774 14013 4808
rect 14047 4774 14059 4808
rect 14093 4837 15162 4879
rect 14093 4803 14111 4837
rect 14145 4803 15111 4837
rect 15145 4803 15162 4837
rect 14093 4792 15162 4803
rect 15409 4821 15475 4879
rect 14001 4715 14059 4774
rect 14001 4681 14013 4715
rect 14047 4681 14059 4715
rect 14001 4646 14059 4681
rect 13725 4557 13745 4591
rect 13779 4557 13855 4591
rect 13889 4557 13967 4591
rect 14410 4627 14478 4644
rect 14410 4593 14427 4627
rect 14461 4593 14478 4627
rect 13173 4475 13225 4504
rect 13264 4479 13397 4513
rect 13173 4471 13191 4475
rect 13173 4437 13185 4471
rect 13363 4458 13397 4479
rect 13219 4437 13225 4441
rect 13173 4403 13225 4437
rect 13261 4411 13277 4445
rect 13311 4411 13327 4445
rect 13261 4369 13327 4411
rect 13363 4403 13397 4424
rect 13449 4464 13967 4523
rect 13449 4430 13467 4464
rect 13501 4430 13915 4464
rect 13949 4430 13967 4464
rect 13449 4369 13967 4430
rect 14001 4497 14059 4514
rect 14001 4463 14013 4497
rect 14047 4463 14059 4497
rect 14410 4478 14478 4593
rect 14774 4591 14844 4792
rect 15409 4787 15425 4821
rect 15459 4787 15475 4821
rect 15409 4753 15475 4787
rect 15234 4701 15312 4720
rect 15409 4719 15425 4753
rect 15459 4719 15475 4753
rect 15509 4837 15616 4845
rect 15509 4803 15525 4837
rect 15559 4803 15616 4837
rect 15509 4769 15616 4803
rect 15509 4735 15525 4769
rect 15559 4735 15616 4769
rect 15509 4721 15616 4735
rect 15234 4667 15256 4701
rect 15290 4685 15312 4701
rect 15290 4667 15519 4685
rect 15234 4651 15519 4667
rect 14774 4557 14791 4591
rect 14825 4557 14844 4591
rect 14774 4542 14844 4557
rect 15209 4607 15280 4617
rect 15243 4601 15280 4607
rect 15243 4573 15246 4601
rect 15209 4567 15246 4573
rect 15209 4505 15280 4567
rect 14001 4369 14059 4463
rect 14093 4464 15162 4478
rect 15314 4471 15348 4651
rect 15382 4601 15435 4617
rect 15416 4567 15435 4601
rect 15382 4539 15435 4567
rect 15485 4601 15519 4651
rect 15485 4551 15519 4567
rect 15382 4505 15393 4539
rect 15427 4505 15435 4539
rect 15553 4539 15616 4721
rect 15657 4837 15991 4879
rect 15657 4803 15675 4837
rect 15709 4803 15939 4837
rect 15973 4803 15991 4837
rect 15657 4735 15991 4803
rect 15657 4701 15675 4735
rect 15709 4701 15939 4735
rect 15973 4701 15991 4735
rect 15657 4661 15991 4701
rect 15553 4517 15577 4539
rect 15493 4515 15577 4517
rect 15493 4481 15509 4515
rect 15543 4505 15577 4515
rect 15611 4505 15616 4539
rect 15543 4481 15616 4505
rect 14093 4430 14111 4464
rect 14145 4430 15111 4464
rect 15145 4430 15162 4464
rect 14093 4369 15162 4430
rect 15230 4455 15278 4471
rect 15230 4421 15244 4455
rect 15230 4369 15278 4421
rect 15314 4455 15370 4471
rect 15314 4421 15328 4455
rect 15362 4421 15370 4455
rect 15314 4405 15370 4421
rect 15416 4455 15459 4471
rect 15416 4421 15424 4455
rect 15458 4421 15459 4455
rect 15416 4369 15459 4421
rect 15493 4447 15616 4481
rect 15493 4413 15509 4447
rect 15543 4413 15616 4447
rect 15493 4403 15616 4413
rect 15657 4593 15677 4627
rect 15711 4593 15807 4627
rect 15657 4523 15807 4593
rect 15841 4591 15991 4661
rect 15841 4557 15937 4591
rect 15971 4557 15991 4591
rect 16025 4829 16079 4845
rect 16025 4795 16043 4829
rect 16077 4795 16079 4829
rect 16025 4748 16079 4795
rect 16025 4714 16043 4748
rect 16077 4714 16079 4748
rect 16113 4829 16179 4879
rect 16113 4795 16129 4829
rect 16163 4795 16179 4829
rect 16113 4761 16179 4795
rect 16113 4727 16129 4761
rect 16163 4727 16179 4761
rect 16215 4829 16249 4845
rect 16215 4761 16249 4795
rect 16025 4664 16079 4714
rect 16215 4693 16249 4727
rect 15657 4471 15991 4523
rect 15657 4437 15675 4471
rect 15709 4437 15939 4471
rect 15973 4437 15991 4471
rect 15657 4369 15991 4437
rect 16025 4504 16059 4664
rect 16116 4659 16249 4693
rect 16301 4837 16635 4879
rect 16301 4803 16319 4837
rect 16353 4803 16583 4837
rect 16617 4803 16635 4837
rect 16301 4735 16635 4803
rect 16301 4701 16319 4735
rect 16353 4701 16583 4735
rect 16617 4701 16635 4735
rect 16301 4661 16635 4701
rect 16116 4630 16150 4659
rect 16093 4614 16150 4630
rect 16127 4580 16150 4614
rect 16093 4564 16150 4580
rect 16116 4513 16150 4564
rect 16197 4607 16263 4623
rect 16197 4601 16221 4607
rect 16197 4567 16213 4601
rect 16255 4573 16263 4607
rect 16247 4567 16263 4573
rect 16197 4549 16263 4567
rect 16301 4593 16321 4627
rect 16355 4593 16451 4627
rect 16301 4523 16451 4593
rect 16485 4591 16635 4661
rect 16485 4557 16581 4591
rect 16615 4557 16635 4591
rect 16669 4829 16723 4845
rect 16669 4795 16687 4829
rect 16721 4795 16723 4829
rect 16669 4748 16723 4795
rect 16669 4714 16687 4748
rect 16721 4714 16723 4748
rect 16757 4829 16823 4879
rect 16757 4795 16773 4829
rect 16807 4795 16823 4829
rect 16757 4761 16823 4795
rect 16757 4727 16773 4761
rect 16807 4727 16823 4761
rect 16859 4829 16893 4845
rect 16859 4761 16893 4795
rect 16945 4837 18014 4879
rect 16945 4803 16963 4837
rect 16997 4803 17963 4837
rect 17997 4803 18014 4837
rect 16945 4792 18014 4803
rect 18049 4837 18567 4879
rect 18049 4803 18067 4837
rect 18101 4803 18515 4837
rect 18549 4803 18567 4837
rect 16669 4664 16723 4714
rect 16859 4693 16893 4727
rect 16025 4475 16077 4504
rect 16116 4479 16249 4513
rect 16025 4471 16043 4475
rect 16025 4437 16037 4471
rect 16215 4458 16249 4479
rect 16071 4437 16077 4441
rect 16025 4403 16077 4437
rect 16113 4411 16129 4445
rect 16163 4411 16179 4445
rect 16113 4369 16179 4411
rect 16215 4403 16249 4424
rect 16301 4471 16635 4523
rect 16301 4437 16319 4471
rect 16353 4437 16583 4471
rect 16617 4437 16635 4471
rect 16301 4369 16635 4437
rect 16669 4504 16703 4664
rect 16760 4659 16893 4693
rect 16760 4630 16794 4659
rect 16737 4614 16794 4630
rect 17262 4627 17330 4644
rect 16771 4580 16794 4614
rect 16737 4564 16794 4580
rect 16760 4513 16794 4564
rect 16841 4607 16907 4623
rect 16841 4601 16865 4607
rect 16841 4567 16857 4601
rect 16899 4573 16907 4607
rect 16891 4567 16907 4573
rect 16841 4549 16907 4567
rect 17262 4593 17279 4627
rect 17313 4593 17330 4627
rect 16669 4475 16721 4504
rect 16760 4479 16893 4513
rect 16669 4471 16687 4475
rect 16669 4437 16681 4471
rect 16859 4458 16893 4479
rect 17262 4478 17330 4593
rect 17626 4591 17696 4792
rect 18049 4735 18567 4803
rect 18049 4701 18067 4735
rect 18101 4701 18515 4735
rect 18549 4701 18567 4735
rect 18049 4661 18567 4701
rect 17626 4557 17643 4591
rect 17677 4557 17696 4591
rect 17626 4542 17696 4557
rect 18049 4593 18127 4627
rect 18161 4593 18237 4627
rect 18271 4593 18291 4627
rect 18049 4523 18291 4593
rect 18325 4591 18567 4661
rect 18325 4557 18345 4591
rect 18379 4557 18455 4591
rect 18489 4557 18567 4591
rect 18601 4837 18843 4879
rect 18601 4803 18619 4837
rect 18653 4803 18791 4837
rect 18825 4803 18843 4837
rect 18601 4742 18843 4803
rect 18601 4708 18619 4742
rect 18653 4708 18791 4742
rect 18825 4708 18843 4742
rect 18601 4661 18843 4708
rect 18601 4587 18705 4661
rect 18601 4553 18651 4587
rect 18685 4553 18705 4587
rect 18739 4593 18759 4627
rect 18793 4593 18843 4627
rect 16715 4437 16721 4441
rect 16669 4403 16721 4437
rect 16757 4411 16773 4445
rect 16807 4411 16823 4445
rect 16757 4369 16823 4411
rect 16859 4403 16893 4424
rect 16945 4464 18014 4478
rect 16945 4430 16963 4464
rect 16997 4430 17963 4464
rect 17997 4430 18014 4464
rect 16945 4369 18014 4430
rect 18049 4464 18567 4523
rect 18739 4519 18843 4593
rect 18049 4430 18067 4464
rect 18101 4430 18515 4464
rect 18549 4430 18567 4464
rect 18049 4369 18567 4430
rect 18601 4466 18843 4519
rect 18601 4432 18619 4466
rect 18653 4432 18791 4466
rect 18825 4432 18843 4466
rect 18601 4369 18843 4432
rect 1104 4335 1133 4369
rect 1167 4335 1225 4369
rect 1259 4335 1317 4369
rect 1351 4335 1409 4369
rect 1443 4335 1501 4369
rect 1535 4335 1593 4369
rect 1627 4335 1685 4369
rect 1719 4335 1777 4369
rect 1811 4335 1869 4369
rect 1903 4335 1961 4369
rect 1995 4335 2053 4369
rect 2087 4335 2145 4369
rect 2179 4335 2237 4369
rect 2271 4335 2329 4369
rect 2363 4335 2421 4369
rect 2455 4335 2513 4369
rect 2547 4335 2605 4369
rect 2639 4335 2697 4369
rect 2731 4335 2789 4369
rect 2823 4335 2881 4369
rect 2915 4335 2973 4369
rect 3007 4335 3065 4369
rect 3099 4335 3157 4369
rect 3191 4335 3249 4369
rect 3283 4335 3341 4369
rect 3375 4335 3433 4369
rect 3467 4335 3525 4369
rect 3559 4335 3617 4369
rect 3651 4335 3709 4369
rect 3743 4335 3801 4369
rect 3835 4335 3893 4369
rect 3927 4335 3985 4369
rect 4019 4335 4077 4369
rect 4111 4335 4169 4369
rect 4203 4335 4261 4369
rect 4295 4335 4353 4369
rect 4387 4335 4445 4369
rect 4479 4335 4537 4369
rect 4571 4335 4629 4369
rect 4663 4335 4721 4369
rect 4755 4335 4813 4369
rect 4847 4335 4905 4369
rect 4939 4335 4997 4369
rect 5031 4335 5089 4369
rect 5123 4335 5181 4369
rect 5215 4335 5273 4369
rect 5307 4335 5365 4369
rect 5399 4335 5457 4369
rect 5491 4335 5549 4369
rect 5583 4335 5641 4369
rect 5675 4335 5733 4369
rect 5767 4335 5825 4369
rect 5859 4335 5917 4369
rect 5951 4335 6009 4369
rect 6043 4335 6101 4369
rect 6135 4335 6193 4369
rect 6227 4335 6285 4369
rect 6319 4335 6377 4369
rect 6411 4335 6469 4369
rect 6503 4335 6561 4369
rect 6595 4335 6653 4369
rect 6687 4335 6745 4369
rect 6779 4335 6837 4369
rect 6871 4335 6929 4369
rect 6963 4335 7021 4369
rect 7055 4335 7113 4369
rect 7147 4335 7205 4369
rect 7239 4335 7297 4369
rect 7331 4335 7389 4369
rect 7423 4335 7481 4369
rect 7515 4335 7573 4369
rect 7607 4335 7665 4369
rect 7699 4335 7757 4369
rect 7791 4335 7849 4369
rect 7883 4335 7941 4369
rect 7975 4335 8033 4369
rect 8067 4335 8125 4369
rect 8159 4335 8217 4369
rect 8251 4335 8309 4369
rect 8343 4335 8401 4369
rect 8435 4335 8493 4369
rect 8527 4335 8585 4369
rect 8619 4335 8677 4369
rect 8711 4335 8769 4369
rect 8803 4335 8861 4369
rect 8895 4335 8953 4369
rect 8987 4335 9045 4369
rect 9079 4335 9137 4369
rect 9171 4335 9229 4369
rect 9263 4335 9321 4369
rect 9355 4335 9413 4369
rect 9447 4335 9505 4369
rect 9539 4335 9597 4369
rect 9631 4335 9689 4369
rect 9723 4335 9781 4369
rect 9815 4335 9873 4369
rect 9907 4335 9965 4369
rect 9999 4335 10057 4369
rect 10091 4335 10149 4369
rect 10183 4335 10241 4369
rect 10275 4335 10333 4369
rect 10367 4335 10425 4369
rect 10459 4335 10517 4369
rect 10551 4335 10609 4369
rect 10643 4335 10701 4369
rect 10735 4335 10793 4369
rect 10827 4335 10885 4369
rect 10919 4335 10977 4369
rect 11011 4335 11069 4369
rect 11103 4335 11161 4369
rect 11195 4335 11253 4369
rect 11287 4335 11345 4369
rect 11379 4335 11437 4369
rect 11471 4335 11529 4369
rect 11563 4335 11621 4369
rect 11655 4335 11713 4369
rect 11747 4335 11805 4369
rect 11839 4335 11897 4369
rect 11931 4335 11989 4369
rect 12023 4335 12081 4369
rect 12115 4335 12173 4369
rect 12207 4335 12265 4369
rect 12299 4335 12357 4369
rect 12391 4335 12449 4369
rect 12483 4335 12541 4369
rect 12575 4335 12633 4369
rect 12667 4335 12725 4369
rect 12759 4335 12817 4369
rect 12851 4335 12909 4369
rect 12943 4335 13001 4369
rect 13035 4335 13093 4369
rect 13127 4335 13185 4369
rect 13219 4335 13277 4369
rect 13311 4335 13369 4369
rect 13403 4335 13461 4369
rect 13495 4335 13553 4369
rect 13587 4335 13645 4369
rect 13679 4335 13737 4369
rect 13771 4335 13829 4369
rect 13863 4335 13921 4369
rect 13955 4335 14013 4369
rect 14047 4335 14105 4369
rect 14139 4335 14197 4369
rect 14231 4335 14289 4369
rect 14323 4335 14381 4369
rect 14415 4335 14473 4369
rect 14507 4335 14565 4369
rect 14599 4335 14657 4369
rect 14691 4335 14749 4369
rect 14783 4335 14841 4369
rect 14875 4335 14933 4369
rect 14967 4335 15025 4369
rect 15059 4335 15117 4369
rect 15151 4335 15209 4369
rect 15243 4335 15301 4369
rect 15335 4335 15393 4369
rect 15427 4335 15485 4369
rect 15519 4335 15577 4369
rect 15611 4335 15669 4369
rect 15703 4335 15761 4369
rect 15795 4335 15853 4369
rect 15887 4335 15945 4369
rect 15979 4335 16037 4369
rect 16071 4335 16129 4369
rect 16163 4335 16221 4369
rect 16255 4335 16313 4369
rect 16347 4335 16405 4369
rect 16439 4335 16497 4369
rect 16531 4335 16589 4369
rect 16623 4335 16681 4369
rect 16715 4335 16773 4369
rect 16807 4335 16865 4369
rect 16899 4335 16957 4369
rect 16991 4335 17049 4369
rect 17083 4335 17141 4369
rect 17175 4335 17233 4369
rect 17267 4335 17325 4369
rect 17359 4335 17417 4369
rect 17451 4335 17509 4369
rect 17543 4335 17601 4369
rect 17635 4335 17693 4369
rect 17727 4335 17785 4369
rect 17819 4335 17877 4369
rect 17911 4335 17969 4369
rect 18003 4335 18061 4369
rect 18095 4335 18153 4369
rect 18187 4335 18245 4369
rect 18279 4335 18337 4369
rect 18371 4335 18429 4369
rect 18463 4335 18521 4369
rect 18555 4335 18613 4369
rect 18647 4335 18705 4369
rect 18739 4335 18797 4369
rect 18831 4335 18860 4369
rect 1121 4272 1363 4335
rect 1121 4238 1139 4272
rect 1173 4238 1311 4272
rect 1345 4238 1363 4272
rect 1121 4185 1363 4238
rect 1397 4274 2099 4335
rect 1397 4240 1415 4274
rect 1449 4240 2047 4274
rect 2081 4240 2099 4274
rect 1121 4111 1225 4185
rect 1397 4181 2099 4240
rect 2243 4280 2277 4301
rect 2313 4293 2379 4335
rect 2313 4259 2329 4293
rect 2363 4259 2379 4293
rect 2415 4267 2467 4301
rect 2415 4263 2421 4267
rect 2243 4225 2277 4246
rect 2455 4233 2467 4267
rect 2449 4229 2467 4233
rect 2243 4191 2376 4225
rect 2415 4200 2467 4229
rect 1121 4077 1171 4111
rect 1205 4077 1225 4111
rect 1259 4117 1279 4151
rect 1313 4117 1363 4151
rect 1259 4043 1363 4117
rect 1397 4111 1727 4181
rect 1397 4077 1475 4111
rect 1509 4077 1574 4111
rect 1608 4077 1673 4111
rect 1707 4077 1727 4111
rect 1761 4113 1781 4147
rect 1815 4113 1884 4147
rect 1918 4113 1987 4147
rect 2021 4113 2099 4147
rect 1761 4043 2099 4113
rect 2229 4137 2295 4155
rect 2229 4131 2245 4137
rect 2229 4097 2237 4131
rect 2279 4103 2295 4137
rect 2271 4097 2295 4103
rect 2229 4081 2295 4097
rect 2342 4140 2376 4191
rect 2342 4124 2399 4140
rect 2342 4090 2365 4124
rect 2342 4074 2399 4090
rect 2342 4045 2376 4074
rect 1121 3996 1363 4043
rect 1121 3962 1139 3996
rect 1173 3962 1311 3996
rect 1345 3962 1363 3996
rect 1121 3901 1363 3962
rect 1121 3867 1139 3901
rect 1173 3867 1311 3901
rect 1345 3867 1363 3901
rect 1121 3825 1363 3867
rect 1397 4003 2099 4043
rect 1397 3969 1415 4003
rect 1449 3969 2047 4003
rect 2081 3969 2099 4003
rect 1397 3901 2099 3969
rect 1397 3867 1415 3901
rect 1449 3867 2047 3901
rect 2081 3867 2099 3901
rect 1397 3825 2099 3867
rect 2243 4011 2376 4045
rect 2433 4040 2467 4200
rect 2501 4267 2835 4335
rect 2955 4293 3021 4335
rect 2501 4233 2519 4267
rect 2553 4233 2783 4267
rect 2817 4233 2835 4267
rect 2501 4181 2835 4233
rect 2870 4267 2921 4283
rect 2870 4233 2887 4267
rect 2955 4259 2971 4293
rect 3005 4259 3021 4293
rect 3161 4297 3227 4335
rect 3055 4267 3089 4283
rect 2870 4225 2921 4233
rect 3161 4263 3177 4297
rect 3211 4263 3227 4297
rect 3747 4293 3813 4335
rect 2870 4191 3020 4225
rect 2501 4111 2651 4181
rect 2501 4077 2521 4111
rect 2555 4077 2651 4111
rect 2685 4113 2781 4147
rect 2815 4113 2835 4147
rect 2685 4043 2835 4113
rect 2243 3977 2277 4011
rect 2413 3990 2467 4040
rect 2243 3909 2277 3943
rect 2243 3859 2277 3875
rect 2313 3943 2329 3977
rect 2363 3943 2379 3977
rect 2313 3909 2379 3943
rect 2313 3875 2329 3909
rect 2363 3875 2379 3909
rect 2313 3825 2379 3875
rect 2413 3956 2415 3990
rect 2449 3956 2467 3990
rect 2413 3909 2467 3956
rect 2413 3875 2415 3909
rect 2449 3875 2467 3909
rect 2413 3859 2467 3875
rect 2501 4003 2835 4043
rect 2870 4137 2940 4157
rect 2870 4103 2884 4137
rect 2918 4103 2940 4137
rect 2870 4063 2940 4103
rect 2870 4029 2881 4063
rect 2915 4029 2940 4063
rect 2870 4027 2940 4029
rect 2974 4131 3020 4191
rect 3008 4122 3020 4131
rect 2974 4088 2986 4097
rect 2501 3969 2519 4003
rect 2553 3969 2783 4003
rect 2817 3969 2835 4003
rect 2974 3993 3020 4088
rect 2501 3901 2835 3969
rect 2501 3867 2519 3901
rect 2553 3867 2783 3901
rect 2817 3867 2835 3901
rect 2501 3825 2835 3867
rect 2870 3977 3020 3993
rect 2870 3943 2887 3977
rect 2921 3959 3020 3977
rect 3055 3995 3089 4233
rect 3261 4257 3310 4291
rect 3344 4257 3360 4291
rect 3401 4257 3417 4291
rect 3451 4257 3572 4291
rect 3135 4076 3227 4229
rect 3135 4063 3193 4076
rect 3135 4029 3157 4063
rect 3191 4042 3193 4063
rect 3191 4029 3227 4042
rect 3135 4019 3227 4029
rect 2870 3909 2921 3943
rect 2870 3875 2887 3909
rect 2870 3859 2921 3875
rect 2955 3891 2971 3925
rect 3005 3891 3021 3925
rect 2955 3825 3021 3891
rect 3055 3909 3089 3943
rect 3055 3859 3089 3875
rect 3123 3862 3188 4019
rect 3261 3985 3295 4257
rect 3329 4183 3399 4199
rect 3329 4149 3352 4183
rect 3386 4149 3399 4183
rect 3329 4131 3399 4149
rect 3329 4097 3341 4131
rect 3375 4097 3399 4131
rect 3329 4075 3399 4097
rect 3433 4189 3504 4199
rect 3433 4155 3454 4189
rect 3488 4155 3504 4189
rect 3433 4037 3467 4155
rect 3538 4115 3572 4257
rect 3747 4259 3763 4293
rect 3797 4259 3813 4293
rect 3747 4243 3813 4259
rect 3855 4263 3875 4297
rect 3909 4263 3925 4297
rect 3969 4293 4159 4301
rect 3647 4165 3685 4199
rect 3719 4183 3771 4199
rect 3855 4185 3907 4263
rect 3969 4259 3985 4293
rect 4019 4259 4159 4293
rect 3969 4245 4159 4259
rect 4193 4297 4231 4335
rect 4193 4263 4197 4297
rect 4528 4293 4589 4335
rect 4193 4247 4231 4263
rect 4265 4277 4479 4293
rect 4265 4259 4415 4277
rect 3613 4149 3709 4165
rect 3743 4149 3771 4183
rect 3805 4135 3839 4151
rect 3374 4021 3467 4037
rect 3408 3995 3467 4021
rect 3408 3987 3433 3995
rect 3261 3951 3340 3985
rect 3374 3961 3433 3987
rect 3374 3959 3467 3961
rect 3501 4101 3805 4115
rect 3501 4081 3839 4101
rect 3306 3925 3340 3951
rect 3501 3925 3535 4081
rect 3873 4047 3907 4185
rect 3607 4013 3623 4047
rect 3657 4013 3907 4047
rect 3945 4195 3987 4211
rect 3945 4161 3953 4195
rect 3945 4053 3987 4161
rect 4021 4147 4091 4211
rect 4021 4113 4049 4147
rect 4083 4131 4091 4147
rect 4021 4097 4057 4113
rect 4021 4087 4091 4097
rect 4125 4089 4159 4245
rect 4265 4213 4299 4259
rect 4449 4243 4479 4277
rect 4528 4259 4539 4293
rect 4573 4259 4589 4293
rect 4528 4243 4589 4259
rect 4623 4243 4674 4299
rect 4193 4179 4299 4213
rect 4333 4199 4381 4225
rect 4193 4173 4237 4179
rect 4227 4139 4237 4173
rect 4367 4165 4381 4199
rect 4333 4145 4381 4165
rect 4193 4123 4237 4139
rect 4273 4136 4289 4145
rect 4323 4111 4381 4145
rect 4307 4102 4381 4111
rect 4125 4055 4206 4089
rect 4273 4071 4381 4102
rect 4415 4188 4479 4243
rect 4657 4209 4674 4243
rect 4623 4193 4674 4209
rect 4415 4153 4480 4188
rect 4415 4137 4598 4153
rect 4415 4103 4564 4137
rect 4415 4093 4598 4103
rect 4450 4087 4598 4093
rect 3945 4021 4080 4053
rect 4172 4037 4206 4055
rect 3945 4019 4088 4021
rect 3873 3985 3907 4013
rect 4046 3995 4088 4019
rect 3222 3901 3272 3917
rect 3222 3867 3238 3901
rect 3222 3825 3272 3867
rect 3306 3909 3356 3925
rect 3306 3875 3322 3909
rect 3306 3859 3356 3875
rect 3399 3903 3535 3925
rect 3399 3869 3415 3903
rect 3449 3869 3535 3903
rect 3569 3945 3784 3979
rect 3873 3951 3985 3985
rect 4046 3961 4057 3995
rect 4122 3987 4138 4021
rect 4091 3961 4138 3987
rect 4172 4003 4366 4037
rect 4400 4003 4416 4037
rect 3569 3927 3603 3945
rect 3750 3927 3784 3945
rect 3569 3877 3603 3893
rect 3650 3877 3666 3911
rect 3700 3877 3716 3911
rect 3750 3877 3784 3893
rect 3843 3901 3917 3917
rect 3399 3859 3535 3869
rect 3650 3825 3716 3877
rect 3843 3867 3863 3901
rect 3897 3867 3917 3901
rect 3843 3825 3917 3867
rect 3951 3909 3985 3951
rect 4172 3927 4206 4003
rect 4450 3969 4484 4087
rect 4632 4063 4674 4193
rect 4709 4267 5043 4335
rect 4709 4233 4727 4267
rect 4761 4233 4991 4267
rect 5025 4233 5043 4267
rect 4709 4181 5043 4233
rect 5113 4305 5181 4335
rect 5113 4271 5131 4305
rect 5165 4271 5181 4305
rect 5113 4237 5181 4271
rect 5113 4203 5131 4237
rect 5165 4203 5181 4237
rect 5215 4267 5231 4301
rect 5265 4267 5319 4301
rect 5215 4233 5319 4267
rect 5215 4199 5231 4233
rect 5265 4199 5319 4233
rect 4709 4111 4859 4181
rect 4709 4077 4729 4111
rect 4763 4077 4859 4111
rect 4893 4113 4989 4147
rect 5023 4113 5043 4147
rect 3951 3859 3985 3875
rect 4032 3902 4206 3927
rect 4324 3935 4484 3969
rect 4528 3969 4589 4053
rect 4528 3935 4539 3969
rect 4573 3935 4589 3969
rect 4324 3927 4358 3935
rect 4032 3868 4048 3902
rect 4082 3868 4206 3902
rect 4032 3859 4206 3868
rect 4240 3901 4290 3917
rect 4274 3867 4290 3901
rect 4528 3901 4589 3935
rect 4324 3877 4358 3893
rect 4240 3825 4290 3867
rect 4394 3867 4410 3901
rect 4444 3867 4460 3901
rect 4394 3825 4460 3867
rect 4528 3867 4539 3901
rect 4573 3867 4589 3901
rect 4623 4005 4674 4063
rect 4893 4043 5043 4113
rect 4657 3971 4674 4005
rect 4623 3937 4674 3971
rect 4657 3927 4674 3937
rect 4623 3893 4629 3903
rect 4663 3893 4674 3927
rect 4623 3887 4674 3893
rect 4709 4003 5043 4043
rect 4709 3969 4727 4003
rect 4761 3969 4991 4003
rect 5025 3969 5043 4003
rect 4709 3901 5043 3969
rect 4528 3825 4589 3867
rect 4709 3867 4727 3901
rect 4761 3867 4991 3901
rect 5025 3867 5043 3901
rect 4709 3825 5043 3867
rect 5077 3995 5181 4169
rect 5215 4004 5319 4199
rect 5353 4274 6055 4335
rect 5353 4240 5371 4274
rect 5405 4240 6003 4274
rect 6037 4240 6055 4274
rect 5353 4181 6055 4240
rect 6273 4241 6331 4335
rect 6273 4207 6285 4241
rect 6319 4207 6331 4241
rect 6273 4190 6331 4207
rect 6365 4272 6607 4335
rect 6365 4238 6383 4272
rect 6417 4238 6555 4272
rect 6589 4238 6607 4272
rect 6365 4185 6607 4238
rect 6641 4263 6693 4301
rect 6641 4229 6659 4263
rect 6729 4293 6795 4335
rect 6729 4259 6745 4293
rect 6779 4259 6795 4293
rect 6831 4280 6865 4301
rect 6641 4200 6693 4229
rect 6831 4225 6865 4246
rect 5353 4111 5683 4181
rect 5353 4077 5431 4111
rect 5465 4077 5530 4111
rect 5564 4077 5629 4111
rect 5663 4077 5683 4111
rect 5717 4113 5737 4147
rect 5771 4113 5840 4147
rect 5874 4113 5943 4147
rect 5977 4113 6055 4147
rect 5717 4043 6055 4113
rect 6365 4111 6469 4185
rect 6365 4077 6415 4111
rect 6449 4077 6469 4111
rect 6503 4117 6523 4151
rect 6557 4117 6607 4151
rect 5077 3961 5089 3995
rect 5123 3970 5181 3995
rect 5353 4003 6055 4043
rect 5123 3961 5131 3970
rect 5077 3936 5131 3961
rect 5165 3936 5181 3970
rect 5077 3902 5181 3936
rect 5077 3868 5131 3902
rect 5165 3868 5181 3902
rect 5077 3859 5181 3868
rect 5215 3936 5231 3970
rect 5265 3936 5281 3970
rect 5215 3902 5281 3936
rect 5215 3868 5231 3902
rect 5265 3868 5281 3902
rect 5215 3825 5281 3868
rect 5353 3969 5371 4003
rect 5405 3969 6003 4003
rect 6037 3969 6055 4003
rect 5353 3901 6055 3969
rect 5353 3867 5371 3901
rect 5405 3867 6003 3901
rect 6037 3867 6055 3901
rect 5353 3825 6055 3867
rect 6273 4023 6331 4058
rect 6503 4043 6607 4117
rect 6273 3989 6285 4023
rect 6319 3989 6331 4023
rect 6273 3930 6331 3989
rect 6273 3896 6285 3930
rect 6319 3896 6331 3930
rect 6273 3825 6331 3896
rect 6365 3996 6607 4043
rect 6365 3962 6383 3996
rect 6417 3962 6555 3996
rect 6589 3962 6607 3996
rect 6365 3901 6607 3962
rect 6365 3867 6383 3901
rect 6417 3867 6555 3901
rect 6589 3867 6607 3901
rect 6365 3825 6607 3867
rect 6641 4040 6675 4200
rect 6732 4191 6865 4225
rect 6917 4274 7619 4335
rect 6917 4240 6935 4274
rect 6969 4240 7567 4274
rect 7601 4240 7619 4274
rect 6732 4140 6766 4191
rect 6917 4181 7619 4240
rect 7708 4278 7757 4294
rect 7708 4244 7717 4278
rect 7751 4244 7757 4278
rect 6709 4124 6766 4140
rect 6743 4090 6766 4124
rect 6709 4074 6766 4090
rect 6813 4137 6879 4155
rect 6813 4103 6829 4137
rect 6863 4131 6879 4137
rect 6813 4097 6837 4103
rect 6871 4097 6879 4131
rect 6813 4081 6879 4097
rect 6917 4111 7247 4181
rect 7708 4173 7757 4244
rect 7801 4278 7903 4335
rect 7835 4244 7869 4278
rect 7801 4228 7903 4244
rect 6917 4077 6995 4111
rect 7029 4077 7094 4111
rect 7128 4077 7193 4111
rect 7227 4077 7247 4111
rect 7281 4113 7301 4147
rect 7335 4113 7404 4147
rect 7438 4113 7507 4147
rect 7541 4113 7619 4147
rect 6732 4045 6766 4074
rect 6641 3995 6695 4040
rect 6732 4011 6865 4045
rect 7281 4043 7619 4113
rect 6641 3961 6653 3995
rect 6687 3990 6695 3995
rect 6641 3956 6659 3961
rect 6693 3956 6695 3990
rect 6831 3977 6865 4011
rect 6641 3909 6695 3956
rect 6641 3875 6659 3909
rect 6693 3875 6695 3909
rect 6641 3859 6695 3875
rect 6729 3943 6745 3977
rect 6779 3943 6795 3977
rect 6729 3909 6795 3943
rect 6729 3875 6745 3909
rect 6779 3875 6795 3909
rect 6729 3825 6795 3875
rect 6831 3909 6865 3943
rect 6831 3859 6865 3875
rect 6917 4003 7619 4043
rect 6917 3969 6935 4003
rect 6969 3969 7567 4003
rect 7601 3969 7619 4003
rect 6917 3901 7619 3969
rect 6917 3867 6935 3901
rect 6969 3867 7567 3901
rect 7601 3867 7619 3901
rect 7653 4139 7849 4173
rect 7883 4139 7899 4173
rect 7653 3977 7721 4139
rect 7755 4063 7905 4064
rect 7755 4029 7757 4063
rect 7791 4060 7905 4063
rect 7755 4026 7771 4029
rect 7805 4026 7905 4060
rect 7653 3961 7756 3977
rect 7653 3927 7717 3961
rect 7751 3927 7756 3961
rect 7653 3895 7756 3927
rect 7803 3961 7837 3977
rect 6917 3825 7619 3867
rect 7803 3825 7837 3927
rect 7871 3893 7905 4026
rect 7939 4063 7977 4301
rect 8011 4267 8066 4301
rect 8104 4278 8210 4301
rect 8011 4233 8033 4267
rect 8138 4244 8210 4278
rect 8295 4293 8361 4335
rect 8295 4259 8311 4293
rect 8345 4259 8361 4293
rect 8295 4255 8361 4259
rect 8395 4274 8446 4301
rect 8429 4267 8446 4274
rect 8011 4173 8066 4233
rect 8104 4228 8210 4244
rect 8175 4221 8210 4228
rect 8395 4233 8401 4240
rect 8435 4233 8446 4267
rect 8045 4139 8066 4173
rect 8011 4069 8066 4139
rect 8107 4173 8141 4189
rect 7939 4060 7941 4063
rect 7975 4029 7977 4063
rect 8107 4029 8141 4139
rect 7973 4026 8141 4029
rect 7939 3995 8141 4026
rect 8175 4187 8361 4221
rect 8395 4187 8446 4233
rect 8175 3961 8209 4187
rect 8327 4153 8361 4187
rect 7984 3927 8000 3961
rect 8034 3927 8075 3961
rect 8109 3927 8209 3961
rect 8243 4137 8282 4153
rect 8243 4103 8248 4137
rect 8243 4087 8282 4103
rect 8327 4137 8378 4153
rect 8327 4103 8344 4137
rect 8327 4087 8378 4103
rect 8243 3893 8277 4087
rect 8412 4053 8446 4187
rect 8481 4267 8815 4335
rect 8481 4233 8499 4267
rect 8533 4233 8763 4267
rect 8797 4233 8815 4267
rect 8941 4293 9002 4335
rect 8941 4259 8959 4293
rect 8993 4259 9002 4293
rect 8941 4233 9002 4259
rect 9038 4280 9088 4299
rect 9038 4246 9045 4280
rect 9079 4246 9088 4280
rect 8481 4181 8815 4233
rect 8481 4111 8631 4181
rect 8941 4165 8955 4199
rect 8989 4165 9004 4199
rect 8481 4077 8501 4111
rect 8535 4077 8631 4111
rect 8665 4113 8761 4147
rect 8795 4113 8815 4147
rect 7871 3859 8277 3893
rect 8311 4037 8345 4053
rect 8311 3969 8345 4003
rect 8311 3901 8345 3935
rect 8311 3825 8345 3867
rect 8379 4037 8446 4053
rect 8665 4043 8815 4113
rect 8941 4137 9004 4165
rect 8941 4103 8961 4137
rect 8995 4103 9004 4137
rect 8941 4087 9004 4103
rect 9038 4137 9088 4246
rect 9122 4280 9174 4335
rect 9122 4246 9131 4280
rect 9165 4246 9174 4280
rect 9122 4230 9174 4246
rect 9210 4280 9260 4299
rect 9210 4246 9217 4280
rect 9251 4246 9260 4280
rect 9210 4137 9260 4246
rect 9294 4280 9346 4335
rect 9294 4246 9303 4280
rect 9337 4246 9346 4280
rect 9294 4223 9346 4246
rect 9380 4280 9432 4296
rect 9380 4246 9389 4280
rect 9423 4246 9432 4280
rect 9380 4205 9432 4246
rect 9466 4289 9518 4335
rect 9466 4255 9475 4289
rect 9509 4255 9518 4289
rect 9466 4239 9518 4255
rect 9552 4280 9604 4296
rect 9552 4246 9561 4280
rect 9595 4246 9604 4280
rect 9552 4205 9604 4246
rect 9638 4289 9690 4335
rect 9638 4255 9647 4289
rect 9681 4255 9690 4289
rect 9638 4239 9690 4255
rect 9724 4280 9776 4296
rect 9724 4246 9733 4280
rect 9767 4246 9776 4280
rect 9724 4205 9776 4246
rect 9810 4289 9859 4335
rect 9810 4255 9819 4289
rect 9853 4255 9859 4289
rect 9810 4239 9859 4255
rect 9893 4280 9948 4296
rect 9893 4246 9905 4280
rect 9939 4246 9948 4280
rect 9893 4205 9948 4246
rect 9982 4289 10031 4335
rect 9982 4255 9991 4289
rect 10025 4255 10031 4289
rect 9982 4239 10031 4255
rect 10065 4280 10117 4296
rect 10065 4246 10076 4280
rect 10110 4246 10117 4280
rect 10065 4205 10117 4246
rect 10153 4289 10203 4335
rect 10153 4255 10162 4289
rect 10196 4255 10203 4289
rect 10153 4239 10203 4255
rect 10237 4280 10289 4296
rect 10237 4246 10248 4280
rect 10282 4246 10289 4280
rect 10237 4205 10289 4246
rect 10325 4289 10375 4335
rect 10325 4255 10334 4289
rect 10368 4255 10375 4289
rect 10325 4239 10375 4255
rect 10409 4280 10461 4296
rect 10409 4246 10420 4280
rect 10454 4246 10461 4280
rect 10409 4205 10461 4246
rect 10497 4289 10549 4335
rect 10497 4255 10506 4289
rect 10540 4255 10549 4289
rect 10497 4239 10549 4255
rect 10583 4280 10635 4296
rect 10583 4246 10592 4280
rect 10626 4246 10635 4280
rect 10583 4205 10635 4246
rect 10669 4289 10729 4335
rect 10669 4255 10678 4289
rect 10712 4255 10729 4289
rect 10669 4239 10729 4255
rect 10781 4274 11299 4335
rect 10781 4240 10799 4274
rect 10833 4240 11247 4274
rect 11281 4240 11299 4274
rect 9380 4171 10729 4205
rect 9038 4103 9388 4137
rect 9422 4103 9456 4137
rect 9490 4103 9524 4137
rect 9558 4103 9592 4137
rect 9626 4103 9660 4137
rect 9694 4103 9728 4137
rect 9762 4103 9796 4137
rect 9830 4103 9864 4137
rect 9898 4103 9932 4137
rect 9966 4103 10000 4137
rect 10034 4103 10068 4137
rect 10102 4103 10136 4137
rect 10170 4103 10204 4137
rect 10238 4103 10272 4137
rect 10306 4103 10340 4137
rect 10374 4103 10408 4137
rect 10442 4103 10462 4137
rect 9038 4087 10462 4103
rect 8379 4003 8395 4037
rect 8429 4003 8446 4037
rect 8379 3969 8446 4003
rect 8379 3935 8395 3969
rect 8429 3935 8446 3969
rect 8379 3901 8446 3935
rect 8379 3867 8395 3901
rect 8429 3867 8446 3901
rect 8379 3859 8446 3867
rect 8481 4003 8815 4043
rect 8481 3969 8499 4003
rect 8533 3969 8763 4003
rect 8797 3969 8815 4003
rect 8481 3901 8815 3969
rect 8481 3867 8499 3901
rect 8533 3867 8763 3901
rect 8797 3867 8815 3901
rect 8481 3825 8815 3867
rect 8943 3969 9002 3987
rect 8943 3935 8959 3969
rect 8993 3935 9002 3969
rect 8943 3901 9002 3935
rect 8943 3867 8959 3901
rect 8993 3867 9002 3901
rect 8943 3825 9002 3867
rect 9038 3977 9087 4087
rect 9038 3943 9045 3977
rect 9079 3943 9087 3977
rect 9038 3909 9087 3943
rect 9038 3875 9045 3909
rect 9079 3875 9087 3909
rect 9038 3859 9087 3875
rect 9122 3969 9174 3987
rect 9122 3935 9131 3969
rect 9165 3935 9174 3969
rect 9122 3901 9174 3935
rect 9122 3867 9131 3901
rect 9165 3867 9174 3901
rect 9122 3825 9174 3867
rect 9210 3985 9260 4087
rect 10496 4053 10729 4171
rect 10781 4181 11299 4240
rect 11425 4241 11483 4335
rect 11425 4207 11437 4241
rect 11471 4207 11483 4241
rect 11425 4190 11483 4207
rect 11702 4267 11753 4299
rect 11702 4233 11713 4267
rect 11747 4243 11753 4267
rect 11787 4293 11848 4335
rect 12145 4297 12183 4335
rect 11787 4259 11803 4293
rect 11837 4259 11848 4293
rect 11787 4243 11848 4259
rect 11897 4277 12111 4293
rect 11897 4243 11927 4277
rect 11961 4259 12111 4277
rect 11702 4209 11719 4233
rect 11702 4193 11753 4209
rect 10781 4111 11023 4181
rect 10781 4077 10859 4111
rect 10893 4077 10969 4111
rect 11003 4077 11023 4111
rect 11057 4113 11077 4147
rect 11111 4113 11187 4147
rect 11221 4113 11299 4147
rect 9380 4031 10729 4053
rect 11057 4043 11299 4113
rect 11702 4063 11744 4193
rect 11897 4188 11961 4243
rect 11896 4153 11961 4188
rect 11778 4137 11961 4153
rect 11812 4103 11961 4137
rect 11778 4093 11961 4103
rect 11995 4199 12043 4225
rect 11995 4165 12009 4199
rect 12077 4213 12111 4259
rect 12179 4263 12183 4297
rect 12145 4247 12183 4263
rect 12217 4293 12407 4301
rect 12217 4259 12357 4293
rect 12391 4259 12407 4293
rect 12451 4263 12467 4297
rect 12501 4263 12521 4297
rect 12217 4245 12407 4259
rect 12077 4179 12183 4213
rect 11995 4145 12043 4165
rect 12139 4173 12183 4179
rect 11995 4111 12053 4145
rect 12087 4136 12103 4145
rect 12139 4139 12149 4173
rect 12139 4123 12183 4139
rect 11995 4102 12069 4111
rect 11778 4087 11926 4093
rect 9380 3997 9389 4031
rect 9423 4005 9561 4031
rect 9423 3997 9432 4005
rect 9210 3951 9217 3985
rect 9251 3951 9260 3985
rect 9210 3917 9260 3951
rect 9210 3883 9217 3917
rect 9251 3883 9260 3917
rect 9210 3860 9260 3883
rect 9294 3969 9346 3985
rect 9294 3935 9303 3969
rect 9337 3935 9346 3969
rect 9294 3901 9346 3935
rect 9294 3867 9303 3901
rect 9337 3867 9346 3901
rect 9294 3826 9346 3867
rect 9380 3945 9432 3997
rect 9552 3997 9561 4005
rect 9595 4005 9733 4031
rect 9595 3997 9604 4005
rect 9380 3911 9389 3945
rect 9423 3911 9432 3945
rect 9380 3860 9432 3911
rect 9466 3925 9518 3971
rect 9466 3891 9475 3925
rect 9509 3891 9518 3925
rect 9466 3826 9518 3891
rect 9552 3945 9604 3997
rect 9724 3997 9733 4005
rect 9767 4005 9905 4031
rect 9767 3997 9776 4005
rect 9552 3911 9561 3945
rect 9595 3911 9604 3945
rect 9552 3860 9604 3911
rect 9638 3925 9690 3971
rect 9638 3891 9647 3925
rect 9681 3891 9690 3925
rect 9638 3826 9690 3891
rect 9724 3945 9776 3997
rect 9896 3997 9905 4005
rect 9939 4005 10076 4031
rect 9939 3997 9948 4005
rect 9724 3911 9733 3945
rect 9767 3911 9776 3945
rect 9724 3860 9776 3911
rect 9810 3925 9862 3971
rect 9810 3891 9819 3925
rect 9853 3891 9862 3925
rect 9810 3826 9862 3891
rect 9896 3945 9948 3997
rect 10065 3997 10076 4005
rect 10110 4005 10248 4031
rect 10110 3997 10117 4005
rect 9896 3911 9905 3945
rect 9939 3911 9948 3945
rect 9896 3860 9948 3911
rect 9982 3925 10031 3971
rect 9982 3891 9991 3925
rect 10025 3891 10031 3925
rect 9982 3826 10031 3891
rect 10065 3945 10117 3997
rect 10237 3997 10248 4005
rect 10282 4005 10420 4031
rect 10282 3997 10289 4005
rect 10065 3911 10076 3945
rect 10110 3911 10117 3945
rect 10065 3860 10117 3911
rect 10154 3925 10203 3971
rect 10154 3891 10162 3925
rect 10196 3891 10203 3925
rect 10154 3826 10203 3891
rect 10237 3945 10289 3997
rect 10409 3997 10420 4005
rect 10454 4008 10592 4031
rect 10454 3997 10461 4008
rect 10237 3927 10248 3945
rect 10237 3893 10241 3927
rect 10282 3911 10289 3945
rect 10275 3893 10289 3911
rect 10237 3860 10289 3893
rect 10326 3925 10375 3971
rect 10326 3891 10334 3925
rect 10368 3891 10375 3925
rect 10326 3826 10375 3891
rect 10409 3945 10461 3997
rect 10583 3997 10592 4008
rect 10626 4008 10729 4031
rect 10626 3997 10641 4008
rect 10409 3911 10420 3945
rect 10454 3911 10461 3945
rect 10409 3860 10461 3911
rect 10498 3925 10549 3971
rect 10498 3891 10506 3925
rect 10540 3891 10549 3925
rect 10498 3826 10549 3891
rect 10583 3945 10641 3997
rect 10781 4003 11299 4043
rect 10583 3911 10592 3945
rect 10626 3911 10641 3945
rect 10583 3860 10641 3911
rect 10675 3925 10729 3974
rect 10675 3891 10678 3925
rect 10712 3891 10729 3925
rect 9294 3825 10549 3826
rect 10675 3825 10729 3891
rect 10781 3969 10799 4003
rect 10833 3969 11247 4003
rect 11281 3969 11299 4003
rect 10781 3901 11299 3969
rect 10781 3867 10799 3901
rect 10833 3867 11247 3901
rect 11281 3867 11299 3901
rect 10781 3825 11299 3867
rect 11425 4023 11483 4058
rect 11425 3989 11437 4023
rect 11471 3989 11483 4023
rect 11425 3930 11483 3989
rect 11425 3896 11437 3930
rect 11471 3896 11483 3930
rect 11425 3825 11483 3896
rect 11702 4005 11753 4063
rect 11702 3971 11719 4005
rect 11702 3937 11753 3971
rect 11702 3903 11719 3937
rect 11702 3887 11753 3903
rect 11787 3969 11848 4053
rect 11787 3935 11803 3969
rect 11837 3935 11848 3969
rect 11892 3969 11926 4087
rect 11995 4071 12103 4102
rect 12217 4089 12251 4245
rect 12170 4055 12251 4089
rect 12285 4147 12355 4211
rect 12285 4131 12293 4147
rect 12327 4113 12355 4147
rect 12319 4097 12355 4113
rect 12285 4087 12355 4097
rect 12389 4195 12431 4211
rect 12423 4161 12431 4195
rect 12170 4037 12204 4055
rect 12389 4053 12431 4161
rect 11960 4003 11976 4037
rect 12010 4003 12204 4037
rect 12296 4021 12431 4053
rect 11892 3935 12052 3969
rect 11787 3901 11848 3935
rect 12018 3927 12052 3935
rect 11787 3867 11803 3901
rect 11837 3867 11848 3901
rect 11787 3825 11848 3867
rect 11916 3867 11932 3901
rect 11966 3867 11982 3901
rect 12170 3927 12204 4003
rect 12238 3987 12254 4021
rect 12288 4019 12431 4021
rect 12469 4185 12521 4263
rect 12563 4293 12629 4335
rect 12563 4259 12579 4293
rect 12613 4259 12629 4293
rect 13149 4297 13215 4335
rect 12563 4243 12629 4259
rect 12804 4257 12925 4291
rect 12959 4257 12975 4291
rect 13016 4257 13032 4291
rect 13066 4257 13115 4291
rect 13149 4263 13165 4297
rect 13199 4263 13215 4297
rect 13355 4293 13421 4335
rect 13287 4267 13321 4283
rect 12469 4047 12503 4185
rect 12605 4183 12657 4199
rect 12537 4135 12571 4151
rect 12605 4149 12633 4183
rect 12691 4165 12729 4199
rect 12667 4149 12763 4165
rect 12804 4115 12838 4257
rect 12872 4189 12943 4199
rect 12872 4155 12888 4189
rect 12922 4155 12943 4189
rect 12571 4101 12875 4115
rect 12537 4081 12875 4101
rect 12288 3995 12330 4019
rect 12238 3961 12285 3987
rect 12319 3961 12330 3995
rect 12469 4013 12719 4047
rect 12753 4013 12769 4047
rect 12469 3985 12503 4013
rect 12391 3951 12503 3985
rect 12018 3877 12052 3893
rect 12086 3901 12136 3917
rect 11916 3825 11982 3867
rect 12086 3867 12102 3901
rect 12086 3825 12136 3867
rect 12170 3902 12344 3927
rect 12170 3868 12294 3902
rect 12328 3868 12344 3902
rect 12170 3859 12344 3868
rect 12391 3909 12425 3951
rect 12592 3945 12807 3979
rect 12592 3927 12626 3945
rect 12391 3859 12425 3875
rect 12459 3901 12533 3917
rect 12459 3867 12479 3901
rect 12513 3867 12533 3901
rect 12773 3927 12807 3945
rect 12592 3877 12626 3893
rect 12660 3877 12676 3911
rect 12710 3877 12726 3911
rect 12773 3877 12807 3893
rect 12841 3925 12875 4081
rect 12909 4037 12943 4155
rect 12977 4183 13047 4199
rect 12977 4149 12990 4183
rect 13024 4149 13047 4183
rect 12977 4131 13047 4149
rect 12977 4097 13001 4131
rect 13035 4097 13047 4131
rect 12977 4075 13047 4097
rect 12909 4021 13002 4037
rect 12909 3995 12968 4021
rect 12943 3987 12968 3995
rect 12943 3961 13002 3987
rect 13081 3985 13115 4257
rect 13355 4259 13371 4293
rect 13405 4259 13421 4293
rect 13455 4267 13506 4283
rect 13149 4076 13241 4229
rect 13183 4063 13241 4076
rect 13183 4042 13185 4063
rect 13149 4029 13185 4042
rect 13219 4029 13241 4063
rect 13149 4019 13241 4029
rect 12909 3959 13002 3961
rect 13036 3951 13115 3985
rect 13036 3925 13070 3951
rect 12841 3903 12977 3925
rect 12459 3825 12533 3867
rect 12660 3825 12726 3877
rect 12841 3869 12927 3903
rect 12961 3869 12977 3903
rect 12841 3859 12977 3869
rect 13020 3909 13070 3925
rect 13054 3875 13070 3909
rect 13020 3859 13070 3875
rect 13104 3901 13154 3917
rect 13138 3867 13154 3901
rect 13104 3825 13154 3867
rect 13188 3862 13253 4019
rect 13287 3995 13321 4233
rect 13489 4233 13506 4267
rect 13455 4225 13506 4233
rect 13356 4191 13506 4225
rect 13541 4267 13875 4335
rect 13995 4293 14061 4335
rect 13541 4233 13559 4267
rect 13593 4233 13823 4267
rect 13857 4233 13875 4267
rect 13356 4131 13402 4191
rect 13541 4181 13875 4233
rect 13910 4267 13961 4283
rect 13910 4233 13927 4267
rect 13995 4259 14011 4293
rect 14045 4259 14061 4293
rect 14201 4297 14267 4335
rect 14095 4267 14129 4283
rect 13910 4225 13961 4233
rect 14201 4263 14217 4297
rect 14251 4263 14267 4297
rect 14787 4293 14853 4335
rect 13910 4191 14060 4225
rect 13356 4122 13368 4131
rect 13390 4088 13402 4097
rect 13356 3993 13402 4088
rect 13436 4137 13506 4157
rect 13436 4103 13458 4137
rect 13492 4103 13506 4137
rect 13436 4063 13506 4103
rect 13541 4111 13691 4181
rect 13541 4077 13561 4111
rect 13595 4077 13691 4111
rect 13725 4113 13821 4147
rect 13855 4113 13875 4147
rect 13436 4029 13461 4063
rect 13495 4029 13506 4063
rect 13725 4043 13875 4113
rect 13436 4027 13506 4029
rect 13541 4003 13875 4043
rect 13910 4137 13980 4157
rect 13910 4103 13924 4137
rect 13958 4103 13980 4137
rect 13910 4063 13980 4103
rect 13910 4029 13921 4063
rect 13955 4029 13980 4063
rect 13910 4027 13980 4029
rect 14014 4131 14060 4191
rect 14048 4122 14060 4131
rect 14014 4088 14026 4097
rect 13356 3977 13506 3993
rect 13356 3959 13455 3977
rect 13287 3909 13321 3943
rect 13489 3943 13506 3977
rect 13287 3859 13321 3875
rect 13355 3891 13371 3925
rect 13405 3891 13421 3925
rect 13355 3825 13421 3891
rect 13455 3909 13506 3943
rect 13489 3875 13506 3909
rect 13455 3859 13506 3875
rect 13541 3969 13559 4003
rect 13593 3969 13823 4003
rect 13857 3969 13875 4003
rect 14014 3993 14060 4088
rect 13541 3901 13875 3969
rect 13541 3867 13559 3901
rect 13593 3867 13823 3901
rect 13857 3867 13875 3901
rect 13541 3825 13875 3867
rect 13910 3977 14060 3993
rect 13910 3943 13927 3977
rect 13961 3959 14060 3977
rect 14095 3995 14129 4233
rect 14301 4257 14350 4291
rect 14384 4257 14400 4291
rect 14441 4257 14457 4291
rect 14491 4257 14612 4291
rect 14175 4076 14267 4229
rect 14175 4063 14233 4076
rect 14175 4029 14197 4063
rect 14231 4042 14233 4063
rect 14231 4029 14267 4042
rect 14175 4019 14267 4029
rect 13910 3909 13961 3943
rect 13910 3875 13927 3909
rect 13910 3859 13961 3875
rect 13995 3891 14011 3925
rect 14045 3891 14061 3925
rect 13995 3825 14061 3891
rect 14095 3909 14129 3943
rect 14095 3859 14129 3875
rect 14163 3862 14228 4019
rect 14301 3985 14335 4257
rect 14369 4183 14439 4199
rect 14369 4149 14392 4183
rect 14426 4149 14439 4183
rect 14369 4131 14439 4149
rect 14369 4097 14381 4131
rect 14415 4097 14439 4131
rect 14369 4075 14439 4097
rect 14473 4189 14544 4199
rect 14473 4155 14494 4189
rect 14528 4155 14544 4189
rect 14473 4037 14507 4155
rect 14578 4115 14612 4257
rect 14787 4259 14803 4293
rect 14837 4259 14853 4293
rect 14787 4243 14853 4259
rect 14895 4263 14915 4297
rect 14949 4263 14965 4297
rect 15009 4293 15199 4301
rect 14687 4165 14725 4199
rect 14759 4183 14811 4199
rect 14895 4185 14947 4263
rect 15009 4259 15025 4293
rect 15059 4259 15199 4293
rect 15009 4245 15199 4259
rect 15233 4297 15271 4335
rect 15233 4263 15237 4297
rect 15568 4293 15629 4335
rect 15233 4247 15271 4263
rect 15305 4277 15519 4293
rect 15305 4259 15455 4277
rect 14653 4149 14749 4165
rect 14783 4149 14811 4183
rect 14845 4135 14879 4151
rect 14414 4021 14507 4037
rect 14448 3995 14507 4021
rect 14448 3987 14473 3995
rect 14301 3951 14380 3985
rect 14414 3961 14473 3987
rect 14414 3959 14507 3961
rect 14541 4101 14845 4115
rect 14541 4081 14879 4101
rect 14346 3925 14380 3951
rect 14541 3925 14575 4081
rect 14913 4047 14947 4185
rect 14647 4013 14663 4047
rect 14697 4013 14947 4047
rect 14985 4195 15027 4211
rect 14985 4161 14993 4195
rect 14985 4053 15027 4161
rect 15061 4147 15131 4211
rect 15061 4113 15089 4147
rect 15123 4131 15131 4147
rect 15061 4097 15097 4113
rect 15061 4087 15131 4097
rect 15165 4089 15199 4245
rect 15305 4213 15339 4259
rect 15489 4243 15519 4277
rect 15568 4259 15579 4293
rect 15613 4259 15629 4293
rect 15568 4243 15629 4259
rect 15663 4243 15714 4299
rect 15233 4179 15339 4213
rect 15373 4199 15421 4225
rect 15233 4173 15277 4179
rect 15267 4139 15277 4173
rect 15407 4165 15421 4199
rect 15373 4145 15421 4165
rect 15233 4123 15277 4139
rect 15313 4136 15329 4145
rect 15363 4111 15421 4145
rect 15347 4102 15421 4111
rect 15165 4055 15246 4089
rect 15313 4071 15421 4102
rect 15455 4188 15519 4243
rect 15697 4209 15714 4243
rect 15663 4193 15714 4209
rect 15455 4153 15520 4188
rect 15455 4137 15638 4153
rect 15455 4103 15604 4137
rect 15455 4093 15638 4103
rect 15490 4087 15638 4093
rect 14985 4021 15120 4053
rect 15212 4037 15246 4055
rect 14985 4019 15128 4021
rect 14913 3985 14947 4013
rect 15086 3995 15128 4019
rect 14262 3901 14312 3917
rect 14262 3867 14278 3901
rect 14262 3825 14312 3867
rect 14346 3909 14396 3925
rect 14346 3875 14362 3909
rect 14346 3859 14396 3875
rect 14439 3903 14575 3925
rect 14439 3869 14455 3903
rect 14489 3869 14575 3903
rect 14609 3945 14824 3979
rect 14913 3951 15025 3985
rect 15086 3961 15097 3995
rect 15162 3987 15178 4021
rect 15131 3961 15178 3987
rect 15212 4003 15406 4037
rect 15440 4003 15456 4037
rect 14609 3927 14643 3945
rect 14790 3927 14824 3945
rect 14609 3877 14643 3893
rect 14690 3877 14706 3911
rect 14740 3877 14756 3911
rect 14790 3877 14824 3893
rect 14883 3901 14957 3917
rect 14439 3859 14575 3869
rect 14690 3825 14756 3877
rect 14883 3867 14903 3901
rect 14937 3867 14957 3901
rect 14883 3825 14957 3867
rect 14991 3909 15025 3951
rect 15212 3927 15246 4003
rect 15490 3969 15524 4087
rect 15672 4063 15714 4193
rect 15749 4274 16451 4335
rect 15749 4240 15767 4274
rect 15801 4240 16399 4274
rect 16433 4240 16451 4274
rect 15749 4181 16451 4240
rect 16577 4241 16635 4335
rect 16577 4207 16589 4241
rect 16623 4207 16635 4241
rect 16669 4274 17738 4335
rect 16669 4240 16687 4274
rect 16721 4240 17687 4274
rect 17721 4240 17738 4274
rect 16669 4226 17738 4240
rect 17773 4274 18475 4335
rect 17773 4240 17791 4274
rect 17825 4240 18423 4274
rect 18457 4240 18475 4274
rect 16577 4190 16635 4207
rect 15749 4111 16079 4181
rect 15749 4077 15827 4111
rect 15861 4077 15926 4111
rect 15960 4077 16025 4111
rect 16059 4077 16079 4111
rect 16113 4113 16133 4147
rect 16167 4113 16236 4147
rect 16270 4113 16339 4147
rect 16373 4113 16451 4147
rect 14991 3859 15025 3875
rect 15072 3902 15246 3927
rect 15364 3935 15524 3969
rect 15568 3969 15629 4053
rect 15568 3935 15579 3969
rect 15613 3935 15629 3969
rect 15364 3927 15398 3935
rect 15072 3868 15088 3902
rect 15122 3868 15246 3902
rect 15072 3859 15246 3868
rect 15280 3901 15330 3917
rect 15314 3867 15330 3901
rect 15568 3901 15629 3935
rect 15364 3877 15398 3893
rect 15280 3825 15330 3867
rect 15434 3867 15450 3901
rect 15484 3867 15500 3901
rect 15434 3825 15500 3867
rect 15568 3867 15579 3901
rect 15613 3867 15629 3901
rect 15663 4005 15714 4063
rect 16113 4043 16451 4113
rect 16986 4111 17054 4226
rect 17773 4181 18475 4240
rect 18601 4272 18843 4335
rect 18601 4238 18619 4272
rect 18653 4238 18791 4272
rect 18825 4238 18843 4272
rect 18601 4185 18843 4238
rect 16986 4077 17003 4111
rect 17037 4077 17054 4111
rect 16986 4060 17054 4077
rect 17350 4147 17420 4162
rect 17350 4113 17367 4147
rect 17401 4113 17420 4147
rect 15697 3971 15714 4005
rect 15663 3937 15714 3971
rect 15697 3927 15714 3937
rect 15663 3893 15669 3903
rect 15703 3893 15714 3927
rect 15663 3887 15714 3893
rect 15749 4003 16451 4043
rect 15749 3969 15767 4003
rect 15801 3969 16399 4003
rect 16433 3969 16451 4003
rect 15749 3901 16451 3969
rect 15568 3825 15629 3867
rect 15749 3867 15767 3901
rect 15801 3867 16399 3901
rect 16433 3867 16451 3901
rect 15749 3825 16451 3867
rect 16577 4023 16635 4058
rect 16577 3989 16589 4023
rect 16623 3989 16635 4023
rect 16577 3930 16635 3989
rect 16577 3896 16589 3930
rect 16623 3896 16635 3930
rect 17350 3912 17420 4113
rect 17773 4111 18103 4181
rect 17773 4077 17851 4111
rect 17885 4077 17950 4111
rect 17984 4077 18049 4111
rect 18083 4077 18103 4111
rect 18137 4113 18157 4147
rect 18191 4113 18260 4147
rect 18294 4113 18363 4147
rect 18397 4113 18475 4147
rect 18137 4043 18475 4113
rect 17773 4003 18475 4043
rect 17773 3969 17791 4003
rect 17825 3969 18423 4003
rect 18457 3969 18475 4003
rect 16577 3825 16635 3896
rect 16669 3901 17738 3912
rect 16669 3867 16687 3901
rect 16721 3867 17687 3901
rect 17721 3867 17738 3901
rect 16669 3825 17738 3867
rect 17773 3901 18475 3969
rect 17773 3867 17791 3901
rect 17825 3867 18423 3901
rect 18457 3867 18475 3901
rect 17773 3825 18475 3867
rect 18601 4117 18651 4151
rect 18685 4117 18705 4151
rect 18601 4043 18705 4117
rect 18739 4111 18843 4185
rect 18739 4077 18759 4111
rect 18793 4077 18843 4111
rect 18601 3996 18843 4043
rect 18601 3962 18619 3996
rect 18653 3962 18791 3996
rect 18825 3962 18843 3996
rect 18601 3901 18843 3962
rect 18601 3867 18619 3901
rect 18653 3867 18791 3901
rect 18825 3867 18843 3901
rect 18601 3825 18843 3867
rect 1104 3791 1133 3825
rect 1167 3791 1225 3825
rect 1259 3791 1317 3825
rect 1351 3791 1409 3825
rect 1443 3791 1501 3825
rect 1535 3791 1593 3825
rect 1627 3791 1685 3825
rect 1719 3791 1777 3825
rect 1811 3791 1869 3825
rect 1903 3791 1961 3825
rect 1995 3791 2053 3825
rect 2087 3791 2145 3825
rect 2179 3791 2237 3825
rect 2271 3791 2329 3825
rect 2363 3791 2421 3825
rect 2455 3791 2513 3825
rect 2547 3791 2605 3825
rect 2639 3791 2697 3825
rect 2731 3791 2789 3825
rect 2823 3791 2881 3825
rect 2915 3791 2973 3825
rect 3007 3791 3065 3825
rect 3099 3791 3157 3825
rect 3191 3791 3249 3825
rect 3283 3791 3341 3825
rect 3375 3791 3433 3825
rect 3467 3791 3525 3825
rect 3559 3791 3617 3825
rect 3651 3791 3709 3825
rect 3743 3791 3801 3825
rect 3835 3791 3893 3825
rect 3927 3791 3985 3825
rect 4019 3791 4077 3825
rect 4111 3791 4169 3825
rect 4203 3791 4261 3825
rect 4295 3791 4353 3825
rect 4387 3791 4445 3825
rect 4479 3791 4537 3825
rect 4571 3791 4629 3825
rect 4663 3791 4721 3825
rect 4755 3791 4813 3825
rect 4847 3791 4905 3825
rect 4939 3791 4997 3825
rect 5031 3791 5089 3825
rect 5123 3791 5181 3825
rect 5215 3791 5273 3825
rect 5307 3791 5365 3825
rect 5399 3791 5457 3825
rect 5491 3791 5549 3825
rect 5583 3791 5641 3825
rect 5675 3791 5733 3825
rect 5767 3791 5825 3825
rect 5859 3791 5917 3825
rect 5951 3791 6009 3825
rect 6043 3791 6101 3825
rect 6135 3791 6193 3825
rect 6227 3791 6285 3825
rect 6319 3791 6377 3825
rect 6411 3791 6469 3825
rect 6503 3791 6561 3825
rect 6595 3791 6653 3825
rect 6687 3791 6745 3825
rect 6779 3791 6837 3825
rect 6871 3791 6929 3825
rect 6963 3791 7021 3825
rect 7055 3791 7113 3825
rect 7147 3791 7205 3825
rect 7239 3791 7297 3825
rect 7331 3791 7389 3825
rect 7423 3791 7481 3825
rect 7515 3791 7573 3825
rect 7607 3791 7665 3825
rect 7699 3791 7757 3825
rect 7791 3791 7849 3825
rect 7883 3791 7941 3825
rect 7975 3791 8033 3825
rect 8067 3791 8125 3825
rect 8159 3791 8217 3825
rect 8251 3791 8309 3825
rect 8343 3791 8401 3825
rect 8435 3791 8493 3825
rect 8527 3791 8585 3825
rect 8619 3791 8677 3825
rect 8711 3791 8769 3825
rect 8803 3791 8861 3825
rect 8895 3791 8953 3825
rect 8987 3791 9045 3825
rect 9079 3791 9137 3825
rect 9171 3791 9229 3825
rect 9263 3791 9321 3825
rect 9355 3791 9413 3825
rect 9447 3791 9505 3825
rect 9539 3791 9597 3825
rect 9631 3791 9689 3825
rect 9723 3791 9781 3825
rect 9815 3791 9873 3825
rect 9907 3791 9965 3825
rect 9999 3791 10057 3825
rect 10091 3791 10149 3825
rect 10183 3791 10241 3825
rect 10275 3791 10333 3825
rect 10367 3791 10425 3825
rect 10459 3791 10517 3825
rect 10551 3791 10609 3825
rect 10643 3791 10701 3825
rect 10735 3791 10793 3825
rect 10827 3791 10885 3825
rect 10919 3791 10977 3825
rect 11011 3791 11069 3825
rect 11103 3791 11161 3825
rect 11195 3791 11253 3825
rect 11287 3791 11345 3825
rect 11379 3791 11437 3825
rect 11471 3791 11529 3825
rect 11563 3791 11621 3825
rect 11655 3791 11713 3825
rect 11747 3791 11805 3825
rect 11839 3791 11897 3825
rect 11931 3791 11989 3825
rect 12023 3791 12081 3825
rect 12115 3791 12173 3825
rect 12207 3791 12265 3825
rect 12299 3791 12357 3825
rect 12391 3791 12449 3825
rect 12483 3791 12541 3825
rect 12575 3791 12633 3825
rect 12667 3791 12725 3825
rect 12759 3791 12817 3825
rect 12851 3791 12909 3825
rect 12943 3791 13001 3825
rect 13035 3791 13093 3825
rect 13127 3791 13185 3825
rect 13219 3791 13277 3825
rect 13311 3791 13369 3825
rect 13403 3791 13461 3825
rect 13495 3791 13553 3825
rect 13587 3791 13645 3825
rect 13679 3791 13737 3825
rect 13771 3791 13829 3825
rect 13863 3791 13921 3825
rect 13955 3791 14013 3825
rect 14047 3791 14105 3825
rect 14139 3791 14197 3825
rect 14231 3791 14289 3825
rect 14323 3791 14381 3825
rect 14415 3791 14473 3825
rect 14507 3791 14565 3825
rect 14599 3791 14657 3825
rect 14691 3791 14749 3825
rect 14783 3791 14841 3825
rect 14875 3791 14933 3825
rect 14967 3791 15025 3825
rect 15059 3791 15117 3825
rect 15151 3791 15209 3825
rect 15243 3791 15301 3825
rect 15335 3791 15393 3825
rect 15427 3791 15485 3825
rect 15519 3791 15577 3825
rect 15611 3791 15669 3825
rect 15703 3791 15761 3825
rect 15795 3791 15853 3825
rect 15887 3791 15945 3825
rect 15979 3791 16037 3825
rect 16071 3791 16129 3825
rect 16163 3791 16221 3825
rect 16255 3791 16313 3825
rect 16347 3791 16405 3825
rect 16439 3791 16497 3825
rect 16531 3791 16589 3825
rect 16623 3791 16681 3825
rect 16715 3791 16773 3825
rect 16807 3791 16865 3825
rect 16899 3791 16957 3825
rect 16991 3791 17049 3825
rect 17083 3791 17141 3825
rect 17175 3791 17233 3825
rect 17267 3791 17325 3825
rect 17359 3791 17417 3825
rect 17451 3791 17509 3825
rect 17543 3791 17601 3825
rect 17635 3791 17693 3825
rect 17727 3791 17785 3825
rect 17819 3791 17877 3825
rect 17911 3791 17969 3825
rect 18003 3791 18061 3825
rect 18095 3791 18153 3825
rect 18187 3791 18245 3825
rect 18279 3791 18337 3825
rect 18371 3791 18429 3825
rect 18463 3791 18521 3825
rect 18555 3791 18613 3825
rect 18647 3791 18705 3825
rect 18739 3791 18797 3825
rect 18831 3791 18860 3825
rect 1121 3749 1363 3791
rect 1121 3715 1139 3749
rect 1173 3715 1311 3749
rect 1345 3715 1363 3749
rect 1121 3654 1363 3715
rect 1121 3620 1139 3654
rect 1173 3620 1311 3654
rect 1345 3620 1363 3654
rect 1121 3573 1363 3620
rect 1397 3749 1639 3791
rect 1397 3715 1415 3749
rect 1449 3715 1587 3749
rect 1621 3715 1639 3749
rect 1397 3654 1639 3715
rect 1397 3620 1415 3654
rect 1449 3620 1587 3654
rect 1621 3620 1639 3654
rect 1674 3741 1725 3757
rect 1674 3707 1691 3741
rect 1674 3673 1725 3707
rect 1759 3725 1825 3791
rect 1759 3691 1775 3725
rect 1809 3691 1825 3725
rect 1859 3741 1893 3757
rect 1674 3639 1691 3673
rect 1859 3673 1893 3707
rect 1725 3639 1824 3657
rect 1674 3623 1824 3639
rect 1397 3573 1639 3620
rect 1121 3505 1171 3539
rect 1205 3505 1225 3539
rect 1121 3431 1225 3505
rect 1259 3499 1363 3573
rect 1259 3465 1279 3499
rect 1313 3465 1363 3499
rect 1397 3505 1447 3539
rect 1481 3505 1501 3539
rect 1397 3431 1501 3505
rect 1535 3499 1639 3573
rect 1535 3465 1555 3499
rect 1589 3465 1639 3499
rect 1674 3587 1744 3589
rect 1674 3553 1685 3587
rect 1719 3553 1744 3587
rect 1674 3513 1744 3553
rect 1674 3479 1688 3513
rect 1722 3479 1744 3513
rect 1674 3459 1744 3479
rect 1778 3528 1824 3623
rect 1778 3519 1790 3528
rect 1812 3485 1824 3494
rect 1121 3378 1363 3431
rect 1121 3344 1139 3378
rect 1173 3344 1311 3378
rect 1345 3344 1363 3378
rect 1121 3281 1363 3344
rect 1397 3378 1639 3431
rect 1778 3425 1824 3485
rect 1397 3344 1415 3378
rect 1449 3344 1587 3378
rect 1621 3344 1639 3378
rect 1397 3281 1639 3344
rect 1674 3391 1824 3425
rect 1674 3383 1725 3391
rect 1674 3349 1691 3383
rect 1859 3383 1893 3621
rect 1927 3723 1992 3754
rect 1927 3689 1948 3723
rect 1982 3689 1992 3723
rect 2026 3749 2076 3791
rect 2026 3715 2042 3749
rect 2026 3699 2076 3715
rect 2110 3741 2160 3757
rect 2110 3707 2126 3741
rect 1927 3597 1992 3689
rect 2110 3691 2160 3707
rect 2203 3747 2339 3757
rect 2203 3713 2219 3747
rect 2253 3713 2339 3747
rect 2454 3739 2520 3791
rect 2647 3749 2721 3791
rect 2203 3691 2339 3713
rect 2110 3665 2144 3691
rect 2065 3631 2144 3665
rect 2178 3655 2271 3657
rect 1939 3574 2031 3597
rect 1939 3540 1997 3574
rect 1939 3387 2031 3540
rect 1674 3333 1725 3349
rect 1759 3323 1775 3357
rect 1809 3323 1825 3357
rect 2065 3359 2099 3631
rect 2178 3629 2237 3655
rect 2212 3621 2237 3629
rect 2212 3595 2271 3621
rect 2178 3579 2271 3595
rect 2133 3519 2203 3541
rect 2133 3485 2145 3519
rect 2179 3485 2203 3519
rect 2133 3467 2203 3485
rect 2133 3433 2156 3467
rect 2190 3433 2203 3467
rect 2133 3417 2203 3433
rect 2237 3461 2271 3579
rect 2305 3535 2339 3691
rect 2373 3723 2407 3739
rect 2454 3705 2470 3739
rect 2504 3705 2520 3739
rect 2554 3723 2588 3739
rect 2373 3671 2407 3689
rect 2647 3715 2667 3749
rect 2701 3715 2721 3749
rect 2647 3699 2721 3715
rect 2755 3741 2789 3757
rect 2554 3671 2588 3689
rect 2373 3637 2588 3671
rect 2755 3665 2789 3707
rect 2836 3748 3010 3757
rect 2836 3714 2852 3748
rect 2886 3714 3010 3748
rect 2836 3689 3010 3714
rect 3044 3749 3094 3791
rect 3078 3715 3094 3749
rect 3198 3749 3264 3791
rect 3044 3699 3094 3715
rect 3128 3723 3162 3739
rect 2677 3631 2789 3665
rect 2677 3603 2711 3631
rect 2411 3569 2427 3603
rect 2461 3569 2711 3603
rect 2850 3621 2861 3655
rect 2895 3629 2942 3655
rect 2850 3597 2892 3621
rect 2305 3515 2643 3535
rect 2305 3501 2609 3515
rect 2237 3427 2258 3461
rect 2292 3427 2308 3461
rect 2237 3417 2308 3427
rect 2342 3359 2376 3501
rect 2417 3451 2513 3467
rect 2451 3417 2489 3451
rect 2547 3433 2575 3467
rect 2609 3465 2643 3481
rect 2523 3417 2575 3433
rect 2677 3431 2711 3569
rect 1859 3333 1893 3349
rect 1759 3281 1825 3323
rect 1965 3319 1981 3353
rect 2015 3319 2031 3353
rect 2065 3325 2114 3359
rect 2148 3325 2164 3359
rect 2205 3325 2221 3359
rect 2255 3325 2376 3359
rect 2551 3357 2617 3373
rect 1965 3281 2031 3319
rect 2551 3323 2567 3357
rect 2601 3323 2617 3357
rect 2551 3281 2617 3323
rect 2659 3353 2711 3431
rect 2749 3595 2892 3597
rect 2926 3595 2942 3629
rect 2976 3613 3010 3689
rect 3198 3715 3214 3749
rect 3248 3715 3264 3749
rect 3332 3749 3393 3791
rect 3332 3715 3343 3749
rect 3377 3715 3393 3749
rect 3128 3681 3162 3689
rect 3332 3681 3393 3715
rect 3128 3647 3288 3681
rect 2749 3563 2884 3595
rect 2976 3579 3170 3613
rect 3204 3579 3220 3613
rect 2749 3455 2791 3563
rect 2976 3561 3010 3579
rect 2749 3421 2757 3455
rect 2749 3405 2791 3421
rect 2825 3519 2895 3529
rect 2825 3503 2861 3519
rect 2825 3469 2853 3503
rect 2887 3469 2895 3485
rect 2825 3405 2895 3469
rect 2929 3527 3010 3561
rect 2929 3371 2963 3527
rect 3077 3514 3185 3545
rect 3254 3529 3288 3647
rect 3332 3647 3343 3681
rect 3377 3647 3393 3681
rect 3332 3563 3393 3647
rect 3427 3713 3478 3729
rect 3461 3679 3478 3713
rect 3427 3645 3478 3679
rect 3461 3611 3478 3645
rect 3427 3553 3478 3611
rect 3697 3720 3755 3791
rect 3697 3686 3709 3720
rect 3743 3686 3755 3720
rect 3697 3627 3755 3686
rect 3697 3593 3709 3627
rect 3743 3593 3755 3627
rect 3697 3558 3755 3593
rect 3789 3749 4491 3791
rect 3789 3715 3807 3749
rect 3841 3715 4439 3749
rect 4473 3715 4491 3749
rect 3789 3647 4491 3715
rect 3789 3613 3807 3647
rect 3841 3613 4439 3647
rect 4473 3613 4491 3647
rect 4543 3725 4597 3791
rect 4723 3790 5978 3791
rect 4543 3691 4560 3725
rect 4594 3691 4597 3725
rect 4543 3642 4597 3691
rect 4631 3705 4689 3756
rect 4631 3671 4646 3705
rect 4680 3671 4689 3705
rect 3789 3573 4491 3613
rect 4631 3619 4689 3671
rect 4723 3725 4774 3790
rect 4723 3691 4732 3725
rect 4766 3691 4774 3725
rect 4723 3645 4774 3691
rect 4811 3705 4863 3756
rect 4811 3671 4818 3705
rect 4852 3671 4863 3705
rect 4631 3608 4646 3619
rect 3254 3523 3402 3529
rect 3111 3505 3185 3514
rect 2997 3477 3041 3493
rect 3031 3443 3041 3477
rect 3077 3471 3093 3480
rect 3127 3471 3185 3505
rect 2997 3437 3041 3443
rect 3137 3451 3185 3471
rect 2997 3403 3103 3437
rect 2773 3357 2963 3371
rect 2659 3319 2679 3353
rect 2713 3319 2729 3353
rect 2773 3323 2789 3357
rect 2823 3323 2963 3357
rect 2773 3315 2963 3323
rect 2997 3353 3035 3369
rect 2997 3319 3001 3353
rect 3069 3357 3103 3403
rect 3171 3417 3185 3451
rect 3137 3391 3185 3417
rect 3219 3513 3402 3523
rect 3219 3479 3368 3513
rect 3219 3463 3402 3479
rect 3219 3428 3284 3463
rect 3219 3373 3283 3428
rect 3436 3423 3478 3553
rect 3789 3505 3867 3539
rect 3901 3505 3966 3539
rect 4000 3505 4065 3539
rect 4099 3505 4119 3539
rect 3789 3435 4119 3505
rect 4153 3503 4491 3573
rect 4153 3469 4173 3503
rect 4207 3469 4276 3503
rect 4310 3469 4379 3503
rect 4413 3469 4491 3503
rect 4543 3585 4646 3608
rect 4680 3608 4689 3619
rect 4811 3619 4863 3671
rect 4897 3725 4946 3790
rect 4897 3691 4904 3725
rect 4938 3691 4946 3725
rect 4897 3645 4946 3691
rect 4983 3723 5035 3756
rect 4983 3705 4997 3723
rect 4983 3671 4990 3705
rect 5031 3689 5035 3723
rect 5024 3671 5035 3689
rect 4811 3608 4818 3619
rect 4680 3585 4818 3608
rect 4852 3611 4863 3619
rect 4983 3619 5035 3671
rect 5069 3725 5118 3790
rect 5069 3691 5076 3725
rect 5110 3691 5118 3725
rect 5069 3645 5118 3691
rect 5155 3705 5207 3756
rect 5155 3671 5162 3705
rect 5196 3671 5207 3705
rect 4983 3611 4990 3619
rect 4852 3585 4990 3611
rect 5024 3611 5035 3619
rect 5155 3619 5207 3671
rect 5241 3725 5290 3790
rect 5241 3691 5247 3725
rect 5281 3691 5290 3725
rect 5241 3645 5290 3691
rect 5324 3705 5376 3756
rect 5324 3671 5333 3705
rect 5367 3671 5376 3705
rect 5155 3611 5162 3619
rect 5024 3585 5162 3611
rect 5196 3611 5207 3619
rect 5324 3619 5376 3671
rect 5410 3725 5462 3790
rect 5410 3691 5419 3725
rect 5453 3691 5462 3725
rect 5410 3645 5462 3691
rect 5496 3705 5548 3756
rect 5496 3671 5505 3705
rect 5539 3671 5548 3705
rect 5324 3611 5333 3619
rect 5196 3585 5333 3611
rect 5367 3611 5376 3619
rect 5496 3619 5548 3671
rect 5582 3725 5634 3790
rect 5582 3691 5591 3725
rect 5625 3691 5634 3725
rect 5582 3645 5634 3691
rect 5668 3705 5720 3756
rect 5668 3671 5677 3705
rect 5711 3671 5720 3705
rect 5496 3611 5505 3619
rect 5367 3585 5505 3611
rect 5539 3611 5548 3619
rect 5668 3619 5720 3671
rect 5754 3725 5806 3790
rect 5754 3691 5763 3725
rect 5797 3691 5806 3725
rect 5754 3645 5806 3691
rect 5840 3705 5892 3756
rect 5840 3671 5849 3705
rect 5883 3671 5892 3705
rect 5668 3611 5677 3619
rect 5539 3585 5677 3611
rect 5711 3611 5720 3619
rect 5840 3619 5892 3671
rect 5926 3749 5978 3790
rect 5926 3715 5935 3749
rect 5969 3715 5978 3749
rect 5926 3681 5978 3715
rect 5926 3647 5935 3681
rect 5969 3647 5978 3681
rect 5926 3631 5978 3647
rect 6012 3733 6062 3756
rect 6012 3699 6021 3733
rect 6055 3699 6062 3733
rect 6012 3665 6062 3699
rect 6012 3631 6021 3665
rect 6055 3631 6062 3665
rect 5840 3611 5849 3619
rect 5711 3585 5849 3611
rect 5883 3585 5892 3619
rect 4543 3563 5892 3585
rect 4543 3445 4776 3563
rect 6012 3529 6062 3631
rect 6098 3749 6150 3791
rect 6098 3715 6107 3749
rect 6141 3715 6150 3749
rect 6098 3681 6150 3715
rect 6098 3647 6107 3681
rect 6141 3647 6150 3681
rect 6098 3629 6150 3647
rect 6185 3741 6234 3757
rect 6185 3707 6193 3741
rect 6227 3707 6234 3741
rect 6185 3673 6234 3707
rect 6185 3639 6193 3673
rect 6227 3639 6234 3673
rect 6185 3529 6234 3639
rect 6270 3749 6329 3791
rect 6270 3715 6279 3749
rect 6313 3715 6329 3749
rect 6270 3681 6329 3715
rect 6270 3647 6279 3681
rect 6313 3647 6329 3681
rect 6270 3629 6329 3647
rect 6365 3749 6699 3791
rect 6365 3715 6383 3749
rect 6417 3715 6647 3749
rect 6681 3715 6699 3749
rect 6365 3647 6699 3715
rect 6365 3613 6383 3647
rect 6417 3613 6647 3647
rect 6681 3613 6699 3647
rect 6734 3741 6785 3757
rect 6734 3707 6751 3741
rect 6734 3673 6785 3707
rect 6819 3725 6885 3791
rect 6819 3691 6835 3725
rect 6869 3691 6885 3725
rect 6919 3741 6953 3757
rect 6734 3639 6751 3673
rect 6919 3673 6953 3707
rect 6785 3639 6884 3657
rect 6734 3623 6884 3639
rect 6365 3573 6699 3613
rect 4810 3513 6234 3529
rect 4810 3479 4830 3513
rect 4864 3479 4898 3513
rect 4932 3479 4966 3513
rect 5000 3479 5034 3513
rect 5068 3479 5102 3513
rect 5136 3479 5170 3513
rect 5204 3479 5238 3513
rect 5272 3479 5306 3513
rect 5340 3479 5374 3513
rect 5408 3479 5442 3513
rect 5476 3479 5510 3513
rect 5544 3479 5578 3513
rect 5612 3479 5646 3513
rect 5680 3479 5714 3513
rect 5748 3479 5782 3513
rect 5816 3479 5850 3513
rect 5884 3479 6234 3513
rect 3427 3407 3478 3423
rect 3461 3383 3478 3407
rect 3069 3339 3219 3357
rect 3253 3339 3283 3373
rect 3069 3323 3283 3339
rect 3332 3357 3393 3373
rect 3332 3323 3343 3357
rect 3377 3323 3393 3357
rect 2997 3281 3035 3319
rect 3332 3281 3393 3323
rect 3427 3349 3433 3373
rect 3467 3349 3478 3383
rect 3427 3317 3478 3349
rect 3697 3409 3755 3426
rect 3697 3375 3709 3409
rect 3743 3375 3755 3409
rect 3697 3281 3755 3375
rect 3789 3376 4491 3435
rect 4543 3411 5892 3445
rect 3789 3342 3807 3376
rect 3841 3342 4439 3376
rect 4473 3342 4491 3376
rect 3789 3281 4491 3342
rect 4543 3361 4603 3377
rect 4543 3327 4560 3361
rect 4594 3327 4603 3361
rect 4543 3281 4603 3327
rect 4637 3370 4689 3411
rect 4637 3336 4646 3370
rect 4680 3336 4689 3370
rect 4637 3320 4689 3336
rect 4723 3361 4775 3377
rect 4723 3327 4732 3361
rect 4766 3327 4775 3361
rect 4723 3281 4775 3327
rect 4811 3370 4863 3411
rect 4811 3336 4818 3370
rect 4852 3336 4863 3370
rect 4811 3320 4863 3336
rect 4897 3361 4947 3377
rect 4897 3327 4904 3361
rect 4938 3327 4947 3361
rect 4897 3281 4947 3327
rect 4983 3370 5035 3411
rect 4983 3336 4990 3370
rect 5024 3336 5035 3370
rect 4983 3320 5035 3336
rect 5069 3361 5119 3377
rect 5069 3327 5076 3361
rect 5110 3327 5119 3361
rect 5069 3281 5119 3327
rect 5155 3370 5207 3411
rect 5155 3336 5162 3370
rect 5196 3336 5207 3370
rect 5155 3320 5207 3336
rect 5241 3361 5290 3377
rect 5241 3327 5247 3361
rect 5281 3327 5290 3361
rect 5241 3281 5290 3327
rect 5324 3370 5379 3411
rect 5324 3336 5333 3370
rect 5367 3336 5379 3370
rect 5324 3320 5379 3336
rect 5413 3361 5462 3377
rect 5413 3327 5419 3361
rect 5453 3327 5462 3361
rect 5413 3281 5462 3327
rect 5496 3370 5548 3411
rect 5496 3336 5505 3370
rect 5539 3336 5548 3370
rect 5496 3320 5548 3336
rect 5582 3361 5634 3377
rect 5582 3327 5591 3361
rect 5625 3327 5634 3361
rect 5582 3281 5634 3327
rect 5668 3370 5720 3411
rect 5668 3336 5677 3370
rect 5711 3336 5720 3370
rect 5668 3320 5720 3336
rect 5754 3361 5806 3377
rect 5754 3327 5763 3361
rect 5797 3327 5806 3361
rect 5754 3281 5806 3327
rect 5840 3370 5892 3411
rect 5840 3336 5849 3370
rect 5883 3336 5892 3370
rect 5840 3320 5892 3336
rect 5926 3370 5978 3393
rect 5926 3336 5935 3370
rect 5969 3336 5978 3370
rect 5926 3281 5978 3336
rect 6012 3370 6062 3479
rect 6012 3336 6021 3370
rect 6055 3336 6062 3370
rect 6012 3317 6062 3336
rect 6098 3370 6150 3386
rect 6098 3336 6107 3370
rect 6141 3336 6150 3370
rect 6098 3281 6150 3336
rect 6184 3370 6234 3479
rect 6268 3519 6331 3529
rect 6268 3513 6285 3519
rect 6268 3479 6277 3513
rect 6319 3485 6331 3519
rect 6311 3479 6331 3485
rect 6268 3417 6331 3479
rect 6365 3505 6385 3539
rect 6419 3505 6515 3539
rect 6365 3435 6515 3505
rect 6549 3503 6699 3573
rect 6549 3469 6645 3503
rect 6679 3469 6699 3503
rect 6734 3519 6804 3589
rect 6734 3485 6745 3519
rect 6779 3513 6804 3519
rect 6734 3479 6748 3485
rect 6782 3479 6804 3513
rect 6734 3459 6804 3479
rect 6838 3528 6884 3623
rect 6838 3519 6850 3528
rect 6872 3485 6884 3494
rect 6365 3383 6699 3435
rect 6838 3425 6884 3485
rect 6184 3336 6193 3370
rect 6227 3336 6234 3370
rect 6184 3317 6234 3336
rect 6270 3357 6331 3383
rect 6270 3323 6279 3357
rect 6313 3323 6331 3357
rect 6270 3281 6331 3323
rect 6365 3349 6383 3383
rect 6417 3349 6647 3383
rect 6681 3349 6699 3383
rect 6365 3281 6699 3349
rect 6734 3391 6884 3425
rect 6734 3383 6785 3391
rect 6734 3349 6751 3383
rect 6919 3383 6953 3621
rect 6987 3597 7052 3754
rect 7086 3749 7136 3791
rect 7086 3715 7102 3749
rect 7086 3699 7136 3715
rect 7170 3741 7220 3757
rect 7170 3707 7186 3741
rect 7170 3691 7220 3707
rect 7263 3747 7399 3757
rect 7263 3713 7279 3747
rect 7313 3713 7399 3747
rect 7514 3739 7580 3791
rect 7707 3749 7781 3791
rect 7263 3691 7399 3713
rect 7170 3665 7204 3691
rect 7125 3631 7204 3665
rect 7238 3655 7331 3657
rect 6999 3574 7091 3597
rect 6999 3540 7057 3574
rect 6999 3451 7091 3540
rect 6999 3417 7021 3451
rect 7055 3417 7091 3451
rect 6999 3387 7091 3417
rect 6734 3333 6785 3349
rect 6819 3323 6835 3357
rect 6869 3323 6885 3357
rect 7125 3359 7159 3631
rect 7238 3629 7297 3655
rect 7272 3621 7297 3629
rect 7272 3595 7331 3621
rect 7238 3579 7331 3595
rect 7193 3519 7263 3541
rect 7193 3485 7205 3519
rect 7239 3485 7263 3519
rect 7193 3467 7263 3485
rect 7193 3433 7216 3467
rect 7250 3433 7263 3467
rect 7193 3417 7263 3433
rect 7297 3461 7331 3579
rect 7365 3535 7399 3691
rect 7433 3723 7467 3739
rect 7514 3705 7530 3739
rect 7564 3705 7580 3739
rect 7614 3723 7648 3739
rect 7433 3671 7467 3689
rect 7707 3715 7727 3749
rect 7761 3715 7781 3749
rect 7707 3699 7781 3715
rect 7815 3741 7849 3757
rect 7614 3671 7648 3689
rect 7433 3637 7648 3671
rect 7815 3665 7849 3707
rect 7896 3748 8070 3757
rect 7896 3714 7912 3748
rect 7946 3714 8070 3748
rect 7896 3689 8070 3714
rect 8104 3749 8154 3791
rect 8138 3715 8154 3749
rect 8258 3749 8324 3791
rect 8104 3699 8154 3715
rect 8188 3723 8222 3739
rect 7737 3631 7849 3665
rect 7737 3603 7771 3631
rect 7471 3569 7487 3603
rect 7521 3569 7771 3603
rect 7910 3621 7921 3655
rect 7955 3629 8002 3655
rect 7910 3597 7952 3621
rect 7365 3515 7703 3535
rect 7365 3501 7669 3515
rect 7297 3427 7318 3461
rect 7352 3427 7368 3461
rect 7297 3417 7368 3427
rect 7402 3359 7436 3501
rect 7477 3451 7573 3467
rect 7511 3417 7549 3451
rect 7607 3433 7635 3467
rect 7669 3465 7703 3481
rect 7583 3417 7635 3433
rect 7737 3431 7771 3569
rect 6919 3333 6953 3349
rect 6819 3281 6885 3323
rect 7025 3319 7041 3353
rect 7075 3319 7091 3353
rect 7125 3325 7174 3359
rect 7208 3325 7224 3359
rect 7265 3325 7281 3359
rect 7315 3325 7436 3359
rect 7611 3357 7677 3373
rect 7025 3281 7091 3319
rect 7611 3323 7627 3357
rect 7661 3323 7677 3357
rect 7611 3281 7677 3323
rect 7719 3353 7771 3431
rect 7809 3595 7952 3597
rect 7986 3595 8002 3629
rect 8036 3613 8070 3689
rect 8258 3715 8274 3749
rect 8308 3715 8324 3749
rect 8392 3749 8453 3791
rect 8392 3715 8403 3749
rect 8437 3715 8453 3749
rect 8573 3749 8815 3791
rect 8188 3681 8222 3689
rect 8392 3681 8453 3715
rect 8188 3647 8348 3681
rect 7809 3563 7944 3595
rect 8036 3579 8230 3613
rect 8264 3579 8280 3613
rect 7809 3455 7851 3563
rect 8036 3561 8070 3579
rect 7809 3421 7817 3455
rect 7809 3405 7851 3421
rect 7885 3519 7955 3529
rect 7885 3503 7921 3519
rect 7885 3469 7913 3503
rect 7947 3469 7955 3485
rect 7885 3405 7955 3469
rect 7989 3527 8070 3561
rect 7989 3371 8023 3527
rect 8137 3514 8245 3545
rect 8314 3529 8348 3647
rect 8392 3647 8403 3681
rect 8437 3647 8453 3681
rect 8392 3563 8453 3647
rect 8487 3713 8538 3729
rect 8521 3679 8538 3713
rect 8487 3655 8538 3679
rect 8487 3645 8493 3655
rect 8527 3621 8538 3655
rect 8521 3611 8538 3621
rect 8487 3553 8538 3611
rect 8573 3715 8591 3749
rect 8625 3715 8763 3749
rect 8797 3715 8815 3749
rect 8573 3654 8815 3715
rect 8573 3620 8591 3654
rect 8625 3620 8763 3654
rect 8797 3620 8815 3654
rect 8573 3573 8815 3620
rect 8314 3523 8462 3529
rect 8171 3505 8245 3514
rect 8057 3477 8101 3493
rect 8091 3443 8101 3477
rect 8137 3471 8153 3480
rect 8187 3471 8245 3505
rect 8057 3437 8101 3443
rect 8197 3451 8245 3471
rect 8057 3403 8163 3437
rect 7833 3357 8023 3371
rect 7719 3319 7739 3353
rect 7773 3319 7789 3353
rect 7833 3323 7849 3357
rect 7883 3323 8023 3357
rect 7833 3315 8023 3323
rect 8057 3353 8095 3369
rect 8057 3319 8061 3353
rect 8129 3357 8163 3403
rect 8231 3417 8245 3451
rect 8197 3391 8245 3417
rect 8279 3513 8462 3523
rect 8279 3479 8428 3513
rect 8279 3463 8462 3479
rect 8279 3428 8344 3463
rect 8279 3373 8343 3428
rect 8496 3423 8538 3553
rect 8487 3407 8538 3423
rect 8521 3373 8538 3407
rect 8129 3339 8279 3357
rect 8313 3339 8343 3373
rect 8129 3323 8343 3339
rect 8392 3357 8453 3373
rect 8392 3323 8403 3357
rect 8437 3323 8453 3357
rect 8057 3281 8095 3319
rect 8392 3281 8453 3323
rect 8487 3317 8538 3373
rect 8573 3505 8623 3539
rect 8657 3505 8677 3539
rect 8573 3431 8677 3505
rect 8711 3499 8815 3573
rect 8849 3720 8907 3791
rect 8849 3686 8861 3720
rect 8895 3686 8907 3720
rect 8849 3627 8907 3686
rect 8849 3593 8861 3627
rect 8895 3593 8907 3627
rect 8849 3558 8907 3593
rect 9143 3741 9177 3757
rect 9143 3673 9177 3707
rect 9220 3741 9286 3791
rect 9220 3707 9236 3741
rect 9270 3707 9286 3741
rect 9220 3673 9286 3707
rect 9220 3639 9236 3673
rect 9270 3639 9286 3673
rect 9320 3725 9371 3757
rect 9320 3691 9322 3725
rect 9356 3691 9371 3725
rect 9320 3655 9371 3691
rect 9143 3605 9177 3639
rect 9320 3621 9321 3655
rect 9355 3644 9371 3655
rect 9320 3610 9322 3621
rect 9356 3610 9371 3644
rect 9143 3571 9286 3605
rect 9320 3576 9371 3610
rect 8711 3465 8731 3499
rect 8765 3465 8815 3499
rect 9125 3519 9196 3535
rect 9125 3485 9137 3519
rect 9171 3513 9196 3519
rect 9125 3479 9145 3485
rect 9179 3479 9196 3513
rect 9125 3461 9196 3479
rect 9252 3529 9286 3571
rect 9252 3513 9303 3529
rect 9252 3479 9269 3513
rect 9252 3463 9303 3479
rect 8573 3378 8815 3431
rect 8573 3344 8591 3378
rect 8625 3344 8763 3378
rect 8797 3344 8815 3378
rect 8573 3281 8815 3344
rect 8849 3409 8907 3426
rect 9252 3425 9286 3463
rect 9337 3430 9371 3576
rect 9406 3749 9458 3791
rect 9440 3715 9458 3749
rect 9406 3681 9458 3715
rect 9440 3647 9458 3681
rect 9406 3613 9458 3647
rect 9440 3579 9458 3613
rect 9406 3561 9458 3579
rect 9493 3749 10011 3791
rect 9493 3715 9511 3749
rect 9545 3715 9959 3749
rect 9993 3715 10011 3749
rect 9493 3647 10011 3715
rect 9493 3613 9511 3647
rect 9545 3613 9959 3647
rect 9993 3613 10011 3647
rect 9493 3573 10011 3613
rect 9493 3505 9571 3539
rect 9605 3505 9681 3539
rect 9715 3505 9735 3539
rect 8849 3375 8861 3409
rect 8895 3375 8907 3409
rect 8849 3281 8907 3375
rect 9143 3391 9286 3425
rect 9143 3370 9177 3391
rect 9320 3387 9371 3430
rect 9143 3315 9177 3336
rect 9220 3323 9236 3357
rect 9270 3323 9286 3357
rect 9220 3281 9286 3323
rect 9320 3353 9322 3387
rect 9356 3353 9371 3387
rect 9320 3315 9371 3353
rect 9406 3429 9458 3449
rect 9440 3395 9458 3429
rect 9406 3361 9458 3395
rect 9440 3327 9458 3361
rect 9406 3281 9458 3327
rect 9493 3435 9735 3505
rect 9769 3503 10011 3573
rect 9769 3469 9789 3503
rect 9823 3469 9899 3503
rect 9933 3469 10011 3503
rect 10045 3741 10099 3757
rect 10045 3707 10063 3741
rect 10097 3707 10099 3741
rect 10045 3660 10099 3707
rect 10045 3626 10063 3660
rect 10097 3626 10099 3660
rect 10133 3741 10199 3791
rect 10133 3707 10149 3741
rect 10183 3707 10199 3741
rect 10133 3673 10199 3707
rect 10133 3639 10149 3673
rect 10183 3639 10199 3673
rect 10235 3741 10269 3757
rect 10235 3673 10269 3707
rect 10045 3576 10099 3626
rect 10235 3605 10269 3639
rect 9493 3376 10011 3435
rect 9493 3342 9511 3376
rect 9545 3342 9959 3376
rect 9993 3342 10011 3376
rect 9493 3281 10011 3342
rect 10045 3416 10079 3576
rect 10136 3571 10269 3605
rect 10321 3749 10839 3791
rect 10321 3715 10339 3749
rect 10373 3715 10787 3749
rect 10821 3715 10839 3749
rect 10321 3647 10839 3715
rect 10321 3613 10339 3647
rect 10373 3613 10787 3647
rect 10821 3613 10839 3647
rect 10321 3573 10839 3613
rect 10136 3542 10170 3571
rect 10113 3526 10170 3542
rect 10147 3492 10170 3526
rect 10113 3476 10170 3492
rect 10136 3425 10170 3476
rect 10217 3519 10283 3535
rect 10217 3513 10241 3519
rect 10217 3479 10233 3513
rect 10275 3485 10283 3519
rect 10267 3479 10283 3485
rect 10217 3461 10283 3479
rect 10321 3505 10399 3539
rect 10433 3505 10509 3539
rect 10543 3505 10563 3539
rect 10321 3435 10563 3505
rect 10597 3503 10839 3573
rect 10983 3741 11017 3757
rect 10983 3673 11017 3707
rect 11053 3741 11119 3791
rect 11053 3707 11069 3741
rect 11103 3707 11119 3741
rect 11053 3673 11119 3707
rect 11053 3639 11069 3673
rect 11103 3639 11119 3673
rect 11153 3741 11207 3757
rect 11153 3707 11155 3741
rect 11189 3707 11207 3741
rect 11153 3660 11207 3707
rect 10983 3605 11017 3639
rect 11153 3626 11155 3660
rect 11189 3655 11207 3660
rect 11153 3621 11161 3626
rect 11195 3621 11207 3655
rect 10983 3571 11116 3605
rect 11153 3576 11207 3621
rect 11082 3542 11116 3571
rect 10597 3469 10617 3503
rect 10651 3469 10727 3503
rect 10761 3469 10839 3503
rect 10969 3519 11035 3535
rect 10969 3485 10977 3519
rect 11011 3513 11035 3519
rect 10969 3479 10985 3485
rect 11019 3479 11035 3513
rect 10969 3461 11035 3479
rect 11082 3526 11139 3542
rect 11082 3492 11105 3526
rect 11082 3476 11139 3492
rect 10045 3387 10097 3416
rect 10136 3391 10269 3425
rect 10045 3383 10063 3387
rect 10045 3349 10057 3383
rect 10235 3370 10269 3391
rect 10091 3349 10097 3353
rect 10045 3315 10097 3349
rect 10133 3323 10149 3357
rect 10183 3323 10199 3357
rect 10133 3281 10199 3323
rect 10235 3315 10269 3336
rect 10321 3376 10839 3435
rect 11082 3425 11116 3476
rect 10321 3342 10339 3376
rect 10373 3342 10787 3376
rect 10821 3342 10839 3376
rect 10321 3281 10839 3342
rect 10983 3391 11116 3425
rect 11173 3416 11207 3576
rect 11241 3749 11943 3791
rect 11241 3715 11259 3749
rect 11293 3715 11891 3749
rect 11925 3715 11943 3749
rect 12063 3749 12124 3791
rect 11241 3647 11943 3715
rect 11241 3613 11259 3647
rect 11293 3613 11891 3647
rect 11925 3613 11943 3647
rect 11241 3573 11943 3613
rect 10983 3370 11017 3391
rect 11155 3387 11207 3416
rect 10983 3315 11017 3336
rect 11053 3323 11069 3357
rect 11103 3323 11119 3357
rect 11053 3281 11119 3323
rect 11189 3353 11207 3387
rect 11155 3315 11207 3353
rect 11241 3505 11319 3539
rect 11353 3505 11418 3539
rect 11452 3505 11517 3539
rect 11551 3505 11571 3539
rect 11241 3435 11571 3505
rect 11605 3503 11943 3573
rect 11605 3469 11625 3503
rect 11659 3469 11728 3503
rect 11762 3469 11831 3503
rect 11865 3469 11943 3503
rect 11978 3713 12029 3729
rect 11978 3679 11995 3713
rect 11978 3655 12029 3679
rect 11978 3621 11989 3655
rect 12023 3645 12029 3655
rect 11978 3611 11995 3621
rect 11978 3553 12029 3611
rect 12063 3715 12079 3749
rect 12113 3715 12124 3749
rect 12192 3749 12258 3791
rect 12192 3715 12208 3749
rect 12242 3715 12258 3749
rect 12362 3749 12412 3791
rect 12294 3723 12328 3739
rect 12063 3681 12124 3715
rect 12362 3715 12378 3749
rect 12362 3699 12412 3715
rect 12446 3748 12620 3757
rect 12446 3714 12570 3748
rect 12604 3714 12620 3748
rect 12294 3681 12328 3689
rect 12063 3647 12079 3681
rect 12113 3647 12124 3681
rect 12063 3563 12124 3647
rect 12168 3647 12328 3681
rect 12446 3689 12620 3714
rect 12667 3741 12701 3757
rect 11241 3376 11943 3435
rect 11241 3342 11259 3376
rect 11293 3342 11891 3376
rect 11925 3342 11943 3376
rect 11241 3281 11943 3342
rect 11978 3423 12020 3553
rect 12168 3529 12202 3647
rect 12446 3613 12480 3689
rect 12667 3665 12701 3707
rect 12735 3749 12809 3791
rect 12735 3715 12755 3749
rect 12789 3715 12809 3749
rect 12936 3739 13002 3791
rect 13117 3747 13253 3757
rect 12735 3699 12809 3715
rect 12868 3723 12902 3739
rect 12936 3705 12952 3739
rect 12986 3705 13002 3739
rect 13049 3723 13083 3739
rect 12868 3671 12902 3689
rect 13049 3671 13083 3689
rect 12236 3579 12252 3613
rect 12286 3579 12480 3613
rect 12514 3629 12561 3655
rect 12514 3595 12530 3629
rect 12595 3621 12606 3655
rect 12667 3631 12779 3665
rect 12868 3637 13083 3671
rect 13117 3713 13203 3747
rect 13237 3713 13253 3747
rect 13117 3691 13253 3713
rect 13296 3741 13346 3757
rect 13330 3707 13346 3741
rect 13296 3691 13346 3707
rect 13380 3749 13430 3791
rect 13414 3715 13430 3749
rect 13380 3699 13430 3715
rect 12564 3597 12606 3621
rect 12745 3603 12779 3631
rect 12564 3595 12707 3597
rect 12446 3561 12480 3579
rect 12572 3563 12707 3595
rect 12054 3523 12202 3529
rect 12054 3513 12237 3523
rect 12088 3479 12237 3513
rect 12054 3463 12237 3479
rect 12172 3428 12237 3463
rect 11978 3407 12029 3423
rect 11978 3373 11995 3407
rect 12173 3373 12237 3428
rect 12271 3514 12379 3545
rect 12446 3527 12527 3561
rect 12271 3505 12345 3514
rect 12271 3471 12329 3505
rect 12363 3471 12379 3480
rect 12415 3477 12459 3493
rect 12271 3451 12319 3471
rect 12271 3417 12285 3451
rect 12415 3443 12425 3477
rect 12415 3437 12459 3443
rect 12271 3391 12319 3417
rect 12353 3403 12459 3437
rect 11978 3317 12029 3373
rect 12063 3357 12124 3373
rect 12063 3323 12079 3357
rect 12113 3323 12124 3357
rect 12173 3339 12203 3373
rect 12353 3357 12387 3403
rect 12493 3371 12527 3527
rect 12561 3519 12631 3529
rect 12595 3503 12631 3519
rect 12561 3469 12569 3485
rect 12603 3469 12631 3503
rect 12561 3405 12631 3469
rect 12665 3455 12707 3563
rect 12699 3421 12707 3455
rect 12665 3405 12707 3421
rect 12745 3569 12995 3603
rect 13029 3569 13045 3603
rect 12745 3431 12779 3569
rect 13117 3535 13151 3691
rect 13312 3665 13346 3691
rect 12813 3515 13151 3535
rect 12847 3501 13151 3515
rect 13185 3655 13278 3657
rect 13219 3629 13278 3655
rect 13312 3631 13391 3665
rect 13219 3621 13244 3629
rect 13185 3595 13244 3621
rect 13185 3579 13278 3595
rect 12813 3465 12847 3481
rect 12881 3433 12909 3467
rect 12943 3451 13039 3467
rect 12237 3339 12387 3357
rect 12173 3323 12387 3339
rect 12421 3353 12459 3369
rect 12063 3281 12124 3323
rect 12455 3319 12459 3353
rect 12421 3281 12459 3319
rect 12493 3357 12683 3371
rect 12493 3323 12633 3357
rect 12667 3323 12683 3357
rect 12745 3353 12797 3431
rect 12881 3417 12933 3433
rect 12967 3417 13005 3451
rect 12493 3315 12683 3323
rect 12727 3319 12743 3353
rect 12777 3319 12797 3353
rect 12839 3357 12905 3373
rect 12839 3323 12855 3357
rect 12889 3323 12905 3357
rect 13080 3359 13114 3501
rect 13185 3461 13219 3579
rect 13148 3427 13164 3461
rect 13198 3427 13219 3461
rect 13148 3417 13219 3427
rect 13253 3519 13323 3541
rect 13253 3485 13277 3519
rect 13311 3485 13323 3519
rect 13253 3467 13323 3485
rect 13253 3433 13266 3467
rect 13300 3433 13323 3467
rect 13253 3417 13323 3433
rect 13357 3359 13391 3631
rect 13464 3597 13529 3754
rect 13563 3741 13597 3757
rect 13563 3673 13597 3707
rect 13631 3725 13697 3791
rect 13631 3691 13647 3725
rect 13681 3691 13697 3725
rect 13731 3741 13782 3757
rect 13765 3707 13782 3741
rect 13731 3673 13782 3707
rect 13425 3574 13517 3597
rect 13459 3540 13517 3574
rect 13425 3451 13517 3540
rect 13425 3417 13461 3451
rect 13495 3417 13517 3451
rect 13425 3387 13517 3417
rect 13080 3325 13201 3359
rect 13235 3325 13251 3359
rect 13292 3325 13308 3359
rect 13342 3325 13391 3359
rect 13563 3383 13597 3621
rect 13632 3639 13731 3657
rect 13765 3639 13782 3673
rect 13632 3623 13782 3639
rect 14001 3720 14059 3791
rect 14001 3686 14013 3720
rect 14047 3686 14059 3720
rect 14093 3749 15162 3791
rect 14093 3715 14111 3749
rect 14145 3715 15111 3749
rect 15145 3715 15162 3749
rect 14093 3704 15162 3715
rect 15197 3749 16266 3791
rect 15197 3715 15215 3749
rect 15249 3715 16215 3749
rect 16249 3715 16266 3749
rect 15197 3704 16266 3715
rect 16301 3749 17370 3791
rect 16301 3715 16319 3749
rect 16353 3715 17319 3749
rect 17353 3715 17370 3749
rect 16301 3704 17370 3715
rect 17405 3749 18474 3791
rect 17405 3715 17423 3749
rect 17457 3715 18423 3749
rect 18457 3715 18474 3749
rect 17405 3704 18474 3715
rect 18601 3749 18843 3791
rect 18601 3715 18619 3749
rect 18653 3715 18791 3749
rect 18825 3715 18843 3749
rect 14001 3627 14059 3686
rect 13632 3528 13678 3623
rect 14001 3593 14013 3627
rect 14047 3593 14059 3627
rect 13666 3519 13678 3528
rect 13632 3485 13644 3494
rect 13632 3425 13678 3485
rect 13712 3587 13782 3589
rect 13712 3553 13737 3587
rect 13771 3553 13782 3587
rect 14001 3558 14059 3593
rect 13712 3513 13782 3553
rect 13712 3479 13734 3513
rect 13768 3479 13782 3513
rect 13712 3459 13782 3479
rect 14410 3539 14478 3556
rect 14410 3505 14427 3539
rect 14461 3505 14478 3539
rect 13632 3391 13782 3425
rect 12839 3281 12905 3323
rect 13425 3319 13441 3353
rect 13475 3319 13491 3353
rect 13731 3383 13782 3391
rect 13563 3333 13597 3349
rect 13425 3281 13491 3319
rect 13631 3323 13647 3357
rect 13681 3323 13697 3357
rect 13765 3349 13782 3383
rect 13731 3333 13782 3349
rect 14001 3409 14059 3426
rect 14001 3375 14013 3409
rect 14047 3375 14059 3409
rect 14410 3390 14478 3505
rect 14774 3503 14844 3704
rect 14774 3469 14791 3503
rect 14825 3469 14844 3503
rect 14774 3454 14844 3469
rect 15514 3539 15582 3556
rect 15514 3505 15531 3539
rect 15565 3505 15582 3539
rect 15514 3390 15582 3505
rect 15878 3503 15948 3704
rect 15878 3469 15895 3503
rect 15929 3469 15948 3503
rect 15878 3454 15948 3469
rect 16618 3539 16686 3556
rect 16618 3505 16635 3539
rect 16669 3505 16686 3539
rect 16618 3390 16686 3505
rect 16982 3503 17052 3704
rect 16982 3469 16999 3503
rect 17033 3469 17052 3503
rect 16982 3454 17052 3469
rect 17722 3539 17790 3556
rect 17722 3505 17739 3539
rect 17773 3505 17790 3539
rect 17722 3390 17790 3505
rect 18086 3503 18156 3704
rect 18086 3469 18103 3503
rect 18137 3469 18156 3503
rect 18086 3454 18156 3469
rect 18601 3654 18843 3715
rect 18601 3620 18619 3654
rect 18653 3620 18791 3654
rect 18825 3620 18843 3654
rect 18601 3573 18843 3620
rect 18601 3499 18705 3573
rect 18601 3465 18651 3499
rect 18685 3465 18705 3499
rect 18739 3505 18759 3539
rect 18793 3505 18843 3539
rect 18739 3431 18843 3505
rect 13631 3281 13697 3323
rect 14001 3281 14059 3375
rect 14093 3376 15162 3390
rect 14093 3342 14111 3376
rect 14145 3342 15111 3376
rect 15145 3342 15162 3376
rect 14093 3281 15162 3342
rect 15197 3376 16266 3390
rect 15197 3342 15215 3376
rect 15249 3342 16215 3376
rect 16249 3342 16266 3376
rect 15197 3281 16266 3342
rect 16301 3376 17370 3390
rect 16301 3342 16319 3376
rect 16353 3342 17319 3376
rect 17353 3342 17370 3376
rect 16301 3281 17370 3342
rect 17405 3376 18474 3390
rect 17405 3342 17423 3376
rect 17457 3342 18423 3376
rect 18457 3342 18474 3376
rect 17405 3281 18474 3342
rect 18601 3378 18843 3431
rect 18601 3344 18619 3378
rect 18653 3344 18791 3378
rect 18825 3344 18843 3378
rect 18601 3281 18843 3344
rect 1104 3247 1133 3281
rect 1167 3247 1225 3281
rect 1259 3247 1317 3281
rect 1351 3247 1409 3281
rect 1443 3247 1501 3281
rect 1535 3247 1593 3281
rect 1627 3247 1685 3281
rect 1719 3247 1777 3281
rect 1811 3247 1869 3281
rect 1903 3247 1961 3281
rect 1995 3247 2053 3281
rect 2087 3247 2145 3281
rect 2179 3247 2237 3281
rect 2271 3247 2329 3281
rect 2363 3247 2421 3281
rect 2455 3247 2513 3281
rect 2547 3247 2605 3281
rect 2639 3247 2697 3281
rect 2731 3247 2789 3281
rect 2823 3247 2881 3281
rect 2915 3247 2973 3281
rect 3007 3247 3065 3281
rect 3099 3247 3157 3281
rect 3191 3247 3249 3281
rect 3283 3247 3341 3281
rect 3375 3247 3433 3281
rect 3467 3247 3525 3281
rect 3559 3247 3617 3281
rect 3651 3247 3709 3281
rect 3743 3247 3801 3281
rect 3835 3247 3893 3281
rect 3927 3247 3985 3281
rect 4019 3247 4077 3281
rect 4111 3247 4169 3281
rect 4203 3247 4261 3281
rect 4295 3247 4353 3281
rect 4387 3247 4445 3281
rect 4479 3247 4537 3281
rect 4571 3247 4629 3281
rect 4663 3247 4721 3281
rect 4755 3247 4813 3281
rect 4847 3247 4905 3281
rect 4939 3247 4997 3281
rect 5031 3247 5089 3281
rect 5123 3247 5181 3281
rect 5215 3247 5273 3281
rect 5307 3247 5365 3281
rect 5399 3247 5457 3281
rect 5491 3247 5549 3281
rect 5583 3247 5641 3281
rect 5675 3247 5733 3281
rect 5767 3247 5825 3281
rect 5859 3247 5917 3281
rect 5951 3247 6009 3281
rect 6043 3247 6101 3281
rect 6135 3247 6193 3281
rect 6227 3247 6285 3281
rect 6319 3247 6377 3281
rect 6411 3247 6469 3281
rect 6503 3247 6561 3281
rect 6595 3247 6653 3281
rect 6687 3247 6745 3281
rect 6779 3247 6837 3281
rect 6871 3247 6929 3281
rect 6963 3247 7021 3281
rect 7055 3247 7113 3281
rect 7147 3247 7205 3281
rect 7239 3247 7297 3281
rect 7331 3247 7389 3281
rect 7423 3247 7481 3281
rect 7515 3247 7573 3281
rect 7607 3247 7665 3281
rect 7699 3247 7757 3281
rect 7791 3247 7849 3281
rect 7883 3247 7941 3281
rect 7975 3247 8033 3281
rect 8067 3247 8125 3281
rect 8159 3247 8217 3281
rect 8251 3247 8309 3281
rect 8343 3247 8401 3281
rect 8435 3247 8493 3281
rect 8527 3247 8585 3281
rect 8619 3247 8677 3281
rect 8711 3247 8769 3281
rect 8803 3247 8861 3281
rect 8895 3247 8953 3281
rect 8987 3247 9045 3281
rect 9079 3247 9137 3281
rect 9171 3247 9229 3281
rect 9263 3247 9321 3281
rect 9355 3247 9413 3281
rect 9447 3247 9505 3281
rect 9539 3247 9597 3281
rect 9631 3247 9689 3281
rect 9723 3247 9781 3281
rect 9815 3247 9873 3281
rect 9907 3247 9965 3281
rect 9999 3247 10057 3281
rect 10091 3247 10149 3281
rect 10183 3247 10241 3281
rect 10275 3247 10333 3281
rect 10367 3247 10425 3281
rect 10459 3247 10517 3281
rect 10551 3247 10609 3281
rect 10643 3247 10701 3281
rect 10735 3247 10793 3281
rect 10827 3247 10885 3281
rect 10919 3247 10977 3281
rect 11011 3247 11069 3281
rect 11103 3247 11161 3281
rect 11195 3247 11253 3281
rect 11287 3247 11345 3281
rect 11379 3247 11437 3281
rect 11471 3247 11529 3281
rect 11563 3247 11621 3281
rect 11655 3247 11713 3281
rect 11747 3247 11805 3281
rect 11839 3247 11897 3281
rect 11931 3247 11989 3281
rect 12023 3247 12081 3281
rect 12115 3247 12173 3281
rect 12207 3247 12265 3281
rect 12299 3247 12357 3281
rect 12391 3247 12449 3281
rect 12483 3247 12541 3281
rect 12575 3247 12633 3281
rect 12667 3247 12725 3281
rect 12759 3247 12817 3281
rect 12851 3247 12909 3281
rect 12943 3247 13001 3281
rect 13035 3247 13093 3281
rect 13127 3247 13185 3281
rect 13219 3247 13277 3281
rect 13311 3247 13369 3281
rect 13403 3247 13461 3281
rect 13495 3247 13553 3281
rect 13587 3247 13645 3281
rect 13679 3247 13737 3281
rect 13771 3247 13829 3281
rect 13863 3247 13921 3281
rect 13955 3247 14013 3281
rect 14047 3247 14105 3281
rect 14139 3247 14197 3281
rect 14231 3247 14289 3281
rect 14323 3247 14381 3281
rect 14415 3247 14473 3281
rect 14507 3247 14565 3281
rect 14599 3247 14657 3281
rect 14691 3247 14749 3281
rect 14783 3247 14841 3281
rect 14875 3247 14933 3281
rect 14967 3247 15025 3281
rect 15059 3247 15117 3281
rect 15151 3247 15209 3281
rect 15243 3247 15301 3281
rect 15335 3247 15393 3281
rect 15427 3247 15485 3281
rect 15519 3247 15577 3281
rect 15611 3247 15669 3281
rect 15703 3247 15761 3281
rect 15795 3247 15853 3281
rect 15887 3247 15945 3281
rect 15979 3247 16037 3281
rect 16071 3247 16129 3281
rect 16163 3247 16221 3281
rect 16255 3247 16313 3281
rect 16347 3247 16405 3281
rect 16439 3247 16497 3281
rect 16531 3247 16589 3281
rect 16623 3247 16681 3281
rect 16715 3247 16773 3281
rect 16807 3247 16865 3281
rect 16899 3247 16957 3281
rect 16991 3247 17049 3281
rect 17083 3247 17141 3281
rect 17175 3247 17233 3281
rect 17267 3247 17325 3281
rect 17359 3247 17417 3281
rect 17451 3247 17509 3281
rect 17543 3247 17601 3281
rect 17635 3247 17693 3281
rect 17727 3247 17785 3281
rect 17819 3247 17877 3281
rect 17911 3247 17969 3281
rect 18003 3247 18061 3281
rect 18095 3247 18153 3281
rect 18187 3247 18245 3281
rect 18279 3247 18337 3281
rect 18371 3247 18429 3281
rect 18463 3247 18521 3281
rect 18555 3247 18613 3281
rect 18647 3247 18705 3281
rect 18739 3247 18797 3281
rect 18831 3247 18860 3281
rect 1121 3184 1363 3247
rect 1121 3150 1139 3184
rect 1173 3150 1311 3184
rect 1345 3150 1363 3184
rect 1121 3097 1363 3150
rect 1397 3186 1915 3247
rect 1397 3152 1415 3186
rect 1449 3152 1863 3186
rect 1897 3152 1915 3186
rect 1121 3023 1225 3097
rect 1397 3093 1915 3152
rect 1950 3179 2001 3211
rect 1950 3145 1961 3179
rect 1995 3155 2001 3179
rect 2035 3205 2096 3247
rect 2393 3209 2431 3247
rect 2035 3171 2051 3205
rect 2085 3171 2096 3205
rect 2035 3155 2096 3171
rect 2145 3189 2359 3205
rect 2145 3155 2175 3189
rect 2209 3171 2359 3189
rect 1950 3121 1967 3145
rect 1950 3105 2001 3121
rect 1121 2989 1171 3023
rect 1205 2989 1225 3023
rect 1259 3029 1279 3063
rect 1313 3029 1363 3063
rect 1259 2955 1363 3029
rect 1397 3023 1639 3093
rect 1397 2989 1475 3023
rect 1509 2989 1585 3023
rect 1619 2989 1639 3023
rect 1673 3025 1693 3059
rect 1727 3025 1803 3059
rect 1837 3025 1915 3059
rect 1673 2955 1915 3025
rect 1121 2908 1363 2955
rect 1121 2874 1139 2908
rect 1173 2874 1311 2908
rect 1345 2874 1363 2908
rect 1121 2813 1363 2874
rect 1121 2779 1139 2813
rect 1173 2779 1311 2813
rect 1345 2779 1363 2813
rect 1121 2737 1363 2779
rect 1397 2915 1915 2955
rect 1397 2881 1415 2915
rect 1449 2881 1863 2915
rect 1897 2881 1915 2915
rect 1397 2813 1915 2881
rect 1397 2779 1415 2813
rect 1449 2779 1863 2813
rect 1897 2779 1915 2813
rect 1950 2975 1992 3105
rect 2145 3100 2209 3155
rect 2144 3065 2209 3100
rect 2026 3049 2209 3065
rect 2060 3015 2209 3049
rect 2026 3005 2209 3015
rect 2243 3111 2291 3137
rect 2243 3077 2257 3111
rect 2325 3125 2359 3171
rect 2427 3175 2431 3209
rect 2393 3159 2431 3175
rect 2465 3205 2655 3213
rect 2465 3171 2605 3205
rect 2639 3171 2655 3205
rect 2699 3175 2715 3209
rect 2749 3175 2769 3209
rect 2465 3157 2655 3171
rect 2325 3091 2431 3125
rect 2243 3057 2291 3077
rect 2387 3085 2431 3091
rect 2243 3023 2301 3057
rect 2335 3048 2351 3057
rect 2387 3051 2397 3085
rect 2387 3035 2431 3051
rect 2243 3014 2317 3023
rect 2026 2999 2174 3005
rect 1950 2917 2001 2975
rect 1950 2883 1967 2917
rect 1950 2849 2001 2883
rect 1950 2815 1967 2849
rect 1950 2799 2001 2815
rect 2035 2881 2096 2965
rect 2035 2847 2051 2881
rect 2085 2847 2096 2881
rect 2140 2881 2174 2999
rect 2243 2983 2351 3014
rect 2465 3001 2499 3157
rect 2418 2967 2499 3001
rect 2533 3059 2603 3123
rect 2533 3043 2541 3059
rect 2575 3025 2603 3059
rect 2567 3009 2603 3025
rect 2533 2999 2603 3009
rect 2637 3107 2679 3123
rect 2671 3073 2679 3107
rect 2418 2949 2452 2967
rect 2637 2965 2679 3073
rect 2208 2915 2224 2949
rect 2258 2915 2452 2949
rect 2544 2933 2679 2965
rect 2140 2847 2300 2881
rect 2035 2813 2096 2847
rect 2266 2839 2300 2847
rect 1397 2737 1915 2779
rect 2035 2779 2051 2813
rect 2085 2779 2096 2813
rect 2035 2737 2096 2779
rect 2164 2779 2180 2813
rect 2214 2779 2230 2813
rect 2418 2839 2452 2915
rect 2486 2899 2502 2933
rect 2536 2931 2679 2933
rect 2717 3097 2769 3175
rect 2811 3205 2877 3247
rect 2811 3171 2827 3205
rect 2861 3171 2877 3205
rect 3397 3209 3463 3247
rect 2811 3155 2877 3171
rect 3052 3169 3173 3203
rect 3207 3169 3223 3203
rect 3264 3169 3280 3203
rect 3314 3169 3363 3203
rect 3397 3175 3413 3209
rect 3447 3175 3463 3209
rect 3603 3205 3669 3247
rect 3535 3179 3569 3195
rect 2717 2959 2751 3097
rect 2853 3095 2905 3111
rect 2785 3047 2819 3063
rect 2853 3061 2881 3095
rect 2939 3077 2977 3111
rect 2915 3061 3011 3077
rect 3052 3027 3086 3169
rect 3120 3101 3191 3111
rect 3120 3067 3136 3101
rect 3170 3067 3191 3101
rect 2819 3013 3123 3027
rect 2785 2993 3123 3013
rect 2536 2907 2578 2931
rect 2486 2873 2533 2899
rect 2567 2873 2578 2907
rect 2717 2925 2967 2959
rect 3001 2925 3017 2959
rect 2717 2897 2751 2925
rect 2639 2863 2751 2897
rect 2266 2789 2300 2805
rect 2334 2813 2384 2829
rect 2164 2737 2230 2779
rect 2334 2779 2350 2813
rect 2334 2737 2384 2779
rect 2418 2814 2592 2839
rect 2418 2780 2542 2814
rect 2576 2780 2592 2814
rect 2418 2771 2592 2780
rect 2639 2821 2673 2863
rect 2840 2857 3055 2891
rect 2840 2839 2874 2857
rect 2639 2771 2673 2787
rect 2707 2813 2781 2829
rect 2707 2779 2727 2813
rect 2761 2779 2781 2813
rect 3021 2839 3055 2857
rect 2840 2789 2874 2805
rect 2908 2789 2924 2823
rect 2958 2789 2974 2823
rect 3021 2789 3055 2805
rect 3089 2837 3123 2993
rect 3157 2949 3191 3067
rect 3225 3095 3295 3111
rect 3225 3061 3238 3095
rect 3272 3061 3295 3095
rect 3225 3043 3295 3061
rect 3225 3009 3249 3043
rect 3283 3009 3295 3043
rect 3225 2987 3295 3009
rect 3157 2933 3250 2949
rect 3157 2907 3216 2933
rect 3191 2899 3216 2907
rect 3191 2873 3250 2899
rect 3329 2897 3363 3169
rect 3603 3171 3619 3205
rect 3653 3171 3669 3205
rect 3703 3179 3754 3195
rect 3397 3111 3489 3141
rect 3397 3077 3433 3111
rect 3467 3077 3489 3111
rect 3397 2988 3489 3077
rect 3431 2954 3489 2988
rect 3397 2931 3489 2954
rect 3157 2871 3250 2873
rect 3284 2863 3363 2897
rect 3284 2837 3318 2863
rect 3089 2815 3225 2837
rect 2707 2737 2781 2779
rect 2908 2737 2974 2789
rect 3089 2781 3175 2815
rect 3209 2781 3225 2815
rect 3089 2771 3225 2781
rect 3268 2821 3318 2837
rect 3302 2787 3318 2821
rect 3268 2771 3318 2787
rect 3352 2813 3402 2829
rect 3386 2779 3402 2813
rect 3352 2737 3402 2779
rect 3436 2774 3501 2931
rect 3535 2907 3569 3145
rect 3737 3145 3754 3179
rect 3703 3137 3754 3145
rect 3604 3103 3754 3137
rect 3789 3179 4123 3247
rect 4243 3205 4309 3247
rect 3789 3145 3807 3179
rect 3841 3145 4071 3179
rect 4105 3145 4123 3179
rect 3604 3043 3650 3103
rect 3789 3093 4123 3145
rect 4175 3179 4209 3195
rect 4243 3171 4259 3205
rect 4293 3171 4309 3205
rect 4431 3205 4497 3247
rect 4343 3179 4388 3195
rect 4175 3137 4209 3145
rect 4377 3145 4388 3179
rect 4431 3171 4447 3205
rect 4481 3171 4497 3205
rect 4625 3205 4828 3211
rect 4531 3187 4565 3203
rect 4175 3103 4308 3137
rect 3604 3034 3616 3043
rect 3638 3000 3650 3009
rect 3604 2905 3650 3000
rect 3684 3049 3754 3069
rect 3684 3015 3706 3049
rect 3740 3043 3754 3049
rect 3684 3009 3709 3015
rect 3743 3009 3754 3043
rect 3684 2939 3754 3009
rect 3789 3023 3939 3093
rect 3789 2989 3809 3023
rect 3843 2989 3939 3023
rect 3973 3025 4069 3059
rect 4103 3025 4123 3059
rect 3973 2955 4123 3025
rect 3789 2915 4123 2955
rect 4158 3043 4228 3069
rect 4158 3009 4169 3043
rect 4203 3034 4228 3043
rect 4158 3000 4172 3009
rect 4206 3000 4228 3034
rect 4158 2939 4228 3000
rect 4262 3034 4308 3103
rect 4262 3000 4274 3034
rect 3604 2889 3754 2905
rect 3604 2871 3703 2889
rect 3535 2821 3569 2855
rect 3737 2855 3754 2889
rect 3535 2771 3569 2787
rect 3603 2803 3619 2837
rect 3653 2803 3669 2837
rect 3603 2737 3669 2803
rect 3703 2821 3754 2855
rect 3737 2787 3754 2821
rect 3703 2771 3754 2787
rect 3789 2881 3807 2915
rect 3841 2881 4071 2915
rect 4105 2881 4123 2915
rect 4262 2907 4308 3000
rect 3789 2813 4123 2881
rect 3789 2779 3807 2813
rect 3841 2779 4071 2813
rect 4105 2779 4123 2813
rect 3789 2737 4123 2779
rect 4175 2889 4262 2905
rect 4209 2873 4262 2889
rect 4296 2873 4308 2907
rect 4209 2871 4308 2873
rect 4343 3111 4388 3145
rect 4625 3171 4641 3205
rect 4675 3171 4828 3205
rect 4531 3137 4565 3153
rect 4343 3077 4354 3111
rect 4343 2889 4388 3077
rect 4175 2821 4209 2855
rect 4377 2855 4388 2889
rect 4426 3099 4565 3137
rect 4610 3107 4654 3123
rect 4426 2905 4460 3099
rect 4644 3073 4654 3107
rect 4494 3047 4576 3063
rect 4528 3043 4576 3047
rect 4528 3013 4537 3043
rect 4494 3009 4537 3013
rect 4571 3009 4576 3043
rect 4494 2939 4576 3009
rect 4610 2949 4654 3073
rect 4690 3111 4760 3135
rect 4690 3095 4726 3111
rect 4690 3061 4706 3095
rect 4740 3061 4760 3077
rect 4794 3025 4828 3171
rect 4862 3209 4944 3247
rect 4896 3175 4944 3209
rect 5092 3205 5156 3247
rect 4862 3159 4944 3175
rect 5002 3189 5052 3205
rect 5002 3155 5018 3189
rect 5092 3171 5122 3205
rect 5092 3155 5156 3171
rect 5268 3169 5284 3203
rect 5318 3169 5438 3203
rect 5002 3119 5052 3155
rect 4862 3111 4944 3117
rect 4862 3085 4910 3111
rect 4862 3051 4878 3085
rect 4912 3051 4944 3077
rect 5002 3051 5086 3119
rect 4744 3017 4828 3025
rect 4744 3001 5014 3017
rect 4744 2983 4980 3001
rect 4610 2933 4710 2949
rect 4610 2907 4676 2933
rect 4426 2889 4565 2905
rect 4426 2871 4531 2889
rect 4175 2771 4209 2787
rect 4243 2803 4259 2837
rect 4293 2803 4309 2837
rect 4243 2737 4309 2803
rect 4343 2821 4388 2855
rect 4610 2873 4634 2907
rect 4668 2899 4676 2907
rect 4668 2873 4710 2899
rect 4377 2787 4388 2821
rect 4343 2771 4388 2787
rect 4431 2803 4447 2837
rect 4481 2803 4497 2837
rect 4431 2737 4497 2803
rect 4531 2821 4565 2855
rect 4744 2814 4778 2983
rect 4964 2967 4980 2983
rect 4964 2951 5014 2967
rect 4812 2933 4862 2949
rect 4846 2899 4862 2933
rect 4812 2897 4862 2899
rect 5048 2897 5086 3051
rect 4812 2847 5086 2897
rect 5120 3095 5370 3119
rect 5120 3085 5320 3095
rect 5120 2933 5154 3085
rect 5304 3061 5320 3085
rect 5354 3061 5370 3095
rect 5188 3043 5224 3051
rect 5188 2995 5190 3043
rect 5404 3017 5438 3169
rect 5478 3185 5610 3247
rect 5836 3205 5893 3247
rect 5478 3151 5542 3185
rect 5576 3151 5610 3185
rect 5646 3178 5710 3194
rect 5680 3144 5710 3178
rect 5646 3128 5710 3144
rect 5476 3111 5608 3117
rect 5476 3085 5562 3111
rect 5476 3051 5492 3085
rect 5526 3077 5562 3085
rect 5596 3077 5608 3111
rect 5526 3063 5608 3077
rect 5526 3051 5542 3063
rect 5572 3017 5588 3029
rect 5188 2969 5224 2995
rect 5258 2995 5588 3017
rect 5622 2995 5638 3029
rect 5258 2983 5638 2995
rect 5120 2899 5158 2933
rect 5192 2907 5224 2933
rect 5120 2873 5190 2899
rect 5120 2871 5224 2873
rect 5258 2881 5292 2983
rect 5672 2949 5710 3128
rect 5326 2915 5342 2949
rect 5376 2915 5710 2949
rect 5646 2911 5710 2915
rect 5750 3179 5800 3195
rect 5784 3145 5800 3179
rect 5836 3171 5845 3205
rect 5879 3171 5893 3205
rect 5836 3155 5893 3171
rect 5929 3155 5980 3211
rect 5750 3065 5800 3145
rect 5963 3121 5980 3155
rect 5929 3105 5980 3121
rect 5750 3049 5910 3065
rect 5750 3015 5876 3049
rect 5750 2999 5910 3015
rect 5646 2907 5680 2911
rect 5258 2847 5500 2881
rect 4531 2771 4565 2787
rect 4612 2780 4628 2814
rect 4662 2780 4778 2814
rect 4938 2839 4972 2847
rect 4826 2779 4842 2813
rect 4876 2779 4902 2813
rect 5258 2831 5292 2847
rect 5166 2815 5292 2831
rect 4938 2789 4972 2805
rect 4826 2737 4902 2779
rect 5006 2779 5022 2813
rect 5056 2779 5072 2813
rect 5166 2781 5182 2815
rect 5216 2781 5292 2815
rect 5452 2839 5500 2847
rect 5006 2737 5072 2779
rect 5328 2779 5362 2813
rect 5396 2779 5412 2813
rect 5452 2805 5466 2839
rect 5452 2789 5500 2805
rect 5546 2839 5612 2875
rect 5546 2805 5562 2839
rect 5596 2805 5612 2839
rect 5328 2737 5412 2779
rect 5546 2737 5612 2805
rect 5750 2881 5800 2999
rect 5944 2975 5980 3105
rect 6273 3153 6331 3247
rect 6273 3119 6285 3153
rect 6319 3119 6331 3153
rect 6273 3102 6331 3119
rect 6365 3186 7067 3247
rect 6365 3152 6383 3186
rect 6417 3152 7015 3186
rect 7049 3152 7067 3186
rect 6365 3093 7067 3152
rect 7194 3179 7245 3211
rect 7194 3145 7205 3179
rect 7239 3155 7245 3179
rect 7279 3205 7340 3247
rect 7637 3209 7675 3247
rect 7279 3171 7295 3205
rect 7329 3171 7340 3205
rect 7279 3155 7340 3171
rect 7389 3189 7603 3205
rect 7389 3155 7419 3189
rect 7453 3171 7603 3189
rect 7194 3121 7211 3145
rect 7194 3105 7245 3121
rect 6365 3023 6695 3093
rect 6365 2989 6443 3023
rect 6477 2989 6542 3023
rect 6576 2989 6641 3023
rect 6675 2989 6695 3023
rect 6729 3025 6749 3059
rect 6783 3025 6852 3059
rect 6886 3025 6955 3059
rect 6989 3025 7067 3059
rect 5944 2941 5963 2975
rect 5944 2933 5980 2941
rect 5929 2917 5980 2933
rect 5646 2839 5680 2873
rect 5646 2789 5680 2805
rect 5734 2847 5750 2881
rect 5784 2847 5800 2881
rect 5734 2813 5800 2847
rect 5734 2779 5750 2813
rect 5784 2779 5800 2813
rect 5836 2881 5893 2897
rect 5836 2847 5845 2881
rect 5879 2847 5893 2881
rect 5836 2813 5893 2847
rect 5836 2779 5845 2813
rect 5879 2779 5893 2813
rect 5963 2883 5980 2917
rect 5929 2849 5980 2883
rect 5963 2815 5980 2849
rect 5929 2799 5980 2815
rect 6273 2935 6331 2970
rect 6729 2955 7067 3025
rect 6273 2901 6285 2935
rect 6319 2901 6331 2935
rect 6273 2842 6331 2901
rect 6273 2808 6285 2842
rect 6319 2808 6331 2842
rect 5836 2737 5893 2779
rect 6273 2737 6331 2808
rect 6365 2915 7067 2955
rect 6365 2881 6383 2915
rect 6417 2881 7015 2915
rect 7049 2881 7067 2915
rect 6365 2813 7067 2881
rect 6365 2779 6383 2813
rect 6417 2779 7015 2813
rect 7049 2779 7067 2813
rect 7194 2975 7236 3105
rect 7389 3100 7453 3155
rect 7388 3065 7453 3100
rect 7270 3049 7453 3065
rect 7304 3015 7453 3049
rect 7270 3005 7453 3015
rect 7487 3111 7535 3137
rect 7487 3077 7501 3111
rect 7569 3125 7603 3171
rect 7671 3175 7675 3209
rect 7637 3159 7675 3175
rect 7709 3205 7899 3213
rect 7709 3171 7849 3205
rect 7883 3171 7899 3205
rect 7943 3175 7959 3209
rect 7993 3175 8013 3209
rect 7709 3157 7899 3171
rect 7569 3091 7675 3125
rect 7487 3057 7535 3077
rect 7631 3085 7675 3091
rect 7487 3023 7545 3057
rect 7579 3048 7595 3057
rect 7631 3051 7641 3085
rect 7631 3035 7675 3051
rect 7487 3014 7561 3023
rect 7270 2999 7418 3005
rect 7194 2917 7245 2975
rect 7194 2883 7211 2917
rect 7194 2849 7245 2883
rect 7194 2815 7211 2849
rect 7194 2799 7245 2815
rect 7279 2881 7340 2965
rect 7279 2847 7295 2881
rect 7329 2847 7340 2881
rect 7384 2881 7418 2999
rect 7487 2983 7595 3014
rect 7709 3001 7743 3157
rect 7662 2967 7743 3001
rect 7777 3059 7847 3123
rect 7777 3043 7785 3059
rect 7819 3025 7847 3059
rect 7811 3009 7847 3025
rect 7777 2999 7847 3009
rect 7881 3107 7923 3123
rect 7915 3073 7923 3107
rect 7662 2949 7696 2967
rect 7881 2965 7923 3073
rect 7452 2915 7468 2949
rect 7502 2915 7696 2949
rect 7788 2933 7923 2965
rect 7384 2847 7544 2881
rect 7279 2813 7340 2847
rect 7510 2839 7544 2847
rect 6365 2737 7067 2779
rect 7279 2779 7295 2813
rect 7329 2779 7340 2813
rect 7279 2737 7340 2779
rect 7408 2779 7424 2813
rect 7458 2779 7474 2813
rect 7662 2839 7696 2915
rect 7730 2899 7746 2933
rect 7780 2931 7923 2933
rect 7961 3097 8013 3175
rect 8055 3205 8121 3247
rect 8055 3171 8071 3205
rect 8105 3171 8121 3205
rect 8641 3209 8707 3247
rect 8055 3155 8121 3171
rect 8296 3169 8417 3203
rect 8451 3169 8467 3203
rect 8508 3169 8524 3203
rect 8558 3169 8607 3203
rect 8641 3175 8657 3209
rect 8691 3175 8707 3209
rect 8847 3205 8913 3247
rect 8779 3179 8813 3195
rect 7961 2959 7995 3097
rect 8097 3095 8149 3111
rect 8029 3047 8063 3063
rect 8097 3061 8125 3095
rect 8183 3077 8221 3111
rect 8159 3061 8255 3077
rect 8296 3027 8330 3169
rect 8364 3101 8435 3111
rect 8364 3067 8380 3101
rect 8414 3067 8435 3101
rect 8063 3013 8367 3027
rect 8029 2993 8367 3013
rect 7780 2907 7822 2931
rect 7730 2873 7777 2899
rect 7811 2873 7822 2907
rect 7961 2925 8211 2959
rect 8245 2925 8261 2959
rect 7961 2897 7995 2925
rect 7883 2863 7995 2897
rect 7510 2789 7544 2805
rect 7578 2813 7628 2829
rect 7408 2737 7474 2779
rect 7578 2779 7594 2813
rect 7578 2737 7628 2779
rect 7662 2814 7836 2839
rect 7662 2780 7786 2814
rect 7820 2780 7836 2814
rect 7662 2771 7836 2780
rect 7883 2821 7917 2863
rect 8084 2857 8299 2891
rect 8084 2839 8118 2857
rect 7883 2771 7917 2787
rect 7951 2813 8025 2829
rect 7951 2779 7971 2813
rect 8005 2779 8025 2813
rect 8265 2839 8299 2857
rect 8084 2789 8118 2805
rect 8152 2789 8168 2823
rect 8202 2789 8218 2823
rect 8265 2789 8299 2805
rect 8333 2837 8367 2993
rect 8401 2949 8435 3067
rect 8469 3095 8539 3111
rect 8469 3061 8482 3095
rect 8516 3061 8539 3095
rect 8469 3043 8539 3061
rect 8469 3009 8493 3043
rect 8527 3009 8539 3043
rect 8469 2987 8539 3009
rect 8401 2933 8494 2949
rect 8401 2907 8460 2933
rect 8435 2899 8460 2907
rect 8435 2873 8494 2899
rect 8573 2897 8607 3169
rect 8847 3171 8863 3205
rect 8897 3171 8913 3205
rect 8947 3179 8998 3195
rect 8641 3111 8733 3141
rect 8641 3077 8689 3111
rect 8723 3077 8733 3111
rect 8641 2988 8733 3077
rect 8675 2954 8733 2988
rect 8641 2931 8733 2954
rect 8401 2871 8494 2873
rect 8528 2863 8607 2897
rect 8528 2837 8562 2863
rect 8333 2815 8469 2837
rect 7951 2737 8025 2779
rect 8152 2737 8218 2789
rect 8333 2781 8419 2815
rect 8453 2781 8469 2815
rect 8333 2771 8469 2781
rect 8512 2821 8562 2837
rect 8546 2787 8562 2821
rect 8512 2771 8562 2787
rect 8596 2813 8646 2829
rect 8630 2779 8646 2813
rect 8596 2737 8646 2779
rect 8680 2774 8745 2931
rect 8779 2907 8813 3145
rect 8981 3145 8998 3179
rect 8947 3137 8998 3145
rect 8848 3103 8998 3137
rect 9033 3179 9367 3247
rect 9033 3145 9051 3179
rect 9085 3145 9315 3179
rect 9349 3145 9367 3179
rect 9401 3205 9462 3247
rect 9401 3171 9419 3205
rect 9453 3171 9462 3205
rect 9401 3145 9462 3171
rect 9498 3192 9548 3211
rect 9498 3158 9505 3192
rect 9539 3158 9548 3192
rect 8848 3043 8894 3103
rect 9033 3093 9367 3145
rect 8848 3034 8860 3043
rect 8882 3000 8894 3009
rect 8848 2905 8894 3000
rect 8928 3049 8998 3069
rect 8928 3015 8950 3049
rect 8984 3015 8998 3049
rect 8928 2975 8998 3015
rect 9033 3023 9183 3093
rect 9401 3077 9413 3111
rect 9447 3077 9464 3111
rect 9033 2989 9053 3023
rect 9087 2989 9183 3023
rect 9217 3025 9313 3059
rect 9347 3025 9367 3059
rect 8928 2941 8953 2975
rect 8987 2941 8998 2975
rect 9217 2955 9367 3025
rect 9401 3049 9464 3077
rect 9401 3015 9421 3049
rect 9455 3015 9464 3049
rect 9401 2999 9464 3015
rect 9498 3049 9548 3158
rect 9582 3192 9634 3247
rect 9582 3158 9591 3192
rect 9625 3158 9634 3192
rect 9582 3142 9634 3158
rect 9670 3192 9720 3211
rect 9670 3158 9677 3192
rect 9711 3158 9720 3192
rect 9670 3049 9720 3158
rect 9754 3192 9806 3247
rect 9754 3158 9763 3192
rect 9797 3158 9806 3192
rect 9754 3135 9806 3158
rect 9840 3192 9892 3208
rect 9840 3158 9849 3192
rect 9883 3158 9892 3192
rect 9840 3117 9892 3158
rect 9926 3201 9978 3247
rect 9926 3167 9935 3201
rect 9969 3167 9978 3201
rect 9926 3151 9978 3167
rect 10012 3192 10064 3208
rect 10012 3158 10021 3192
rect 10055 3158 10064 3192
rect 10012 3117 10064 3158
rect 10098 3201 10150 3247
rect 10098 3167 10107 3201
rect 10141 3167 10150 3201
rect 10098 3151 10150 3167
rect 10184 3192 10236 3208
rect 10184 3158 10193 3192
rect 10227 3158 10236 3192
rect 10184 3117 10236 3158
rect 10270 3201 10319 3247
rect 10270 3167 10279 3201
rect 10313 3167 10319 3201
rect 10270 3151 10319 3167
rect 10353 3192 10408 3208
rect 10353 3158 10365 3192
rect 10399 3158 10408 3192
rect 10353 3117 10408 3158
rect 10442 3201 10491 3247
rect 10442 3167 10451 3201
rect 10485 3167 10491 3201
rect 10442 3151 10491 3167
rect 10525 3192 10577 3208
rect 10525 3158 10536 3192
rect 10570 3158 10577 3192
rect 10525 3117 10577 3158
rect 10613 3201 10663 3247
rect 10613 3167 10622 3201
rect 10656 3167 10663 3201
rect 10613 3151 10663 3167
rect 10697 3192 10749 3208
rect 10697 3158 10708 3192
rect 10742 3158 10749 3192
rect 10697 3117 10749 3158
rect 10785 3201 10835 3247
rect 10785 3167 10794 3201
rect 10828 3167 10835 3201
rect 10785 3151 10835 3167
rect 10869 3192 10921 3208
rect 10869 3158 10880 3192
rect 10914 3158 10921 3192
rect 10869 3117 10921 3158
rect 10957 3201 11009 3247
rect 10957 3167 10966 3201
rect 11000 3167 11009 3201
rect 10957 3151 11009 3167
rect 11043 3192 11095 3208
rect 11043 3158 11052 3192
rect 11086 3158 11095 3192
rect 11043 3117 11095 3158
rect 11129 3201 11189 3247
rect 11129 3167 11138 3201
rect 11172 3167 11189 3201
rect 11129 3151 11189 3167
rect 11425 3153 11483 3247
rect 11425 3119 11437 3153
rect 11471 3119 11483 3153
rect 9840 3083 11189 3117
rect 11425 3102 11483 3119
rect 11702 3155 11753 3211
rect 11787 3205 11848 3247
rect 12145 3209 12183 3247
rect 11787 3171 11803 3205
rect 11837 3171 11848 3205
rect 11787 3155 11848 3171
rect 11897 3189 12111 3205
rect 11897 3155 11927 3189
rect 11961 3171 12111 3189
rect 11702 3121 11719 3155
rect 11702 3105 11753 3121
rect 9498 3015 9848 3049
rect 9882 3015 9916 3049
rect 9950 3015 9984 3049
rect 10018 3015 10052 3049
rect 10086 3015 10120 3049
rect 10154 3015 10188 3049
rect 10222 3015 10256 3049
rect 10290 3015 10324 3049
rect 10358 3015 10392 3049
rect 10426 3015 10460 3049
rect 10494 3015 10528 3049
rect 10562 3015 10596 3049
rect 10630 3015 10664 3049
rect 10698 3015 10732 3049
rect 10766 3015 10800 3049
rect 10834 3015 10868 3049
rect 10902 3015 10922 3049
rect 9498 2999 10922 3015
rect 8928 2939 8998 2941
rect 9033 2915 9367 2955
rect 8848 2889 8998 2905
rect 8848 2871 8947 2889
rect 8779 2821 8813 2855
rect 8981 2855 8998 2889
rect 8779 2771 8813 2787
rect 8847 2803 8863 2837
rect 8897 2803 8913 2837
rect 8847 2737 8913 2803
rect 8947 2821 8998 2855
rect 8981 2787 8998 2821
rect 8947 2771 8998 2787
rect 9033 2881 9051 2915
rect 9085 2881 9315 2915
rect 9349 2881 9367 2915
rect 9033 2813 9367 2881
rect 9033 2779 9051 2813
rect 9085 2779 9315 2813
rect 9349 2779 9367 2813
rect 9033 2737 9367 2779
rect 9403 2881 9462 2899
rect 9403 2847 9419 2881
rect 9453 2847 9462 2881
rect 9403 2813 9462 2847
rect 9403 2779 9419 2813
rect 9453 2779 9462 2813
rect 9403 2737 9462 2779
rect 9498 2889 9547 2999
rect 9498 2855 9505 2889
rect 9539 2855 9547 2889
rect 9498 2821 9547 2855
rect 9498 2787 9505 2821
rect 9539 2787 9547 2821
rect 9498 2771 9547 2787
rect 9582 2881 9634 2899
rect 9582 2847 9591 2881
rect 9625 2847 9634 2881
rect 9582 2813 9634 2847
rect 9582 2779 9591 2813
rect 9625 2779 9634 2813
rect 9582 2737 9634 2779
rect 9670 2897 9720 2999
rect 10956 2965 11189 3083
rect 11702 2975 11744 3105
rect 11897 3100 11961 3155
rect 11896 3065 11961 3100
rect 11778 3049 11961 3065
rect 11812 3015 11961 3049
rect 11778 3005 11961 3015
rect 11995 3111 12043 3137
rect 11995 3077 12009 3111
rect 12077 3125 12111 3171
rect 12179 3175 12183 3209
rect 12145 3159 12183 3175
rect 12217 3205 12407 3213
rect 12217 3171 12357 3205
rect 12391 3171 12407 3205
rect 12451 3175 12467 3209
rect 12501 3175 12521 3209
rect 12217 3157 12407 3171
rect 12077 3091 12183 3125
rect 11995 3057 12043 3077
rect 12139 3085 12183 3091
rect 11995 3023 12053 3057
rect 12087 3048 12103 3057
rect 12139 3051 12149 3085
rect 12139 3035 12183 3051
rect 11995 3014 12069 3023
rect 11778 2999 11926 3005
rect 9840 2943 11189 2965
rect 9840 2909 9849 2943
rect 9883 2917 10021 2943
rect 9883 2909 9892 2917
rect 9670 2863 9677 2897
rect 9711 2863 9720 2897
rect 9670 2829 9720 2863
rect 9670 2795 9677 2829
rect 9711 2795 9720 2829
rect 9670 2772 9720 2795
rect 9754 2881 9806 2897
rect 9754 2847 9763 2881
rect 9797 2847 9806 2881
rect 9754 2813 9806 2847
rect 9754 2779 9763 2813
rect 9797 2779 9806 2813
rect 9754 2738 9806 2779
rect 9840 2857 9892 2909
rect 10012 2909 10021 2917
rect 10055 2917 10193 2943
rect 10055 2909 10064 2917
rect 9840 2823 9849 2857
rect 9883 2823 9892 2857
rect 9840 2772 9892 2823
rect 9926 2837 9978 2883
rect 9926 2803 9935 2837
rect 9969 2803 9978 2837
rect 9926 2738 9978 2803
rect 10012 2857 10064 2909
rect 10184 2909 10193 2917
rect 10227 2917 10365 2943
rect 10227 2909 10236 2917
rect 10012 2823 10021 2857
rect 10055 2823 10064 2857
rect 10012 2772 10064 2823
rect 10098 2837 10150 2883
rect 10098 2803 10107 2837
rect 10141 2803 10150 2837
rect 10098 2738 10150 2803
rect 10184 2857 10236 2909
rect 10356 2909 10365 2917
rect 10399 2917 10536 2943
rect 10399 2909 10408 2917
rect 10184 2823 10193 2857
rect 10227 2823 10236 2857
rect 10184 2772 10236 2823
rect 10270 2837 10322 2883
rect 10270 2803 10279 2837
rect 10313 2803 10322 2837
rect 10270 2738 10322 2803
rect 10356 2857 10408 2909
rect 10525 2909 10536 2917
rect 10570 2917 10708 2943
rect 10570 2909 10577 2917
rect 10356 2823 10365 2857
rect 10399 2823 10408 2857
rect 10356 2772 10408 2823
rect 10442 2837 10491 2883
rect 10442 2803 10451 2837
rect 10485 2803 10491 2837
rect 10442 2738 10491 2803
rect 10525 2857 10577 2909
rect 10697 2909 10708 2917
rect 10742 2917 10880 2943
rect 10742 2909 10749 2917
rect 10697 2907 10749 2909
rect 10525 2823 10536 2857
rect 10570 2823 10577 2857
rect 10525 2772 10577 2823
rect 10614 2837 10663 2883
rect 10614 2803 10622 2837
rect 10656 2803 10663 2837
rect 10614 2738 10663 2803
rect 10697 2873 10701 2907
rect 10735 2873 10749 2907
rect 10869 2909 10880 2917
rect 10914 2920 11052 2943
rect 10914 2909 10921 2920
rect 10697 2857 10749 2873
rect 10697 2823 10708 2857
rect 10742 2823 10749 2857
rect 10697 2772 10749 2823
rect 10786 2837 10835 2883
rect 10786 2803 10794 2837
rect 10828 2803 10835 2837
rect 10786 2738 10835 2803
rect 10869 2857 10921 2909
rect 11043 2909 11052 2920
rect 11086 2920 11189 2943
rect 11425 2935 11483 2970
rect 11086 2909 11101 2920
rect 10869 2823 10880 2857
rect 10914 2823 10921 2857
rect 10869 2772 10921 2823
rect 10958 2837 11009 2883
rect 10958 2803 10966 2837
rect 11000 2803 11009 2837
rect 10958 2738 11009 2803
rect 11043 2857 11101 2909
rect 11425 2901 11437 2935
rect 11471 2901 11483 2935
rect 11043 2823 11052 2857
rect 11086 2823 11101 2857
rect 11043 2772 11101 2823
rect 11135 2837 11189 2886
rect 11135 2803 11138 2837
rect 11172 2803 11189 2837
rect 9754 2737 11009 2738
rect 11135 2737 11189 2803
rect 11425 2842 11483 2901
rect 11425 2808 11437 2842
rect 11471 2808 11483 2842
rect 11425 2737 11483 2808
rect 11702 2917 11753 2975
rect 11702 2907 11719 2917
rect 11702 2873 11713 2907
rect 11747 2873 11753 2883
rect 11702 2849 11753 2873
rect 11702 2815 11719 2849
rect 11702 2799 11753 2815
rect 11787 2881 11848 2965
rect 11787 2847 11803 2881
rect 11837 2847 11848 2881
rect 11892 2881 11926 2999
rect 11995 2983 12103 3014
rect 12217 3001 12251 3157
rect 12170 2967 12251 3001
rect 12285 3059 12355 3123
rect 12285 3043 12293 3059
rect 12327 3025 12355 3059
rect 12319 3009 12355 3025
rect 12285 2999 12355 3009
rect 12389 3107 12431 3123
rect 12423 3073 12431 3107
rect 12170 2949 12204 2967
rect 12389 2965 12431 3073
rect 11960 2915 11976 2949
rect 12010 2915 12204 2949
rect 12296 2933 12431 2965
rect 11892 2847 12052 2881
rect 11787 2813 11848 2847
rect 12018 2839 12052 2847
rect 11787 2779 11803 2813
rect 11837 2779 11848 2813
rect 11787 2737 11848 2779
rect 11916 2779 11932 2813
rect 11966 2779 11982 2813
rect 12170 2839 12204 2915
rect 12238 2899 12254 2933
rect 12288 2931 12431 2933
rect 12469 3097 12521 3175
rect 12563 3205 12629 3247
rect 12563 3171 12579 3205
rect 12613 3171 12629 3205
rect 13149 3209 13215 3247
rect 12563 3155 12629 3171
rect 12804 3169 12925 3203
rect 12959 3169 12975 3203
rect 13016 3169 13032 3203
rect 13066 3169 13115 3203
rect 13149 3175 13165 3209
rect 13199 3175 13215 3209
rect 13355 3205 13421 3247
rect 13287 3179 13321 3195
rect 12469 2959 12503 3097
rect 12605 3095 12657 3111
rect 12537 3047 12571 3063
rect 12605 3061 12633 3095
rect 12691 3077 12729 3111
rect 12667 3061 12763 3077
rect 12804 3027 12838 3169
rect 12872 3101 12943 3111
rect 12872 3067 12888 3101
rect 12922 3067 12943 3101
rect 12571 3013 12875 3027
rect 12537 2993 12875 3013
rect 12288 2907 12330 2931
rect 12238 2873 12285 2899
rect 12319 2873 12330 2907
rect 12469 2925 12719 2959
rect 12753 2925 12769 2959
rect 12469 2897 12503 2925
rect 12391 2863 12503 2897
rect 12018 2789 12052 2805
rect 12086 2813 12136 2829
rect 11916 2737 11982 2779
rect 12086 2779 12102 2813
rect 12086 2737 12136 2779
rect 12170 2814 12344 2839
rect 12170 2780 12294 2814
rect 12328 2780 12344 2814
rect 12170 2771 12344 2780
rect 12391 2821 12425 2863
rect 12592 2857 12807 2891
rect 12592 2839 12626 2857
rect 12391 2771 12425 2787
rect 12459 2813 12533 2829
rect 12459 2779 12479 2813
rect 12513 2779 12533 2813
rect 12773 2839 12807 2857
rect 12592 2789 12626 2805
rect 12660 2789 12676 2823
rect 12710 2789 12726 2823
rect 12773 2789 12807 2805
rect 12841 2837 12875 2993
rect 12909 2949 12943 3067
rect 12977 3095 13047 3111
rect 12977 3061 12990 3095
rect 13024 3061 13047 3095
rect 12977 3043 13047 3061
rect 12977 3009 13001 3043
rect 13035 3009 13047 3043
rect 12977 2987 13047 3009
rect 12909 2933 13002 2949
rect 12909 2907 12968 2933
rect 12943 2899 12968 2907
rect 12943 2873 13002 2899
rect 13081 2897 13115 3169
rect 13355 3171 13371 3205
rect 13405 3171 13421 3205
rect 13455 3179 13506 3195
rect 13149 3111 13241 3141
rect 13149 3077 13185 3111
rect 13219 3077 13241 3111
rect 13149 2988 13241 3077
rect 13183 2954 13241 2988
rect 13149 2931 13241 2954
rect 12909 2871 13002 2873
rect 13036 2863 13115 2897
rect 13036 2837 13070 2863
rect 12841 2815 12977 2837
rect 12459 2737 12533 2779
rect 12660 2737 12726 2789
rect 12841 2781 12927 2815
rect 12961 2781 12977 2815
rect 12841 2771 12977 2781
rect 13020 2821 13070 2837
rect 13054 2787 13070 2821
rect 13020 2771 13070 2787
rect 13104 2813 13154 2829
rect 13138 2779 13154 2813
rect 13104 2737 13154 2779
rect 13188 2774 13253 2931
rect 13287 2907 13321 3145
rect 13489 3145 13506 3179
rect 13455 3137 13506 3145
rect 13356 3103 13506 3137
rect 13541 3179 13875 3247
rect 13541 3145 13559 3179
rect 13593 3145 13823 3179
rect 13857 3145 13875 3179
rect 13356 3043 13402 3103
rect 13541 3093 13875 3145
rect 13927 3192 13961 3213
rect 14004 3205 14070 3247
rect 14004 3171 14020 3205
rect 14054 3171 14070 3205
rect 14104 3175 14155 3213
rect 13927 3137 13961 3158
rect 14104 3141 14106 3175
rect 14140 3141 14155 3175
rect 13927 3103 14070 3137
rect 13356 3034 13368 3043
rect 13390 3000 13402 3009
rect 13356 2905 13402 3000
rect 13436 3049 13506 3069
rect 13436 3015 13458 3049
rect 13492 3015 13506 3049
rect 13436 2975 13506 3015
rect 13541 3023 13691 3093
rect 13541 2989 13561 3023
rect 13595 2989 13691 3023
rect 13725 3025 13821 3059
rect 13855 3025 13875 3059
rect 13436 2941 13461 2975
rect 13495 2941 13506 2975
rect 13725 2955 13875 3025
rect 13909 3049 13980 3067
rect 13909 3043 13929 3049
rect 13909 3009 13921 3043
rect 13963 3015 13980 3049
rect 13955 3009 13980 3015
rect 13909 2993 13980 3009
rect 14036 3065 14070 3103
rect 14104 3098 14155 3141
rect 14036 3049 14087 3065
rect 14036 3015 14053 3049
rect 14036 2999 14087 3015
rect 14036 2957 14070 2999
rect 13436 2939 13506 2941
rect 13541 2915 13875 2955
rect 13356 2889 13506 2905
rect 13356 2871 13455 2889
rect 13287 2821 13321 2855
rect 13489 2855 13506 2889
rect 13287 2771 13321 2787
rect 13355 2803 13371 2837
rect 13405 2803 13421 2837
rect 13355 2737 13421 2803
rect 13455 2821 13506 2855
rect 13489 2787 13506 2821
rect 13455 2771 13506 2787
rect 13541 2881 13559 2915
rect 13593 2881 13823 2915
rect 13857 2881 13875 2915
rect 13541 2813 13875 2881
rect 13541 2779 13559 2813
rect 13593 2779 13823 2813
rect 13857 2779 13875 2813
rect 13541 2737 13875 2779
rect 13927 2923 14070 2957
rect 14121 2952 14155 3098
rect 14190 3201 14242 3247
rect 14224 3167 14242 3201
rect 14190 3133 14242 3167
rect 14277 3186 15346 3247
rect 14277 3152 14295 3186
rect 14329 3152 15295 3186
rect 15329 3152 15346 3186
rect 14277 3138 15346 3152
rect 15381 3186 16450 3247
rect 15381 3152 15399 3186
rect 15433 3152 16399 3186
rect 16433 3152 16450 3186
rect 15381 3138 16450 3152
rect 16577 3153 16635 3247
rect 14224 3099 14242 3133
rect 14190 3079 14242 3099
rect 14594 3023 14662 3138
rect 14594 2989 14611 3023
rect 14645 2989 14662 3023
rect 14594 2972 14662 2989
rect 14958 3059 15028 3074
rect 14958 3025 14975 3059
rect 15009 3025 15028 3059
rect 13927 2889 13961 2923
rect 14104 2918 14155 2952
rect 13927 2821 13961 2855
rect 13927 2771 13961 2787
rect 14004 2855 14020 2889
rect 14054 2855 14070 2889
rect 14004 2821 14070 2855
rect 14004 2787 14020 2821
rect 14054 2787 14070 2821
rect 14004 2737 14070 2787
rect 14104 2884 14106 2918
rect 14140 2884 14155 2918
rect 14104 2839 14155 2884
rect 14104 2805 14105 2839
rect 14139 2837 14155 2839
rect 14104 2803 14106 2805
rect 14140 2803 14155 2837
rect 14104 2771 14155 2803
rect 14190 2949 14242 2967
rect 14224 2915 14242 2949
rect 14190 2881 14242 2915
rect 14224 2847 14242 2881
rect 14190 2813 14242 2847
rect 14958 2824 15028 3025
rect 15698 3023 15766 3138
rect 16577 3119 16589 3153
rect 16623 3119 16635 3153
rect 16669 3186 17738 3247
rect 16669 3152 16687 3186
rect 16721 3152 17687 3186
rect 17721 3152 17738 3186
rect 16669 3138 17738 3152
rect 17773 3186 18475 3247
rect 17773 3152 17791 3186
rect 17825 3152 18423 3186
rect 18457 3152 18475 3186
rect 16577 3102 16635 3119
rect 15698 2989 15715 3023
rect 15749 2989 15766 3023
rect 15698 2972 15766 2989
rect 16062 3059 16132 3074
rect 16062 3025 16079 3059
rect 16113 3025 16132 3059
rect 16062 2824 16132 3025
rect 16986 3023 17054 3138
rect 17773 3093 18475 3152
rect 18601 3184 18843 3247
rect 18601 3150 18619 3184
rect 18653 3150 18791 3184
rect 18825 3150 18843 3184
rect 18601 3097 18843 3150
rect 16986 2989 17003 3023
rect 17037 2989 17054 3023
rect 16986 2972 17054 2989
rect 17350 3059 17420 3074
rect 17350 3025 17367 3059
rect 17401 3025 17420 3059
rect 16577 2935 16635 2970
rect 16577 2901 16589 2935
rect 16623 2901 16635 2935
rect 16577 2842 16635 2901
rect 14224 2779 14242 2813
rect 14190 2737 14242 2779
rect 14277 2813 15346 2824
rect 14277 2779 14295 2813
rect 14329 2779 15295 2813
rect 15329 2779 15346 2813
rect 14277 2737 15346 2779
rect 15381 2813 16450 2824
rect 15381 2779 15399 2813
rect 15433 2779 16399 2813
rect 16433 2779 16450 2813
rect 15381 2737 16450 2779
rect 16577 2808 16589 2842
rect 16623 2808 16635 2842
rect 17350 2824 17420 3025
rect 17773 3023 18103 3093
rect 17773 2989 17851 3023
rect 17885 2989 17950 3023
rect 17984 2989 18049 3023
rect 18083 2989 18103 3023
rect 18137 3025 18157 3059
rect 18191 3025 18260 3059
rect 18294 3025 18363 3059
rect 18397 3025 18475 3059
rect 18137 2955 18475 3025
rect 17773 2915 18475 2955
rect 17773 2881 17791 2915
rect 17825 2881 18423 2915
rect 18457 2881 18475 2915
rect 16577 2737 16635 2808
rect 16669 2813 17738 2824
rect 16669 2779 16687 2813
rect 16721 2779 17687 2813
rect 17721 2779 17738 2813
rect 16669 2737 17738 2779
rect 17773 2813 18475 2881
rect 17773 2779 17791 2813
rect 17825 2779 18423 2813
rect 18457 2779 18475 2813
rect 17773 2737 18475 2779
rect 18601 3029 18651 3063
rect 18685 3029 18705 3063
rect 18601 2955 18705 3029
rect 18739 3023 18843 3097
rect 18739 2989 18759 3023
rect 18793 2989 18843 3023
rect 18601 2908 18843 2955
rect 18601 2874 18619 2908
rect 18653 2874 18791 2908
rect 18825 2874 18843 2908
rect 18601 2813 18843 2874
rect 18601 2779 18619 2813
rect 18653 2779 18791 2813
rect 18825 2779 18843 2813
rect 18601 2737 18843 2779
rect 1104 2703 1133 2737
rect 1167 2703 1225 2737
rect 1259 2703 1317 2737
rect 1351 2703 1409 2737
rect 1443 2703 1501 2737
rect 1535 2703 1593 2737
rect 1627 2703 1685 2737
rect 1719 2703 1777 2737
rect 1811 2703 1869 2737
rect 1903 2703 1961 2737
rect 1995 2703 2053 2737
rect 2087 2703 2145 2737
rect 2179 2703 2237 2737
rect 2271 2703 2329 2737
rect 2363 2703 2421 2737
rect 2455 2703 2513 2737
rect 2547 2703 2605 2737
rect 2639 2703 2697 2737
rect 2731 2703 2789 2737
rect 2823 2703 2881 2737
rect 2915 2703 2973 2737
rect 3007 2703 3065 2737
rect 3099 2703 3157 2737
rect 3191 2703 3249 2737
rect 3283 2703 3341 2737
rect 3375 2703 3433 2737
rect 3467 2703 3525 2737
rect 3559 2703 3617 2737
rect 3651 2703 3709 2737
rect 3743 2703 3801 2737
rect 3835 2703 3893 2737
rect 3927 2703 3985 2737
rect 4019 2703 4077 2737
rect 4111 2703 4169 2737
rect 4203 2703 4261 2737
rect 4295 2703 4353 2737
rect 4387 2703 4445 2737
rect 4479 2703 4537 2737
rect 4571 2703 4629 2737
rect 4663 2703 4721 2737
rect 4755 2703 4813 2737
rect 4847 2703 4905 2737
rect 4939 2703 4997 2737
rect 5031 2703 5089 2737
rect 5123 2703 5181 2737
rect 5215 2703 5273 2737
rect 5307 2703 5365 2737
rect 5399 2703 5457 2737
rect 5491 2703 5549 2737
rect 5583 2703 5641 2737
rect 5675 2703 5733 2737
rect 5767 2703 5825 2737
rect 5859 2703 5917 2737
rect 5951 2703 6009 2737
rect 6043 2703 6101 2737
rect 6135 2703 6193 2737
rect 6227 2703 6285 2737
rect 6319 2703 6377 2737
rect 6411 2703 6469 2737
rect 6503 2703 6561 2737
rect 6595 2703 6653 2737
rect 6687 2703 6745 2737
rect 6779 2703 6837 2737
rect 6871 2703 6929 2737
rect 6963 2703 7021 2737
rect 7055 2703 7113 2737
rect 7147 2703 7205 2737
rect 7239 2703 7297 2737
rect 7331 2703 7389 2737
rect 7423 2703 7481 2737
rect 7515 2703 7573 2737
rect 7607 2703 7665 2737
rect 7699 2703 7757 2737
rect 7791 2703 7849 2737
rect 7883 2703 7941 2737
rect 7975 2703 8033 2737
rect 8067 2703 8125 2737
rect 8159 2703 8217 2737
rect 8251 2703 8309 2737
rect 8343 2703 8401 2737
rect 8435 2703 8493 2737
rect 8527 2703 8585 2737
rect 8619 2703 8677 2737
rect 8711 2703 8769 2737
rect 8803 2703 8861 2737
rect 8895 2703 8953 2737
rect 8987 2703 9045 2737
rect 9079 2703 9137 2737
rect 9171 2703 9229 2737
rect 9263 2703 9321 2737
rect 9355 2703 9413 2737
rect 9447 2703 9505 2737
rect 9539 2703 9597 2737
rect 9631 2703 9689 2737
rect 9723 2703 9781 2737
rect 9815 2703 9873 2737
rect 9907 2703 9965 2737
rect 9999 2703 10057 2737
rect 10091 2703 10149 2737
rect 10183 2703 10241 2737
rect 10275 2703 10333 2737
rect 10367 2703 10425 2737
rect 10459 2703 10517 2737
rect 10551 2703 10609 2737
rect 10643 2703 10701 2737
rect 10735 2703 10793 2737
rect 10827 2703 10885 2737
rect 10919 2703 10977 2737
rect 11011 2703 11069 2737
rect 11103 2703 11161 2737
rect 11195 2703 11253 2737
rect 11287 2703 11345 2737
rect 11379 2703 11437 2737
rect 11471 2703 11529 2737
rect 11563 2703 11621 2737
rect 11655 2703 11713 2737
rect 11747 2703 11805 2737
rect 11839 2703 11897 2737
rect 11931 2703 11989 2737
rect 12023 2703 12081 2737
rect 12115 2703 12173 2737
rect 12207 2703 12265 2737
rect 12299 2703 12357 2737
rect 12391 2703 12449 2737
rect 12483 2703 12541 2737
rect 12575 2703 12633 2737
rect 12667 2703 12725 2737
rect 12759 2703 12817 2737
rect 12851 2703 12909 2737
rect 12943 2703 13001 2737
rect 13035 2703 13093 2737
rect 13127 2703 13185 2737
rect 13219 2703 13277 2737
rect 13311 2703 13369 2737
rect 13403 2703 13461 2737
rect 13495 2703 13553 2737
rect 13587 2703 13645 2737
rect 13679 2703 13737 2737
rect 13771 2703 13829 2737
rect 13863 2703 13921 2737
rect 13955 2703 14013 2737
rect 14047 2703 14105 2737
rect 14139 2703 14197 2737
rect 14231 2703 14289 2737
rect 14323 2703 14381 2737
rect 14415 2703 14473 2737
rect 14507 2703 14565 2737
rect 14599 2703 14657 2737
rect 14691 2703 14749 2737
rect 14783 2703 14841 2737
rect 14875 2703 14933 2737
rect 14967 2703 15025 2737
rect 15059 2703 15117 2737
rect 15151 2703 15209 2737
rect 15243 2703 15301 2737
rect 15335 2703 15393 2737
rect 15427 2703 15485 2737
rect 15519 2703 15577 2737
rect 15611 2703 15669 2737
rect 15703 2703 15761 2737
rect 15795 2703 15853 2737
rect 15887 2703 15945 2737
rect 15979 2703 16037 2737
rect 16071 2703 16129 2737
rect 16163 2703 16221 2737
rect 16255 2703 16313 2737
rect 16347 2703 16405 2737
rect 16439 2703 16497 2737
rect 16531 2703 16589 2737
rect 16623 2703 16681 2737
rect 16715 2703 16773 2737
rect 16807 2703 16865 2737
rect 16899 2703 16957 2737
rect 16991 2703 17049 2737
rect 17083 2703 17141 2737
rect 17175 2703 17233 2737
rect 17267 2703 17325 2737
rect 17359 2703 17417 2737
rect 17451 2703 17509 2737
rect 17543 2703 17601 2737
rect 17635 2703 17693 2737
rect 17727 2703 17785 2737
rect 17819 2703 17877 2737
rect 17911 2703 17969 2737
rect 18003 2703 18061 2737
rect 18095 2703 18153 2737
rect 18187 2703 18245 2737
rect 18279 2703 18337 2737
rect 18371 2703 18429 2737
rect 18463 2703 18521 2737
rect 18555 2703 18613 2737
rect 18647 2703 18705 2737
rect 18739 2703 18797 2737
rect 18831 2703 18860 2737
rect 1121 2661 1363 2703
rect 1121 2627 1139 2661
rect 1173 2627 1311 2661
rect 1345 2627 1363 2661
rect 1121 2566 1363 2627
rect 1121 2532 1139 2566
rect 1173 2532 1311 2566
rect 1345 2532 1363 2566
rect 1121 2485 1363 2532
rect 1397 2661 1639 2703
rect 1397 2627 1415 2661
rect 1449 2627 1587 2661
rect 1621 2627 1639 2661
rect 1397 2566 1639 2627
rect 1397 2532 1415 2566
rect 1449 2532 1587 2566
rect 1621 2532 1639 2566
rect 1674 2653 1725 2669
rect 1674 2619 1691 2653
rect 1674 2585 1725 2619
rect 1759 2637 1825 2703
rect 1759 2603 1775 2637
rect 1809 2603 1825 2637
rect 1859 2653 1893 2669
rect 1674 2551 1691 2585
rect 1859 2585 1893 2619
rect 1725 2551 1824 2569
rect 1674 2535 1824 2551
rect 1397 2485 1639 2532
rect 1121 2417 1171 2451
rect 1205 2417 1225 2451
rect 1121 2343 1225 2417
rect 1259 2411 1363 2485
rect 1259 2377 1279 2411
rect 1313 2377 1363 2411
rect 1397 2417 1447 2451
rect 1481 2417 1501 2451
rect 1397 2343 1501 2417
rect 1535 2411 1639 2485
rect 1535 2377 1555 2411
rect 1589 2377 1639 2411
rect 1674 2499 1744 2501
rect 1674 2465 1685 2499
rect 1719 2465 1744 2499
rect 1674 2425 1744 2465
rect 1674 2391 1688 2425
rect 1722 2391 1744 2425
rect 1674 2371 1744 2391
rect 1778 2440 1824 2535
rect 1778 2431 1790 2440
rect 1812 2397 1824 2406
rect 1121 2290 1363 2343
rect 1121 2256 1139 2290
rect 1173 2256 1311 2290
rect 1345 2256 1363 2290
rect 1121 2193 1363 2256
rect 1397 2290 1639 2343
rect 1778 2337 1824 2397
rect 1397 2256 1415 2290
rect 1449 2256 1587 2290
rect 1621 2256 1639 2290
rect 1397 2193 1639 2256
rect 1674 2303 1824 2337
rect 1674 2295 1725 2303
rect 1674 2261 1691 2295
rect 1859 2295 1893 2533
rect 1927 2509 1992 2666
rect 2026 2661 2076 2703
rect 2026 2627 2042 2661
rect 2026 2611 2076 2627
rect 2110 2653 2160 2669
rect 2110 2619 2126 2653
rect 2110 2603 2160 2619
rect 2203 2659 2339 2669
rect 2203 2625 2219 2659
rect 2253 2625 2339 2659
rect 2454 2651 2520 2703
rect 2647 2661 2721 2703
rect 2203 2603 2339 2625
rect 2110 2577 2144 2603
rect 2065 2543 2144 2577
rect 2178 2567 2271 2569
rect 1939 2486 2031 2509
rect 1939 2452 1997 2486
rect 1939 2363 2031 2452
rect 1939 2329 1961 2363
rect 1995 2329 2031 2363
rect 1939 2299 2031 2329
rect 1674 2245 1725 2261
rect 1759 2235 1775 2269
rect 1809 2235 1825 2269
rect 2065 2271 2099 2543
rect 2178 2541 2237 2567
rect 2212 2533 2237 2541
rect 2212 2507 2271 2533
rect 2178 2491 2271 2507
rect 2133 2431 2203 2453
rect 2133 2397 2145 2431
rect 2179 2397 2203 2431
rect 2133 2379 2203 2397
rect 2133 2345 2156 2379
rect 2190 2345 2203 2379
rect 2133 2329 2203 2345
rect 2237 2373 2271 2491
rect 2305 2447 2339 2603
rect 2373 2635 2407 2651
rect 2454 2617 2470 2651
rect 2504 2617 2520 2651
rect 2554 2635 2588 2651
rect 2373 2583 2407 2601
rect 2647 2627 2667 2661
rect 2701 2627 2721 2661
rect 2647 2611 2721 2627
rect 2755 2653 2789 2669
rect 2554 2583 2588 2601
rect 2373 2549 2588 2583
rect 2755 2577 2789 2619
rect 2836 2660 3010 2669
rect 2836 2626 2852 2660
rect 2886 2626 3010 2660
rect 2836 2601 3010 2626
rect 3044 2661 3094 2703
rect 3078 2627 3094 2661
rect 3198 2661 3264 2703
rect 3044 2611 3094 2627
rect 3128 2635 3162 2651
rect 2677 2543 2789 2577
rect 2677 2515 2711 2543
rect 2411 2481 2427 2515
rect 2461 2481 2711 2515
rect 2850 2533 2861 2567
rect 2895 2541 2942 2567
rect 2850 2509 2892 2533
rect 2305 2427 2643 2447
rect 2305 2413 2609 2427
rect 2237 2339 2258 2373
rect 2292 2339 2308 2373
rect 2237 2329 2308 2339
rect 2342 2271 2376 2413
rect 2417 2363 2513 2379
rect 2451 2329 2489 2363
rect 2547 2345 2575 2379
rect 2609 2377 2643 2393
rect 2523 2329 2575 2345
rect 2677 2343 2711 2481
rect 1859 2245 1893 2261
rect 1759 2193 1825 2235
rect 1965 2231 1981 2265
rect 2015 2231 2031 2265
rect 2065 2237 2114 2271
rect 2148 2237 2164 2271
rect 2205 2237 2221 2271
rect 2255 2237 2376 2271
rect 2551 2269 2617 2285
rect 1965 2193 2031 2231
rect 2551 2235 2567 2269
rect 2601 2235 2617 2269
rect 2551 2193 2617 2235
rect 2659 2265 2711 2343
rect 2749 2507 2892 2509
rect 2926 2507 2942 2541
rect 2976 2525 3010 2601
rect 3198 2627 3214 2661
rect 3248 2627 3264 2661
rect 3332 2661 3393 2703
rect 3332 2627 3343 2661
rect 3377 2627 3393 2661
rect 3128 2593 3162 2601
rect 3332 2593 3393 2627
rect 3128 2559 3288 2593
rect 2749 2475 2884 2507
rect 2976 2491 3170 2525
rect 3204 2491 3220 2525
rect 2749 2367 2791 2475
rect 2976 2473 3010 2491
rect 2749 2333 2757 2367
rect 2749 2317 2791 2333
rect 2825 2431 2895 2441
rect 2825 2415 2861 2431
rect 2825 2381 2853 2415
rect 2887 2381 2895 2397
rect 2825 2317 2895 2381
rect 2929 2439 3010 2473
rect 2929 2283 2963 2439
rect 3077 2426 3185 2457
rect 3254 2441 3288 2559
rect 3332 2559 3343 2593
rect 3377 2559 3393 2593
rect 3332 2475 3393 2559
rect 3427 2635 3478 2641
rect 3427 2625 3433 2635
rect 3467 2601 3478 2635
rect 3461 2591 3478 2601
rect 3427 2557 3478 2591
rect 3461 2523 3478 2557
rect 3427 2465 3478 2523
rect 3697 2632 3755 2703
rect 3697 2598 3709 2632
rect 3743 2598 3755 2632
rect 3697 2539 3755 2598
rect 3697 2505 3709 2539
rect 3743 2505 3755 2539
rect 3697 2470 3755 2505
rect 3789 2661 4123 2703
rect 3789 2627 3807 2661
rect 3841 2627 4071 2661
rect 4105 2627 4123 2661
rect 3789 2559 4123 2627
rect 3789 2525 3807 2559
rect 3841 2525 4071 2559
rect 4105 2525 4123 2559
rect 4250 2653 4301 2669
rect 4250 2619 4267 2653
rect 4250 2585 4301 2619
rect 4335 2637 4401 2703
rect 4335 2603 4351 2637
rect 4385 2603 4401 2637
rect 4435 2653 4469 2669
rect 4250 2551 4267 2585
rect 4435 2585 4469 2619
rect 4301 2551 4400 2569
rect 4250 2535 4400 2551
rect 3789 2485 4123 2525
rect 3254 2435 3402 2441
rect 3111 2417 3185 2426
rect 2997 2389 3041 2405
rect 3031 2355 3041 2389
rect 3077 2383 3093 2392
rect 3127 2383 3185 2417
rect 2997 2349 3041 2355
rect 3137 2363 3185 2383
rect 2997 2315 3103 2349
rect 2773 2269 2963 2283
rect 2659 2231 2679 2265
rect 2713 2231 2729 2265
rect 2773 2235 2789 2269
rect 2823 2235 2963 2269
rect 2773 2227 2963 2235
rect 2997 2265 3035 2281
rect 2997 2231 3001 2265
rect 3069 2269 3103 2315
rect 3171 2329 3185 2363
rect 3137 2303 3185 2329
rect 3219 2425 3402 2435
rect 3219 2391 3368 2425
rect 3219 2375 3402 2391
rect 3219 2340 3284 2375
rect 3219 2285 3283 2340
rect 3436 2335 3478 2465
rect 3789 2417 3809 2451
rect 3843 2417 3939 2451
rect 3789 2347 3939 2417
rect 3973 2415 4123 2485
rect 3973 2381 4069 2415
rect 4103 2381 4123 2415
rect 4250 2499 4320 2501
rect 4250 2465 4261 2499
rect 4295 2465 4320 2499
rect 4250 2425 4320 2465
rect 4250 2391 4264 2425
rect 4298 2391 4320 2425
rect 4250 2371 4320 2391
rect 4354 2440 4400 2535
rect 4354 2431 4366 2440
rect 4388 2397 4400 2406
rect 3427 2319 3478 2335
rect 3461 2285 3478 2319
rect 3069 2251 3219 2269
rect 3253 2251 3283 2285
rect 3069 2235 3283 2251
rect 3332 2269 3393 2285
rect 3332 2235 3343 2269
rect 3377 2235 3393 2269
rect 2997 2193 3035 2231
rect 3332 2193 3393 2235
rect 3427 2229 3478 2285
rect 3697 2321 3755 2338
rect 3697 2287 3709 2321
rect 3743 2287 3755 2321
rect 3697 2193 3755 2287
rect 3789 2295 4123 2347
rect 4354 2337 4400 2397
rect 3789 2261 3807 2295
rect 3841 2261 4071 2295
rect 4105 2261 4123 2295
rect 3789 2193 4123 2261
rect 4250 2303 4400 2337
rect 4250 2295 4301 2303
rect 4250 2261 4267 2295
rect 4435 2295 4469 2533
rect 4503 2509 4568 2666
rect 4602 2661 4652 2703
rect 4602 2627 4618 2661
rect 4602 2611 4652 2627
rect 4686 2653 4736 2669
rect 4686 2619 4702 2653
rect 4686 2603 4736 2619
rect 4779 2659 4915 2669
rect 4779 2625 4795 2659
rect 4829 2625 4915 2659
rect 5030 2651 5096 2703
rect 5223 2661 5297 2703
rect 4779 2603 4915 2625
rect 4686 2577 4720 2603
rect 4641 2543 4720 2577
rect 4754 2567 4847 2569
rect 4515 2499 4607 2509
rect 4515 2465 4537 2499
rect 4571 2486 4607 2499
rect 4571 2465 4573 2486
rect 4515 2452 4573 2465
rect 4515 2299 4607 2452
rect 4250 2245 4301 2261
rect 4335 2235 4351 2269
rect 4385 2235 4401 2269
rect 4641 2271 4675 2543
rect 4754 2541 4813 2567
rect 4788 2533 4813 2541
rect 4788 2507 4847 2533
rect 4754 2491 4847 2507
rect 4709 2431 4779 2453
rect 4709 2397 4721 2431
rect 4755 2397 4779 2431
rect 4709 2379 4779 2397
rect 4709 2345 4732 2379
rect 4766 2345 4779 2379
rect 4709 2329 4779 2345
rect 4813 2373 4847 2491
rect 4881 2447 4915 2603
rect 4949 2635 4983 2651
rect 5030 2617 5046 2651
rect 5080 2617 5096 2651
rect 5130 2635 5164 2651
rect 4949 2583 4983 2601
rect 5223 2627 5243 2661
rect 5277 2627 5297 2661
rect 5223 2611 5297 2627
rect 5331 2653 5365 2669
rect 5130 2583 5164 2601
rect 4949 2549 5164 2583
rect 5331 2577 5365 2619
rect 5412 2660 5586 2669
rect 5412 2626 5428 2660
rect 5462 2626 5586 2660
rect 5412 2601 5586 2626
rect 5620 2661 5670 2703
rect 5654 2627 5670 2661
rect 5774 2661 5840 2703
rect 5620 2611 5670 2627
rect 5704 2635 5738 2651
rect 5253 2543 5365 2577
rect 5253 2515 5287 2543
rect 4987 2481 5003 2515
rect 5037 2481 5287 2515
rect 5426 2533 5437 2567
rect 5471 2541 5518 2567
rect 5426 2509 5468 2533
rect 4881 2427 5219 2447
rect 4881 2413 5185 2427
rect 4813 2339 4834 2373
rect 4868 2339 4884 2373
rect 4813 2329 4884 2339
rect 4918 2271 4952 2413
rect 4993 2363 5089 2379
rect 5027 2329 5065 2363
rect 5123 2345 5151 2379
rect 5185 2377 5219 2393
rect 5099 2329 5151 2345
rect 5253 2343 5287 2481
rect 4435 2245 4469 2261
rect 4335 2193 4401 2235
rect 4541 2231 4557 2265
rect 4591 2231 4607 2265
rect 4641 2237 4690 2271
rect 4724 2237 4740 2271
rect 4781 2237 4797 2271
rect 4831 2237 4952 2271
rect 5127 2269 5193 2285
rect 4541 2193 4607 2231
rect 5127 2235 5143 2269
rect 5177 2235 5193 2269
rect 5127 2193 5193 2235
rect 5235 2265 5287 2343
rect 5325 2507 5468 2509
rect 5502 2507 5518 2541
rect 5552 2525 5586 2601
rect 5774 2627 5790 2661
rect 5824 2627 5840 2661
rect 5908 2661 5969 2703
rect 5908 2627 5919 2661
rect 5953 2627 5969 2661
rect 5704 2593 5738 2601
rect 5908 2593 5969 2627
rect 5704 2559 5864 2593
rect 5325 2475 5460 2507
rect 5552 2491 5746 2525
rect 5780 2491 5796 2525
rect 5325 2367 5367 2475
rect 5552 2473 5586 2491
rect 5325 2333 5333 2367
rect 5325 2317 5367 2333
rect 5401 2431 5471 2441
rect 5401 2415 5437 2431
rect 5401 2381 5429 2415
rect 5463 2381 5471 2397
rect 5401 2317 5471 2381
rect 5505 2439 5586 2473
rect 5505 2283 5539 2439
rect 5653 2426 5761 2457
rect 5830 2441 5864 2559
rect 5908 2559 5919 2593
rect 5953 2559 5969 2593
rect 5908 2475 5969 2559
rect 6003 2635 6054 2641
rect 6003 2625 6009 2635
rect 6043 2601 6054 2635
rect 6037 2591 6054 2601
rect 6003 2557 6054 2591
rect 6037 2523 6054 2557
rect 6003 2465 6054 2523
rect 6273 2632 6331 2703
rect 6273 2598 6285 2632
rect 6319 2598 6331 2632
rect 6365 2661 7434 2703
rect 6365 2627 6383 2661
rect 6417 2627 7383 2661
rect 7417 2627 7434 2661
rect 6365 2616 7434 2627
rect 7469 2661 8538 2703
rect 7469 2627 7487 2661
rect 7521 2627 8487 2661
rect 8521 2627 8538 2661
rect 7469 2616 8538 2627
rect 8573 2661 8815 2703
rect 8573 2627 8591 2661
rect 8625 2627 8763 2661
rect 8797 2627 8815 2661
rect 6273 2539 6331 2598
rect 6273 2505 6285 2539
rect 6319 2505 6331 2539
rect 6273 2470 6331 2505
rect 5830 2435 5978 2441
rect 5687 2417 5761 2426
rect 5573 2389 5617 2405
rect 5607 2355 5617 2389
rect 5653 2383 5669 2392
rect 5703 2383 5761 2417
rect 5573 2349 5617 2355
rect 5713 2363 5761 2383
rect 5573 2315 5679 2349
rect 5349 2269 5539 2283
rect 5235 2231 5255 2265
rect 5289 2231 5305 2265
rect 5349 2235 5365 2269
rect 5399 2235 5539 2269
rect 5349 2227 5539 2235
rect 5573 2265 5611 2281
rect 5573 2231 5577 2265
rect 5645 2269 5679 2315
rect 5747 2329 5761 2363
rect 5713 2303 5761 2329
rect 5795 2425 5978 2435
rect 5795 2391 5944 2425
rect 5795 2375 5978 2391
rect 5795 2340 5860 2375
rect 5795 2285 5859 2340
rect 6012 2335 6054 2465
rect 6682 2451 6750 2468
rect 6682 2417 6699 2451
rect 6733 2417 6750 2451
rect 6003 2319 6054 2335
rect 6037 2285 6054 2319
rect 5645 2251 5795 2269
rect 5829 2251 5859 2285
rect 5645 2235 5859 2251
rect 5908 2269 5969 2285
rect 5908 2235 5919 2269
rect 5953 2235 5969 2269
rect 5573 2193 5611 2231
rect 5908 2193 5969 2235
rect 6003 2229 6054 2285
rect 6273 2321 6331 2338
rect 6273 2287 6285 2321
rect 6319 2287 6331 2321
rect 6682 2302 6750 2417
rect 7046 2415 7116 2616
rect 7046 2381 7063 2415
rect 7097 2381 7116 2415
rect 7046 2366 7116 2381
rect 7786 2451 7854 2468
rect 7786 2417 7803 2451
rect 7837 2417 7854 2451
rect 7786 2302 7854 2417
rect 8150 2415 8220 2616
rect 8573 2566 8815 2627
rect 8573 2532 8591 2566
rect 8625 2532 8763 2566
rect 8797 2532 8815 2566
rect 8573 2485 8815 2532
rect 8150 2381 8167 2415
rect 8201 2381 8220 2415
rect 8150 2366 8220 2381
rect 8573 2417 8623 2451
rect 8657 2417 8677 2451
rect 8573 2343 8677 2417
rect 8711 2411 8815 2485
rect 8849 2632 8907 2703
rect 9211 2661 9272 2703
rect 8849 2598 8861 2632
rect 8895 2598 8907 2632
rect 8849 2539 8907 2598
rect 8849 2505 8861 2539
rect 8895 2505 8907 2539
rect 8849 2470 8907 2505
rect 9126 2635 9177 2641
rect 9126 2601 9137 2635
rect 9171 2625 9177 2635
rect 9126 2591 9143 2601
rect 9126 2557 9177 2591
rect 9126 2523 9143 2557
rect 8711 2377 8731 2411
rect 8765 2377 8815 2411
rect 9126 2465 9177 2523
rect 9211 2627 9227 2661
rect 9261 2627 9272 2661
rect 9340 2661 9406 2703
rect 9340 2627 9356 2661
rect 9390 2627 9406 2661
rect 9510 2661 9560 2703
rect 9442 2635 9476 2651
rect 9211 2593 9272 2627
rect 9510 2627 9526 2661
rect 9510 2611 9560 2627
rect 9594 2660 9768 2669
rect 9594 2626 9718 2660
rect 9752 2626 9768 2660
rect 9442 2593 9476 2601
rect 9211 2559 9227 2593
rect 9261 2559 9272 2593
rect 9211 2475 9272 2559
rect 9316 2559 9476 2593
rect 9594 2601 9768 2626
rect 9815 2653 9849 2669
rect 6273 2193 6331 2287
rect 6365 2288 7434 2302
rect 6365 2254 6383 2288
rect 6417 2254 7383 2288
rect 7417 2254 7434 2288
rect 6365 2193 7434 2254
rect 7469 2288 8538 2302
rect 7469 2254 7487 2288
rect 7521 2254 8487 2288
rect 8521 2254 8538 2288
rect 7469 2193 8538 2254
rect 8573 2290 8815 2343
rect 8573 2256 8591 2290
rect 8625 2256 8763 2290
rect 8797 2256 8815 2290
rect 8573 2193 8815 2256
rect 8849 2321 8907 2338
rect 8849 2287 8861 2321
rect 8895 2287 8907 2321
rect 8849 2193 8907 2287
rect 9126 2335 9168 2465
rect 9316 2441 9350 2559
rect 9594 2525 9628 2601
rect 9815 2577 9849 2619
rect 9883 2661 9957 2703
rect 9883 2627 9903 2661
rect 9937 2627 9957 2661
rect 10084 2651 10150 2703
rect 10265 2659 10401 2669
rect 9883 2611 9957 2627
rect 10016 2635 10050 2651
rect 10084 2617 10100 2651
rect 10134 2617 10150 2651
rect 10197 2635 10231 2651
rect 10016 2583 10050 2601
rect 10197 2583 10231 2601
rect 9384 2491 9400 2525
rect 9434 2491 9628 2525
rect 9662 2541 9709 2567
rect 9662 2507 9678 2541
rect 9743 2533 9754 2567
rect 9815 2543 9927 2577
rect 10016 2549 10231 2583
rect 10265 2625 10351 2659
rect 10385 2625 10401 2659
rect 10265 2603 10401 2625
rect 10444 2653 10494 2669
rect 10478 2619 10494 2653
rect 10444 2603 10494 2619
rect 10528 2661 10578 2703
rect 10562 2627 10578 2661
rect 10528 2611 10578 2627
rect 9712 2509 9754 2533
rect 9893 2515 9927 2543
rect 9712 2507 9855 2509
rect 9594 2473 9628 2491
rect 9720 2475 9855 2507
rect 9202 2435 9350 2441
rect 9202 2425 9385 2435
rect 9236 2391 9385 2425
rect 9202 2375 9385 2391
rect 9320 2340 9385 2375
rect 9126 2319 9177 2335
rect 9126 2285 9143 2319
rect 9321 2285 9385 2340
rect 9419 2426 9527 2457
rect 9594 2439 9675 2473
rect 9419 2417 9493 2426
rect 9419 2383 9477 2417
rect 9511 2383 9527 2392
rect 9563 2389 9607 2405
rect 9419 2363 9467 2383
rect 9419 2329 9433 2363
rect 9563 2355 9573 2389
rect 9563 2349 9607 2355
rect 9419 2303 9467 2329
rect 9501 2315 9607 2349
rect 9126 2229 9177 2285
rect 9211 2269 9272 2285
rect 9211 2235 9227 2269
rect 9261 2235 9272 2269
rect 9321 2251 9351 2285
rect 9501 2269 9535 2315
rect 9641 2283 9675 2439
rect 9709 2431 9779 2441
rect 9743 2415 9779 2431
rect 9709 2381 9717 2397
rect 9751 2381 9779 2415
rect 9709 2317 9779 2381
rect 9813 2367 9855 2475
rect 9847 2333 9855 2367
rect 9813 2317 9855 2333
rect 9893 2481 10143 2515
rect 10177 2481 10193 2515
rect 9893 2343 9927 2481
rect 10265 2447 10299 2603
rect 10460 2577 10494 2603
rect 9961 2427 10299 2447
rect 9995 2413 10299 2427
rect 10333 2567 10426 2569
rect 10367 2541 10426 2567
rect 10460 2543 10539 2577
rect 10367 2533 10392 2541
rect 10333 2507 10392 2533
rect 10333 2491 10426 2507
rect 9961 2377 9995 2393
rect 10029 2345 10057 2379
rect 10091 2363 10187 2379
rect 9385 2251 9535 2269
rect 9321 2235 9535 2251
rect 9569 2265 9607 2281
rect 9211 2193 9272 2235
rect 9603 2231 9607 2265
rect 9569 2193 9607 2231
rect 9641 2269 9831 2283
rect 9641 2235 9781 2269
rect 9815 2235 9831 2269
rect 9893 2265 9945 2343
rect 10029 2329 10081 2345
rect 10115 2329 10153 2363
rect 9641 2227 9831 2235
rect 9875 2231 9891 2265
rect 9925 2231 9945 2265
rect 9987 2269 10053 2285
rect 9987 2235 10003 2269
rect 10037 2235 10053 2269
rect 10228 2271 10262 2413
rect 10333 2373 10367 2491
rect 10296 2339 10312 2373
rect 10346 2339 10367 2373
rect 10296 2329 10367 2339
rect 10401 2431 10471 2453
rect 10401 2397 10425 2431
rect 10459 2397 10471 2431
rect 10401 2379 10471 2397
rect 10401 2345 10414 2379
rect 10448 2345 10471 2379
rect 10401 2329 10471 2345
rect 10505 2271 10539 2543
rect 10612 2509 10677 2666
rect 10711 2653 10745 2669
rect 10711 2585 10745 2619
rect 10779 2637 10845 2703
rect 10779 2603 10795 2637
rect 10829 2603 10845 2637
rect 10879 2653 10930 2669
rect 10913 2619 10930 2653
rect 10879 2585 10930 2619
rect 10573 2499 10665 2509
rect 10573 2486 10609 2499
rect 10607 2465 10609 2486
rect 10643 2465 10665 2499
rect 10607 2452 10665 2465
rect 10573 2299 10665 2452
rect 10228 2237 10349 2271
rect 10383 2237 10399 2271
rect 10440 2237 10456 2271
rect 10490 2237 10539 2271
rect 10711 2295 10745 2533
rect 10780 2551 10879 2569
rect 10913 2551 10930 2585
rect 10780 2535 10930 2551
rect 10965 2661 11299 2703
rect 10965 2627 10983 2661
rect 11017 2627 11247 2661
rect 11281 2627 11299 2661
rect 10965 2559 11299 2627
rect 10780 2440 10826 2535
rect 10965 2525 10983 2559
rect 11017 2525 11247 2559
rect 11281 2525 11299 2559
rect 10814 2431 10826 2440
rect 10780 2397 10792 2406
rect 10780 2337 10826 2397
rect 10860 2431 10930 2501
rect 10965 2485 11299 2525
rect 10860 2425 10885 2431
rect 10860 2391 10882 2425
rect 10919 2397 10930 2431
rect 10916 2391 10930 2397
rect 10860 2371 10930 2391
rect 10965 2417 10985 2451
rect 11019 2417 11115 2451
rect 10965 2347 11115 2417
rect 11149 2415 11299 2485
rect 11425 2632 11483 2703
rect 11425 2598 11437 2632
rect 11471 2598 11483 2632
rect 11425 2539 11483 2598
rect 11425 2505 11437 2539
rect 11471 2505 11483 2539
rect 11425 2470 11483 2505
rect 11517 2661 11851 2703
rect 11517 2627 11535 2661
rect 11569 2627 11799 2661
rect 11833 2627 11851 2661
rect 12063 2661 12124 2703
rect 11517 2559 11851 2627
rect 11517 2525 11535 2559
rect 11569 2525 11799 2559
rect 11833 2525 11851 2559
rect 11517 2485 11851 2525
rect 11149 2381 11245 2415
rect 11279 2381 11299 2415
rect 11517 2417 11537 2451
rect 11571 2417 11667 2451
rect 11517 2347 11667 2417
rect 11701 2415 11851 2485
rect 11701 2381 11797 2415
rect 11831 2381 11851 2415
rect 11978 2625 12029 2641
rect 11978 2591 11995 2625
rect 11978 2567 12029 2591
rect 11978 2533 11989 2567
rect 12023 2557 12029 2567
rect 11978 2523 11995 2533
rect 11978 2465 12029 2523
rect 12063 2627 12079 2661
rect 12113 2627 12124 2661
rect 12192 2661 12258 2703
rect 12192 2627 12208 2661
rect 12242 2627 12258 2661
rect 12362 2661 12412 2703
rect 12294 2635 12328 2651
rect 12063 2593 12124 2627
rect 12362 2627 12378 2661
rect 12362 2611 12412 2627
rect 12446 2660 12620 2669
rect 12446 2626 12570 2660
rect 12604 2626 12620 2660
rect 12294 2593 12328 2601
rect 12063 2559 12079 2593
rect 12113 2559 12124 2593
rect 12063 2475 12124 2559
rect 12168 2559 12328 2593
rect 12446 2601 12620 2626
rect 12667 2653 12701 2669
rect 10780 2303 10930 2337
rect 9987 2193 10053 2235
rect 10573 2231 10589 2265
rect 10623 2231 10639 2265
rect 10879 2295 10930 2303
rect 10711 2245 10745 2261
rect 10573 2193 10639 2231
rect 10779 2235 10795 2269
rect 10829 2235 10845 2269
rect 10913 2261 10930 2295
rect 10879 2245 10930 2261
rect 10965 2295 11299 2347
rect 10965 2261 10983 2295
rect 11017 2261 11247 2295
rect 11281 2261 11299 2295
rect 10779 2193 10845 2235
rect 10965 2193 11299 2261
rect 11425 2321 11483 2338
rect 11425 2287 11437 2321
rect 11471 2287 11483 2321
rect 11425 2193 11483 2287
rect 11517 2295 11851 2347
rect 11517 2261 11535 2295
rect 11569 2261 11799 2295
rect 11833 2261 11851 2295
rect 11517 2193 11851 2261
rect 11978 2335 12020 2465
rect 12168 2441 12202 2559
rect 12446 2525 12480 2601
rect 12667 2577 12701 2619
rect 12735 2661 12809 2703
rect 12735 2627 12755 2661
rect 12789 2627 12809 2661
rect 12936 2651 13002 2703
rect 13117 2659 13253 2669
rect 12735 2611 12809 2627
rect 12868 2635 12902 2651
rect 12936 2617 12952 2651
rect 12986 2617 13002 2651
rect 13049 2635 13083 2651
rect 12868 2583 12902 2601
rect 13049 2583 13083 2601
rect 12236 2491 12252 2525
rect 12286 2491 12480 2525
rect 12514 2541 12561 2567
rect 12514 2507 12530 2541
rect 12595 2533 12606 2567
rect 12667 2543 12779 2577
rect 12868 2549 13083 2583
rect 13117 2625 13203 2659
rect 13237 2625 13253 2659
rect 13117 2603 13253 2625
rect 13296 2653 13346 2669
rect 13330 2619 13346 2653
rect 13296 2603 13346 2619
rect 13380 2661 13430 2703
rect 13414 2627 13430 2661
rect 13380 2611 13430 2627
rect 12564 2509 12606 2533
rect 12745 2515 12779 2543
rect 12564 2507 12707 2509
rect 12446 2473 12480 2491
rect 12572 2475 12707 2507
rect 12054 2435 12202 2441
rect 12054 2425 12237 2435
rect 12088 2391 12237 2425
rect 12054 2375 12237 2391
rect 12172 2340 12237 2375
rect 11978 2319 12029 2335
rect 11978 2285 11995 2319
rect 12173 2285 12237 2340
rect 12271 2426 12379 2457
rect 12446 2439 12527 2473
rect 12271 2417 12345 2426
rect 12271 2383 12329 2417
rect 12363 2383 12379 2392
rect 12415 2389 12459 2405
rect 12271 2363 12319 2383
rect 12271 2329 12285 2363
rect 12415 2355 12425 2389
rect 12415 2349 12459 2355
rect 12271 2303 12319 2329
rect 12353 2315 12459 2349
rect 11978 2229 12029 2285
rect 12063 2269 12124 2285
rect 12063 2235 12079 2269
rect 12113 2235 12124 2269
rect 12173 2251 12203 2285
rect 12353 2269 12387 2315
rect 12493 2283 12527 2439
rect 12561 2431 12631 2441
rect 12595 2415 12631 2431
rect 12561 2381 12569 2397
rect 12603 2381 12631 2415
rect 12561 2317 12631 2381
rect 12665 2367 12707 2475
rect 12699 2333 12707 2367
rect 12665 2317 12707 2333
rect 12745 2481 12995 2515
rect 13029 2481 13045 2515
rect 12745 2343 12779 2481
rect 13117 2447 13151 2603
rect 13312 2577 13346 2603
rect 12813 2427 13151 2447
rect 12847 2413 13151 2427
rect 13185 2567 13278 2569
rect 13219 2541 13278 2567
rect 13312 2543 13391 2577
rect 13219 2533 13244 2541
rect 13185 2507 13244 2533
rect 13185 2491 13278 2507
rect 12813 2377 12847 2393
rect 12881 2345 12909 2379
rect 12943 2363 13039 2379
rect 12237 2251 12387 2269
rect 12173 2235 12387 2251
rect 12421 2265 12459 2281
rect 12063 2193 12124 2235
rect 12455 2231 12459 2265
rect 12421 2193 12459 2231
rect 12493 2269 12683 2283
rect 12493 2235 12633 2269
rect 12667 2235 12683 2269
rect 12745 2265 12797 2343
rect 12881 2329 12933 2345
rect 12967 2329 13005 2363
rect 12493 2227 12683 2235
rect 12727 2231 12743 2265
rect 12777 2231 12797 2265
rect 12839 2269 12905 2285
rect 12839 2235 12855 2269
rect 12889 2235 12905 2269
rect 13080 2271 13114 2413
rect 13185 2373 13219 2491
rect 13148 2339 13164 2373
rect 13198 2339 13219 2373
rect 13148 2329 13219 2339
rect 13253 2431 13323 2453
rect 13253 2397 13277 2431
rect 13311 2397 13323 2431
rect 13253 2379 13323 2397
rect 13253 2345 13266 2379
rect 13300 2345 13323 2379
rect 13253 2329 13323 2345
rect 13357 2271 13391 2543
rect 13464 2509 13529 2666
rect 13563 2653 13597 2669
rect 13563 2585 13597 2619
rect 13631 2637 13697 2703
rect 13631 2603 13647 2637
rect 13681 2603 13697 2637
rect 13731 2653 13782 2669
rect 13765 2619 13782 2653
rect 13731 2585 13782 2619
rect 13425 2499 13517 2509
rect 13425 2486 13461 2499
rect 13459 2465 13461 2486
rect 13495 2465 13517 2499
rect 13459 2452 13517 2465
rect 13425 2299 13517 2452
rect 13080 2237 13201 2271
rect 13235 2237 13251 2271
rect 13292 2237 13308 2271
rect 13342 2237 13391 2271
rect 13563 2295 13597 2533
rect 13632 2551 13731 2569
rect 13765 2551 13782 2585
rect 13632 2535 13782 2551
rect 14001 2632 14059 2703
rect 14363 2661 14424 2703
rect 14001 2598 14013 2632
rect 14047 2598 14059 2632
rect 14001 2539 14059 2598
rect 13632 2440 13678 2535
rect 14001 2505 14013 2539
rect 14047 2505 14059 2539
rect 13666 2431 13678 2440
rect 13632 2397 13644 2406
rect 13632 2337 13678 2397
rect 13712 2499 13782 2501
rect 13712 2465 13737 2499
rect 13771 2465 13782 2499
rect 14001 2470 14059 2505
rect 14278 2635 14329 2641
rect 14278 2601 14289 2635
rect 14323 2625 14329 2635
rect 14278 2591 14295 2601
rect 14278 2557 14329 2591
rect 14278 2523 14295 2557
rect 13712 2425 13782 2465
rect 13712 2391 13734 2425
rect 13768 2391 13782 2425
rect 13712 2371 13782 2391
rect 14278 2465 14329 2523
rect 14363 2627 14379 2661
rect 14413 2627 14424 2661
rect 14492 2661 14558 2703
rect 14492 2627 14508 2661
rect 14542 2627 14558 2661
rect 14662 2661 14712 2703
rect 14594 2635 14628 2651
rect 14363 2593 14424 2627
rect 14662 2627 14678 2661
rect 14662 2611 14712 2627
rect 14746 2660 14920 2669
rect 14746 2626 14870 2660
rect 14904 2626 14920 2660
rect 14594 2593 14628 2601
rect 14363 2559 14379 2593
rect 14413 2559 14424 2593
rect 14363 2475 14424 2559
rect 14468 2559 14628 2593
rect 14746 2601 14920 2626
rect 14967 2653 15001 2669
rect 13632 2303 13782 2337
rect 12839 2193 12905 2235
rect 13425 2231 13441 2265
rect 13475 2231 13491 2265
rect 13731 2295 13782 2303
rect 13563 2245 13597 2261
rect 13425 2193 13491 2231
rect 13631 2235 13647 2269
rect 13681 2235 13697 2269
rect 13765 2261 13782 2295
rect 13731 2245 13782 2261
rect 14001 2321 14059 2338
rect 14001 2287 14013 2321
rect 14047 2287 14059 2321
rect 13631 2193 13697 2235
rect 14001 2193 14059 2287
rect 14278 2335 14320 2465
rect 14468 2441 14502 2559
rect 14746 2525 14780 2601
rect 14967 2577 15001 2619
rect 15035 2661 15109 2703
rect 15035 2627 15055 2661
rect 15089 2627 15109 2661
rect 15236 2651 15302 2703
rect 15417 2659 15553 2669
rect 15035 2611 15109 2627
rect 15168 2635 15202 2651
rect 15236 2617 15252 2651
rect 15286 2617 15302 2651
rect 15349 2635 15383 2651
rect 15168 2583 15202 2601
rect 15349 2583 15383 2601
rect 14536 2491 14552 2525
rect 14586 2491 14780 2525
rect 14814 2541 14861 2567
rect 14814 2507 14830 2541
rect 14895 2533 14906 2567
rect 14967 2543 15079 2577
rect 15168 2549 15383 2583
rect 15417 2625 15503 2659
rect 15537 2625 15553 2659
rect 15417 2603 15553 2625
rect 15596 2653 15646 2669
rect 15630 2619 15646 2653
rect 15596 2603 15646 2619
rect 15680 2661 15730 2703
rect 15714 2627 15730 2661
rect 15680 2611 15730 2627
rect 14864 2509 14906 2533
rect 15045 2515 15079 2543
rect 14864 2507 15007 2509
rect 14746 2473 14780 2491
rect 14872 2475 15007 2507
rect 14354 2435 14502 2441
rect 14354 2425 14537 2435
rect 14388 2391 14537 2425
rect 14354 2375 14537 2391
rect 14472 2340 14537 2375
rect 14278 2319 14329 2335
rect 14278 2285 14295 2319
rect 14473 2285 14537 2340
rect 14571 2426 14679 2457
rect 14746 2439 14827 2473
rect 14571 2417 14645 2426
rect 14571 2383 14629 2417
rect 14663 2383 14679 2392
rect 14715 2389 14759 2405
rect 14571 2363 14619 2383
rect 14571 2329 14585 2363
rect 14715 2355 14725 2389
rect 14715 2349 14759 2355
rect 14571 2303 14619 2329
rect 14653 2315 14759 2349
rect 14278 2229 14329 2285
rect 14363 2269 14424 2285
rect 14363 2235 14379 2269
rect 14413 2235 14424 2269
rect 14473 2251 14503 2285
rect 14653 2269 14687 2315
rect 14793 2283 14827 2439
rect 14861 2431 14931 2441
rect 14895 2415 14931 2431
rect 14861 2381 14869 2397
rect 14903 2381 14931 2415
rect 14861 2317 14931 2381
rect 14965 2367 15007 2475
rect 14999 2333 15007 2367
rect 14965 2317 15007 2333
rect 15045 2481 15295 2515
rect 15329 2481 15345 2515
rect 15045 2343 15079 2481
rect 15417 2447 15451 2603
rect 15612 2577 15646 2603
rect 15113 2427 15451 2447
rect 15147 2413 15451 2427
rect 15485 2567 15578 2569
rect 15519 2541 15578 2567
rect 15612 2543 15691 2577
rect 15519 2533 15544 2541
rect 15485 2507 15544 2533
rect 15485 2491 15578 2507
rect 15113 2377 15147 2393
rect 15181 2345 15209 2379
rect 15243 2363 15339 2379
rect 14537 2251 14687 2269
rect 14473 2235 14687 2251
rect 14721 2265 14759 2281
rect 14363 2193 14424 2235
rect 14755 2231 14759 2265
rect 14721 2193 14759 2231
rect 14793 2269 14983 2283
rect 14793 2235 14933 2269
rect 14967 2235 14983 2269
rect 15045 2265 15097 2343
rect 15181 2329 15233 2345
rect 15267 2329 15305 2363
rect 14793 2227 14983 2235
rect 15027 2231 15043 2265
rect 15077 2231 15097 2265
rect 15139 2269 15205 2285
rect 15139 2235 15155 2269
rect 15189 2235 15205 2269
rect 15380 2271 15414 2413
rect 15485 2373 15519 2491
rect 15448 2339 15464 2373
rect 15498 2339 15519 2373
rect 15448 2329 15519 2339
rect 15553 2431 15623 2453
rect 15553 2397 15577 2431
rect 15611 2397 15623 2431
rect 15553 2379 15623 2397
rect 15553 2345 15566 2379
rect 15600 2345 15623 2379
rect 15553 2329 15623 2345
rect 15657 2271 15691 2543
rect 15764 2509 15829 2666
rect 15863 2653 15897 2669
rect 15863 2585 15897 2619
rect 15931 2637 15997 2703
rect 15931 2603 15947 2637
rect 15981 2603 15997 2637
rect 16031 2653 16082 2669
rect 16065 2619 16082 2653
rect 16031 2585 16082 2619
rect 15725 2486 15817 2509
rect 15759 2452 15817 2486
rect 15725 2363 15817 2452
rect 15725 2329 15761 2363
rect 15795 2329 15817 2363
rect 15725 2299 15817 2329
rect 15380 2237 15501 2271
rect 15535 2237 15551 2271
rect 15592 2237 15608 2271
rect 15642 2237 15691 2271
rect 15863 2295 15897 2533
rect 15932 2551 16031 2569
rect 16065 2551 16082 2585
rect 15932 2535 16082 2551
rect 16117 2661 16451 2703
rect 16117 2627 16135 2661
rect 16169 2627 16399 2661
rect 16433 2627 16451 2661
rect 16117 2559 16451 2627
rect 15932 2440 15978 2535
rect 16117 2525 16135 2559
rect 16169 2525 16399 2559
rect 16433 2525 16451 2559
rect 15966 2431 15978 2440
rect 15932 2397 15944 2406
rect 15932 2337 15978 2397
rect 16012 2499 16082 2501
rect 16012 2465 16037 2499
rect 16071 2465 16082 2499
rect 16117 2485 16451 2525
rect 16012 2425 16082 2465
rect 16012 2391 16034 2425
rect 16068 2391 16082 2425
rect 16012 2371 16082 2391
rect 16117 2417 16137 2451
rect 16171 2417 16267 2451
rect 16117 2347 16267 2417
rect 16301 2415 16451 2485
rect 16577 2632 16635 2703
rect 16577 2598 16589 2632
rect 16623 2598 16635 2632
rect 16577 2539 16635 2598
rect 16577 2505 16589 2539
rect 16623 2505 16635 2539
rect 16577 2470 16635 2505
rect 16669 2661 17371 2703
rect 16669 2627 16687 2661
rect 16721 2627 17319 2661
rect 17353 2627 17371 2661
rect 16669 2559 17371 2627
rect 16669 2525 16687 2559
rect 16721 2525 17319 2559
rect 17353 2525 17371 2559
rect 16669 2485 17371 2525
rect 16301 2381 16397 2415
rect 16431 2381 16451 2415
rect 16669 2417 16747 2451
rect 16781 2417 16846 2451
rect 16880 2417 16945 2451
rect 16979 2417 16999 2451
rect 16669 2347 16999 2417
rect 17033 2415 17371 2485
rect 17515 2653 17549 2669
rect 17515 2585 17549 2619
rect 17592 2653 17658 2703
rect 17592 2619 17608 2653
rect 17642 2619 17658 2653
rect 17592 2585 17658 2619
rect 17592 2551 17608 2585
rect 17642 2551 17658 2585
rect 17692 2637 17743 2669
rect 17692 2603 17694 2637
rect 17728 2603 17743 2637
rect 17692 2556 17743 2603
rect 17515 2517 17549 2551
rect 17692 2522 17694 2556
rect 17728 2522 17743 2556
rect 17515 2483 17658 2517
rect 17692 2488 17743 2522
rect 17033 2381 17053 2415
rect 17087 2381 17156 2415
rect 17190 2381 17259 2415
rect 17293 2381 17371 2415
rect 17497 2431 17568 2447
rect 17497 2397 17509 2431
rect 17543 2425 17568 2431
rect 17497 2391 17517 2397
rect 17551 2391 17568 2425
rect 17497 2373 17568 2391
rect 17624 2441 17658 2483
rect 17624 2425 17675 2441
rect 17624 2391 17641 2425
rect 17624 2375 17675 2391
rect 15932 2303 16082 2337
rect 15139 2193 15205 2235
rect 15725 2231 15741 2265
rect 15775 2231 15791 2265
rect 16031 2295 16082 2303
rect 15863 2245 15897 2261
rect 15725 2193 15791 2231
rect 15931 2235 15947 2269
rect 15981 2235 15997 2269
rect 16065 2261 16082 2295
rect 16031 2245 16082 2261
rect 16117 2295 16451 2347
rect 16117 2261 16135 2295
rect 16169 2261 16399 2295
rect 16433 2261 16451 2295
rect 15931 2193 15997 2235
rect 16117 2193 16451 2261
rect 16577 2321 16635 2338
rect 16577 2287 16589 2321
rect 16623 2287 16635 2321
rect 16577 2193 16635 2287
rect 16669 2288 17371 2347
rect 17624 2337 17658 2375
rect 17709 2342 17743 2488
rect 17778 2661 17830 2703
rect 17812 2627 17830 2661
rect 17778 2593 17830 2627
rect 17812 2559 17830 2593
rect 17778 2525 17830 2559
rect 17812 2491 17830 2525
rect 17778 2473 17830 2491
rect 17865 2661 18567 2703
rect 17865 2627 17883 2661
rect 17917 2627 18515 2661
rect 18549 2627 18567 2661
rect 17865 2559 18567 2627
rect 17865 2525 17883 2559
rect 17917 2525 18515 2559
rect 18549 2525 18567 2559
rect 17865 2485 18567 2525
rect 17865 2417 17943 2451
rect 17977 2417 18042 2451
rect 18076 2417 18141 2451
rect 18175 2417 18195 2451
rect 16669 2254 16687 2288
rect 16721 2254 17319 2288
rect 17353 2254 17371 2288
rect 16669 2193 17371 2254
rect 17515 2303 17658 2337
rect 17515 2282 17549 2303
rect 17692 2299 17743 2342
rect 17692 2295 17694 2299
rect 17515 2227 17549 2248
rect 17592 2235 17608 2269
rect 17642 2235 17658 2269
rect 17592 2193 17658 2235
rect 17692 2261 17693 2295
rect 17728 2265 17743 2299
rect 17727 2261 17743 2265
rect 17692 2227 17743 2261
rect 17778 2341 17830 2361
rect 17812 2307 17830 2341
rect 17778 2273 17830 2307
rect 17812 2239 17830 2273
rect 17778 2193 17830 2239
rect 17865 2347 18195 2417
rect 18229 2415 18567 2485
rect 18229 2381 18249 2415
rect 18283 2381 18352 2415
rect 18386 2381 18455 2415
rect 18489 2381 18567 2415
rect 18601 2661 18843 2703
rect 18601 2627 18619 2661
rect 18653 2627 18791 2661
rect 18825 2627 18843 2661
rect 18601 2566 18843 2627
rect 18601 2532 18619 2566
rect 18653 2532 18791 2566
rect 18825 2532 18843 2566
rect 18601 2485 18843 2532
rect 18601 2411 18705 2485
rect 18601 2377 18651 2411
rect 18685 2377 18705 2411
rect 18739 2417 18759 2451
rect 18793 2417 18843 2451
rect 17865 2288 18567 2347
rect 18739 2343 18843 2417
rect 17865 2254 17883 2288
rect 17917 2254 18515 2288
rect 18549 2254 18567 2288
rect 17865 2193 18567 2254
rect 18601 2290 18843 2343
rect 18601 2256 18619 2290
rect 18653 2256 18791 2290
rect 18825 2256 18843 2290
rect 18601 2193 18843 2256
rect 1104 2159 1133 2193
rect 1167 2159 1225 2193
rect 1259 2159 1317 2193
rect 1351 2159 1409 2193
rect 1443 2159 1501 2193
rect 1535 2159 1593 2193
rect 1627 2159 1685 2193
rect 1719 2159 1777 2193
rect 1811 2159 1869 2193
rect 1903 2159 1961 2193
rect 1995 2159 2053 2193
rect 2087 2159 2145 2193
rect 2179 2159 2237 2193
rect 2271 2159 2329 2193
rect 2363 2159 2421 2193
rect 2455 2159 2513 2193
rect 2547 2159 2605 2193
rect 2639 2159 2697 2193
rect 2731 2159 2789 2193
rect 2823 2159 2881 2193
rect 2915 2159 2973 2193
rect 3007 2159 3065 2193
rect 3099 2159 3157 2193
rect 3191 2159 3249 2193
rect 3283 2159 3341 2193
rect 3375 2159 3433 2193
rect 3467 2159 3525 2193
rect 3559 2159 3617 2193
rect 3651 2159 3709 2193
rect 3743 2159 3801 2193
rect 3835 2159 3893 2193
rect 3927 2159 3985 2193
rect 4019 2159 4077 2193
rect 4111 2159 4169 2193
rect 4203 2159 4261 2193
rect 4295 2159 4353 2193
rect 4387 2159 4445 2193
rect 4479 2159 4537 2193
rect 4571 2159 4629 2193
rect 4663 2159 4721 2193
rect 4755 2159 4813 2193
rect 4847 2159 4905 2193
rect 4939 2159 4997 2193
rect 5031 2159 5089 2193
rect 5123 2159 5181 2193
rect 5215 2159 5273 2193
rect 5307 2159 5365 2193
rect 5399 2159 5457 2193
rect 5491 2159 5549 2193
rect 5583 2159 5641 2193
rect 5675 2159 5733 2193
rect 5767 2159 5825 2193
rect 5859 2159 5917 2193
rect 5951 2159 6009 2193
rect 6043 2159 6101 2193
rect 6135 2159 6193 2193
rect 6227 2159 6285 2193
rect 6319 2159 6377 2193
rect 6411 2159 6469 2193
rect 6503 2159 6561 2193
rect 6595 2159 6653 2193
rect 6687 2159 6745 2193
rect 6779 2159 6837 2193
rect 6871 2159 6929 2193
rect 6963 2159 7021 2193
rect 7055 2159 7113 2193
rect 7147 2159 7205 2193
rect 7239 2159 7297 2193
rect 7331 2159 7389 2193
rect 7423 2159 7481 2193
rect 7515 2159 7573 2193
rect 7607 2159 7665 2193
rect 7699 2159 7757 2193
rect 7791 2159 7849 2193
rect 7883 2159 7941 2193
rect 7975 2159 8033 2193
rect 8067 2159 8125 2193
rect 8159 2159 8217 2193
rect 8251 2159 8309 2193
rect 8343 2159 8401 2193
rect 8435 2159 8493 2193
rect 8527 2159 8585 2193
rect 8619 2159 8677 2193
rect 8711 2159 8769 2193
rect 8803 2159 8861 2193
rect 8895 2159 8953 2193
rect 8987 2159 9045 2193
rect 9079 2159 9137 2193
rect 9171 2159 9229 2193
rect 9263 2159 9321 2193
rect 9355 2159 9413 2193
rect 9447 2159 9505 2193
rect 9539 2159 9597 2193
rect 9631 2159 9689 2193
rect 9723 2159 9781 2193
rect 9815 2159 9873 2193
rect 9907 2159 9965 2193
rect 9999 2159 10057 2193
rect 10091 2159 10149 2193
rect 10183 2159 10241 2193
rect 10275 2159 10333 2193
rect 10367 2159 10425 2193
rect 10459 2159 10517 2193
rect 10551 2159 10609 2193
rect 10643 2159 10701 2193
rect 10735 2159 10793 2193
rect 10827 2159 10885 2193
rect 10919 2159 10977 2193
rect 11011 2159 11069 2193
rect 11103 2159 11161 2193
rect 11195 2159 11253 2193
rect 11287 2159 11345 2193
rect 11379 2159 11437 2193
rect 11471 2159 11529 2193
rect 11563 2159 11621 2193
rect 11655 2159 11713 2193
rect 11747 2159 11805 2193
rect 11839 2159 11897 2193
rect 11931 2159 11989 2193
rect 12023 2159 12081 2193
rect 12115 2159 12173 2193
rect 12207 2159 12265 2193
rect 12299 2159 12357 2193
rect 12391 2159 12449 2193
rect 12483 2159 12541 2193
rect 12575 2159 12633 2193
rect 12667 2159 12725 2193
rect 12759 2159 12817 2193
rect 12851 2159 12909 2193
rect 12943 2159 13001 2193
rect 13035 2159 13093 2193
rect 13127 2159 13185 2193
rect 13219 2159 13277 2193
rect 13311 2159 13369 2193
rect 13403 2159 13461 2193
rect 13495 2159 13553 2193
rect 13587 2159 13645 2193
rect 13679 2159 13737 2193
rect 13771 2159 13829 2193
rect 13863 2159 13921 2193
rect 13955 2159 14013 2193
rect 14047 2159 14105 2193
rect 14139 2159 14197 2193
rect 14231 2159 14289 2193
rect 14323 2159 14381 2193
rect 14415 2159 14473 2193
rect 14507 2159 14565 2193
rect 14599 2159 14657 2193
rect 14691 2159 14749 2193
rect 14783 2159 14841 2193
rect 14875 2159 14933 2193
rect 14967 2159 15025 2193
rect 15059 2159 15117 2193
rect 15151 2159 15209 2193
rect 15243 2159 15301 2193
rect 15335 2159 15393 2193
rect 15427 2159 15485 2193
rect 15519 2159 15577 2193
rect 15611 2159 15669 2193
rect 15703 2159 15761 2193
rect 15795 2159 15853 2193
rect 15887 2159 15945 2193
rect 15979 2159 16037 2193
rect 16071 2159 16129 2193
rect 16163 2159 16221 2193
rect 16255 2159 16313 2193
rect 16347 2159 16405 2193
rect 16439 2159 16497 2193
rect 16531 2159 16589 2193
rect 16623 2159 16681 2193
rect 16715 2159 16773 2193
rect 16807 2159 16865 2193
rect 16899 2159 16957 2193
rect 16991 2159 17049 2193
rect 17083 2159 17141 2193
rect 17175 2159 17233 2193
rect 17267 2159 17325 2193
rect 17359 2159 17417 2193
rect 17451 2159 17509 2193
rect 17543 2159 17601 2193
rect 17635 2159 17693 2193
rect 17727 2159 17785 2193
rect 17819 2159 17877 2193
rect 17911 2159 17969 2193
rect 18003 2159 18061 2193
rect 18095 2159 18153 2193
rect 18187 2159 18245 2193
rect 18279 2159 18337 2193
rect 18371 2159 18429 2193
rect 18463 2159 18521 2193
rect 18555 2159 18613 2193
rect 18647 2159 18705 2193
rect 18739 2159 18797 2193
rect 18831 2159 18860 2193
<< viali >>
rect 1133 7599 1167 7633
rect 1225 7599 1259 7633
rect 1317 7599 1351 7633
rect 1409 7599 1443 7633
rect 1501 7599 1535 7633
rect 1593 7599 1627 7633
rect 1685 7599 1719 7633
rect 1777 7599 1811 7633
rect 1869 7599 1903 7633
rect 1961 7599 1995 7633
rect 2053 7599 2087 7633
rect 2145 7599 2179 7633
rect 2237 7599 2271 7633
rect 2329 7599 2363 7633
rect 2421 7599 2455 7633
rect 2513 7599 2547 7633
rect 2605 7599 2639 7633
rect 2697 7599 2731 7633
rect 2789 7599 2823 7633
rect 2881 7599 2915 7633
rect 2973 7599 3007 7633
rect 3065 7599 3099 7633
rect 3157 7599 3191 7633
rect 3249 7599 3283 7633
rect 3341 7599 3375 7633
rect 3433 7599 3467 7633
rect 3525 7599 3559 7633
rect 3617 7599 3651 7633
rect 3709 7599 3743 7633
rect 3801 7599 3835 7633
rect 3893 7599 3927 7633
rect 3985 7599 4019 7633
rect 4077 7599 4111 7633
rect 4169 7599 4203 7633
rect 4261 7599 4295 7633
rect 4353 7599 4387 7633
rect 4445 7599 4479 7633
rect 4537 7599 4571 7633
rect 4629 7599 4663 7633
rect 4721 7599 4755 7633
rect 4813 7599 4847 7633
rect 4905 7599 4939 7633
rect 4997 7599 5031 7633
rect 5089 7599 5123 7633
rect 5181 7599 5215 7633
rect 5273 7599 5307 7633
rect 5365 7599 5399 7633
rect 5457 7599 5491 7633
rect 5549 7599 5583 7633
rect 5641 7599 5675 7633
rect 5733 7599 5767 7633
rect 5825 7599 5859 7633
rect 5917 7599 5951 7633
rect 6009 7599 6043 7633
rect 6101 7599 6135 7633
rect 6193 7599 6227 7633
rect 6285 7599 6319 7633
rect 6377 7599 6411 7633
rect 6469 7599 6503 7633
rect 6561 7599 6595 7633
rect 6653 7599 6687 7633
rect 6745 7599 6779 7633
rect 6837 7599 6871 7633
rect 6929 7599 6963 7633
rect 7021 7599 7055 7633
rect 7113 7599 7147 7633
rect 7205 7599 7239 7633
rect 7297 7599 7331 7633
rect 7389 7599 7423 7633
rect 7481 7599 7515 7633
rect 7573 7599 7607 7633
rect 7665 7599 7699 7633
rect 7757 7599 7791 7633
rect 7849 7599 7883 7633
rect 7941 7599 7975 7633
rect 8033 7599 8067 7633
rect 8125 7599 8159 7633
rect 8217 7599 8251 7633
rect 8309 7599 8343 7633
rect 8401 7599 8435 7633
rect 8493 7599 8527 7633
rect 8585 7599 8619 7633
rect 8677 7599 8711 7633
rect 8769 7599 8803 7633
rect 8861 7599 8895 7633
rect 8953 7599 8987 7633
rect 9045 7599 9079 7633
rect 9137 7599 9171 7633
rect 9229 7599 9263 7633
rect 9321 7599 9355 7633
rect 9413 7599 9447 7633
rect 9505 7599 9539 7633
rect 9597 7599 9631 7633
rect 9689 7599 9723 7633
rect 9781 7599 9815 7633
rect 9873 7599 9907 7633
rect 9965 7599 9999 7633
rect 10057 7599 10091 7633
rect 10149 7599 10183 7633
rect 10241 7599 10275 7633
rect 10333 7599 10367 7633
rect 10425 7599 10459 7633
rect 10517 7599 10551 7633
rect 10609 7599 10643 7633
rect 10701 7599 10735 7633
rect 10793 7599 10827 7633
rect 10885 7599 10919 7633
rect 10977 7599 11011 7633
rect 11069 7599 11103 7633
rect 11161 7599 11195 7633
rect 11253 7599 11287 7633
rect 11345 7599 11379 7633
rect 11437 7599 11471 7633
rect 11529 7599 11563 7633
rect 11621 7599 11655 7633
rect 11713 7599 11747 7633
rect 11805 7599 11839 7633
rect 11897 7599 11931 7633
rect 11989 7599 12023 7633
rect 12081 7599 12115 7633
rect 12173 7599 12207 7633
rect 12265 7599 12299 7633
rect 12357 7599 12391 7633
rect 12449 7599 12483 7633
rect 12541 7599 12575 7633
rect 12633 7599 12667 7633
rect 12725 7599 12759 7633
rect 12817 7599 12851 7633
rect 12909 7599 12943 7633
rect 13001 7599 13035 7633
rect 13093 7599 13127 7633
rect 13185 7599 13219 7633
rect 13277 7599 13311 7633
rect 13369 7599 13403 7633
rect 13461 7599 13495 7633
rect 13553 7599 13587 7633
rect 13645 7599 13679 7633
rect 13737 7599 13771 7633
rect 13829 7599 13863 7633
rect 13921 7599 13955 7633
rect 14013 7599 14047 7633
rect 14105 7599 14139 7633
rect 14197 7599 14231 7633
rect 14289 7599 14323 7633
rect 14381 7599 14415 7633
rect 14473 7599 14507 7633
rect 14565 7599 14599 7633
rect 14657 7599 14691 7633
rect 14749 7599 14783 7633
rect 14841 7599 14875 7633
rect 14933 7599 14967 7633
rect 15025 7599 15059 7633
rect 15117 7599 15151 7633
rect 15209 7599 15243 7633
rect 15301 7599 15335 7633
rect 15393 7599 15427 7633
rect 15485 7599 15519 7633
rect 15577 7599 15611 7633
rect 15669 7599 15703 7633
rect 15761 7599 15795 7633
rect 15853 7599 15887 7633
rect 15945 7599 15979 7633
rect 16037 7599 16071 7633
rect 16129 7599 16163 7633
rect 16221 7599 16255 7633
rect 16313 7599 16347 7633
rect 16405 7599 16439 7633
rect 16497 7599 16531 7633
rect 16589 7599 16623 7633
rect 16681 7599 16715 7633
rect 16773 7599 16807 7633
rect 16865 7599 16899 7633
rect 16957 7599 16991 7633
rect 17049 7599 17083 7633
rect 17141 7599 17175 7633
rect 17233 7599 17267 7633
rect 17325 7599 17359 7633
rect 17417 7599 17451 7633
rect 17509 7599 17543 7633
rect 17601 7599 17635 7633
rect 17693 7599 17727 7633
rect 17785 7599 17819 7633
rect 17877 7599 17911 7633
rect 17969 7599 18003 7633
rect 18061 7599 18095 7633
rect 18153 7599 18187 7633
rect 18245 7599 18279 7633
rect 18337 7599 18371 7633
rect 18429 7599 18463 7633
rect 18521 7599 18555 7633
rect 18613 7599 18647 7633
rect 18705 7599 18739 7633
rect 18797 7599 18831 7633
rect 1685 7527 1719 7531
rect 1685 7497 1718 7527
rect 1718 7497 1719 7527
rect 1869 7367 1895 7395
rect 1895 7367 1903 7395
rect 1869 7361 1903 7367
rect 4077 7527 4111 7531
rect 4077 7497 4110 7527
rect 4110 7497 4111 7527
rect 4261 7367 4287 7395
rect 4287 7367 4295 7395
rect 4261 7361 4295 7367
rect 5733 7527 5767 7531
rect 5733 7497 5766 7527
rect 5766 7497 5767 7527
rect 5917 7367 5943 7395
rect 5943 7367 5951 7395
rect 5917 7361 5951 7367
rect 7941 7527 7975 7531
rect 7941 7497 7974 7527
rect 7974 7497 7975 7527
rect 9597 7457 9620 7463
rect 9620 7457 9631 7463
rect 8125 7367 8151 7395
rect 8151 7367 8159 7395
rect 8125 7361 8159 7367
rect 9597 7429 9631 7457
rect 10149 7429 10183 7463
rect 12449 7527 12483 7531
rect 12449 7497 12450 7527
rect 12450 7497 12483 7527
rect 10333 7225 10367 7259
rect 12265 7367 12273 7395
rect 12273 7367 12299 7395
rect 12265 7361 12299 7367
rect 14657 7527 14691 7531
rect 14657 7497 14658 7527
rect 14658 7497 14691 7527
rect 14473 7367 14481 7395
rect 14481 7367 14507 7395
rect 14473 7361 14507 7367
rect 17049 7527 17083 7531
rect 17049 7497 17050 7527
rect 17050 7497 17083 7527
rect 16865 7367 16873 7395
rect 16873 7367 16899 7395
rect 16865 7361 16899 7367
rect 18245 7527 18279 7531
rect 18245 7497 18246 7527
rect 18246 7497 18279 7527
rect 18061 7367 18069 7395
rect 18069 7367 18095 7395
rect 18061 7361 18095 7367
rect 1133 7055 1167 7089
rect 1225 7055 1259 7089
rect 1317 7055 1351 7089
rect 1409 7055 1443 7089
rect 1501 7055 1535 7089
rect 1593 7055 1627 7089
rect 1685 7055 1719 7089
rect 1777 7055 1811 7089
rect 1869 7055 1903 7089
rect 1961 7055 1995 7089
rect 2053 7055 2087 7089
rect 2145 7055 2179 7089
rect 2237 7055 2271 7089
rect 2329 7055 2363 7089
rect 2421 7055 2455 7089
rect 2513 7055 2547 7089
rect 2605 7055 2639 7089
rect 2697 7055 2731 7089
rect 2789 7055 2823 7089
rect 2881 7055 2915 7089
rect 2973 7055 3007 7089
rect 3065 7055 3099 7089
rect 3157 7055 3191 7089
rect 3249 7055 3283 7089
rect 3341 7055 3375 7089
rect 3433 7055 3467 7089
rect 3525 7055 3559 7089
rect 3617 7055 3651 7089
rect 3709 7055 3743 7089
rect 3801 7055 3835 7089
rect 3893 7055 3927 7089
rect 3985 7055 4019 7089
rect 4077 7055 4111 7089
rect 4169 7055 4203 7089
rect 4261 7055 4295 7089
rect 4353 7055 4387 7089
rect 4445 7055 4479 7089
rect 4537 7055 4571 7089
rect 4629 7055 4663 7089
rect 4721 7055 4755 7089
rect 4813 7055 4847 7089
rect 4905 7055 4939 7089
rect 4997 7055 5031 7089
rect 5089 7055 5123 7089
rect 5181 7055 5215 7089
rect 5273 7055 5307 7089
rect 5365 7055 5399 7089
rect 5457 7055 5491 7089
rect 5549 7055 5583 7089
rect 5641 7055 5675 7089
rect 5733 7055 5767 7089
rect 5825 7055 5859 7089
rect 5917 7055 5951 7089
rect 6009 7055 6043 7089
rect 6101 7055 6135 7089
rect 6193 7055 6227 7089
rect 6285 7055 6319 7089
rect 6377 7055 6411 7089
rect 6469 7055 6503 7089
rect 6561 7055 6595 7089
rect 6653 7055 6687 7089
rect 6745 7055 6779 7089
rect 6837 7055 6871 7089
rect 6929 7055 6963 7089
rect 7021 7055 7055 7089
rect 7113 7055 7147 7089
rect 7205 7055 7239 7089
rect 7297 7055 7331 7089
rect 7389 7055 7423 7089
rect 7481 7055 7515 7089
rect 7573 7055 7607 7089
rect 7665 7055 7699 7089
rect 7757 7055 7791 7089
rect 7849 7055 7883 7089
rect 7941 7055 7975 7089
rect 8033 7055 8067 7089
rect 8125 7055 8159 7089
rect 8217 7055 8251 7089
rect 8309 7055 8343 7089
rect 8401 7055 8435 7089
rect 8493 7055 8527 7089
rect 8585 7055 8619 7089
rect 8677 7055 8711 7089
rect 8769 7055 8803 7089
rect 8861 7055 8895 7089
rect 8953 7055 8987 7089
rect 9045 7055 9079 7089
rect 9137 7055 9171 7089
rect 9229 7055 9263 7089
rect 9321 7055 9355 7089
rect 9413 7055 9447 7089
rect 9505 7055 9539 7089
rect 9597 7055 9631 7089
rect 9689 7055 9723 7089
rect 9781 7055 9815 7089
rect 9873 7055 9907 7089
rect 9965 7055 9999 7089
rect 10057 7055 10091 7089
rect 10149 7055 10183 7089
rect 10241 7055 10275 7089
rect 10333 7055 10367 7089
rect 10425 7055 10459 7089
rect 10517 7055 10551 7089
rect 10609 7055 10643 7089
rect 10701 7055 10735 7089
rect 10793 7055 10827 7089
rect 10885 7055 10919 7089
rect 10977 7055 11011 7089
rect 11069 7055 11103 7089
rect 11161 7055 11195 7089
rect 11253 7055 11287 7089
rect 11345 7055 11379 7089
rect 11437 7055 11471 7089
rect 11529 7055 11563 7089
rect 11621 7055 11655 7089
rect 11713 7055 11747 7089
rect 11805 7055 11839 7089
rect 11897 7055 11931 7089
rect 11989 7055 12023 7089
rect 12081 7055 12115 7089
rect 12173 7055 12207 7089
rect 12265 7055 12299 7089
rect 12357 7055 12391 7089
rect 12449 7055 12483 7089
rect 12541 7055 12575 7089
rect 12633 7055 12667 7089
rect 12725 7055 12759 7089
rect 12817 7055 12851 7089
rect 12909 7055 12943 7089
rect 13001 7055 13035 7089
rect 13093 7055 13127 7089
rect 13185 7055 13219 7089
rect 13277 7055 13311 7089
rect 13369 7055 13403 7089
rect 13461 7055 13495 7089
rect 13553 7055 13587 7089
rect 13645 7055 13679 7089
rect 13737 7055 13771 7089
rect 13829 7055 13863 7089
rect 13921 7055 13955 7089
rect 14013 7055 14047 7089
rect 14105 7055 14139 7089
rect 14197 7055 14231 7089
rect 14289 7055 14323 7089
rect 14381 7055 14415 7089
rect 14473 7055 14507 7089
rect 14565 7055 14599 7089
rect 14657 7055 14691 7089
rect 14749 7055 14783 7089
rect 14841 7055 14875 7089
rect 14933 7055 14967 7089
rect 15025 7055 15059 7089
rect 15117 7055 15151 7089
rect 15209 7055 15243 7089
rect 15301 7055 15335 7089
rect 15393 7055 15427 7089
rect 15485 7055 15519 7089
rect 15577 7055 15611 7089
rect 15669 7055 15703 7089
rect 15761 7055 15795 7089
rect 15853 7055 15887 7089
rect 15945 7055 15979 7089
rect 16037 7055 16071 7089
rect 16129 7055 16163 7089
rect 16221 7055 16255 7089
rect 16313 7055 16347 7089
rect 16405 7055 16439 7089
rect 16497 7055 16531 7089
rect 16589 7055 16623 7089
rect 16681 7055 16715 7089
rect 16773 7055 16807 7089
rect 16865 7055 16899 7089
rect 16957 7055 16991 7089
rect 17049 7055 17083 7089
rect 17141 7055 17175 7089
rect 17233 7055 17267 7089
rect 17325 7055 17359 7089
rect 17417 7055 17451 7089
rect 17509 7055 17543 7089
rect 17601 7055 17635 7089
rect 17693 7055 17727 7089
rect 17785 7055 17819 7089
rect 17877 7055 17911 7089
rect 17969 7055 18003 7089
rect 18061 7055 18095 7089
rect 18153 7055 18187 7089
rect 18245 7055 18279 7089
rect 18337 7055 18371 7089
rect 18429 7055 18463 7089
rect 18521 7055 18555 7089
rect 18613 7055 18647 7089
rect 18705 7055 18739 7089
rect 18797 7055 18831 7089
rect 1133 6511 1167 6545
rect 1225 6511 1259 6545
rect 1317 6511 1351 6545
rect 1409 6511 1443 6545
rect 1501 6511 1535 6545
rect 1593 6511 1627 6545
rect 1685 6511 1719 6545
rect 1777 6511 1811 6545
rect 1869 6511 1903 6545
rect 1961 6511 1995 6545
rect 2053 6511 2087 6545
rect 2145 6511 2179 6545
rect 2237 6511 2271 6545
rect 2329 6511 2363 6545
rect 2421 6511 2455 6545
rect 2513 6511 2547 6545
rect 2605 6511 2639 6545
rect 2697 6511 2731 6545
rect 2789 6511 2823 6545
rect 2881 6511 2915 6545
rect 2973 6511 3007 6545
rect 3065 6511 3099 6545
rect 3157 6511 3191 6545
rect 3249 6511 3283 6545
rect 3341 6511 3375 6545
rect 3433 6511 3467 6545
rect 3525 6511 3559 6545
rect 3617 6511 3651 6545
rect 3709 6511 3743 6545
rect 3801 6511 3835 6545
rect 3893 6511 3927 6545
rect 3985 6511 4019 6545
rect 4077 6511 4111 6545
rect 4169 6511 4203 6545
rect 4261 6511 4295 6545
rect 4353 6511 4387 6545
rect 4445 6511 4479 6545
rect 4537 6511 4571 6545
rect 4629 6511 4663 6545
rect 4721 6511 4755 6545
rect 4813 6511 4847 6545
rect 4905 6511 4939 6545
rect 4997 6511 5031 6545
rect 5089 6511 5123 6545
rect 5181 6511 5215 6545
rect 5273 6511 5307 6545
rect 5365 6511 5399 6545
rect 5457 6511 5491 6545
rect 5549 6511 5583 6545
rect 5641 6511 5675 6545
rect 5733 6511 5767 6545
rect 5825 6511 5859 6545
rect 5917 6511 5951 6545
rect 6009 6511 6043 6545
rect 6101 6511 6135 6545
rect 6193 6511 6227 6545
rect 6285 6511 6319 6545
rect 6377 6511 6411 6545
rect 6469 6511 6503 6545
rect 6561 6511 6595 6545
rect 6653 6511 6687 6545
rect 6745 6511 6779 6545
rect 6837 6511 6871 6545
rect 6929 6511 6963 6545
rect 7021 6511 7055 6545
rect 7113 6511 7147 6545
rect 7205 6511 7239 6545
rect 7297 6511 7331 6545
rect 7389 6511 7423 6545
rect 7481 6511 7515 6545
rect 7573 6511 7607 6545
rect 7665 6511 7699 6545
rect 7757 6511 7791 6545
rect 7849 6511 7883 6545
rect 7941 6511 7975 6545
rect 8033 6511 8067 6545
rect 8125 6511 8159 6545
rect 8217 6511 8251 6545
rect 8309 6511 8343 6545
rect 8401 6511 8435 6545
rect 8493 6511 8527 6545
rect 8585 6511 8619 6545
rect 8677 6511 8711 6545
rect 8769 6511 8803 6545
rect 8861 6511 8895 6545
rect 8953 6511 8987 6545
rect 9045 6511 9079 6545
rect 9137 6511 9171 6545
rect 9229 6511 9263 6545
rect 9321 6511 9355 6545
rect 9413 6511 9447 6545
rect 9505 6511 9539 6545
rect 9597 6511 9631 6545
rect 9689 6511 9723 6545
rect 9781 6511 9815 6545
rect 9873 6511 9907 6545
rect 9965 6511 9999 6545
rect 10057 6511 10091 6545
rect 10149 6511 10183 6545
rect 10241 6511 10275 6545
rect 10333 6511 10367 6545
rect 10425 6511 10459 6545
rect 10517 6511 10551 6545
rect 10609 6511 10643 6545
rect 10701 6511 10735 6545
rect 10793 6511 10827 6545
rect 10885 6511 10919 6545
rect 10977 6511 11011 6545
rect 11069 6511 11103 6545
rect 11161 6511 11195 6545
rect 11253 6511 11287 6545
rect 11345 6511 11379 6545
rect 11437 6511 11471 6545
rect 11529 6511 11563 6545
rect 11621 6511 11655 6545
rect 11713 6511 11747 6545
rect 11805 6511 11839 6545
rect 11897 6511 11931 6545
rect 11989 6511 12023 6545
rect 12081 6511 12115 6545
rect 12173 6511 12207 6545
rect 12265 6511 12299 6545
rect 12357 6511 12391 6545
rect 12449 6511 12483 6545
rect 12541 6511 12575 6545
rect 12633 6511 12667 6545
rect 12725 6511 12759 6545
rect 12817 6511 12851 6545
rect 12909 6511 12943 6545
rect 13001 6511 13035 6545
rect 13093 6511 13127 6545
rect 13185 6511 13219 6545
rect 13277 6511 13311 6545
rect 13369 6511 13403 6545
rect 13461 6511 13495 6545
rect 13553 6511 13587 6545
rect 13645 6511 13679 6545
rect 13737 6511 13771 6545
rect 13829 6511 13863 6545
rect 13921 6511 13955 6545
rect 14013 6511 14047 6545
rect 14105 6511 14139 6545
rect 14197 6511 14231 6545
rect 14289 6511 14323 6545
rect 14381 6511 14415 6545
rect 14473 6511 14507 6545
rect 14565 6511 14599 6545
rect 14657 6511 14691 6545
rect 14749 6511 14783 6545
rect 14841 6511 14875 6545
rect 14933 6511 14967 6545
rect 15025 6511 15059 6545
rect 15117 6511 15151 6545
rect 15209 6511 15243 6545
rect 15301 6511 15335 6545
rect 15393 6511 15427 6545
rect 15485 6511 15519 6545
rect 15577 6511 15611 6545
rect 15669 6511 15703 6545
rect 15761 6511 15795 6545
rect 15853 6511 15887 6545
rect 15945 6511 15979 6545
rect 16037 6511 16071 6545
rect 16129 6511 16163 6545
rect 16221 6511 16255 6545
rect 16313 6511 16347 6545
rect 16405 6511 16439 6545
rect 16497 6511 16531 6545
rect 16589 6511 16623 6545
rect 16681 6511 16715 6545
rect 16773 6511 16807 6545
rect 16865 6511 16899 6545
rect 16957 6511 16991 6545
rect 17049 6511 17083 6545
rect 17141 6511 17175 6545
rect 17233 6511 17267 6545
rect 17325 6511 17359 6545
rect 17417 6511 17451 6545
rect 17509 6511 17543 6545
rect 17601 6511 17635 6545
rect 17693 6511 17727 6545
rect 17785 6511 17819 6545
rect 17877 6511 17911 6545
rect 17969 6511 18003 6545
rect 18061 6511 18095 6545
rect 18153 6511 18187 6545
rect 18245 6511 18279 6545
rect 18337 6511 18371 6545
rect 18429 6511 18463 6545
rect 18521 6511 18555 6545
rect 18613 6511 18647 6545
rect 18705 6511 18739 6545
rect 18797 6511 18831 6545
rect 8033 6273 8067 6307
rect 8217 6279 8240 6307
rect 8240 6279 8251 6307
rect 8217 6273 8251 6279
rect 8401 6069 8435 6103
rect 1133 5967 1167 6001
rect 1225 5967 1259 6001
rect 1317 5967 1351 6001
rect 1409 5967 1443 6001
rect 1501 5967 1535 6001
rect 1593 5967 1627 6001
rect 1685 5967 1719 6001
rect 1777 5967 1811 6001
rect 1869 5967 1903 6001
rect 1961 5967 1995 6001
rect 2053 5967 2087 6001
rect 2145 5967 2179 6001
rect 2237 5967 2271 6001
rect 2329 5967 2363 6001
rect 2421 5967 2455 6001
rect 2513 5967 2547 6001
rect 2605 5967 2639 6001
rect 2697 5967 2731 6001
rect 2789 5967 2823 6001
rect 2881 5967 2915 6001
rect 2973 5967 3007 6001
rect 3065 5967 3099 6001
rect 3157 5967 3191 6001
rect 3249 5967 3283 6001
rect 3341 5967 3375 6001
rect 3433 5967 3467 6001
rect 3525 5967 3559 6001
rect 3617 5967 3651 6001
rect 3709 5967 3743 6001
rect 3801 5967 3835 6001
rect 3893 5967 3927 6001
rect 3985 5967 4019 6001
rect 4077 5967 4111 6001
rect 4169 5967 4203 6001
rect 4261 5967 4295 6001
rect 4353 5967 4387 6001
rect 4445 5967 4479 6001
rect 4537 5967 4571 6001
rect 4629 5967 4663 6001
rect 4721 5967 4755 6001
rect 4813 5967 4847 6001
rect 4905 5967 4939 6001
rect 4997 5967 5031 6001
rect 5089 5967 5123 6001
rect 5181 5967 5215 6001
rect 5273 5967 5307 6001
rect 5365 5967 5399 6001
rect 5457 5967 5491 6001
rect 5549 5967 5583 6001
rect 5641 5967 5675 6001
rect 5733 5967 5767 6001
rect 5825 5967 5859 6001
rect 5917 5967 5951 6001
rect 6009 5967 6043 6001
rect 6101 5967 6135 6001
rect 6193 5967 6227 6001
rect 6285 5967 6319 6001
rect 6377 5967 6411 6001
rect 6469 5967 6503 6001
rect 6561 5967 6595 6001
rect 6653 5967 6687 6001
rect 6745 5967 6779 6001
rect 6837 5967 6871 6001
rect 6929 5967 6963 6001
rect 7021 5967 7055 6001
rect 7113 5967 7147 6001
rect 7205 5967 7239 6001
rect 7297 5967 7331 6001
rect 7389 5967 7423 6001
rect 7481 5967 7515 6001
rect 7573 5967 7607 6001
rect 7665 5967 7699 6001
rect 7757 5967 7791 6001
rect 7849 5967 7883 6001
rect 7941 5967 7975 6001
rect 8033 5967 8067 6001
rect 8125 5967 8159 6001
rect 8217 5967 8251 6001
rect 8309 5967 8343 6001
rect 8401 5967 8435 6001
rect 8493 5967 8527 6001
rect 8585 5967 8619 6001
rect 8677 5967 8711 6001
rect 8769 5967 8803 6001
rect 8861 5967 8895 6001
rect 8953 5967 8987 6001
rect 9045 5967 9079 6001
rect 9137 5967 9171 6001
rect 9229 5967 9263 6001
rect 9321 5967 9355 6001
rect 9413 5967 9447 6001
rect 9505 5967 9539 6001
rect 9597 5967 9631 6001
rect 9689 5967 9723 6001
rect 9781 5967 9815 6001
rect 9873 5967 9907 6001
rect 9965 5967 9999 6001
rect 10057 5967 10091 6001
rect 10149 5967 10183 6001
rect 10241 5967 10275 6001
rect 10333 5967 10367 6001
rect 10425 5967 10459 6001
rect 10517 5967 10551 6001
rect 10609 5967 10643 6001
rect 10701 5967 10735 6001
rect 10793 5967 10827 6001
rect 10885 5967 10919 6001
rect 10977 5967 11011 6001
rect 11069 5967 11103 6001
rect 11161 5967 11195 6001
rect 11253 5967 11287 6001
rect 11345 5967 11379 6001
rect 11437 5967 11471 6001
rect 11529 5967 11563 6001
rect 11621 5967 11655 6001
rect 11713 5967 11747 6001
rect 11805 5967 11839 6001
rect 11897 5967 11931 6001
rect 11989 5967 12023 6001
rect 12081 5967 12115 6001
rect 12173 5967 12207 6001
rect 12265 5967 12299 6001
rect 12357 5967 12391 6001
rect 12449 5967 12483 6001
rect 12541 5967 12575 6001
rect 12633 5967 12667 6001
rect 12725 5967 12759 6001
rect 12817 5967 12851 6001
rect 12909 5967 12943 6001
rect 13001 5967 13035 6001
rect 13093 5967 13127 6001
rect 13185 5967 13219 6001
rect 13277 5967 13311 6001
rect 13369 5967 13403 6001
rect 13461 5967 13495 6001
rect 13553 5967 13587 6001
rect 13645 5967 13679 6001
rect 13737 5967 13771 6001
rect 13829 5967 13863 6001
rect 13921 5967 13955 6001
rect 14013 5967 14047 6001
rect 14105 5967 14139 6001
rect 14197 5967 14231 6001
rect 14289 5967 14323 6001
rect 14381 5967 14415 6001
rect 14473 5967 14507 6001
rect 14565 5967 14599 6001
rect 14657 5967 14691 6001
rect 14749 5967 14783 6001
rect 14841 5967 14875 6001
rect 14933 5967 14967 6001
rect 15025 5967 15059 6001
rect 15117 5967 15151 6001
rect 15209 5967 15243 6001
rect 15301 5967 15335 6001
rect 15393 5967 15427 6001
rect 15485 5967 15519 6001
rect 15577 5967 15611 6001
rect 15669 5967 15703 6001
rect 15761 5967 15795 6001
rect 15853 5967 15887 6001
rect 15945 5967 15979 6001
rect 16037 5967 16071 6001
rect 16129 5967 16163 6001
rect 16221 5967 16255 6001
rect 16313 5967 16347 6001
rect 16405 5967 16439 6001
rect 16497 5967 16531 6001
rect 16589 5967 16623 6001
rect 16681 5967 16715 6001
rect 16773 5967 16807 6001
rect 16865 5967 16899 6001
rect 16957 5967 16991 6001
rect 17049 5967 17083 6001
rect 17141 5967 17175 6001
rect 17233 5967 17267 6001
rect 17325 5967 17359 6001
rect 17417 5967 17451 6001
rect 17509 5967 17543 6001
rect 17601 5967 17635 6001
rect 17693 5967 17727 6001
rect 17785 5967 17819 6001
rect 17877 5967 17911 6001
rect 17969 5967 18003 6001
rect 18061 5967 18095 6001
rect 18153 5967 18187 6001
rect 18245 5967 18279 6001
rect 18337 5967 18371 6001
rect 18429 5967 18463 6001
rect 18521 5967 18555 6001
rect 18613 5967 18647 6001
rect 18705 5967 18739 6001
rect 18797 5967 18831 6001
rect 6929 5689 6963 5695
rect 6929 5661 6955 5689
rect 6955 5661 6963 5689
rect 7757 5729 7791 5763
rect 6745 5529 6751 5559
rect 6751 5529 6779 5559
rect 6745 5525 6779 5529
rect 7849 5525 7883 5559
rect 7941 5619 7953 5627
rect 7953 5619 7975 5627
rect 7941 5593 7975 5619
rect 8309 5891 8337 5899
rect 8337 5891 8343 5899
rect 8309 5865 8343 5891
rect 11529 5593 11563 5627
rect 11713 5593 11747 5627
rect 11897 5525 11931 5559
rect 12817 5593 12851 5627
rect 13001 5593 13035 5627
rect 13185 5525 13219 5559
rect 1133 5423 1167 5457
rect 1225 5423 1259 5457
rect 1317 5423 1351 5457
rect 1409 5423 1443 5457
rect 1501 5423 1535 5457
rect 1593 5423 1627 5457
rect 1685 5423 1719 5457
rect 1777 5423 1811 5457
rect 1869 5423 1903 5457
rect 1961 5423 1995 5457
rect 2053 5423 2087 5457
rect 2145 5423 2179 5457
rect 2237 5423 2271 5457
rect 2329 5423 2363 5457
rect 2421 5423 2455 5457
rect 2513 5423 2547 5457
rect 2605 5423 2639 5457
rect 2697 5423 2731 5457
rect 2789 5423 2823 5457
rect 2881 5423 2915 5457
rect 2973 5423 3007 5457
rect 3065 5423 3099 5457
rect 3157 5423 3191 5457
rect 3249 5423 3283 5457
rect 3341 5423 3375 5457
rect 3433 5423 3467 5457
rect 3525 5423 3559 5457
rect 3617 5423 3651 5457
rect 3709 5423 3743 5457
rect 3801 5423 3835 5457
rect 3893 5423 3927 5457
rect 3985 5423 4019 5457
rect 4077 5423 4111 5457
rect 4169 5423 4203 5457
rect 4261 5423 4295 5457
rect 4353 5423 4387 5457
rect 4445 5423 4479 5457
rect 4537 5423 4571 5457
rect 4629 5423 4663 5457
rect 4721 5423 4755 5457
rect 4813 5423 4847 5457
rect 4905 5423 4939 5457
rect 4997 5423 5031 5457
rect 5089 5423 5123 5457
rect 5181 5423 5215 5457
rect 5273 5423 5307 5457
rect 5365 5423 5399 5457
rect 5457 5423 5491 5457
rect 5549 5423 5583 5457
rect 5641 5423 5675 5457
rect 5733 5423 5767 5457
rect 5825 5423 5859 5457
rect 5917 5423 5951 5457
rect 6009 5423 6043 5457
rect 6101 5423 6135 5457
rect 6193 5423 6227 5457
rect 6285 5423 6319 5457
rect 6377 5423 6411 5457
rect 6469 5423 6503 5457
rect 6561 5423 6595 5457
rect 6653 5423 6687 5457
rect 6745 5423 6779 5457
rect 6837 5423 6871 5457
rect 6929 5423 6963 5457
rect 7021 5423 7055 5457
rect 7113 5423 7147 5457
rect 7205 5423 7239 5457
rect 7297 5423 7331 5457
rect 7389 5423 7423 5457
rect 7481 5423 7515 5457
rect 7573 5423 7607 5457
rect 7665 5423 7699 5457
rect 7757 5423 7791 5457
rect 7849 5423 7883 5457
rect 7941 5423 7975 5457
rect 8033 5423 8067 5457
rect 8125 5423 8159 5457
rect 8217 5423 8251 5457
rect 8309 5423 8343 5457
rect 8401 5423 8435 5457
rect 8493 5423 8527 5457
rect 8585 5423 8619 5457
rect 8677 5423 8711 5457
rect 8769 5423 8803 5457
rect 8861 5423 8895 5457
rect 8953 5423 8987 5457
rect 9045 5423 9079 5457
rect 9137 5423 9171 5457
rect 9229 5423 9263 5457
rect 9321 5423 9355 5457
rect 9413 5423 9447 5457
rect 9505 5423 9539 5457
rect 9597 5423 9631 5457
rect 9689 5423 9723 5457
rect 9781 5423 9815 5457
rect 9873 5423 9907 5457
rect 9965 5423 9999 5457
rect 10057 5423 10091 5457
rect 10149 5423 10183 5457
rect 10241 5423 10275 5457
rect 10333 5423 10367 5457
rect 10425 5423 10459 5457
rect 10517 5423 10551 5457
rect 10609 5423 10643 5457
rect 10701 5423 10735 5457
rect 10793 5423 10827 5457
rect 10885 5423 10919 5457
rect 10977 5423 11011 5457
rect 11069 5423 11103 5457
rect 11161 5423 11195 5457
rect 11253 5423 11287 5457
rect 11345 5423 11379 5457
rect 11437 5423 11471 5457
rect 11529 5423 11563 5457
rect 11621 5423 11655 5457
rect 11713 5423 11747 5457
rect 11805 5423 11839 5457
rect 11897 5423 11931 5457
rect 11989 5423 12023 5457
rect 12081 5423 12115 5457
rect 12173 5423 12207 5457
rect 12265 5423 12299 5457
rect 12357 5423 12391 5457
rect 12449 5423 12483 5457
rect 12541 5423 12575 5457
rect 12633 5423 12667 5457
rect 12725 5423 12759 5457
rect 12817 5423 12851 5457
rect 12909 5423 12943 5457
rect 13001 5423 13035 5457
rect 13093 5423 13127 5457
rect 13185 5423 13219 5457
rect 13277 5423 13311 5457
rect 13369 5423 13403 5457
rect 13461 5423 13495 5457
rect 13553 5423 13587 5457
rect 13645 5423 13679 5457
rect 13737 5423 13771 5457
rect 13829 5423 13863 5457
rect 13921 5423 13955 5457
rect 14013 5423 14047 5457
rect 14105 5423 14139 5457
rect 14197 5423 14231 5457
rect 14289 5423 14323 5457
rect 14381 5423 14415 5457
rect 14473 5423 14507 5457
rect 14565 5423 14599 5457
rect 14657 5423 14691 5457
rect 14749 5423 14783 5457
rect 14841 5423 14875 5457
rect 14933 5423 14967 5457
rect 15025 5423 15059 5457
rect 15117 5423 15151 5457
rect 15209 5423 15243 5457
rect 15301 5423 15335 5457
rect 15393 5423 15427 5457
rect 15485 5423 15519 5457
rect 15577 5423 15611 5457
rect 15669 5423 15703 5457
rect 15761 5423 15795 5457
rect 15853 5423 15887 5457
rect 15945 5423 15979 5457
rect 16037 5423 16071 5457
rect 16129 5423 16163 5457
rect 16221 5423 16255 5457
rect 16313 5423 16347 5457
rect 16405 5423 16439 5457
rect 16497 5423 16531 5457
rect 16589 5423 16623 5457
rect 16681 5423 16715 5457
rect 16773 5423 16807 5457
rect 16865 5423 16899 5457
rect 16957 5423 16991 5457
rect 17049 5423 17083 5457
rect 17141 5423 17175 5457
rect 17233 5423 17267 5457
rect 17325 5423 17359 5457
rect 17417 5423 17451 5457
rect 17509 5423 17543 5457
rect 17601 5423 17635 5457
rect 17693 5423 17727 5457
rect 17785 5423 17819 5457
rect 17877 5423 17911 5457
rect 17969 5423 18003 5457
rect 18061 5423 18095 5457
rect 18153 5423 18187 5457
rect 18245 5423 18279 5457
rect 18337 5423 18371 5457
rect 18429 5423 18463 5457
rect 18521 5423 18555 5457
rect 18613 5423 18647 5457
rect 18705 5423 18739 5457
rect 18797 5423 18831 5457
rect 2789 5117 2823 5151
rect 2882 5210 2916 5219
rect 2882 5185 2894 5210
rect 2894 5185 2916 5210
rect 3065 5117 3099 5151
rect 2963 5065 2997 5083
rect 2963 5049 2997 5065
rect 3249 5185 3283 5219
rect 3521 5253 3555 5287
rect 3593 5271 3627 5287
rect 3593 5253 3617 5271
rect 3617 5253 3627 5271
rect 3341 5049 3375 5083
rect 3965 5201 3991 5219
rect 3991 5201 3999 5219
rect 3965 5185 3999 5201
rect 4537 5331 4571 5355
rect 4241 5253 4275 5287
rect 4181 5199 4197 5224
rect 4197 5199 4215 5224
rect 4181 5190 4215 5199
rect 4537 5321 4565 5331
rect 4565 5321 4571 5331
rect 3965 5075 3996 5083
rect 3996 5075 3999 5083
rect 3965 5049 3999 5075
rect 7021 5321 7055 5355
rect 6653 4989 6687 5015
rect 6653 4981 6659 4989
rect 6659 4981 6687 4989
rect 7113 5321 7147 5355
rect 7205 5117 7239 5151
rect 7849 5117 7883 5151
rect 7942 5210 7976 5219
rect 7942 5185 7954 5210
rect 7954 5185 7976 5210
rect 8125 5117 8159 5151
rect 8023 5065 8057 5083
rect 8023 5049 8057 5065
rect 8309 5185 8343 5219
rect 8581 5253 8615 5287
rect 8653 5271 8687 5287
rect 8653 5253 8677 5271
rect 8677 5253 8687 5271
rect 8401 5049 8435 5083
rect 9025 5201 9051 5219
rect 9051 5201 9059 5219
rect 9025 5185 9059 5201
rect 9301 5253 9335 5287
rect 9241 5199 9257 5224
rect 9257 5199 9275 5224
rect 9241 5190 9275 5199
rect 9025 5075 9056 5083
rect 9056 5075 9059 5083
rect 9025 5049 9059 5075
rect 9597 4991 9625 5015
rect 9625 4991 9631 5015
rect 9597 4981 9631 4991
rect 10333 5253 10367 5287
rect 10149 5148 10183 5151
rect 10149 5117 10163 5148
rect 10163 5117 10183 5148
rect 10425 5321 10459 5355
rect 11713 5328 11719 5355
rect 11719 5328 11747 5355
rect 11713 5321 11747 5328
rect 10793 4989 10827 5015
rect 10793 4981 10821 4989
rect 10821 4981 10827 4989
rect 12081 5261 12115 5287
rect 12081 5253 12103 5261
rect 12103 5253 12115 5261
rect 12173 5321 12207 5355
rect 12265 5117 12299 5151
rect 13185 5321 13219 5355
rect 13093 5117 13127 5151
rect 13277 5185 13311 5219
rect 13645 4989 13679 5015
rect 13645 4981 13673 4989
rect 13673 4981 13679 4989
rect 1133 4879 1167 4913
rect 1225 4879 1259 4913
rect 1317 4879 1351 4913
rect 1409 4879 1443 4913
rect 1501 4879 1535 4913
rect 1593 4879 1627 4913
rect 1685 4879 1719 4913
rect 1777 4879 1811 4913
rect 1869 4879 1903 4913
rect 1961 4879 1995 4913
rect 2053 4879 2087 4913
rect 2145 4879 2179 4913
rect 2237 4879 2271 4913
rect 2329 4879 2363 4913
rect 2421 4879 2455 4913
rect 2513 4879 2547 4913
rect 2605 4879 2639 4913
rect 2697 4879 2731 4913
rect 2789 4879 2823 4913
rect 2881 4879 2915 4913
rect 2973 4879 3007 4913
rect 3065 4879 3099 4913
rect 3157 4879 3191 4913
rect 3249 4879 3283 4913
rect 3341 4879 3375 4913
rect 3433 4879 3467 4913
rect 3525 4879 3559 4913
rect 3617 4879 3651 4913
rect 3709 4879 3743 4913
rect 3801 4879 3835 4913
rect 3893 4879 3927 4913
rect 3985 4879 4019 4913
rect 4077 4879 4111 4913
rect 4169 4879 4203 4913
rect 4261 4879 4295 4913
rect 4353 4879 4387 4913
rect 4445 4879 4479 4913
rect 4537 4879 4571 4913
rect 4629 4879 4663 4913
rect 4721 4879 4755 4913
rect 4813 4879 4847 4913
rect 4905 4879 4939 4913
rect 4997 4879 5031 4913
rect 5089 4879 5123 4913
rect 5181 4879 5215 4913
rect 5273 4879 5307 4913
rect 5365 4879 5399 4913
rect 5457 4879 5491 4913
rect 5549 4879 5583 4913
rect 5641 4879 5675 4913
rect 5733 4879 5767 4913
rect 5825 4879 5859 4913
rect 5917 4879 5951 4913
rect 6009 4879 6043 4913
rect 6101 4879 6135 4913
rect 6193 4879 6227 4913
rect 6285 4879 6319 4913
rect 6377 4879 6411 4913
rect 6469 4879 6503 4913
rect 6561 4879 6595 4913
rect 6653 4879 6687 4913
rect 6745 4879 6779 4913
rect 6837 4879 6871 4913
rect 6929 4879 6963 4913
rect 7021 4879 7055 4913
rect 7113 4879 7147 4913
rect 7205 4879 7239 4913
rect 7297 4879 7331 4913
rect 7389 4879 7423 4913
rect 7481 4879 7515 4913
rect 7573 4879 7607 4913
rect 7665 4879 7699 4913
rect 7757 4879 7791 4913
rect 7849 4879 7883 4913
rect 7941 4879 7975 4913
rect 8033 4879 8067 4913
rect 8125 4879 8159 4913
rect 8217 4879 8251 4913
rect 8309 4879 8343 4913
rect 8401 4879 8435 4913
rect 8493 4879 8527 4913
rect 8585 4879 8619 4913
rect 8677 4879 8711 4913
rect 8769 4879 8803 4913
rect 8861 4879 8895 4913
rect 8953 4879 8987 4913
rect 9045 4879 9079 4913
rect 9137 4879 9171 4913
rect 9229 4879 9263 4913
rect 9321 4879 9355 4913
rect 9413 4879 9447 4913
rect 9505 4879 9539 4913
rect 9597 4879 9631 4913
rect 9689 4879 9723 4913
rect 9781 4879 9815 4913
rect 9873 4879 9907 4913
rect 9965 4879 9999 4913
rect 10057 4879 10091 4913
rect 10149 4879 10183 4913
rect 10241 4879 10275 4913
rect 10333 4879 10367 4913
rect 10425 4879 10459 4913
rect 10517 4879 10551 4913
rect 10609 4879 10643 4913
rect 10701 4879 10735 4913
rect 10793 4879 10827 4913
rect 10885 4879 10919 4913
rect 10977 4879 11011 4913
rect 11069 4879 11103 4913
rect 11161 4879 11195 4913
rect 11253 4879 11287 4913
rect 11345 4879 11379 4913
rect 11437 4879 11471 4913
rect 11529 4879 11563 4913
rect 11621 4879 11655 4913
rect 11713 4879 11747 4913
rect 11805 4879 11839 4913
rect 11897 4879 11931 4913
rect 11989 4879 12023 4913
rect 12081 4879 12115 4913
rect 12173 4879 12207 4913
rect 12265 4879 12299 4913
rect 12357 4879 12391 4913
rect 12449 4879 12483 4913
rect 12541 4879 12575 4913
rect 12633 4879 12667 4913
rect 12725 4879 12759 4913
rect 12817 4879 12851 4913
rect 12909 4879 12943 4913
rect 13001 4879 13035 4913
rect 13093 4879 13127 4913
rect 13185 4879 13219 4913
rect 13277 4879 13311 4913
rect 13369 4879 13403 4913
rect 13461 4879 13495 4913
rect 13553 4879 13587 4913
rect 13645 4879 13679 4913
rect 13737 4879 13771 4913
rect 13829 4879 13863 4913
rect 13921 4879 13955 4913
rect 14013 4879 14047 4913
rect 14105 4879 14139 4913
rect 14197 4879 14231 4913
rect 14289 4879 14323 4913
rect 14381 4879 14415 4913
rect 14473 4879 14507 4913
rect 14565 4879 14599 4913
rect 14657 4879 14691 4913
rect 14749 4879 14783 4913
rect 14841 4879 14875 4913
rect 14933 4879 14967 4913
rect 15025 4879 15059 4913
rect 15117 4879 15151 4913
rect 15209 4879 15243 4913
rect 15301 4879 15335 4913
rect 15393 4879 15427 4913
rect 15485 4879 15519 4913
rect 15577 4879 15611 4913
rect 15669 4879 15703 4913
rect 15761 4879 15795 4913
rect 15853 4879 15887 4913
rect 15945 4879 15979 4913
rect 16037 4879 16071 4913
rect 16129 4879 16163 4913
rect 16221 4879 16255 4913
rect 16313 4879 16347 4913
rect 16405 4879 16439 4913
rect 16497 4879 16531 4913
rect 16589 4879 16623 4913
rect 16681 4879 16715 4913
rect 16773 4879 16807 4913
rect 16865 4879 16899 4913
rect 16957 4879 16991 4913
rect 17049 4879 17083 4913
rect 17141 4879 17175 4913
rect 17233 4879 17267 4913
rect 17325 4879 17359 4913
rect 17417 4879 17451 4913
rect 17509 4879 17543 4913
rect 17601 4879 17635 4913
rect 17693 4879 17727 4913
rect 17785 4879 17819 4913
rect 17877 4879 17911 4913
rect 17969 4879 18003 4913
rect 18061 4879 18095 4913
rect 18153 4879 18187 4913
rect 18245 4879 18279 4913
rect 18337 4879 18371 4913
rect 18429 4879 18463 4913
rect 18521 4879 18555 4913
rect 18613 4879 18647 4913
rect 18705 4879 18739 4913
rect 18797 4879 18831 4913
rect 2421 4437 2446 4471
rect 2446 4437 2455 4471
rect 3065 4573 3099 4607
rect 4353 4505 4387 4539
rect 4077 4437 4084 4471
rect 4084 4437 4111 4471
rect 4905 4573 4939 4607
rect 6193 4505 6227 4539
rect 6377 4573 6411 4607
rect 7205 4777 7239 4811
rect 6837 4573 6871 4607
rect 7021 4505 7055 4539
rect 6009 4437 6043 4471
rect 7849 4735 7855 4743
rect 7855 4735 7883 4743
rect 7849 4709 7883 4735
rect 8217 4437 8251 4471
rect 8401 4641 8435 4675
rect 8309 4573 8343 4607
rect 9137 4505 9171 4539
rect 9321 4505 9355 4539
rect 9505 4437 9539 4471
rect 9965 4573 9999 4607
rect 10517 4573 10551 4607
rect 10701 4505 10735 4539
rect 10885 4437 10919 4471
rect 11529 4714 11557 4743
rect 11557 4714 11563 4743
rect 11529 4709 11563 4714
rect 11345 4601 11379 4607
rect 11345 4573 11353 4601
rect 11353 4573 11379 4601
rect 12081 4644 12095 4675
rect 12095 4644 12115 4675
rect 12081 4641 12115 4644
rect 12265 4644 12297 4675
rect 12297 4644 12299 4675
rect 12265 4641 12299 4644
rect 12725 4803 12753 4811
rect 12753 4803 12759 4811
rect 12725 4777 12759 4803
rect 12357 4437 12391 4471
rect 13369 4601 13403 4607
rect 13369 4573 13395 4601
rect 13395 4573 13403 4601
rect 13185 4441 13191 4471
rect 13191 4441 13219 4471
rect 13185 4437 13219 4441
rect 15209 4573 15243 4607
rect 15393 4505 15427 4539
rect 15577 4505 15611 4539
rect 16221 4601 16255 4607
rect 16221 4573 16247 4601
rect 16247 4573 16255 4601
rect 16037 4441 16043 4471
rect 16043 4441 16071 4471
rect 16037 4437 16071 4441
rect 16865 4601 16899 4607
rect 16865 4573 16891 4601
rect 16891 4573 16899 4601
rect 16681 4441 16687 4471
rect 16687 4441 16715 4471
rect 16681 4437 16715 4441
rect 1133 4335 1167 4369
rect 1225 4335 1259 4369
rect 1317 4335 1351 4369
rect 1409 4335 1443 4369
rect 1501 4335 1535 4369
rect 1593 4335 1627 4369
rect 1685 4335 1719 4369
rect 1777 4335 1811 4369
rect 1869 4335 1903 4369
rect 1961 4335 1995 4369
rect 2053 4335 2087 4369
rect 2145 4335 2179 4369
rect 2237 4335 2271 4369
rect 2329 4335 2363 4369
rect 2421 4335 2455 4369
rect 2513 4335 2547 4369
rect 2605 4335 2639 4369
rect 2697 4335 2731 4369
rect 2789 4335 2823 4369
rect 2881 4335 2915 4369
rect 2973 4335 3007 4369
rect 3065 4335 3099 4369
rect 3157 4335 3191 4369
rect 3249 4335 3283 4369
rect 3341 4335 3375 4369
rect 3433 4335 3467 4369
rect 3525 4335 3559 4369
rect 3617 4335 3651 4369
rect 3709 4335 3743 4369
rect 3801 4335 3835 4369
rect 3893 4335 3927 4369
rect 3985 4335 4019 4369
rect 4077 4335 4111 4369
rect 4169 4335 4203 4369
rect 4261 4335 4295 4369
rect 4353 4335 4387 4369
rect 4445 4335 4479 4369
rect 4537 4335 4571 4369
rect 4629 4335 4663 4369
rect 4721 4335 4755 4369
rect 4813 4335 4847 4369
rect 4905 4335 4939 4369
rect 4997 4335 5031 4369
rect 5089 4335 5123 4369
rect 5181 4335 5215 4369
rect 5273 4335 5307 4369
rect 5365 4335 5399 4369
rect 5457 4335 5491 4369
rect 5549 4335 5583 4369
rect 5641 4335 5675 4369
rect 5733 4335 5767 4369
rect 5825 4335 5859 4369
rect 5917 4335 5951 4369
rect 6009 4335 6043 4369
rect 6101 4335 6135 4369
rect 6193 4335 6227 4369
rect 6285 4335 6319 4369
rect 6377 4335 6411 4369
rect 6469 4335 6503 4369
rect 6561 4335 6595 4369
rect 6653 4335 6687 4369
rect 6745 4335 6779 4369
rect 6837 4335 6871 4369
rect 6929 4335 6963 4369
rect 7021 4335 7055 4369
rect 7113 4335 7147 4369
rect 7205 4335 7239 4369
rect 7297 4335 7331 4369
rect 7389 4335 7423 4369
rect 7481 4335 7515 4369
rect 7573 4335 7607 4369
rect 7665 4335 7699 4369
rect 7757 4335 7791 4369
rect 7849 4335 7883 4369
rect 7941 4335 7975 4369
rect 8033 4335 8067 4369
rect 8125 4335 8159 4369
rect 8217 4335 8251 4369
rect 8309 4335 8343 4369
rect 8401 4335 8435 4369
rect 8493 4335 8527 4369
rect 8585 4335 8619 4369
rect 8677 4335 8711 4369
rect 8769 4335 8803 4369
rect 8861 4335 8895 4369
rect 8953 4335 8987 4369
rect 9045 4335 9079 4369
rect 9137 4335 9171 4369
rect 9229 4335 9263 4369
rect 9321 4335 9355 4369
rect 9413 4335 9447 4369
rect 9505 4335 9539 4369
rect 9597 4335 9631 4369
rect 9689 4335 9723 4369
rect 9781 4335 9815 4369
rect 9873 4335 9907 4369
rect 9965 4335 9999 4369
rect 10057 4335 10091 4369
rect 10149 4335 10183 4369
rect 10241 4335 10275 4369
rect 10333 4335 10367 4369
rect 10425 4335 10459 4369
rect 10517 4335 10551 4369
rect 10609 4335 10643 4369
rect 10701 4335 10735 4369
rect 10793 4335 10827 4369
rect 10885 4335 10919 4369
rect 10977 4335 11011 4369
rect 11069 4335 11103 4369
rect 11161 4335 11195 4369
rect 11253 4335 11287 4369
rect 11345 4335 11379 4369
rect 11437 4335 11471 4369
rect 11529 4335 11563 4369
rect 11621 4335 11655 4369
rect 11713 4335 11747 4369
rect 11805 4335 11839 4369
rect 11897 4335 11931 4369
rect 11989 4335 12023 4369
rect 12081 4335 12115 4369
rect 12173 4335 12207 4369
rect 12265 4335 12299 4369
rect 12357 4335 12391 4369
rect 12449 4335 12483 4369
rect 12541 4335 12575 4369
rect 12633 4335 12667 4369
rect 12725 4335 12759 4369
rect 12817 4335 12851 4369
rect 12909 4335 12943 4369
rect 13001 4335 13035 4369
rect 13093 4335 13127 4369
rect 13185 4335 13219 4369
rect 13277 4335 13311 4369
rect 13369 4335 13403 4369
rect 13461 4335 13495 4369
rect 13553 4335 13587 4369
rect 13645 4335 13679 4369
rect 13737 4335 13771 4369
rect 13829 4335 13863 4369
rect 13921 4335 13955 4369
rect 14013 4335 14047 4369
rect 14105 4335 14139 4369
rect 14197 4335 14231 4369
rect 14289 4335 14323 4369
rect 14381 4335 14415 4369
rect 14473 4335 14507 4369
rect 14565 4335 14599 4369
rect 14657 4335 14691 4369
rect 14749 4335 14783 4369
rect 14841 4335 14875 4369
rect 14933 4335 14967 4369
rect 15025 4335 15059 4369
rect 15117 4335 15151 4369
rect 15209 4335 15243 4369
rect 15301 4335 15335 4369
rect 15393 4335 15427 4369
rect 15485 4335 15519 4369
rect 15577 4335 15611 4369
rect 15669 4335 15703 4369
rect 15761 4335 15795 4369
rect 15853 4335 15887 4369
rect 15945 4335 15979 4369
rect 16037 4335 16071 4369
rect 16129 4335 16163 4369
rect 16221 4335 16255 4369
rect 16313 4335 16347 4369
rect 16405 4335 16439 4369
rect 16497 4335 16531 4369
rect 16589 4335 16623 4369
rect 16681 4335 16715 4369
rect 16773 4335 16807 4369
rect 16865 4335 16899 4369
rect 16957 4335 16991 4369
rect 17049 4335 17083 4369
rect 17141 4335 17175 4369
rect 17233 4335 17267 4369
rect 17325 4335 17359 4369
rect 17417 4335 17451 4369
rect 17509 4335 17543 4369
rect 17601 4335 17635 4369
rect 17693 4335 17727 4369
rect 17785 4335 17819 4369
rect 17877 4335 17911 4369
rect 17969 4335 18003 4369
rect 18061 4335 18095 4369
rect 18153 4335 18187 4369
rect 18245 4335 18279 4369
rect 18337 4335 18371 4369
rect 18429 4335 18463 4369
rect 18521 4335 18555 4369
rect 18613 4335 18647 4369
rect 18705 4335 18739 4369
rect 18797 4335 18831 4369
rect 2421 4263 2455 4267
rect 2421 4233 2449 4263
rect 2449 4233 2455 4263
rect 2237 4103 2245 4131
rect 2245 4103 2271 4131
rect 2237 4097 2271 4103
rect 2881 4029 2915 4063
rect 2974 4122 3008 4131
rect 2974 4097 2986 4122
rect 2986 4097 3008 4122
rect 3157 4029 3191 4063
rect 3055 3977 3089 3995
rect 3055 3961 3089 3977
rect 3341 4097 3375 4131
rect 3613 4165 3647 4199
rect 3685 4183 3719 4199
rect 3685 4165 3709 4183
rect 3709 4165 3719 4183
rect 3433 3961 3467 3995
rect 4057 4113 4083 4131
rect 4083 4113 4091 4131
rect 4057 4097 4091 4113
rect 4333 4165 4367 4199
rect 4273 4111 4289 4136
rect 4289 4111 4307 4136
rect 4273 4102 4307 4111
rect 4057 3987 4088 3995
rect 4088 3987 4091 3995
rect 4057 3961 4091 3987
rect 4629 3903 4657 3927
rect 4657 3903 4663 3927
rect 4629 3893 4663 3903
rect 5089 3961 5123 3995
rect 6837 4103 6863 4131
rect 6863 4103 6871 4131
rect 6837 4097 6871 4103
rect 6653 3990 6687 3995
rect 6653 3961 6659 3990
rect 6659 3961 6687 3990
rect 7757 4060 7791 4063
rect 7757 4029 7771 4060
rect 7771 4029 7791 4060
rect 8033 4233 8067 4267
rect 8401 4240 8429 4267
rect 8429 4240 8435 4267
rect 8401 4233 8435 4240
rect 7941 4060 7975 4063
rect 7941 4029 7973 4060
rect 7973 4029 7975 4060
rect 8955 4165 8989 4199
rect 11713 4243 11747 4267
rect 11713 4233 11719 4243
rect 11719 4233 11747 4243
rect 12009 4165 12043 4199
rect 12069 4111 12087 4136
rect 12087 4111 12103 4136
rect 12069 4102 12103 4111
rect 10241 3911 10248 3927
rect 10248 3911 10275 3927
rect 10241 3893 10275 3911
rect 12285 4113 12293 4131
rect 12293 4113 12319 4131
rect 12285 4097 12319 4113
rect 12657 4183 12691 4199
rect 12657 4165 12667 4183
rect 12667 4165 12691 4183
rect 12729 4165 12763 4199
rect 12285 3987 12288 3995
rect 12288 3987 12319 3995
rect 12285 3961 12319 3987
rect 13001 4097 13035 4131
rect 12909 3961 12943 3995
rect 13185 4029 13219 4063
rect 13287 3977 13321 3995
rect 13287 3961 13321 3977
rect 13368 4122 13402 4131
rect 13368 4097 13390 4122
rect 13390 4097 13402 4122
rect 13461 4029 13495 4063
rect 13921 4029 13955 4063
rect 14014 4122 14048 4131
rect 14014 4097 14026 4122
rect 14026 4097 14048 4122
rect 14197 4029 14231 4063
rect 14095 3977 14129 3995
rect 14095 3961 14129 3977
rect 14381 4097 14415 4131
rect 14653 4165 14687 4199
rect 14725 4183 14759 4199
rect 14725 4165 14749 4183
rect 14749 4165 14759 4183
rect 14473 3961 14507 3995
rect 15097 4113 15123 4131
rect 15123 4113 15131 4131
rect 15097 4097 15131 4113
rect 15373 4165 15407 4199
rect 15313 4111 15329 4136
rect 15329 4111 15347 4136
rect 15313 4102 15347 4111
rect 15097 3987 15128 3995
rect 15128 3987 15131 3995
rect 15097 3961 15131 3987
rect 15669 3903 15697 3927
rect 15697 3903 15703 3927
rect 15669 3893 15703 3903
rect 1133 3791 1167 3825
rect 1225 3791 1259 3825
rect 1317 3791 1351 3825
rect 1409 3791 1443 3825
rect 1501 3791 1535 3825
rect 1593 3791 1627 3825
rect 1685 3791 1719 3825
rect 1777 3791 1811 3825
rect 1869 3791 1903 3825
rect 1961 3791 1995 3825
rect 2053 3791 2087 3825
rect 2145 3791 2179 3825
rect 2237 3791 2271 3825
rect 2329 3791 2363 3825
rect 2421 3791 2455 3825
rect 2513 3791 2547 3825
rect 2605 3791 2639 3825
rect 2697 3791 2731 3825
rect 2789 3791 2823 3825
rect 2881 3791 2915 3825
rect 2973 3791 3007 3825
rect 3065 3791 3099 3825
rect 3157 3791 3191 3825
rect 3249 3791 3283 3825
rect 3341 3791 3375 3825
rect 3433 3791 3467 3825
rect 3525 3791 3559 3825
rect 3617 3791 3651 3825
rect 3709 3791 3743 3825
rect 3801 3791 3835 3825
rect 3893 3791 3927 3825
rect 3985 3791 4019 3825
rect 4077 3791 4111 3825
rect 4169 3791 4203 3825
rect 4261 3791 4295 3825
rect 4353 3791 4387 3825
rect 4445 3791 4479 3825
rect 4537 3791 4571 3825
rect 4629 3791 4663 3825
rect 4721 3791 4755 3825
rect 4813 3791 4847 3825
rect 4905 3791 4939 3825
rect 4997 3791 5031 3825
rect 5089 3791 5123 3825
rect 5181 3791 5215 3825
rect 5273 3791 5307 3825
rect 5365 3791 5399 3825
rect 5457 3791 5491 3825
rect 5549 3791 5583 3825
rect 5641 3791 5675 3825
rect 5733 3791 5767 3825
rect 5825 3791 5859 3825
rect 5917 3791 5951 3825
rect 6009 3791 6043 3825
rect 6101 3791 6135 3825
rect 6193 3791 6227 3825
rect 6285 3791 6319 3825
rect 6377 3791 6411 3825
rect 6469 3791 6503 3825
rect 6561 3791 6595 3825
rect 6653 3791 6687 3825
rect 6745 3791 6779 3825
rect 6837 3791 6871 3825
rect 6929 3791 6963 3825
rect 7021 3791 7055 3825
rect 7113 3791 7147 3825
rect 7205 3791 7239 3825
rect 7297 3791 7331 3825
rect 7389 3791 7423 3825
rect 7481 3791 7515 3825
rect 7573 3791 7607 3825
rect 7665 3791 7699 3825
rect 7757 3791 7791 3825
rect 7849 3791 7883 3825
rect 7941 3791 7975 3825
rect 8033 3791 8067 3825
rect 8125 3791 8159 3825
rect 8217 3791 8251 3825
rect 8309 3791 8343 3825
rect 8401 3791 8435 3825
rect 8493 3791 8527 3825
rect 8585 3791 8619 3825
rect 8677 3791 8711 3825
rect 8769 3791 8803 3825
rect 8861 3791 8895 3825
rect 8953 3791 8987 3825
rect 9045 3791 9079 3825
rect 9137 3791 9171 3825
rect 9229 3791 9263 3825
rect 9321 3791 9355 3825
rect 9413 3791 9447 3825
rect 9505 3791 9539 3825
rect 9597 3791 9631 3825
rect 9689 3791 9723 3825
rect 9781 3791 9815 3825
rect 9873 3791 9907 3825
rect 9965 3791 9999 3825
rect 10057 3791 10091 3825
rect 10149 3791 10183 3825
rect 10241 3791 10275 3825
rect 10333 3791 10367 3825
rect 10425 3791 10459 3825
rect 10517 3791 10551 3825
rect 10609 3791 10643 3825
rect 10701 3791 10735 3825
rect 10793 3791 10827 3825
rect 10885 3791 10919 3825
rect 10977 3791 11011 3825
rect 11069 3791 11103 3825
rect 11161 3791 11195 3825
rect 11253 3791 11287 3825
rect 11345 3791 11379 3825
rect 11437 3791 11471 3825
rect 11529 3791 11563 3825
rect 11621 3791 11655 3825
rect 11713 3791 11747 3825
rect 11805 3791 11839 3825
rect 11897 3791 11931 3825
rect 11989 3791 12023 3825
rect 12081 3791 12115 3825
rect 12173 3791 12207 3825
rect 12265 3791 12299 3825
rect 12357 3791 12391 3825
rect 12449 3791 12483 3825
rect 12541 3791 12575 3825
rect 12633 3791 12667 3825
rect 12725 3791 12759 3825
rect 12817 3791 12851 3825
rect 12909 3791 12943 3825
rect 13001 3791 13035 3825
rect 13093 3791 13127 3825
rect 13185 3791 13219 3825
rect 13277 3791 13311 3825
rect 13369 3791 13403 3825
rect 13461 3791 13495 3825
rect 13553 3791 13587 3825
rect 13645 3791 13679 3825
rect 13737 3791 13771 3825
rect 13829 3791 13863 3825
rect 13921 3791 13955 3825
rect 14013 3791 14047 3825
rect 14105 3791 14139 3825
rect 14197 3791 14231 3825
rect 14289 3791 14323 3825
rect 14381 3791 14415 3825
rect 14473 3791 14507 3825
rect 14565 3791 14599 3825
rect 14657 3791 14691 3825
rect 14749 3791 14783 3825
rect 14841 3791 14875 3825
rect 14933 3791 14967 3825
rect 15025 3791 15059 3825
rect 15117 3791 15151 3825
rect 15209 3791 15243 3825
rect 15301 3791 15335 3825
rect 15393 3791 15427 3825
rect 15485 3791 15519 3825
rect 15577 3791 15611 3825
rect 15669 3791 15703 3825
rect 15761 3791 15795 3825
rect 15853 3791 15887 3825
rect 15945 3791 15979 3825
rect 16037 3791 16071 3825
rect 16129 3791 16163 3825
rect 16221 3791 16255 3825
rect 16313 3791 16347 3825
rect 16405 3791 16439 3825
rect 16497 3791 16531 3825
rect 16589 3791 16623 3825
rect 16681 3791 16715 3825
rect 16773 3791 16807 3825
rect 16865 3791 16899 3825
rect 16957 3791 16991 3825
rect 17049 3791 17083 3825
rect 17141 3791 17175 3825
rect 17233 3791 17267 3825
rect 17325 3791 17359 3825
rect 17417 3791 17451 3825
rect 17509 3791 17543 3825
rect 17601 3791 17635 3825
rect 17693 3791 17727 3825
rect 17785 3791 17819 3825
rect 17877 3791 17911 3825
rect 17969 3791 18003 3825
rect 18061 3791 18095 3825
rect 18153 3791 18187 3825
rect 18245 3791 18279 3825
rect 18337 3791 18371 3825
rect 18429 3791 18463 3825
rect 18521 3791 18555 3825
rect 18613 3791 18647 3825
rect 18705 3791 18739 3825
rect 18797 3791 18831 3825
rect 1685 3553 1719 3587
rect 1778 3494 1790 3519
rect 1790 3494 1812 3519
rect 1778 3485 1812 3494
rect 1859 3639 1893 3655
rect 1859 3621 1893 3639
rect 1948 3689 1982 3723
rect 2237 3621 2271 3655
rect 2145 3485 2179 3519
rect 2861 3629 2895 3655
rect 2861 3621 2892 3629
rect 2892 3621 2895 3629
rect 2417 3417 2451 3451
rect 2489 3433 2513 3451
rect 2513 3433 2523 3451
rect 2489 3417 2523 3433
rect 2861 3503 2895 3519
rect 2861 3485 2887 3503
rect 2887 3485 2895 3503
rect 3077 3505 3111 3514
rect 3077 3480 3093 3505
rect 3093 3480 3111 3505
rect 3137 3417 3171 3451
rect 4997 3705 5031 3723
rect 4997 3689 5024 3705
rect 5024 3689 5031 3705
rect 3433 3373 3461 3383
rect 3461 3373 3467 3383
rect 3433 3349 3467 3373
rect 6285 3513 6319 3519
rect 6285 3485 6311 3513
rect 6311 3485 6319 3513
rect 6745 3513 6779 3519
rect 6745 3485 6748 3513
rect 6748 3485 6779 3513
rect 6838 3494 6850 3519
rect 6850 3494 6872 3519
rect 6838 3485 6872 3494
rect 6919 3639 6953 3655
rect 6919 3621 6953 3639
rect 7021 3417 7055 3451
rect 7297 3621 7331 3655
rect 7205 3485 7239 3519
rect 7921 3629 7955 3655
rect 7921 3621 7952 3629
rect 7952 3621 7955 3629
rect 7477 3417 7511 3451
rect 7549 3433 7573 3451
rect 7573 3433 7583 3451
rect 7549 3417 7583 3433
rect 7921 3503 7955 3519
rect 7921 3485 7947 3503
rect 7947 3485 7955 3503
rect 8493 3645 8527 3655
rect 8493 3621 8521 3645
rect 8521 3621 8527 3645
rect 8137 3505 8171 3514
rect 8137 3480 8153 3505
rect 8153 3480 8171 3505
rect 8197 3417 8231 3451
rect 9321 3644 9355 3655
rect 9321 3621 9322 3644
rect 9322 3621 9355 3644
rect 9137 3513 9171 3519
rect 9137 3485 9145 3513
rect 9145 3485 9171 3513
rect 10241 3513 10275 3519
rect 10241 3485 10267 3513
rect 10267 3485 10275 3513
rect 11161 3626 11189 3655
rect 11189 3626 11195 3655
rect 11161 3621 11195 3626
rect 10977 3513 11011 3519
rect 10977 3485 10985 3513
rect 10985 3485 11011 3513
rect 10057 3353 10063 3383
rect 10063 3353 10091 3383
rect 10057 3349 10091 3353
rect 11989 3645 12023 3655
rect 11989 3621 11995 3645
rect 11995 3621 12023 3645
rect 12561 3629 12595 3655
rect 12561 3621 12564 3629
rect 12564 3621 12595 3629
rect 12345 3505 12379 3514
rect 12345 3480 12363 3505
rect 12363 3480 12379 3505
rect 12285 3417 12319 3451
rect 12561 3503 12595 3519
rect 12561 3485 12569 3503
rect 12569 3485 12595 3503
rect 13185 3621 13219 3655
rect 12933 3433 12943 3451
rect 12943 3433 12967 3451
rect 12933 3417 12967 3433
rect 13005 3417 13039 3451
rect 13277 3485 13311 3519
rect 13563 3639 13597 3655
rect 13563 3621 13597 3639
rect 13461 3417 13495 3451
rect 13644 3494 13666 3519
rect 13666 3494 13678 3519
rect 13644 3485 13678 3494
rect 13737 3553 13771 3587
rect 1133 3247 1167 3281
rect 1225 3247 1259 3281
rect 1317 3247 1351 3281
rect 1409 3247 1443 3281
rect 1501 3247 1535 3281
rect 1593 3247 1627 3281
rect 1685 3247 1719 3281
rect 1777 3247 1811 3281
rect 1869 3247 1903 3281
rect 1961 3247 1995 3281
rect 2053 3247 2087 3281
rect 2145 3247 2179 3281
rect 2237 3247 2271 3281
rect 2329 3247 2363 3281
rect 2421 3247 2455 3281
rect 2513 3247 2547 3281
rect 2605 3247 2639 3281
rect 2697 3247 2731 3281
rect 2789 3247 2823 3281
rect 2881 3247 2915 3281
rect 2973 3247 3007 3281
rect 3065 3247 3099 3281
rect 3157 3247 3191 3281
rect 3249 3247 3283 3281
rect 3341 3247 3375 3281
rect 3433 3247 3467 3281
rect 3525 3247 3559 3281
rect 3617 3247 3651 3281
rect 3709 3247 3743 3281
rect 3801 3247 3835 3281
rect 3893 3247 3927 3281
rect 3985 3247 4019 3281
rect 4077 3247 4111 3281
rect 4169 3247 4203 3281
rect 4261 3247 4295 3281
rect 4353 3247 4387 3281
rect 4445 3247 4479 3281
rect 4537 3247 4571 3281
rect 4629 3247 4663 3281
rect 4721 3247 4755 3281
rect 4813 3247 4847 3281
rect 4905 3247 4939 3281
rect 4997 3247 5031 3281
rect 5089 3247 5123 3281
rect 5181 3247 5215 3281
rect 5273 3247 5307 3281
rect 5365 3247 5399 3281
rect 5457 3247 5491 3281
rect 5549 3247 5583 3281
rect 5641 3247 5675 3281
rect 5733 3247 5767 3281
rect 5825 3247 5859 3281
rect 5917 3247 5951 3281
rect 6009 3247 6043 3281
rect 6101 3247 6135 3281
rect 6193 3247 6227 3281
rect 6285 3247 6319 3281
rect 6377 3247 6411 3281
rect 6469 3247 6503 3281
rect 6561 3247 6595 3281
rect 6653 3247 6687 3281
rect 6745 3247 6779 3281
rect 6837 3247 6871 3281
rect 6929 3247 6963 3281
rect 7021 3247 7055 3281
rect 7113 3247 7147 3281
rect 7205 3247 7239 3281
rect 7297 3247 7331 3281
rect 7389 3247 7423 3281
rect 7481 3247 7515 3281
rect 7573 3247 7607 3281
rect 7665 3247 7699 3281
rect 7757 3247 7791 3281
rect 7849 3247 7883 3281
rect 7941 3247 7975 3281
rect 8033 3247 8067 3281
rect 8125 3247 8159 3281
rect 8217 3247 8251 3281
rect 8309 3247 8343 3281
rect 8401 3247 8435 3281
rect 8493 3247 8527 3281
rect 8585 3247 8619 3281
rect 8677 3247 8711 3281
rect 8769 3247 8803 3281
rect 8861 3247 8895 3281
rect 8953 3247 8987 3281
rect 9045 3247 9079 3281
rect 9137 3247 9171 3281
rect 9229 3247 9263 3281
rect 9321 3247 9355 3281
rect 9413 3247 9447 3281
rect 9505 3247 9539 3281
rect 9597 3247 9631 3281
rect 9689 3247 9723 3281
rect 9781 3247 9815 3281
rect 9873 3247 9907 3281
rect 9965 3247 9999 3281
rect 10057 3247 10091 3281
rect 10149 3247 10183 3281
rect 10241 3247 10275 3281
rect 10333 3247 10367 3281
rect 10425 3247 10459 3281
rect 10517 3247 10551 3281
rect 10609 3247 10643 3281
rect 10701 3247 10735 3281
rect 10793 3247 10827 3281
rect 10885 3247 10919 3281
rect 10977 3247 11011 3281
rect 11069 3247 11103 3281
rect 11161 3247 11195 3281
rect 11253 3247 11287 3281
rect 11345 3247 11379 3281
rect 11437 3247 11471 3281
rect 11529 3247 11563 3281
rect 11621 3247 11655 3281
rect 11713 3247 11747 3281
rect 11805 3247 11839 3281
rect 11897 3247 11931 3281
rect 11989 3247 12023 3281
rect 12081 3247 12115 3281
rect 12173 3247 12207 3281
rect 12265 3247 12299 3281
rect 12357 3247 12391 3281
rect 12449 3247 12483 3281
rect 12541 3247 12575 3281
rect 12633 3247 12667 3281
rect 12725 3247 12759 3281
rect 12817 3247 12851 3281
rect 12909 3247 12943 3281
rect 13001 3247 13035 3281
rect 13093 3247 13127 3281
rect 13185 3247 13219 3281
rect 13277 3247 13311 3281
rect 13369 3247 13403 3281
rect 13461 3247 13495 3281
rect 13553 3247 13587 3281
rect 13645 3247 13679 3281
rect 13737 3247 13771 3281
rect 13829 3247 13863 3281
rect 13921 3247 13955 3281
rect 14013 3247 14047 3281
rect 14105 3247 14139 3281
rect 14197 3247 14231 3281
rect 14289 3247 14323 3281
rect 14381 3247 14415 3281
rect 14473 3247 14507 3281
rect 14565 3247 14599 3281
rect 14657 3247 14691 3281
rect 14749 3247 14783 3281
rect 14841 3247 14875 3281
rect 14933 3247 14967 3281
rect 15025 3247 15059 3281
rect 15117 3247 15151 3281
rect 15209 3247 15243 3281
rect 15301 3247 15335 3281
rect 15393 3247 15427 3281
rect 15485 3247 15519 3281
rect 15577 3247 15611 3281
rect 15669 3247 15703 3281
rect 15761 3247 15795 3281
rect 15853 3247 15887 3281
rect 15945 3247 15979 3281
rect 16037 3247 16071 3281
rect 16129 3247 16163 3281
rect 16221 3247 16255 3281
rect 16313 3247 16347 3281
rect 16405 3247 16439 3281
rect 16497 3247 16531 3281
rect 16589 3247 16623 3281
rect 16681 3247 16715 3281
rect 16773 3247 16807 3281
rect 16865 3247 16899 3281
rect 16957 3247 16991 3281
rect 17049 3247 17083 3281
rect 17141 3247 17175 3281
rect 17233 3247 17267 3281
rect 17325 3247 17359 3281
rect 17417 3247 17451 3281
rect 17509 3247 17543 3281
rect 17601 3247 17635 3281
rect 17693 3247 17727 3281
rect 17785 3247 17819 3281
rect 17877 3247 17911 3281
rect 17969 3247 18003 3281
rect 18061 3247 18095 3281
rect 18153 3247 18187 3281
rect 18245 3247 18279 3281
rect 18337 3247 18371 3281
rect 18429 3247 18463 3281
rect 18521 3247 18555 3281
rect 18613 3247 18647 3281
rect 18705 3247 18739 3281
rect 18797 3247 18831 3281
rect 1961 3155 1995 3179
rect 1961 3145 1967 3155
rect 1967 3145 1995 3155
rect 2257 3077 2291 3111
rect 2317 3023 2335 3048
rect 2335 3023 2351 3048
rect 2317 3014 2351 3023
rect 2533 3025 2541 3043
rect 2541 3025 2567 3043
rect 2533 3009 2567 3025
rect 2905 3095 2939 3111
rect 2905 3077 2915 3095
rect 2915 3077 2939 3095
rect 2977 3077 3011 3111
rect 2533 2899 2536 2907
rect 2536 2899 2567 2907
rect 2533 2873 2567 2899
rect 3249 3009 3283 3043
rect 3157 2873 3191 2907
rect 3433 3077 3467 3111
rect 3535 2889 3569 2907
rect 3535 2873 3569 2889
rect 3616 3034 3650 3043
rect 3616 3009 3638 3034
rect 3638 3009 3650 3034
rect 3709 3015 3740 3043
rect 3740 3015 3743 3043
rect 3709 3009 3743 3015
rect 4169 3034 4203 3043
rect 4169 3009 4172 3034
rect 4172 3009 4203 3034
rect 4262 2873 4296 2907
rect 4354 3077 4388 3111
rect 4537 3009 4571 3043
rect 4726 3095 4760 3111
rect 4726 3077 4740 3095
rect 4740 3077 4760 3095
rect 4910 3085 4944 3111
rect 4910 3077 4912 3085
rect 4912 3077 4944 3085
rect 4634 2873 4668 2907
rect 5190 3029 5224 3043
rect 5190 3009 5224 3029
rect 5562 3077 5596 3111
rect 5190 2899 5192 2907
rect 5192 2899 5224 2907
rect 5190 2873 5224 2899
rect 7205 3155 7239 3179
rect 7205 3145 7211 3155
rect 7211 3145 7239 3155
rect 5963 2941 5997 2975
rect 7501 3077 7535 3111
rect 7561 3023 7579 3048
rect 7579 3023 7595 3048
rect 7561 3014 7595 3023
rect 7777 3025 7785 3043
rect 7785 3025 7811 3043
rect 7777 3009 7811 3025
rect 8149 3095 8183 3111
rect 8149 3077 8159 3095
rect 8159 3077 8183 3095
rect 8221 3077 8255 3111
rect 7777 2899 7780 2907
rect 7780 2899 7811 2907
rect 7777 2873 7811 2899
rect 8493 3009 8527 3043
rect 8401 2873 8435 2907
rect 8689 3077 8723 3111
rect 8779 2889 8813 2907
rect 8779 2873 8813 2889
rect 8860 3034 8894 3043
rect 8860 3009 8882 3034
rect 8882 3009 8894 3034
rect 9413 3077 9447 3111
rect 8953 2941 8987 2975
rect 12009 3077 12043 3111
rect 12069 3023 12087 3048
rect 12087 3023 12103 3048
rect 12069 3014 12103 3023
rect 10701 2873 10735 2907
rect 11713 2883 11719 2907
rect 11719 2883 11747 2907
rect 11713 2873 11747 2883
rect 12285 3025 12293 3043
rect 12293 3025 12319 3043
rect 12285 3009 12319 3025
rect 12657 3095 12691 3111
rect 12657 3077 12667 3095
rect 12667 3077 12691 3095
rect 12729 3077 12763 3111
rect 12285 2899 12288 2907
rect 12288 2899 12319 2907
rect 12285 2873 12319 2899
rect 13001 3009 13035 3043
rect 12909 2873 12943 2907
rect 13185 3077 13219 3111
rect 13287 2889 13321 2907
rect 13287 2873 13321 2889
rect 13368 3034 13402 3043
rect 13368 3009 13390 3034
rect 13390 3009 13402 3034
rect 13461 2941 13495 2975
rect 13921 3015 13929 3043
rect 13929 3015 13955 3043
rect 13921 3009 13955 3015
rect 14105 2837 14139 2839
rect 14105 2805 14106 2837
rect 14106 2805 14139 2837
rect 1133 2703 1167 2737
rect 1225 2703 1259 2737
rect 1317 2703 1351 2737
rect 1409 2703 1443 2737
rect 1501 2703 1535 2737
rect 1593 2703 1627 2737
rect 1685 2703 1719 2737
rect 1777 2703 1811 2737
rect 1869 2703 1903 2737
rect 1961 2703 1995 2737
rect 2053 2703 2087 2737
rect 2145 2703 2179 2737
rect 2237 2703 2271 2737
rect 2329 2703 2363 2737
rect 2421 2703 2455 2737
rect 2513 2703 2547 2737
rect 2605 2703 2639 2737
rect 2697 2703 2731 2737
rect 2789 2703 2823 2737
rect 2881 2703 2915 2737
rect 2973 2703 3007 2737
rect 3065 2703 3099 2737
rect 3157 2703 3191 2737
rect 3249 2703 3283 2737
rect 3341 2703 3375 2737
rect 3433 2703 3467 2737
rect 3525 2703 3559 2737
rect 3617 2703 3651 2737
rect 3709 2703 3743 2737
rect 3801 2703 3835 2737
rect 3893 2703 3927 2737
rect 3985 2703 4019 2737
rect 4077 2703 4111 2737
rect 4169 2703 4203 2737
rect 4261 2703 4295 2737
rect 4353 2703 4387 2737
rect 4445 2703 4479 2737
rect 4537 2703 4571 2737
rect 4629 2703 4663 2737
rect 4721 2703 4755 2737
rect 4813 2703 4847 2737
rect 4905 2703 4939 2737
rect 4997 2703 5031 2737
rect 5089 2703 5123 2737
rect 5181 2703 5215 2737
rect 5273 2703 5307 2737
rect 5365 2703 5399 2737
rect 5457 2703 5491 2737
rect 5549 2703 5583 2737
rect 5641 2703 5675 2737
rect 5733 2703 5767 2737
rect 5825 2703 5859 2737
rect 5917 2703 5951 2737
rect 6009 2703 6043 2737
rect 6101 2703 6135 2737
rect 6193 2703 6227 2737
rect 6285 2703 6319 2737
rect 6377 2703 6411 2737
rect 6469 2703 6503 2737
rect 6561 2703 6595 2737
rect 6653 2703 6687 2737
rect 6745 2703 6779 2737
rect 6837 2703 6871 2737
rect 6929 2703 6963 2737
rect 7021 2703 7055 2737
rect 7113 2703 7147 2737
rect 7205 2703 7239 2737
rect 7297 2703 7331 2737
rect 7389 2703 7423 2737
rect 7481 2703 7515 2737
rect 7573 2703 7607 2737
rect 7665 2703 7699 2737
rect 7757 2703 7791 2737
rect 7849 2703 7883 2737
rect 7941 2703 7975 2737
rect 8033 2703 8067 2737
rect 8125 2703 8159 2737
rect 8217 2703 8251 2737
rect 8309 2703 8343 2737
rect 8401 2703 8435 2737
rect 8493 2703 8527 2737
rect 8585 2703 8619 2737
rect 8677 2703 8711 2737
rect 8769 2703 8803 2737
rect 8861 2703 8895 2737
rect 8953 2703 8987 2737
rect 9045 2703 9079 2737
rect 9137 2703 9171 2737
rect 9229 2703 9263 2737
rect 9321 2703 9355 2737
rect 9413 2703 9447 2737
rect 9505 2703 9539 2737
rect 9597 2703 9631 2737
rect 9689 2703 9723 2737
rect 9781 2703 9815 2737
rect 9873 2703 9907 2737
rect 9965 2703 9999 2737
rect 10057 2703 10091 2737
rect 10149 2703 10183 2737
rect 10241 2703 10275 2737
rect 10333 2703 10367 2737
rect 10425 2703 10459 2737
rect 10517 2703 10551 2737
rect 10609 2703 10643 2737
rect 10701 2703 10735 2737
rect 10793 2703 10827 2737
rect 10885 2703 10919 2737
rect 10977 2703 11011 2737
rect 11069 2703 11103 2737
rect 11161 2703 11195 2737
rect 11253 2703 11287 2737
rect 11345 2703 11379 2737
rect 11437 2703 11471 2737
rect 11529 2703 11563 2737
rect 11621 2703 11655 2737
rect 11713 2703 11747 2737
rect 11805 2703 11839 2737
rect 11897 2703 11931 2737
rect 11989 2703 12023 2737
rect 12081 2703 12115 2737
rect 12173 2703 12207 2737
rect 12265 2703 12299 2737
rect 12357 2703 12391 2737
rect 12449 2703 12483 2737
rect 12541 2703 12575 2737
rect 12633 2703 12667 2737
rect 12725 2703 12759 2737
rect 12817 2703 12851 2737
rect 12909 2703 12943 2737
rect 13001 2703 13035 2737
rect 13093 2703 13127 2737
rect 13185 2703 13219 2737
rect 13277 2703 13311 2737
rect 13369 2703 13403 2737
rect 13461 2703 13495 2737
rect 13553 2703 13587 2737
rect 13645 2703 13679 2737
rect 13737 2703 13771 2737
rect 13829 2703 13863 2737
rect 13921 2703 13955 2737
rect 14013 2703 14047 2737
rect 14105 2703 14139 2737
rect 14197 2703 14231 2737
rect 14289 2703 14323 2737
rect 14381 2703 14415 2737
rect 14473 2703 14507 2737
rect 14565 2703 14599 2737
rect 14657 2703 14691 2737
rect 14749 2703 14783 2737
rect 14841 2703 14875 2737
rect 14933 2703 14967 2737
rect 15025 2703 15059 2737
rect 15117 2703 15151 2737
rect 15209 2703 15243 2737
rect 15301 2703 15335 2737
rect 15393 2703 15427 2737
rect 15485 2703 15519 2737
rect 15577 2703 15611 2737
rect 15669 2703 15703 2737
rect 15761 2703 15795 2737
rect 15853 2703 15887 2737
rect 15945 2703 15979 2737
rect 16037 2703 16071 2737
rect 16129 2703 16163 2737
rect 16221 2703 16255 2737
rect 16313 2703 16347 2737
rect 16405 2703 16439 2737
rect 16497 2703 16531 2737
rect 16589 2703 16623 2737
rect 16681 2703 16715 2737
rect 16773 2703 16807 2737
rect 16865 2703 16899 2737
rect 16957 2703 16991 2737
rect 17049 2703 17083 2737
rect 17141 2703 17175 2737
rect 17233 2703 17267 2737
rect 17325 2703 17359 2737
rect 17417 2703 17451 2737
rect 17509 2703 17543 2737
rect 17601 2703 17635 2737
rect 17693 2703 17727 2737
rect 17785 2703 17819 2737
rect 17877 2703 17911 2737
rect 17969 2703 18003 2737
rect 18061 2703 18095 2737
rect 18153 2703 18187 2737
rect 18245 2703 18279 2737
rect 18337 2703 18371 2737
rect 18429 2703 18463 2737
rect 18521 2703 18555 2737
rect 18613 2703 18647 2737
rect 18705 2703 18739 2737
rect 18797 2703 18831 2737
rect 1685 2465 1719 2499
rect 1778 2406 1790 2431
rect 1790 2406 1812 2431
rect 1778 2397 1812 2406
rect 1859 2551 1893 2567
rect 1859 2533 1893 2551
rect 1961 2329 1995 2363
rect 2237 2533 2271 2567
rect 2145 2397 2179 2431
rect 2861 2541 2895 2567
rect 2861 2533 2892 2541
rect 2892 2533 2895 2541
rect 2417 2329 2451 2363
rect 2489 2345 2513 2363
rect 2513 2345 2523 2363
rect 2489 2329 2523 2345
rect 2861 2415 2895 2431
rect 2861 2397 2887 2415
rect 2887 2397 2895 2415
rect 3433 2625 3467 2635
rect 3433 2601 3461 2625
rect 3461 2601 3467 2625
rect 3077 2417 3111 2426
rect 3077 2392 3093 2417
rect 3093 2392 3111 2417
rect 3137 2329 3171 2363
rect 4261 2465 4295 2499
rect 4354 2406 4366 2431
rect 4366 2406 4388 2431
rect 4354 2397 4388 2406
rect 4435 2551 4469 2567
rect 4435 2533 4469 2551
rect 4537 2465 4571 2499
rect 4813 2533 4847 2567
rect 4721 2397 4755 2431
rect 5437 2541 5471 2567
rect 5437 2533 5468 2541
rect 5468 2533 5471 2541
rect 4993 2329 5027 2363
rect 5065 2345 5089 2363
rect 5089 2345 5099 2363
rect 5065 2329 5099 2345
rect 5437 2415 5471 2431
rect 5437 2397 5463 2415
rect 5463 2397 5471 2415
rect 6009 2625 6043 2635
rect 6009 2601 6037 2625
rect 6037 2601 6043 2625
rect 5653 2417 5687 2426
rect 5653 2392 5669 2417
rect 5669 2392 5687 2417
rect 5713 2329 5747 2363
rect 9137 2625 9171 2635
rect 9137 2601 9143 2625
rect 9143 2601 9171 2625
rect 9709 2541 9743 2567
rect 9709 2533 9712 2541
rect 9712 2533 9743 2541
rect 9493 2417 9527 2426
rect 9493 2392 9511 2417
rect 9511 2392 9527 2417
rect 9433 2329 9467 2363
rect 9709 2415 9743 2431
rect 9709 2397 9717 2415
rect 9717 2397 9743 2415
rect 10333 2533 10367 2567
rect 10081 2345 10091 2363
rect 10091 2345 10115 2363
rect 10081 2329 10115 2345
rect 10153 2329 10187 2363
rect 10425 2397 10459 2431
rect 10711 2551 10745 2567
rect 10711 2533 10745 2551
rect 10609 2465 10643 2499
rect 10792 2406 10814 2431
rect 10814 2406 10826 2431
rect 10792 2397 10826 2406
rect 10885 2425 10919 2431
rect 10885 2397 10916 2425
rect 10916 2397 10919 2425
rect 11989 2557 12023 2567
rect 11989 2533 11995 2557
rect 11995 2533 12023 2557
rect 12561 2541 12595 2567
rect 12561 2533 12564 2541
rect 12564 2533 12595 2541
rect 12345 2417 12379 2426
rect 12345 2392 12363 2417
rect 12363 2392 12379 2417
rect 12285 2329 12319 2363
rect 12561 2415 12595 2431
rect 12561 2397 12569 2415
rect 12569 2397 12595 2415
rect 13185 2533 13219 2567
rect 12933 2345 12943 2363
rect 12943 2345 12967 2363
rect 12933 2329 12967 2345
rect 13005 2329 13039 2363
rect 13277 2397 13311 2431
rect 13563 2551 13597 2567
rect 13563 2533 13597 2551
rect 13461 2465 13495 2499
rect 13644 2406 13666 2431
rect 13666 2406 13678 2431
rect 13644 2397 13678 2406
rect 13737 2465 13771 2499
rect 14289 2625 14323 2635
rect 14289 2601 14295 2625
rect 14295 2601 14323 2625
rect 14861 2541 14895 2567
rect 14861 2533 14864 2541
rect 14864 2533 14895 2541
rect 14645 2417 14679 2426
rect 14645 2392 14663 2417
rect 14663 2392 14679 2417
rect 14585 2329 14619 2363
rect 14861 2415 14895 2431
rect 14861 2397 14869 2415
rect 14869 2397 14895 2415
rect 15485 2533 15519 2567
rect 15233 2345 15243 2363
rect 15243 2345 15267 2363
rect 15233 2329 15267 2345
rect 15305 2329 15339 2363
rect 15577 2397 15611 2431
rect 15863 2551 15897 2567
rect 15863 2533 15897 2551
rect 15761 2329 15795 2363
rect 15944 2406 15966 2431
rect 15966 2406 15978 2431
rect 15944 2397 15978 2406
rect 16037 2465 16071 2499
rect 17509 2425 17543 2431
rect 17509 2397 17517 2425
rect 17517 2397 17543 2425
rect 17693 2265 17694 2295
rect 17694 2265 17727 2295
rect 17693 2261 17727 2265
rect 1133 2159 1167 2193
rect 1225 2159 1259 2193
rect 1317 2159 1351 2193
rect 1409 2159 1443 2193
rect 1501 2159 1535 2193
rect 1593 2159 1627 2193
rect 1685 2159 1719 2193
rect 1777 2159 1811 2193
rect 1869 2159 1903 2193
rect 1961 2159 1995 2193
rect 2053 2159 2087 2193
rect 2145 2159 2179 2193
rect 2237 2159 2271 2193
rect 2329 2159 2363 2193
rect 2421 2159 2455 2193
rect 2513 2159 2547 2193
rect 2605 2159 2639 2193
rect 2697 2159 2731 2193
rect 2789 2159 2823 2193
rect 2881 2159 2915 2193
rect 2973 2159 3007 2193
rect 3065 2159 3099 2193
rect 3157 2159 3191 2193
rect 3249 2159 3283 2193
rect 3341 2159 3375 2193
rect 3433 2159 3467 2193
rect 3525 2159 3559 2193
rect 3617 2159 3651 2193
rect 3709 2159 3743 2193
rect 3801 2159 3835 2193
rect 3893 2159 3927 2193
rect 3985 2159 4019 2193
rect 4077 2159 4111 2193
rect 4169 2159 4203 2193
rect 4261 2159 4295 2193
rect 4353 2159 4387 2193
rect 4445 2159 4479 2193
rect 4537 2159 4571 2193
rect 4629 2159 4663 2193
rect 4721 2159 4755 2193
rect 4813 2159 4847 2193
rect 4905 2159 4939 2193
rect 4997 2159 5031 2193
rect 5089 2159 5123 2193
rect 5181 2159 5215 2193
rect 5273 2159 5307 2193
rect 5365 2159 5399 2193
rect 5457 2159 5491 2193
rect 5549 2159 5583 2193
rect 5641 2159 5675 2193
rect 5733 2159 5767 2193
rect 5825 2159 5859 2193
rect 5917 2159 5951 2193
rect 6009 2159 6043 2193
rect 6101 2159 6135 2193
rect 6193 2159 6227 2193
rect 6285 2159 6319 2193
rect 6377 2159 6411 2193
rect 6469 2159 6503 2193
rect 6561 2159 6595 2193
rect 6653 2159 6687 2193
rect 6745 2159 6779 2193
rect 6837 2159 6871 2193
rect 6929 2159 6963 2193
rect 7021 2159 7055 2193
rect 7113 2159 7147 2193
rect 7205 2159 7239 2193
rect 7297 2159 7331 2193
rect 7389 2159 7423 2193
rect 7481 2159 7515 2193
rect 7573 2159 7607 2193
rect 7665 2159 7699 2193
rect 7757 2159 7791 2193
rect 7849 2159 7883 2193
rect 7941 2159 7975 2193
rect 8033 2159 8067 2193
rect 8125 2159 8159 2193
rect 8217 2159 8251 2193
rect 8309 2159 8343 2193
rect 8401 2159 8435 2193
rect 8493 2159 8527 2193
rect 8585 2159 8619 2193
rect 8677 2159 8711 2193
rect 8769 2159 8803 2193
rect 8861 2159 8895 2193
rect 8953 2159 8987 2193
rect 9045 2159 9079 2193
rect 9137 2159 9171 2193
rect 9229 2159 9263 2193
rect 9321 2159 9355 2193
rect 9413 2159 9447 2193
rect 9505 2159 9539 2193
rect 9597 2159 9631 2193
rect 9689 2159 9723 2193
rect 9781 2159 9815 2193
rect 9873 2159 9907 2193
rect 9965 2159 9999 2193
rect 10057 2159 10091 2193
rect 10149 2159 10183 2193
rect 10241 2159 10275 2193
rect 10333 2159 10367 2193
rect 10425 2159 10459 2193
rect 10517 2159 10551 2193
rect 10609 2159 10643 2193
rect 10701 2159 10735 2193
rect 10793 2159 10827 2193
rect 10885 2159 10919 2193
rect 10977 2159 11011 2193
rect 11069 2159 11103 2193
rect 11161 2159 11195 2193
rect 11253 2159 11287 2193
rect 11345 2159 11379 2193
rect 11437 2159 11471 2193
rect 11529 2159 11563 2193
rect 11621 2159 11655 2193
rect 11713 2159 11747 2193
rect 11805 2159 11839 2193
rect 11897 2159 11931 2193
rect 11989 2159 12023 2193
rect 12081 2159 12115 2193
rect 12173 2159 12207 2193
rect 12265 2159 12299 2193
rect 12357 2159 12391 2193
rect 12449 2159 12483 2193
rect 12541 2159 12575 2193
rect 12633 2159 12667 2193
rect 12725 2159 12759 2193
rect 12817 2159 12851 2193
rect 12909 2159 12943 2193
rect 13001 2159 13035 2193
rect 13093 2159 13127 2193
rect 13185 2159 13219 2193
rect 13277 2159 13311 2193
rect 13369 2159 13403 2193
rect 13461 2159 13495 2193
rect 13553 2159 13587 2193
rect 13645 2159 13679 2193
rect 13737 2159 13771 2193
rect 13829 2159 13863 2193
rect 13921 2159 13955 2193
rect 14013 2159 14047 2193
rect 14105 2159 14139 2193
rect 14197 2159 14231 2193
rect 14289 2159 14323 2193
rect 14381 2159 14415 2193
rect 14473 2159 14507 2193
rect 14565 2159 14599 2193
rect 14657 2159 14691 2193
rect 14749 2159 14783 2193
rect 14841 2159 14875 2193
rect 14933 2159 14967 2193
rect 15025 2159 15059 2193
rect 15117 2159 15151 2193
rect 15209 2159 15243 2193
rect 15301 2159 15335 2193
rect 15393 2159 15427 2193
rect 15485 2159 15519 2193
rect 15577 2159 15611 2193
rect 15669 2159 15703 2193
rect 15761 2159 15795 2193
rect 15853 2159 15887 2193
rect 15945 2159 15979 2193
rect 16037 2159 16071 2193
rect 16129 2159 16163 2193
rect 16221 2159 16255 2193
rect 16313 2159 16347 2193
rect 16405 2159 16439 2193
rect 16497 2159 16531 2193
rect 16589 2159 16623 2193
rect 16681 2159 16715 2193
rect 16773 2159 16807 2193
rect 16865 2159 16899 2193
rect 16957 2159 16991 2193
rect 17049 2159 17083 2193
rect 17141 2159 17175 2193
rect 17233 2159 17267 2193
rect 17325 2159 17359 2193
rect 17417 2159 17451 2193
rect 17509 2159 17543 2193
rect 17601 2159 17635 2193
rect 17693 2159 17727 2193
rect 17785 2159 17819 2193
rect 17877 2159 17911 2193
rect 17969 2159 18003 2193
rect 18061 2159 18095 2193
rect 18153 2159 18187 2193
rect 18245 2159 18279 2193
rect 18337 2159 18371 2193
rect 18429 2159 18463 2193
rect 18521 2159 18555 2193
rect 18613 2159 18647 2193
rect 18705 2159 18739 2193
rect 18797 2159 18831 2193
<< metal1 >>
rect 1104 7642 19019 7664
rect 1104 7633 5388 7642
rect 1104 7599 1133 7633
rect 1167 7599 1225 7633
rect 1259 7599 1317 7633
rect 1351 7599 1409 7633
rect 1443 7599 1501 7633
rect 1535 7599 1593 7633
rect 1627 7599 1685 7633
rect 1719 7599 1777 7633
rect 1811 7599 1869 7633
rect 1903 7599 1961 7633
rect 1995 7599 2053 7633
rect 2087 7599 2145 7633
rect 2179 7599 2237 7633
rect 2271 7599 2329 7633
rect 2363 7599 2421 7633
rect 2455 7599 2513 7633
rect 2547 7599 2605 7633
rect 2639 7599 2697 7633
rect 2731 7599 2789 7633
rect 2823 7599 2881 7633
rect 2915 7599 2973 7633
rect 3007 7599 3065 7633
rect 3099 7599 3157 7633
rect 3191 7599 3249 7633
rect 3283 7599 3341 7633
rect 3375 7599 3433 7633
rect 3467 7599 3525 7633
rect 3559 7599 3617 7633
rect 3651 7599 3709 7633
rect 3743 7599 3801 7633
rect 3835 7599 3893 7633
rect 3927 7599 3985 7633
rect 4019 7599 4077 7633
rect 4111 7599 4169 7633
rect 4203 7599 4261 7633
rect 4295 7599 4353 7633
rect 4387 7599 4445 7633
rect 4479 7599 4537 7633
rect 4571 7599 4629 7633
rect 4663 7599 4721 7633
rect 4755 7599 4813 7633
rect 4847 7599 4905 7633
rect 4939 7599 4997 7633
rect 5031 7599 5089 7633
rect 5123 7599 5181 7633
rect 5215 7599 5273 7633
rect 5307 7599 5365 7633
rect 1104 7590 5388 7599
rect 5440 7590 5452 7642
rect 5504 7590 5516 7642
rect 5568 7633 5580 7642
rect 5632 7633 5644 7642
rect 5696 7633 9827 7642
rect 9879 7633 9891 7642
rect 5632 7599 5641 7633
rect 5696 7599 5733 7633
rect 5767 7599 5825 7633
rect 5859 7599 5917 7633
rect 5951 7599 6009 7633
rect 6043 7599 6101 7633
rect 6135 7599 6193 7633
rect 6227 7599 6285 7633
rect 6319 7599 6377 7633
rect 6411 7599 6469 7633
rect 6503 7599 6561 7633
rect 6595 7599 6653 7633
rect 6687 7599 6745 7633
rect 6779 7599 6837 7633
rect 6871 7599 6929 7633
rect 6963 7599 7021 7633
rect 7055 7599 7113 7633
rect 7147 7599 7205 7633
rect 7239 7599 7297 7633
rect 7331 7599 7389 7633
rect 7423 7599 7481 7633
rect 7515 7599 7573 7633
rect 7607 7599 7665 7633
rect 7699 7599 7757 7633
rect 7791 7599 7849 7633
rect 7883 7599 7941 7633
rect 7975 7599 8033 7633
rect 8067 7599 8125 7633
rect 8159 7599 8217 7633
rect 8251 7599 8309 7633
rect 8343 7599 8401 7633
rect 8435 7599 8493 7633
rect 8527 7599 8585 7633
rect 8619 7599 8677 7633
rect 8711 7599 8769 7633
rect 8803 7599 8861 7633
rect 8895 7599 8953 7633
rect 8987 7599 9045 7633
rect 9079 7599 9137 7633
rect 9171 7599 9229 7633
rect 9263 7599 9321 7633
rect 9355 7599 9413 7633
rect 9447 7599 9505 7633
rect 9539 7599 9597 7633
rect 9631 7599 9689 7633
rect 9723 7599 9781 7633
rect 9815 7599 9827 7633
rect 5568 7590 5580 7599
rect 5632 7590 5644 7599
rect 5696 7590 9827 7599
rect 9879 7590 9891 7599
rect 9943 7590 9955 7642
rect 10007 7590 10019 7642
rect 10071 7633 10083 7642
rect 10135 7633 14266 7642
rect 14318 7633 14330 7642
rect 14382 7633 14394 7642
rect 10135 7599 10149 7633
rect 10183 7599 10241 7633
rect 10275 7599 10333 7633
rect 10367 7599 10425 7633
rect 10459 7599 10517 7633
rect 10551 7599 10609 7633
rect 10643 7599 10701 7633
rect 10735 7599 10793 7633
rect 10827 7599 10885 7633
rect 10919 7599 10977 7633
rect 11011 7599 11069 7633
rect 11103 7599 11161 7633
rect 11195 7599 11253 7633
rect 11287 7599 11345 7633
rect 11379 7599 11437 7633
rect 11471 7599 11529 7633
rect 11563 7599 11621 7633
rect 11655 7599 11713 7633
rect 11747 7599 11805 7633
rect 11839 7599 11897 7633
rect 11931 7599 11989 7633
rect 12023 7599 12081 7633
rect 12115 7599 12173 7633
rect 12207 7599 12265 7633
rect 12299 7599 12357 7633
rect 12391 7599 12449 7633
rect 12483 7599 12541 7633
rect 12575 7599 12633 7633
rect 12667 7599 12725 7633
rect 12759 7599 12817 7633
rect 12851 7599 12909 7633
rect 12943 7599 13001 7633
rect 13035 7599 13093 7633
rect 13127 7599 13185 7633
rect 13219 7599 13277 7633
rect 13311 7599 13369 7633
rect 13403 7599 13461 7633
rect 13495 7599 13553 7633
rect 13587 7599 13645 7633
rect 13679 7599 13737 7633
rect 13771 7599 13829 7633
rect 13863 7599 13921 7633
rect 13955 7599 14013 7633
rect 14047 7599 14105 7633
rect 14139 7599 14197 7633
rect 14231 7599 14266 7633
rect 14323 7599 14330 7633
rect 10071 7590 10083 7599
rect 10135 7590 14266 7599
rect 14318 7590 14330 7599
rect 14382 7590 14394 7599
rect 14446 7590 14458 7642
rect 14510 7590 14522 7642
rect 14574 7633 18705 7642
rect 14599 7599 14657 7633
rect 14691 7599 14749 7633
rect 14783 7599 14841 7633
rect 14875 7599 14933 7633
rect 14967 7599 15025 7633
rect 15059 7599 15117 7633
rect 15151 7599 15209 7633
rect 15243 7599 15301 7633
rect 15335 7599 15393 7633
rect 15427 7599 15485 7633
rect 15519 7599 15577 7633
rect 15611 7599 15669 7633
rect 15703 7599 15761 7633
rect 15795 7599 15853 7633
rect 15887 7599 15945 7633
rect 15979 7599 16037 7633
rect 16071 7599 16129 7633
rect 16163 7599 16221 7633
rect 16255 7599 16313 7633
rect 16347 7599 16405 7633
rect 16439 7599 16497 7633
rect 16531 7599 16589 7633
rect 16623 7599 16681 7633
rect 16715 7599 16773 7633
rect 16807 7599 16865 7633
rect 16899 7599 16957 7633
rect 16991 7599 17049 7633
rect 17083 7599 17141 7633
rect 17175 7599 17233 7633
rect 17267 7599 17325 7633
rect 17359 7599 17417 7633
rect 17451 7599 17509 7633
rect 17543 7599 17601 7633
rect 17635 7599 17693 7633
rect 17727 7599 17785 7633
rect 17819 7599 17877 7633
rect 17911 7599 17969 7633
rect 18003 7599 18061 7633
rect 18095 7599 18153 7633
rect 18187 7599 18245 7633
rect 18279 7599 18337 7633
rect 18371 7599 18429 7633
rect 18463 7599 18521 7633
rect 18555 7599 18613 7633
rect 18647 7599 18705 7633
rect 14574 7590 18705 7599
rect 18757 7590 18769 7642
rect 18821 7633 18833 7642
rect 18831 7599 18833 7633
rect 18821 7590 18833 7599
rect 18885 7590 18897 7642
rect 18949 7590 18961 7642
rect 19013 7590 19019 7642
rect 1104 7568 19019 7590
rect 1118 7488 1124 7540
rect 1176 7528 1182 7540
rect 1673 7531 1731 7537
rect 1673 7528 1685 7531
rect 1176 7500 1685 7528
rect 1176 7488 1182 7500
rect 1673 7497 1685 7500
rect 1719 7497 1731 7531
rect 1673 7491 1731 7497
rect 3326 7488 3332 7540
rect 3384 7528 3390 7540
rect 4065 7531 4123 7537
rect 4065 7528 4077 7531
rect 3384 7500 4077 7528
rect 3384 7488 3390 7500
rect 4065 7497 4077 7500
rect 4111 7497 4123 7531
rect 5718 7528 5724 7540
rect 5679 7500 5724 7528
rect 4065 7491 4123 7497
rect 5718 7488 5724 7500
rect 5776 7488 5782 7540
rect 7926 7528 7932 7540
rect 7887 7500 7932 7528
rect 7926 7488 7932 7500
rect 7984 7488 7990 7540
rect 12434 7528 12440 7540
rect 12395 7500 12440 7528
rect 12434 7488 12440 7500
rect 12492 7488 12498 7540
rect 14642 7528 14648 7540
rect 14603 7500 14648 7528
rect 14642 7488 14648 7500
rect 14700 7488 14706 7540
rect 16574 7488 16580 7540
rect 16632 7528 16638 7540
rect 17037 7531 17095 7537
rect 17037 7528 17049 7531
rect 16632 7500 17049 7528
rect 16632 7488 16638 7500
rect 17037 7497 17049 7500
rect 17083 7497 17095 7531
rect 17037 7491 17095 7497
rect 18233 7531 18291 7537
rect 18233 7497 18245 7531
rect 18279 7528 18291 7531
rect 18414 7528 18420 7540
rect 18279 7500 18420 7528
rect 18279 7497 18291 7500
rect 18233 7491 18291 7497
rect 18414 7488 18420 7500
rect 18472 7488 18478 7540
rect 7282 7420 7288 7472
rect 7340 7460 7346 7472
rect 9585 7463 9643 7469
rect 7340 7432 8248 7460
rect 7340 7420 7346 7432
rect 1857 7395 1915 7401
rect 1857 7361 1869 7395
rect 1903 7361 1915 7395
rect 1857 7355 1915 7361
rect 4249 7395 4307 7401
rect 4249 7361 4261 7395
rect 4295 7361 4307 7395
rect 4249 7355 4307 7361
rect 5905 7395 5963 7401
rect 5905 7361 5917 7395
rect 5951 7392 5963 7395
rect 7006 7392 7012 7404
rect 5951 7364 7012 7392
rect 5951 7361 5963 7364
rect 5905 7355 5963 7361
rect 1872 7324 1900 7355
rect 4264 7324 4292 7355
rect 7006 7352 7012 7364
rect 7064 7352 7070 7404
rect 7466 7352 7472 7404
rect 7524 7392 7530 7404
rect 8113 7395 8171 7401
rect 8113 7392 8125 7395
rect 7524 7364 8125 7392
rect 7524 7352 7530 7364
rect 8113 7361 8125 7364
rect 8159 7361 8171 7395
rect 8220 7392 8248 7432
rect 9585 7429 9597 7463
rect 9631 7460 9643 7463
rect 10137 7463 10195 7469
rect 10137 7460 10149 7463
rect 9631 7432 10149 7460
rect 9631 7429 9643 7432
rect 9585 7423 9643 7429
rect 10137 7429 10149 7432
rect 10183 7460 10195 7463
rect 10226 7460 10232 7472
rect 10183 7432 10232 7460
rect 10183 7429 10195 7432
rect 10137 7423 10195 7429
rect 10226 7420 10232 7432
rect 10284 7420 10290 7472
rect 12253 7395 12311 7401
rect 12253 7392 12265 7395
rect 8220 7364 12265 7392
rect 8113 7355 8171 7361
rect 12253 7361 12265 7364
rect 12299 7361 12311 7395
rect 12253 7355 12311 7361
rect 13814 7352 13820 7404
rect 13872 7392 13878 7404
rect 14461 7395 14519 7401
rect 14461 7392 14473 7395
rect 13872 7364 14473 7392
rect 13872 7352 13878 7364
rect 14461 7361 14473 7364
rect 14507 7361 14519 7395
rect 16850 7392 16856 7404
rect 16811 7364 16856 7392
rect 14461 7355 14519 7361
rect 16850 7352 16856 7364
rect 16908 7352 16914 7404
rect 18049 7395 18107 7401
rect 18049 7361 18061 7395
rect 18095 7361 18107 7395
rect 18049 7355 18107 7361
rect 7926 7324 7932 7336
rect 1872 7296 2774 7324
rect 4264 7296 7932 7324
rect 2746 7188 2774 7296
rect 7926 7284 7932 7296
rect 7984 7284 7990 7336
rect 13354 7284 13360 7336
rect 13412 7324 13418 7336
rect 18064 7324 18092 7355
rect 13412 7296 18092 7324
rect 13412 7284 13418 7296
rect 10318 7256 10324 7268
rect 10279 7228 10324 7256
rect 10318 7216 10324 7228
rect 10376 7216 10382 7268
rect 11054 7188 11060 7200
rect 2746 7160 11060 7188
rect 11054 7148 11060 7160
rect 11112 7148 11118 7200
rect 1104 7098 18860 7120
rect 1104 7089 3169 7098
rect 1104 7055 1133 7089
rect 1167 7055 1225 7089
rect 1259 7055 1317 7089
rect 1351 7055 1409 7089
rect 1443 7055 1501 7089
rect 1535 7055 1593 7089
rect 1627 7055 1685 7089
rect 1719 7055 1777 7089
rect 1811 7055 1869 7089
rect 1903 7055 1961 7089
rect 1995 7055 2053 7089
rect 2087 7055 2145 7089
rect 2179 7055 2237 7089
rect 2271 7055 2329 7089
rect 2363 7055 2421 7089
rect 2455 7055 2513 7089
rect 2547 7055 2605 7089
rect 2639 7055 2697 7089
rect 2731 7055 2789 7089
rect 2823 7055 2881 7089
rect 2915 7055 2973 7089
rect 3007 7055 3065 7089
rect 3099 7055 3157 7089
rect 1104 7046 3169 7055
rect 3221 7046 3233 7098
rect 3285 7046 3297 7098
rect 3349 7089 3361 7098
rect 3349 7046 3361 7055
rect 3413 7046 3425 7098
rect 3477 7089 7608 7098
rect 3477 7055 3525 7089
rect 3559 7055 3617 7089
rect 3651 7055 3709 7089
rect 3743 7055 3801 7089
rect 3835 7055 3893 7089
rect 3927 7055 3985 7089
rect 4019 7055 4077 7089
rect 4111 7055 4169 7089
rect 4203 7055 4261 7089
rect 4295 7055 4353 7089
rect 4387 7055 4445 7089
rect 4479 7055 4537 7089
rect 4571 7055 4629 7089
rect 4663 7055 4721 7089
rect 4755 7055 4813 7089
rect 4847 7055 4905 7089
rect 4939 7055 4997 7089
rect 5031 7055 5089 7089
rect 5123 7055 5181 7089
rect 5215 7055 5273 7089
rect 5307 7055 5365 7089
rect 5399 7055 5457 7089
rect 5491 7055 5549 7089
rect 5583 7055 5641 7089
rect 5675 7055 5733 7089
rect 5767 7055 5825 7089
rect 5859 7055 5917 7089
rect 5951 7055 6009 7089
rect 6043 7055 6101 7089
rect 6135 7055 6193 7089
rect 6227 7055 6285 7089
rect 6319 7055 6377 7089
rect 6411 7055 6469 7089
rect 6503 7055 6561 7089
rect 6595 7055 6653 7089
rect 6687 7055 6745 7089
rect 6779 7055 6837 7089
rect 6871 7055 6929 7089
rect 6963 7055 7021 7089
rect 7055 7055 7113 7089
rect 7147 7055 7205 7089
rect 7239 7055 7297 7089
rect 7331 7055 7389 7089
rect 7423 7055 7481 7089
rect 7515 7055 7573 7089
rect 7607 7055 7608 7089
rect 3477 7046 7608 7055
rect 7660 7089 7672 7098
rect 7660 7055 7665 7089
rect 7660 7046 7672 7055
rect 7724 7046 7736 7098
rect 7788 7089 7800 7098
rect 7852 7089 7864 7098
rect 7916 7089 12047 7098
rect 12099 7089 12111 7098
rect 12163 7089 12175 7098
rect 7791 7055 7800 7089
rect 7916 7055 7941 7089
rect 7975 7055 8033 7089
rect 8067 7055 8125 7089
rect 8159 7055 8217 7089
rect 8251 7055 8309 7089
rect 8343 7055 8401 7089
rect 8435 7055 8493 7089
rect 8527 7055 8585 7089
rect 8619 7055 8677 7089
rect 8711 7055 8769 7089
rect 8803 7055 8861 7089
rect 8895 7055 8953 7089
rect 8987 7055 9045 7089
rect 9079 7055 9137 7089
rect 9171 7055 9229 7089
rect 9263 7055 9321 7089
rect 9355 7055 9413 7089
rect 9447 7055 9505 7089
rect 9539 7055 9597 7089
rect 9631 7055 9689 7089
rect 9723 7055 9781 7089
rect 9815 7055 9873 7089
rect 9907 7055 9965 7089
rect 9999 7055 10057 7089
rect 10091 7055 10149 7089
rect 10183 7055 10241 7089
rect 10275 7055 10333 7089
rect 10367 7055 10425 7089
rect 10459 7055 10517 7089
rect 10551 7055 10609 7089
rect 10643 7055 10701 7089
rect 10735 7055 10793 7089
rect 10827 7055 10885 7089
rect 10919 7055 10977 7089
rect 11011 7055 11069 7089
rect 11103 7055 11161 7089
rect 11195 7055 11253 7089
rect 11287 7055 11345 7089
rect 11379 7055 11437 7089
rect 11471 7055 11529 7089
rect 11563 7055 11621 7089
rect 11655 7055 11713 7089
rect 11747 7055 11805 7089
rect 11839 7055 11897 7089
rect 11931 7055 11989 7089
rect 12023 7055 12047 7089
rect 12163 7055 12173 7089
rect 7788 7046 7800 7055
rect 7852 7046 7864 7055
rect 7916 7046 12047 7055
rect 12099 7046 12111 7055
rect 12163 7046 12175 7055
rect 12227 7046 12239 7098
rect 12291 7089 12303 7098
rect 12299 7055 12303 7089
rect 12291 7046 12303 7055
rect 12355 7089 16486 7098
rect 12355 7055 12357 7089
rect 12391 7055 12449 7089
rect 12483 7055 12541 7089
rect 12575 7055 12633 7089
rect 12667 7055 12725 7089
rect 12759 7055 12817 7089
rect 12851 7055 12909 7089
rect 12943 7055 13001 7089
rect 13035 7055 13093 7089
rect 13127 7055 13185 7089
rect 13219 7055 13277 7089
rect 13311 7055 13369 7089
rect 13403 7055 13461 7089
rect 13495 7055 13553 7089
rect 13587 7055 13645 7089
rect 13679 7055 13737 7089
rect 13771 7055 13829 7089
rect 13863 7055 13921 7089
rect 13955 7055 14013 7089
rect 14047 7055 14105 7089
rect 14139 7055 14197 7089
rect 14231 7055 14289 7089
rect 14323 7055 14381 7089
rect 14415 7055 14473 7089
rect 14507 7055 14565 7089
rect 14599 7055 14657 7089
rect 14691 7055 14749 7089
rect 14783 7055 14841 7089
rect 14875 7055 14933 7089
rect 14967 7055 15025 7089
rect 15059 7055 15117 7089
rect 15151 7055 15209 7089
rect 15243 7055 15301 7089
rect 15335 7055 15393 7089
rect 15427 7055 15485 7089
rect 15519 7055 15577 7089
rect 15611 7055 15669 7089
rect 15703 7055 15761 7089
rect 15795 7055 15853 7089
rect 15887 7055 15945 7089
rect 15979 7055 16037 7089
rect 16071 7055 16129 7089
rect 16163 7055 16221 7089
rect 16255 7055 16313 7089
rect 16347 7055 16405 7089
rect 16439 7055 16486 7089
rect 12355 7046 16486 7055
rect 16538 7046 16550 7098
rect 16602 7089 16614 7098
rect 16602 7046 16614 7055
rect 16666 7046 16678 7098
rect 16730 7046 16742 7098
rect 16794 7089 18860 7098
rect 16807 7055 16865 7089
rect 16899 7055 16957 7089
rect 16991 7055 17049 7089
rect 17083 7055 17141 7089
rect 17175 7055 17233 7089
rect 17267 7055 17325 7089
rect 17359 7055 17417 7089
rect 17451 7055 17509 7089
rect 17543 7055 17601 7089
rect 17635 7055 17693 7089
rect 17727 7055 17785 7089
rect 17819 7055 17877 7089
rect 17911 7055 17969 7089
rect 18003 7055 18061 7089
rect 18095 7055 18153 7089
rect 18187 7055 18245 7089
rect 18279 7055 18337 7089
rect 18371 7055 18429 7089
rect 18463 7055 18521 7089
rect 18555 7055 18613 7089
rect 18647 7055 18705 7089
rect 18739 7055 18797 7089
rect 18831 7055 18860 7089
rect 16794 7046 18860 7055
rect 1104 7024 18860 7046
rect 1104 6554 19019 6576
rect 1104 6545 5388 6554
rect 1104 6511 1133 6545
rect 1167 6511 1225 6545
rect 1259 6511 1317 6545
rect 1351 6511 1409 6545
rect 1443 6511 1501 6545
rect 1535 6511 1593 6545
rect 1627 6511 1685 6545
rect 1719 6511 1777 6545
rect 1811 6511 1869 6545
rect 1903 6511 1961 6545
rect 1995 6511 2053 6545
rect 2087 6511 2145 6545
rect 2179 6511 2237 6545
rect 2271 6511 2329 6545
rect 2363 6511 2421 6545
rect 2455 6511 2513 6545
rect 2547 6511 2605 6545
rect 2639 6511 2697 6545
rect 2731 6511 2789 6545
rect 2823 6511 2881 6545
rect 2915 6511 2973 6545
rect 3007 6511 3065 6545
rect 3099 6511 3157 6545
rect 3191 6511 3249 6545
rect 3283 6511 3341 6545
rect 3375 6511 3433 6545
rect 3467 6511 3525 6545
rect 3559 6511 3617 6545
rect 3651 6511 3709 6545
rect 3743 6511 3801 6545
rect 3835 6511 3893 6545
rect 3927 6511 3985 6545
rect 4019 6511 4077 6545
rect 4111 6511 4169 6545
rect 4203 6511 4261 6545
rect 4295 6511 4353 6545
rect 4387 6511 4445 6545
rect 4479 6511 4537 6545
rect 4571 6511 4629 6545
rect 4663 6511 4721 6545
rect 4755 6511 4813 6545
rect 4847 6511 4905 6545
rect 4939 6511 4997 6545
rect 5031 6511 5089 6545
rect 5123 6511 5181 6545
rect 5215 6511 5273 6545
rect 5307 6511 5365 6545
rect 1104 6502 5388 6511
rect 5440 6502 5452 6554
rect 5504 6502 5516 6554
rect 5568 6545 5580 6554
rect 5632 6545 5644 6554
rect 5696 6545 9827 6554
rect 9879 6545 9891 6554
rect 5632 6511 5641 6545
rect 5696 6511 5733 6545
rect 5767 6511 5825 6545
rect 5859 6511 5917 6545
rect 5951 6511 6009 6545
rect 6043 6511 6101 6545
rect 6135 6511 6193 6545
rect 6227 6511 6285 6545
rect 6319 6511 6377 6545
rect 6411 6511 6469 6545
rect 6503 6511 6561 6545
rect 6595 6511 6653 6545
rect 6687 6511 6745 6545
rect 6779 6511 6837 6545
rect 6871 6511 6929 6545
rect 6963 6511 7021 6545
rect 7055 6511 7113 6545
rect 7147 6511 7205 6545
rect 7239 6511 7297 6545
rect 7331 6511 7389 6545
rect 7423 6511 7481 6545
rect 7515 6511 7573 6545
rect 7607 6511 7665 6545
rect 7699 6511 7757 6545
rect 7791 6511 7849 6545
rect 7883 6511 7941 6545
rect 7975 6511 8033 6545
rect 8067 6511 8125 6545
rect 8159 6511 8217 6545
rect 8251 6511 8309 6545
rect 8343 6511 8401 6545
rect 8435 6511 8493 6545
rect 8527 6511 8585 6545
rect 8619 6511 8677 6545
rect 8711 6511 8769 6545
rect 8803 6511 8861 6545
rect 8895 6511 8953 6545
rect 8987 6511 9045 6545
rect 9079 6511 9137 6545
rect 9171 6511 9229 6545
rect 9263 6511 9321 6545
rect 9355 6511 9413 6545
rect 9447 6511 9505 6545
rect 9539 6511 9597 6545
rect 9631 6511 9689 6545
rect 9723 6511 9781 6545
rect 9815 6511 9827 6545
rect 5568 6502 5580 6511
rect 5632 6502 5644 6511
rect 5696 6502 9827 6511
rect 9879 6502 9891 6511
rect 9943 6502 9955 6554
rect 10007 6502 10019 6554
rect 10071 6545 10083 6554
rect 10135 6545 14266 6554
rect 14318 6545 14330 6554
rect 14382 6545 14394 6554
rect 10135 6511 10149 6545
rect 10183 6511 10241 6545
rect 10275 6511 10333 6545
rect 10367 6511 10425 6545
rect 10459 6511 10517 6545
rect 10551 6511 10609 6545
rect 10643 6511 10701 6545
rect 10735 6511 10793 6545
rect 10827 6511 10885 6545
rect 10919 6511 10977 6545
rect 11011 6511 11069 6545
rect 11103 6511 11161 6545
rect 11195 6511 11253 6545
rect 11287 6511 11345 6545
rect 11379 6511 11437 6545
rect 11471 6511 11529 6545
rect 11563 6511 11621 6545
rect 11655 6511 11713 6545
rect 11747 6511 11805 6545
rect 11839 6511 11897 6545
rect 11931 6511 11989 6545
rect 12023 6511 12081 6545
rect 12115 6511 12173 6545
rect 12207 6511 12265 6545
rect 12299 6511 12357 6545
rect 12391 6511 12449 6545
rect 12483 6511 12541 6545
rect 12575 6511 12633 6545
rect 12667 6511 12725 6545
rect 12759 6511 12817 6545
rect 12851 6511 12909 6545
rect 12943 6511 13001 6545
rect 13035 6511 13093 6545
rect 13127 6511 13185 6545
rect 13219 6511 13277 6545
rect 13311 6511 13369 6545
rect 13403 6511 13461 6545
rect 13495 6511 13553 6545
rect 13587 6511 13645 6545
rect 13679 6511 13737 6545
rect 13771 6511 13829 6545
rect 13863 6511 13921 6545
rect 13955 6511 14013 6545
rect 14047 6511 14105 6545
rect 14139 6511 14197 6545
rect 14231 6511 14266 6545
rect 14323 6511 14330 6545
rect 10071 6502 10083 6511
rect 10135 6502 14266 6511
rect 14318 6502 14330 6511
rect 14382 6502 14394 6511
rect 14446 6502 14458 6554
rect 14510 6502 14522 6554
rect 14574 6545 18705 6554
rect 14599 6511 14657 6545
rect 14691 6511 14749 6545
rect 14783 6511 14841 6545
rect 14875 6511 14933 6545
rect 14967 6511 15025 6545
rect 15059 6511 15117 6545
rect 15151 6511 15209 6545
rect 15243 6511 15301 6545
rect 15335 6511 15393 6545
rect 15427 6511 15485 6545
rect 15519 6511 15577 6545
rect 15611 6511 15669 6545
rect 15703 6511 15761 6545
rect 15795 6511 15853 6545
rect 15887 6511 15945 6545
rect 15979 6511 16037 6545
rect 16071 6511 16129 6545
rect 16163 6511 16221 6545
rect 16255 6511 16313 6545
rect 16347 6511 16405 6545
rect 16439 6511 16497 6545
rect 16531 6511 16589 6545
rect 16623 6511 16681 6545
rect 16715 6511 16773 6545
rect 16807 6511 16865 6545
rect 16899 6511 16957 6545
rect 16991 6511 17049 6545
rect 17083 6511 17141 6545
rect 17175 6511 17233 6545
rect 17267 6511 17325 6545
rect 17359 6511 17417 6545
rect 17451 6511 17509 6545
rect 17543 6511 17601 6545
rect 17635 6511 17693 6545
rect 17727 6511 17785 6545
rect 17819 6511 17877 6545
rect 17911 6511 17969 6545
rect 18003 6511 18061 6545
rect 18095 6511 18153 6545
rect 18187 6511 18245 6545
rect 18279 6511 18337 6545
rect 18371 6511 18429 6545
rect 18463 6511 18521 6545
rect 18555 6511 18613 6545
rect 18647 6511 18705 6545
rect 14574 6502 18705 6511
rect 18757 6502 18769 6554
rect 18821 6545 18833 6554
rect 18831 6511 18833 6545
rect 18821 6502 18833 6511
rect 18885 6502 18897 6554
rect 18949 6502 18961 6554
rect 19013 6502 19019 6554
rect 1104 6480 19019 6502
rect 8018 6304 8024 6316
rect 7979 6276 8024 6304
rect 8018 6264 8024 6276
rect 8076 6264 8082 6316
rect 8202 6304 8208 6316
rect 8163 6276 8208 6304
rect 8202 6264 8208 6276
rect 8260 6264 8266 6316
rect 8389 6103 8447 6109
rect 8389 6069 8401 6103
rect 8435 6100 8447 6103
rect 10962 6100 10968 6112
rect 8435 6072 10968 6100
rect 8435 6069 8447 6072
rect 8389 6063 8447 6069
rect 10962 6060 10968 6072
rect 11020 6060 11026 6112
rect 1104 6010 18860 6032
rect 1104 6001 3169 6010
rect 1104 5967 1133 6001
rect 1167 5967 1225 6001
rect 1259 5967 1317 6001
rect 1351 5967 1409 6001
rect 1443 5967 1501 6001
rect 1535 5967 1593 6001
rect 1627 5967 1685 6001
rect 1719 5967 1777 6001
rect 1811 5967 1869 6001
rect 1903 5967 1961 6001
rect 1995 5967 2053 6001
rect 2087 5967 2145 6001
rect 2179 5967 2237 6001
rect 2271 5967 2329 6001
rect 2363 5967 2421 6001
rect 2455 5967 2513 6001
rect 2547 5967 2605 6001
rect 2639 5967 2697 6001
rect 2731 5967 2789 6001
rect 2823 5967 2881 6001
rect 2915 5967 2973 6001
rect 3007 5967 3065 6001
rect 3099 5967 3157 6001
rect 1104 5958 3169 5967
rect 3221 5958 3233 6010
rect 3285 5958 3297 6010
rect 3349 6001 3361 6010
rect 3349 5958 3361 5967
rect 3413 5958 3425 6010
rect 3477 6001 7608 6010
rect 3477 5967 3525 6001
rect 3559 5967 3617 6001
rect 3651 5967 3709 6001
rect 3743 5967 3801 6001
rect 3835 5967 3893 6001
rect 3927 5967 3985 6001
rect 4019 5967 4077 6001
rect 4111 5967 4169 6001
rect 4203 5967 4261 6001
rect 4295 5967 4353 6001
rect 4387 5967 4445 6001
rect 4479 5967 4537 6001
rect 4571 5967 4629 6001
rect 4663 5967 4721 6001
rect 4755 5967 4813 6001
rect 4847 5967 4905 6001
rect 4939 5967 4997 6001
rect 5031 5967 5089 6001
rect 5123 5967 5181 6001
rect 5215 5967 5273 6001
rect 5307 5967 5365 6001
rect 5399 5967 5457 6001
rect 5491 5967 5549 6001
rect 5583 5967 5641 6001
rect 5675 5967 5733 6001
rect 5767 5967 5825 6001
rect 5859 5967 5917 6001
rect 5951 5967 6009 6001
rect 6043 5967 6101 6001
rect 6135 5967 6193 6001
rect 6227 5967 6285 6001
rect 6319 5967 6377 6001
rect 6411 5967 6469 6001
rect 6503 5967 6561 6001
rect 6595 5967 6653 6001
rect 6687 5967 6745 6001
rect 6779 5967 6837 6001
rect 6871 5967 6929 6001
rect 6963 5967 7021 6001
rect 7055 5967 7113 6001
rect 7147 5967 7205 6001
rect 7239 5967 7297 6001
rect 7331 5967 7389 6001
rect 7423 5967 7481 6001
rect 7515 5967 7573 6001
rect 7607 5967 7608 6001
rect 3477 5958 7608 5967
rect 7660 6001 7672 6010
rect 7660 5967 7665 6001
rect 7660 5958 7672 5967
rect 7724 5958 7736 6010
rect 7788 6001 7800 6010
rect 7852 6001 7864 6010
rect 7916 6001 12047 6010
rect 12099 6001 12111 6010
rect 12163 6001 12175 6010
rect 7791 5967 7800 6001
rect 7916 5967 7941 6001
rect 7975 5967 8033 6001
rect 8067 5967 8125 6001
rect 8159 5967 8217 6001
rect 8251 5967 8309 6001
rect 8343 5967 8401 6001
rect 8435 5967 8493 6001
rect 8527 5967 8585 6001
rect 8619 5967 8677 6001
rect 8711 5967 8769 6001
rect 8803 5967 8861 6001
rect 8895 5967 8953 6001
rect 8987 5967 9045 6001
rect 9079 5967 9137 6001
rect 9171 5967 9229 6001
rect 9263 5967 9321 6001
rect 9355 5967 9413 6001
rect 9447 5967 9505 6001
rect 9539 5967 9597 6001
rect 9631 5967 9689 6001
rect 9723 5967 9781 6001
rect 9815 5967 9873 6001
rect 9907 5967 9965 6001
rect 9999 5967 10057 6001
rect 10091 5967 10149 6001
rect 10183 5967 10241 6001
rect 10275 5967 10333 6001
rect 10367 5967 10425 6001
rect 10459 5967 10517 6001
rect 10551 5967 10609 6001
rect 10643 5967 10701 6001
rect 10735 5967 10793 6001
rect 10827 5967 10885 6001
rect 10919 5967 10977 6001
rect 11011 5967 11069 6001
rect 11103 5967 11161 6001
rect 11195 5967 11253 6001
rect 11287 5967 11345 6001
rect 11379 5967 11437 6001
rect 11471 5967 11529 6001
rect 11563 5967 11621 6001
rect 11655 5967 11713 6001
rect 11747 5967 11805 6001
rect 11839 5967 11897 6001
rect 11931 5967 11989 6001
rect 12023 5967 12047 6001
rect 12163 5967 12173 6001
rect 7788 5958 7800 5967
rect 7852 5958 7864 5967
rect 7916 5958 12047 5967
rect 12099 5958 12111 5967
rect 12163 5958 12175 5967
rect 12227 5958 12239 6010
rect 12291 6001 12303 6010
rect 12299 5967 12303 6001
rect 12291 5958 12303 5967
rect 12355 6001 16486 6010
rect 12355 5967 12357 6001
rect 12391 5967 12449 6001
rect 12483 5967 12541 6001
rect 12575 5967 12633 6001
rect 12667 5967 12725 6001
rect 12759 5967 12817 6001
rect 12851 5967 12909 6001
rect 12943 5967 13001 6001
rect 13035 5967 13093 6001
rect 13127 5967 13185 6001
rect 13219 5967 13277 6001
rect 13311 5967 13369 6001
rect 13403 5967 13461 6001
rect 13495 5967 13553 6001
rect 13587 5967 13645 6001
rect 13679 5967 13737 6001
rect 13771 5967 13829 6001
rect 13863 5967 13921 6001
rect 13955 5967 14013 6001
rect 14047 5967 14105 6001
rect 14139 5967 14197 6001
rect 14231 5967 14289 6001
rect 14323 5967 14381 6001
rect 14415 5967 14473 6001
rect 14507 5967 14565 6001
rect 14599 5967 14657 6001
rect 14691 5967 14749 6001
rect 14783 5967 14841 6001
rect 14875 5967 14933 6001
rect 14967 5967 15025 6001
rect 15059 5967 15117 6001
rect 15151 5967 15209 6001
rect 15243 5967 15301 6001
rect 15335 5967 15393 6001
rect 15427 5967 15485 6001
rect 15519 5967 15577 6001
rect 15611 5967 15669 6001
rect 15703 5967 15761 6001
rect 15795 5967 15853 6001
rect 15887 5967 15945 6001
rect 15979 5967 16037 6001
rect 16071 5967 16129 6001
rect 16163 5967 16221 6001
rect 16255 5967 16313 6001
rect 16347 5967 16405 6001
rect 16439 5967 16486 6001
rect 12355 5958 16486 5967
rect 16538 5958 16550 6010
rect 16602 6001 16614 6010
rect 16602 5958 16614 5967
rect 16666 5958 16678 6010
rect 16730 5958 16742 6010
rect 16794 6001 18860 6010
rect 16807 5967 16865 6001
rect 16899 5967 16957 6001
rect 16991 5967 17049 6001
rect 17083 5967 17141 6001
rect 17175 5967 17233 6001
rect 17267 5967 17325 6001
rect 17359 5967 17417 6001
rect 17451 5967 17509 6001
rect 17543 5967 17601 6001
rect 17635 5967 17693 6001
rect 17727 5967 17785 6001
rect 17819 5967 17877 6001
rect 17911 5967 17969 6001
rect 18003 5967 18061 6001
rect 18095 5967 18153 6001
rect 18187 5967 18245 6001
rect 18279 5967 18337 6001
rect 18371 5967 18429 6001
rect 18463 5967 18521 6001
rect 18555 5967 18613 6001
rect 18647 5967 18705 6001
rect 18739 5967 18797 6001
rect 18831 5967 18860 6001
rect 16794 5958 18860 5967
rect 1104 5936 18860 5958
rect 8018 5856 8024 5908
rect 8076 5896 8082 5908
rect 8297 5899 8355 5905
rect 8297 5896 8309 5899
rect 8076 5868 8309 5896
rect 8076 5856 8082 5868
rect 8297 5865 8309 5868
rect 8343 5865 8355 5899
rect 8297 5859 8355 5865
rect 7745 5763 7803 5769
rect 7745 5729 7757 5763
rect 7791 5760 7803 5763
rect 8110 5760 8116 5772
rect 7791 5732 8116 5760
rect 7791 5729 7803 5732
rect 7745 5723 7803 5729
rect 8110 5720 8116 5732
rect 8168 5720 8174 5772
rect 6914 5692 6920 5704
rect 6875 5664 6920 5692
rect 6914 5652 6920 5664
rect 6972 5652 6978 5704
rect 7466 5584 7472 5636
rect 7524 5624 7530 5636
rect 7929 5627 7987 5633
rect 7929 5624 7941 5627
rect 7524 5596 7941 5624
rect 7524 5584 7530 5596
rect 7929 5593 7941 5596
rect 7975 5593 7987 5627
rect 11514 5624 11520 5636
rect 11475 5596 11520 5624
rect 7929 5587 7987 5593
rect 11514 5584 11520 5596
rect 11572 5584 11578 5636
rect 11698 5624 11704 5636
rect 11659 5596 11704 5624
rect 11698 5584 11704 5596
rect 11756 5584 11762 5636
rect 12802 5624 12808 5636
rect 12763 5596 12808 5624
rect 12802 5584 12808 5596
rect 12860 5584 12866 5636
rect 12894 5584 12900 5636
rect 12952 5624 12958 5636
rect 12989 5627 13047 5633
rect 12989 5624 13001 5627
rect 12952 5596 13001 5624
rect 12952 5584 12958 5596
rect 12989 5593 13001 5596
rect 13035 5593 13047 5627
rect 12989 5587 13047 5593
rect 4614 5516 4620 5568
rect 4672 5556 4678 5568
rect 6733 5559 6791 5565
rect 6733 5556 6745 5559
rect 4672 5528 6745 5556
rect 4672 5516 4678 5528
rect 6733 5525 6745 5528
rect 6779 5525 6791 5559
rect 6733 5519 6791 5525
rect 7374 5516 7380 5568
rect 7432 5556 7438 5568
rect 7837 5559 7895 5565
rect 7837 5556 7849 5559
rect 7432 5528 7849 5556
rect 7432 5516 7438 5528
rect 7837 5525 7849 5528
rect 7883 5525 7895 5559
rect 7837 5519 7895 5525
rect 11885 5559 11943 5565
rect 11885 5525 11897 5559
rect 11931 5556 11943 5559
rect 13078 5556 13084 5568
rect 11931 5528 13084 5556
rect 11931 5525 11943 5528
rect 11885 5519 11943 5525
rect 13078 5516 13084 5528
rect 13136 5516 13142 5568
rect 13173 5559 13231 5565
rect 13173 5525 13185 5559
rect 13219 5556 13231 5559
rect 15102 5556 15108 5568
rect 13219 5528 15108 5556
rect 13219 5525 13231 5528
rect 13173 5519 13231 5525
rect 15102 5516 15108 5528
rect 15160 5516 15166 5568
rect 1104 5466 19019 5488
rect 1104 5457 5388 5466
rect 1104 5423 1133 5457
rect 1167 5423 1225 5457
rect 1259 5423 1317 5457
rect 1351 5423 1409 5457
rect 1443 5423 1501 5457
rect 1535 5423 1593 5457
rect 1627 5423 1685 5457
rect 1719 5423 1777 5457
rect 1811 5423 1869 5457
rect 1903 5423 1961 5457
rect 1995 5423 2053 5457
rect 2087 5423 2145 5457
rect 2179 5423 2237 5457
rect 2271 5423 2329 5457
rect 2363 5423 2421 5457
rect 2455 5423 2513 5457
rect 2547 5423 2605 5457
rect 2639 5423 2697 5457
rect 2731 5423 2789 5457
rect 2823 5423 2881 5457
rect 2915 5423 2973 5457
rect 3007 5423 3065 5457
rect 3099 5423 3157 5457
rect 3191 5423 3249 5457
rect 3283 5423 3341 5457
rect 3375 5423 3433 5457
rect 3467 5423 3525 5457
rect 3559 5423 3617 5457
rect 3651 5423 3709 5457
rect 3743 5423 3801 5457
rect 3835 5423 3893 5457
rect 3927 5423 3985 5457
rect 4019 5423 4077 5457
rect 4111 5423 4169 5457
rect 4203 5423 4261 5457
rect 4295 5423 4353 5457
rect 4387 5423 4445 5457
rect 4479 5423 4537 5457
rect 4571 5423 4629 5457
rect 4663 5423 4721 5457
rect 4755 5423 4813 5457
rect 4847 5423 4905 5457
rect 4939 5423 4997 5457
rect 5031 5423 5089 5457
rect 5123 5423 5181 5457
rect 5215 5423 5273 5457
rect 5307 5423 5365 5457
rect 1104 5414 5388 5423
rect 5440 5414 5452 5466
rect 5504 5414 5516 5466
rect 5568 5457 5580 5466
rect 5632 5457 5644 5466
rect 5696 5457 9827 5466
rect 9879 5457 9891 5466
rect 5632 5423 5641 5457
rect 5696 5423 5733 5457
rect 5767 5423 5825 5457
rect 5859 5423 5917 5457
rect 5951 5423 6009 5457
rect 6043 5423 6101 5457
rect 6135 5423 6193 5457
rect 6227 5423 6285 5457
rect 6319 5423 6377 5457
rect 6411 5423 6469 5457
rect 6503 5423 6561 5457
rect 6595 5423 6653 5457
rect 6687 5423 6745 5457
rect 6779 5423 6837 5457
rect 6871 5423 6929 5457
rect 6963 5423 7021 5457
rect 7055 5423 7113 5457
rect 7147 5423 7205 5457
rect 7239 5423 7297 5457
rect 7331 5423 7389 5457
rect 7423 5423 7481 5457
rect 7515 5423 7573 5457
rect 7607 5423 7665 5457
rect 7699 5423 7757 5457
rect 7791 5423 7849 5457
rect 7883 5423 7941 5457
rect 7975 5423 8033 5457
rect 8067 5423 8125 5457
rect 8159 5423 8217 5457
rect 8251 5423 8309 5457
rect 8343 5423 8401 5457
rect 8435 5423 8493 5457
rect 8527 5423 8585 5457
rect 8619 5423 8677 5457
rect 8711 5423 8769 5457
rect 8803 5423 8861 5457
rect 8895 5423 8953 5457
rect 8987 5423 9045 5457
rect 9079 5423 9137 5457
rect 9171 5423 9229 5457
rect 9263 5423 9321 5457
rect 9355 5423 9413 5457
rect 9447 5423 9505 5457
rect 9539 5423 9597 5457
rect 9631 5423 9689 5457
rect 9723 5423 9781 5457
rect 9815 5423 9827 5457
rect 5568 5414 5580 5423
rect 5632 5414 5644 5423
rect 5696 5414 9827 5423
rect 9879 5414 9891 5423
rect 9943 5414 9955 5466
rect 10007 5414 10019 5466
rect 10071 5457 10083 5466
rect 10135 5457 14266 5466
rect 14318 5457 14330 5466
rect 14382 5457 14394 5466
rect 10135 5423 10149 5457
rect 10183 5423 10241 5457
rect 10275 5423 10333 5457
rect 10367 5423 10425 5457
rect 10459 5423 10517 5457
rect 10551 5423 10609 5457
rect 10643 5423 10701 5457
rect 10735 5423 10793 5457
rect 10827 5423 10885 5457
rect 10919 5423 10977 5457
rect 11011 5423 11069 5457
rect 11103 5423 11161 5457
rect 11195 5423 11253 5457
rect 11287 5423 11345 5457
rect 11379 5423 11437 5457
rect 11471 5423 11529 5457
rect 11563 5423 11621 5457
rect 11655 5423 11713 5457
rect 11747 5423 11805 5457
rect 11839 5423 11897 5457
rect 11931 5423 11989 5457
rect 12023 5423 12081 5457
rect 12115 5423 12173 5457
rect 12207 5423 12265 5457
rect 12299 5423 12357 5457
rect 12391 5423 12449 5457
rect 12483 5423 12541 5457
rect 12575 5423 12633 5457
rect 12667 5423 12725 5457
rect 12759 5423 12817 5457
rect 12851 5423 12909 5457
rect 12943 5423 13001 5457
rect 13035 5423 13093 5457
rect 13127 5423 13185 5457
rect 13219 5423 13277 5457
rect 13311 5423 13369 5457
rect 13403 5423 13461 5457
rect 13495 5423 13553 5457
rect 13587 5423 13645 5457
rect 13679 5423 13737 5457
rect 13771 5423 13829 5457
rect 13863 5423 13921 5457
rect 13955 5423 14013 5457
rect 14047 5423 14105 5457
rect 14139 5423 14197 5457
rect 14231 5423 14266 5457
rect 14323 5423 14330 5457
rect 10071 5414 10083 5423
rect 10135 5414 14266 5423
rect 14318 5414 14330 5423
rect 14382 5414 14394 5423
rect 14446 5414 14458 5466
rect 14510 5414 14522 5466
rect 14574 5457 18705 5466
rect 14599 5423 14657 5457
rect 14691 5423 14749 5457
rect 14783 5423 14841 5457
rect 14875 5423 14933 5457
rect 14967 5423 15025 5457
rect 15059 5423 15117 5457
rect 15151 5423 15209 5457
rect 15243 5423 15301 5457
rect 15335 5423 15393 5457
rect 15427 5423 15485 5457
rect 15519 5423 15577 5457
rect 15611 5423 15669 5457
rect 15703 5423 15761 5457
rect 15795 5423 15853 5457
rect 15887 5423 15945 5457
rect 15979 5423 16037 5457
rect 16071 5423 16129 5457
rect 16163 5423 16221 5457
rect 16255 5423 16313 5457
rect 16347 5423 16405 5457
rect 16439 5423 16497 5457
rect 16531 5423 16589 5457
rect 16623 5423 16681 5457
rect 16715 5423 16773 5457
rect 16807 5423 16865 5457
rect 16899 5423 16957 5457
rect 16991 5423 17049 5457
rect 17083 5423 17141 5457
rect 17175 5423 17233 5457
rect 17267 5423 17325 5457
rect 17359 5423 17417 5457
rect 17451 5423 17509 5457
rect 17543 5423 17601 5457
rect 17635 5423 17693 5457
rect 17727 5423 17785 5457
rect 17819 5423 17877 5457
rect 17911 5423 17969 5457
rect 18003 5423 18061 5457
rect 18095 5423 18153 5457
rect 18187 5423 18245 5457
rect 18279 5423 18337 5457
rect 18371 5423 18429 5457
rect 18463 5423 18521 5457
rect 18555 5423 18613 5457
rect 18647 5423 18705 5457
rect 14574 5414 18705 5423
rect 18757 5414 18769 5466
rect 18821 5457 18833 5466
rect 18831 5423 18833 5457
rect 18821 5414 18833 5423
rect 18885 5414 18897 5466
rect 18949 5414 18961 5466
rect 19013 5414 19019 5466
rect 1104 5392 19019 5414
rect 4525 5355 4583 5361
rect 4525 5321 4537 5355
rect 4571 5321 4583 5355
rect 7006 5352 7012 5364
rect 6967 5324 7012 5352
rect 4525 5315 4583 5321
rect 3509 5287 3639 5293
rect 3509 5253 3521 5287
rect 3555 5253 3593 5287
rect 3627 5284 3639 5287
rect 4229 5287 4287 5293
rect 4229 5284 4241 5287
rect 3627 5256 4241 5284
rect 3627 5253 3639 5256
rect 3509 5247 3639 5253
rect 4169 5253 4241 5256
rect 4275 5284 4287 5287
rect 4430 5284 4436 5296
rect 4275 5256 4436 5284
rect 4275 5253 4287 5256
rect 4169 5247 4287 5253
rect 2870 5219 2928 5225
rect 2870 5185 2882 5219
rect 2916 5216 2928 5219
rect 3237 5219 3295 5225
rect 3237 5216 3249 5219
rect 2916 5188 3249 5216
rect 2916 5185 2928 5188
rect 2870 5179 2928 5185
rect 3237 5185 3249 5188
rect 3283 5216 3295 5219
rect 3953 5219 4011 5225
rect 3953 5216 3965 5219
rect 3283 5188 3965 5216
rect 3283 5185 3295 5188
rect 3237 5179 3295 5185
rect 3953 5185 3965 5188
rect 3999 5185 4011 5219
rect 3953 5179 4011 5185
rect 4169 5224 4227 5247
rect 4430 5244 4436 5256
rect 4488 5244 4494 5296
rect 4540 5284 4568 5315
rect 7006 5312 7012 5324
rect 7064 5312 7070 5364
rect 7101 5355 7159 5361
rect 7101 5321 7113 5355
rect 7147 5352 7159 5355
rect 7374 5352 7380 5364
rect 7147 5324 7380 5352
rect 7147 5321 7159 5324
rect 7101 5315 7159 5321
rect 7374 5312 7380 5324
rect 7432 5312 7438 5364
rect 10413 5355 10471 5361
rect 8496 5324 9720 5352
rect 8496 5284 8524 5324
rect 4540 5256 8524 5284
rect 8569 5287 8699 5293
rect 8569 5253 8581 5287
rect 8615 5253 8653 5287
rect 8687 5284 8699 5287
rect 9289 5287 9347 5293
rect 9289 5284 9301 5287
rect 8687 5256 9301 5284
rect 8687 5253 8699 5256
rect 8569 5247 8699 5253
rect 9229 5253 9301 5256
rect 9335 5253 9347 5287
rect 9229 5247 9347 5253
rect 9229 5228 9287 5247
rect 4169 5190 4181 5224
rect 4215 5190 4227 5224
rect 4169 5184 4227 5190
rect 6730 5176 6736 5228
rect 6788 5216 6794 5228
rect 7930 5219 7988 5225
rect 6788 5188 7880 5216
rect 6788 5176 6794 5188
rect 2777 5151 2835 5157
rect 2777 5117 2789 5151
rect 2823 5148 2835 5151
rect 3050 5148 3056 5160
rect 2823 5120 2912 5148
rect 3011 5120 3056 5148
rect 2823 5117 2835 5120
rect 2777 5111 2835 5117
rect 2884 5012 2912 5120
rect 3050 5108 3056 5120
rect 3108 5108 3114 5160
rect 7852 5157 7880 5188
rect 7930 5185 7942 5219
rect 7976 5216 7988 5219
rect 8297 5219 8355 5225
rect 8297 5216 8309 5219
rect 7976 5188 8309 5216
rect 7976 5185 7988 5188
rect 7930 5179 7988 5185
rect 8297 5185 8309 5188
rect 8343 5216 8355 5219
rect 9013 5219 9071 5225
rect 9013 5216 9025 5219
rect 8343 5188 9025 5216
rect 8343 5185 8355 5188
rect 8297 5179 8355 5185
rect 9013 5185 9025 5188
rect 9059 5185 9071 5219
rect 9013 5179 9071 5185
rect 9214 5176 9220 5228
rect 9272 5224 9287 5228
rect 9275 5190 9287 5224
rect 9272 5184 9287 5190
rect 9692 5216 9720 5324
rect 10413 5321 10425 5355
rect 10459 5352 10471 5355
rect 11054 5352 11060 5364
rect 10459 5324 11060 5352
rect 10459 5321 10471 5324
rect 10413 5315 10471 5321
rect 11054 5312 11060 5324
rect 11112 5312 11118 5364
rect 11514 5312 11520 5364
rect 11572 5352 11578 5364
rect 11701 5355 11759 5361
rect 11701 5352 11713 5355
rect 11572 5324 11713 5352
rect 11572 5312 11578 5324
rect 11701 5321 11713 5324
rect 11747 5321 11759 5355
rect 12161 5355 12219 5361
rect 12161 5352 12173 5355
rect 11701 5315 11759 5321
rect 11808 5324 12173 5352
rect 10318 5284 10324 5296
rect 10231 5256 10324 5284
rect 10318 5244 10324 5256
rect 10376 5284 10382 5296
rect 11808 5284 11836 5324
rect 12161 5321 12173 5324
rect 12207 5352 12219 5355
rect 12434 5352 12440 5364
rect 12207 5324 12440 5352
rect 12207 5321 12219 5324
rect 12161 5315 12219 5321
rect 12434 5312 12440 5324
rect 12492 5352 12498 5364
rect 13173 5355 13231 5361
rect 13173 5352 13185 5355
rect 12492 5324 13185 5352
rect 12492 5312 12498 5324
rect 13173 5321 13185 5324
rect 13219 5321 13231 5355
rect 13173 5315 13231 5321
rect 10376 5256 11836 5284
rect 12069 5287 12127 5293
rect 10376 5244 10382 5256
rect 12069 5253 12081 5287
rect 12115 5253 12127 5287
rect 13814 5284 13820 5296
rect 12069 5247 12127 5253
rect 12406 5256 13820 5284
rect 12084 5216 12112 5247
rect 12406 5216 12434 5256
rect 13814 5244 13820 5256
rect 13872 5244 13878 5296
rect 9692 5188 12434 5216
rect 9272 5176 9278 5184
rect 12986 5176 12992 5228
rect 13044 5216 13050 5228
rect 13265 5219 13323 5225
rect 13265 5216 13277 5219
rect 13044 5188 13277 5216
rect 13044 5176 13050 5188
rect 13265 5185 13277 5188
rect 13311 5216 13323 5219
rect 13354 5216 13360 5228
rect 13311 5188 13360 5216
rect 13311 5185 13323 5188
rect 13265 5179 13323 5185
rect 13354 5176 13360 5188
rect 13412 5176 13418 5228
rect 7193 5151 7251 5157
rect 7193 5117 7205 5151
rect 7239 5117 7251 5151
rect 7193 5111 7251 5117
rect 7837 5151 7895 5157
rect 7837 5117 7849 5151
rect 7883 5117 7895 5151
rect 8110 5148 8116 5160
rect 8071 5120 8116 5148
rect 7837 5111 7895 5117
rect 2951 5083 3009 5089
rect 2951 5049 2963 5083
rect 2997 5080 3009 5083
rect 3329 5083 3387 5089
rect 3329 5080 3341 5083
rect 2997 5052 3341 5080
rect 2997 5049 3009 5052
rect 2951 5043 3009 5049
rect 3329 5049 3341 5052
rect 3375 5080 3387 5083
rect 3953 5083 4011 5089
rect 3953 5080 3965 5083
rect 3375 5052 3965 5080
rect 3375 5049 3387 5052
rect 3329 5043 3387 5049
rect 3953 5049 3965 5052
rect 3999 5049 4011 5083
rect 3953 5043 4011 5049
rect 4246 5040 4252 5092
rect 4304 5080 4310 5092
rect 7208 5080 7236 5111
rect 8110 5108 8116 5120
rect 8168 5108 8174 5160
rect 9674 5108 9680 5160
rect 9732 5148 9738 5160
rect 10137 5151 10195 5157
rect 10137 5148 10149 5151
rect 9732 5120 10149 5148
rect 9732 5108 9738 5120
rect 10137 5117 10149 5120
rect 10183 5117 10195 5151
rect 10137 5111 10195 5117
rect 4304 5052 7236 5080
rect 4304 5040 4310 5052
rect 4154 5012 4160 5024
rect 2884 4984 4160 5012
rect 4154 4972 4160 4984
rect 4212 4972 4218 5024
rect 6641 5015 6699 5021
rect 6641 4981 6653 5015
rect 6687 5012 6699 5015
rect 6822 5012 6828 5024
rect 6687 4984 6828 5012
rect 6687 4981 6699 4984
rect 6641 4975 6699 4981
rect 6822 4972 6828 4984
rect 6880 4972 6886 5024
rect 7208 5012 7236 5052
rect 8011 5083 8069 5089
rect 8011 5049 8023 5083
rect 8057 5080 8069 5083
rect 8389 5083 8447 5089
rect 8389 5080 8401 5083
rect 8057 5052 8401 5080
rect 8057 5049 8069 5052
rect 8011 5043 8069 5049
rect 8389 5049 8401 5052
rect 8435 5080 8447 5083
rect 9013 5083 9071 5089
rect 9013 5080 9025 5083
rect 8435 5052 9025 5080
rect 8435 5049 8447 5052
rect 8389 5043 8447 5049
rect 9013 5049 9025 5052
rect 9059 5049 9071 5083
rect 10152 5080 10180 5111
rect 11882 5108 11888 5160
rect 11940 5148 11946 5160
rect 12253 5151 12311 5157
rect 12253 5148 12265 5151
rect 11940 5120 12265 5148
rect 11940 5108 11946 5120
rect 12253 5117 12265 5120
rect 12299 5117 12311 5151
rect 12253 5111 12311 5117
rect 12894 5108 12900 5160
rect 12952 5148 12958 5160
rect 13081 5151 13139 5157
rect 13081 5148 13093 5151
rect 12952 5120 13093 5148
rect 12952 5108 12958 5120
rect 13081 5117 13093 5120
rect 13127 5117 13139 5151
rect 13081 5111 13139 5117
rect 13906 5080 13912 5092
rect 10152 5052 13912 5080
rect 9013 5043 9071 5049
rect 13906 5040 13912 5052
rect 13964 5040 13970 5092
rect 9306 5012 9312 5024
rect 7208 4984 9312 5012
rect 9306 4972 9312 4984
rect 9364 5012 9370 5024
rect 9585 5015 9643 5021
rect 9585 5012 9597 5015
rect 9364 4984 9597 5012
rect 9364 4972 9370 4984
rect 9585 4981 9597 4984
rect 9631 4981 9643 5015
rect 9585 4975 9643 4981
rect 10502 4972 10508 5024
rect 10560 5012 10566 5024
rect 10781 5015 10839 5021
rect 10781 5012 10793 5015
rect 10560 4984 10793 5012
rect 10560 4972 10566 4984
rect 10781 4981 10793 4984
rect 10827 4981 10839 5015
rect 10781 4975 10839 4981
rect 13633 5015 13691 5021
rect 13633 4981 13645 5015
rect 13679 5012 13691 5015
rect 15194 5012 15200 5024
rect 13679 4984 15200 5012
rect 13679 4981 13691 4984
rect 13633 4975 13691 4981
rect 15194 4972 15200 4984
rect 15252 4972 15258 5024
rect 1104 4922 18860 4944
rect 1104 4913 3169 4922
rect 1104 4879 1133 4913
rect 1167 4879 1225 4913
rect 1259 4879 1317 4913
rect 1351 4879 1409 4913
rect 1443 4879 1501 4913
rect 1535 4879 1593 4913
rect 1627 4879 1685 4913
rect 1719 4879 1777 4913
rect 1811 4879 1869 4913
rect 1903 4879 1961 4913
rect 1995 4879 2053 4913
rect 2087 4879 2145 4913
rect 2179 4879 2237 4913
rect 2271 4879 2329 4913
rect 2363 4879 2421 4913
rect 2455 4879 2513 4913
rect 2547 4879 2605 4913
rect 2639 4879 2697 4913
rect 2731 4879 2789 4913
rect 2823 4879 2881 4913
rect 2915 4879 2973 4913
rect 3007 4879 3065 4913
rect 3099 4879 3157 4913
rect 1104 4870 3169 4879
rect 3221 4870 3233 4922
rect 3285 4870 3297 4922
rect 3349 4913 3361 4922
rect 3349 4870 3361 4879
rect 3413 4870 3425 4922
rect 3477 4913 7608 4922
rect 3477 4879 3525 4913
rect 3559 4879 3617 4913
rect 3651 4879 3709 4913
rect 3743 4879 3801 4913
rect 3835 4879 3893 4913
rect 3927 4879 3985 4913
rect 4019 4879 4077 4913
rect 4111 4879 4169 4913
rect 4203 4879 4261 4913
rect 4295 4879 4353 4913
rect 4387 4879 4445 4913
rect 4479 4879 4537 4913
rect 4571 4879 4629 4913
rect 4663 4879 4721 4913
rect 4755 4879 4813 4913
rect 4847 4879 4905 4913
rect 4939 4879 4997 4913
rect 5031 4879 5089 4913
rect 5123 4879 5181 4913
rect 5215 4879 5273 4913
rect 5307 4879 5365 4913
rect 5399 4879 5457 4913
rect 5491 4879 5549 4913
rect 5583 4879 5641 4913
rect 5675 4879 5733 4913
rect 5767 4879 5825 4913
rect 5859 4879 5917 4913
rect 5951 4879 6009 4913
rect 6043 4879 6101 4913
rect 6135 4879 6193 4913
rect 6227 4879 6285 4913
rect 6319 4879 6377 4913
rect 6411 4879 6469 4913
rect 6503 4879 6561 4913
rect 6595 4879 6653 4913
rect 6687 4879 6745 4913
rect 6779 4879 6837 4913
rect 6871 4879 6929 4913
rect 6963 4879 7021 4913
rect 7055 4879 7113 4913
rect 7147 4879 7205 4913
rect 7239 4879 7297 4913
rect 7331 4879 7389 4913
rect 7423 4879 7481 4913
rect 7515 4879 7573 4913
rect 7607 4879 7608 4913
rect 3477 4870 7608 4879
rect 7660 4913 7672 4922
rect 7660 4879 7665 4913
rect 7660 4870 7672 4879
rect 7724 4870 7736 4922
rect 7788 4913 7800 4922
rect 7852 4913 7864 4922
rect 7916 4913 12047 4922
rect 12099 4913 12111 4922
rect 12163 4913 12175 4922
rect 7791 4879 7800 4913
rect 7916 4879 7941 4913
rect 7975 4879 8033 4913
rect 8067 4879 8125 4913
rect 8159 4879 8217 4913
rect 8251 4879 8309 4913
rect 8343 4879 8401 4913
rect 8435 4879 8493 4913
rect 8527 4879 8585 4913
rect 8619 4879 8677 4913
rect 8711 4879 8769 4913
rect 8803 4879 8861 4913
rect 8895 4879 8953 4913
rect 8987 4879 9045 4913
rect 9079 4879 9137 4913
rect 9171 4879 9229 4913
rect 9263 4879 9321 4913
rect 9355 4879 9413 4913
rect 9447 4879 9505 4913
rect 9539 4879 9597 4913
rect 9631 4879 9689 4913
rect 9723 4879 9781 4913
rect 9815 4879 9873 4913
rect 9907 4879 9965 4913
rect 9999 4879 10057 4913
rect 10091 4879 10149 4913
rect 10183 4879 10241 4913
rect 10275 4879 10333 4913
rect 10367 4879 10425 4913
rect 10459 4879 10517 4913
rect 10551 4879 10609 4913
rect 10643 4879 10701 4913
rect 10735 4879 10793 4913
rect 10827 4879 10885 4913
rect 10919 4879 10977 4913
rect 11011 4879 11069 4913
rect 11103 4879 11161 4913
rect 11195 4879 11253 4913
rect 11287 4879 11345 4913
rect 11379 4879 11437 4913
rect 11471 4879 11529 4913
rect 11563 4879 11621 4913
rect 11655 4879 11713 4913
rect 11747 4879 11805 4913
rect 11839 4879 11897 4913
rect 11931 4879 11989 4913
rect 12023 4879 12047 4913
rect 12163 4879 12173 4913
rect 7788 4870 7800 4879
rect 7852 4870 7864 4879
rect 7916 4870 12047 4879
rect 12099 4870 12111 4879
rect 12163 4870 12175 4879
rect 12227 4870 12239 4922
rect 12291 4913 12303 4922
rect 12299 4879 12303 4913
rect 12291 4870 12303 4879
rect 12355 4913 16486 4922
rect 12355 4879 12357 4913
rect 12391 4879 12449 4913
rect 12483 4879 12541 4913
rect 12575 4879 12633 4913
rect 12667 4879 12725 4913
rect 12759 4879 12817 4913
rect 12851 4879 12909 4913
rect 12943 4879 13001 4913
rect 13035 4879 13093 4913
rect 13127 4879 13185 4913
rect 13219 4879 13277 4913
rect 13311 4879 13369 4913
rect 13403 4879 13461 4913
rect 13495 4879 13553 4913
rect 13587 4879 13645 4913
rect 13679 4879 13737 4913
rect 13771 4879 13829 4913
rect 13863 4879 13921 4913
rect 13955 4879 14013 4913
rect 14047 4879 14105 4913
rect 14139 4879 14197 4913
rect 14231 4879 14289 4913
rect 14323 4879 14381 4913
rect 14415 4879 14473 4913
rect 14507 4879 14565 4913
rect 14599 4879 14657 4913
rect 14691 4879 14749 4913
rect 14783 4879 14841 4913
rect 14875 4879 14933 4913
rect 14967 4879 15025 4913
rect 15059 4879 15117 4913
rect 15151 4879 15209 4913
rect 15243 4879 15301 4913
rect 15335 4879 15393 4913
rect 15427 4879 15485 4913
rect 15519 4879 15577 4913
rect 15611 4879 15669 4913
rect 15703 4879 15761 4913
rect 15795 4879 15853 4913
rect 15887 4879 15945 4913
rect 15979 4879 16037 4913
rect 16071 4879 16129 4913
rect 16163 4879 16221 4913
rect 16255 4879 16313 4913
rect 16347 4879 16405 4913
rect 16439 4879 16486 4913
rect 12355 4870 16486 4879
rect 16538 4870 16550 4922
rect 16602 4913 16614 4922
rect 16602 4870 16614 4879
rect 16666 4870 16678 4922
rect 16730 4870 16742 4922
rect 16794 4913 18860 4922
rect 16807 4879 16865 4913
rect 16899 4879 16957 4913
rect 16991 4879 17049 4913
rect 17083 4879 17141 4913
rect 17175 4879 17233 4913
rect 17267 4879 17325 4913
rect 17359 4879 17417 4913
rect 17451 4879 17509 4913
rect 17543 4879 17601 4913
rect 17635 4879 17693 4913
rect 17727 4879 17785 4913
rect 17819 4879 17877 4913
rect 17911 4879 17969 4913
rect 18003 4879 18061 4913
rect 18095 4879 18153 4913
rect 18187 4879 18245 4913
rect 18279 4879 18337 4913
rect 18371 4879 18429 4913
rect 18463 4879 18521 4913
rect 18555 4879 18613 4913
rect 18647 4879 18705 4913
rect 18739 4879 18797 4913
rect 18831 4879 18860 4913
rect 16794 4870 18860 4879
rect 1104 4848 18860 4870
rect 6914 4768 6920 4820
rect 6972 4808 6978 4820
rect 7193 4811 7251 4817
rect 7193 4808 7205 4811
rect 6972 4780 7205 4808
rect 6972 4768 6978 4780
rect 7193 4777 7205 4780
rect 7239 4777 7251 4811
rect 12713 4811 12771 4817
rect 7193 4771 7251 4777
rect 7760 4780 12204 4808
rect 3050 4700 3056 4752
rect 3108 4740 3114 4752
rect 7760 4740 7788 4780
rect 3108 4712 7788 4740
rect 7837 4743 7895 4749
rect 3108 4700 3114 4712
rect 7837 4709 7849 4743
rect 7883 4709 7895 4743
rect 7837 4703 7895 4709
rect 7852 4672 7880 4703
rect 8294 4700 8300 4752
rect 8352 4740 8358 4752
rect 11517 4743 11575 4749
rect 8352 4712 10824 4740
rect 8352 4700 8358 4712
rect 6380 4644 7880 4672
rect 2774 4564 2780 4616
rect 2832 4604 2838 4616
rect 6380 4613 6408 4644
rect 8018 4632 8024 4684
rect 8076 4672 8082 4684
rect 8202 4672 8208 4684
rect 8076 4644 8208 4672
rect 8076 4632 8082 4644
rect 8202 4632 8208 4644
rect 8260 4672 8266 4684
rect 8389 4675 8447 4681
rect 8389 4672 8401 4675
rect 8260 4644 8401 4672
rect 8260 4632 8266 4644
rect 8389 4641 8401 4644
rect 8435 4641 8447 4675
rect 10318 4672 10324 4684
rect 8389 4635 8447 4641
rect 8496 4644 10324 4672
rect 3053 4607 3111 4613
rect 3053 4604 3065 4607
rect 2832 4576 3065 4604
rect 2832 4564 2838 4576
rect 3053 4573 3065 4576
rect 3099 4604 3111 4607
rect 4893 4607 4951 4613
rect 4893 4604 4905 4607
rect 3099 4576 4905 4604
rect 3099 4573 3111 4576
rect 3053 4567 3111 4573
rect 4893 4573 4905 4576
rect 4939 4573 4951 4607
rect 4893 4567 4951 4573
rect 6365 4607 6423 4613
rect 6365 4573 6377 4607
rect 6411 4573 6423 4607
rect 6822 4604 6828 4616
rect 6783 4576 6828 4604
rect 6365 4567 6423 4573
rect 6822 4564 6828 4576
rect 6880 4564 6886 4616
rect 7374 4564 7380 4616
rect 7432 4604 7438 4616
rect 7834 4604 7840 4616
rect 7432 4576 7840 4604
rect 7432 4564 7438 4576
rect 7834 4564 7840 4576
rect 7892 4604 7898 4616
rect 8297 4607 8355 4613
rect 8297 4604 8309 4607
rect 7892 4576 8309 4604
rect 7892 4564 7898 4576
rect 8297 4573 8309 4576
rect 8343 4604 8355 4607
rect 8496 4604 8524 4644
rect 10318 4632 10324 4644
rect 10376 4632 10382 4684
rect 8343 4576 8524 4604
rect 8343 4573 8355 4576
rect 8297 4567 8355 4573
rect 9030 4564 9036 4616
rect 9088 4604 9094 4616
rect 9582 4604 9588 4616
rect 9088 4576 9588 4604
rect 9088 4564 9094 4576
rect 9582 4564 9588 4576
rect 9640 4604 9646 4616
rect 9953 4607 10011 4613
rect 9953 4604 9965 4607
rect 9640 4576 9965 4604
rect 9640 4564 9646 4576
rect 9953 4573 9965 4576
rect 9999 4573 10011 4607
rect 10502 4604 10508 4616
rect 10463 4576 10508 4604
rect 9953 4567 10011 4573
rect 10502 4564 10508 4576
rect 10560 4564 10566 4616
rect 4341 4539 4399 4545
rect 4341 4505 4353 4539
rect 4387 4536 4399 4539
rect 4982 4536 4988 4548
rect 4387 4508 4988 4536
rect 4387 4505 4399 4508
rect 4341 4499 4399 4505
rect 4982 4496 4988 4508
rect 5040 4496 5046 4548
rect 6178 4536 6184 4548
rect 6139 4508 6184 4536
rect 6178 4496 6184 4508
rect 6236 4496 6242 4548
rect 7009 4539 7067 4545
rect 7009 4505 7021 4539
rect 7055 4536 7067 4539
rect 8110 4536 8116 4548
rect 7055 4508 8116 4536
rect 7055 4505 7067 4508
rect 7009 4499 7067 4505
rect 8110 4496 8116 4508
rect 8168 4496 8174 4548
rect 8386 4496 8392 4548
rect 8444 4536 8450 4548
rect 9125 4539 9183 4545
rect 9125 4536 9137 4539
rect 8444 4508 9137 4536
rect 8444 4496 8450 4508
rect 9125 4505 9137 4508
rect 9171 4505 9183 4539
rect 9306 4536 9312 4548
rect 9267 4508 9312 4536
rect 9125 4499 9183 4505
rect 9306 4496 9312 4508
rect 9364 4496 9370 4548
rect 10686 4536 10692 4548
rect 10647 4508 10692 4536
rect 10686 4496 10692 4508
rect 10744 4496 10750 4548
rect 10796 4536 10824 4712
rect 11517 4709 11529 4743
rect 11563 4740 11575 4743
rect 11974 4740 11980 4752
rect 11563 4712 11980 4740
rect 11563 4709 11575 4712
rect 11517 4703 11575 4709
rect 11974 4700 11980 4712
rect 12032 4700 12038 4752
rect 11698 4632 11704 4684
rect 11756 4672 11762 4684
rect 12069 4675 12127 4681
rect 12069 4672 12081 4675
rect 11756 4644 12081 4672
rect 11756 4632 11762 4644
rect 12069 4641 12081 4644
rect 12115 4641 12127 4675
rect 12069 4635 12127 4641
rect 10962 4564 10968 4616
rect 11020 4604 11026 4616
rect 11333 4607 11391 4613
rect 11333 4604 11345 4607
rect 11020 4576 11345 4604
rect 11020 4564 11026 4576
rect 11333 4573 11345 4576
rect 11379 4573 11391 4607
rect 11333 4567 11391 4573
rect 11882 4536 11888 4548
rect 10796 4508 11888 4536
rect 11882 4496 11888 4508
rect 11940 4496 11946 4548
rect 12176 4536 12204 4780
rect 12713 4777 12725 4811
rect 12759 4808 12771 4811
rect 12802 4808 12808 4820
rect 12759 4780 12808 4808
rect 12759 4777 12771 4780
rect 12713 4771 12771 4777
rect 12802 4768 12808 4780
rect 12860 4768 12866 4820
rect 12342 4700 12348 4752
rect 12400 4740 12406 4752
rect 13722 4740 13728 4752
rect 12400 4712 13728 4740
rect 12400 4700 12406 4712
rect 13722 4700 13728 4712
rect 13780 4700 13786 4752
rect 16850 4740 16856 4752
rect 13832 4712 16856 4740
rect 12253 4675 12311 4681
rect 12253 4641 12265 4675
rect 12299 4672 12311 4675
rect 12434 4672 12440 4684
rect 12299 4644 12440 4672
rect 12299 4641 12311 4644
rect 12253 4635 12311 4641
rect 12434 4632 12440 4644
rect 12492 4632 12498 4684
rect 13832 4672 13860 4712
rect 16850 4700 16856 4712
rect 16908 4700 16914 4752
rect 13004 4644 13860 4672
rect 12342 4564 12348 4616
rect 12400 4604 12406 4616
rect 13004 4604 13032 4644
rect 15102 4632 15108 4684
rect 15160 4672 15166 4684
rect 15160 4644 16252 4672
rect 15160 4632 15166 4644
rect 12400 4576 13032 4604
rect 12400 4564 12406 4576
rect 13078 4564 13084 4616
rect 13136 4604 13142 4616
rect 13357 4607 13415 4613
rect 13357 4604 13369 4607
rect 13136 4576 13369 4604
rect 13136 4564 13142 4576
rect 13357 4573 13369 4576
rect 13403 4573 13415 4607
rect 15194 4604 15200 4616
rect 15155 4576 15200 4604
rect 13357 4567 13415 4573
rect 15194 4564 15200 4576
rect 15252 4564 15258 4616
rect 16224 4613 16252 4644
rect 16209 4607 16267 4613
rect 16209 4573 16221 4607
rect 16255 4573 16267 4607
rect 16853 4607 16911 4613
rect 16853 4604 16865 4607
rect 16209 4567 16267 4573
rect 16546 4576 16865 4604
rect 15378 4536 15384 4548
rect 12176 4508 13216 4536
rect 15339 4508 15384 4536
rect 2222 4428 2228 4480
rect 2280 4468 2286 4480
rect 2409 4471 2467 4477
rect 2409 4468 2421 4471
rect 2280 4440 2421 4468
rect 2280 4428 2286 4440
rect 2409 4437 2421 4440
rect 2455 4437 2467 4471
rect 2409 4431 2467 4437
rect 4065 4471 4123 4477
rect 4065 4437 4077 4471
rect 4111 4468 4123 4471
rect 4430 4468 4436 4480
rect 4111 4440 4436 4468
rect 4111 4437 4123 4440
rect 4065 4431 4123 4437
rect 4430 4428 4436 4440
rect 4488 4428 4494 4480
rect 5997 4471 6055 4477
rect 5997 4437 6009 4471
rect 6043 4468 6055 4471
rect 6822 4468 6828 4480
rect 6043 4440 6828 4468
rect 6043 4437 6055 4440
rect 5997 4431 6055 4437
rect 6822 4428 6828 4440
rect 6880 4428 6886 4480
rect 7282 4428 7288 4480
rect 7340 4468 7346 4480
rect 8205 4471 8263 4477
rect 8205 4468 8217 4471
rect 7340 4440 8217 4468
rect 7340 4428 7346 4440
rect 8205 4437 8217 4440
rect 8251 4437 8263 4471
rect 8205 4431 8263 4437
rect 8846 4428 8852 4480
rect 8904 4468 8910 4480
rect 9398 4468 9404 4480
rect 8904 4440 9404 4468
rect 8904 4428 8910 4440
rect 9398 4428 9404 4440
rect 9456 4428 9462 4480
rect 9493 4471 9551 4477
rect 9493 4437 9505 4471
rect 9539 4468 9551 4471
rect 10226 4468 10232 4480
rect 9539 4440 10232 4468
rect 9539 4437 9551 4440
rect 9493 4431 9551 4437
rect 10226 4428 10232 4440
rect 10284 4428 10290 4480
rect 10873 4471 10931 4477
rect 10873 4437 10885 4471
rect 10919 4468 10931 4471
rect 10962 4468 10968 4480
rect 10919 4440 10968 4468
rect 10919 4437 10931 4440
rect 10873 4431 10931 4437
rect 10962 4428 10968 4440
rect 11020 4428 11026 4480
rect 11054 4428 11060 4480
rect 11112 4468 11118 4480
rect 12342 4468 12348 4480
rect 11112 4440 12348 4468
rect 11112 4428 11118 4440
rect 12342 4428 12348 4440
rect 12400 4428 12406 4480
rect 13188 4477 13216 4508
rect 15378 4496 15384 4508
rect 15436 4496 15442 4548
rect 15565 4539 15623 4545
rect 15565 4505 15577 4539
rect 15611 4536 15623 4539
rect 16546 4536 16574 4576
rect 16853 4573 16865 4576
rect 16899 4573 16911 4607
rect 16853 4567 16911 4573
rect 15611 4508 16574 4536
rect 15611 4505 15623 4508
rect 15565 4499 15623 4505
rect 13173 4471 13231 4477
rect 13173 4437 13185 4471
rect 13219 4437 13231 4471
rect 16022 4468 16028 4480
rect 15983 4440 16028 4468
rect 13173 4431 13231 4437
rect 16022 4428 16028 4440
rect 16080 4428 16086 4480
rect 16669 4471 16727 4477
rect 16669 4437 16681 4471
rect 16715 4468 16727 4471
rect 16850 4468 16856 4480
rect 16715 4440 16856 4468
rect 16715 4437 16727 4440
rect 16669 4431 16727 4437
rect 16850 4428 16856 4440
rect 16908 4428 16914 4480
rect 1104 4378 19019 4400
rect 1104 4369 5388 4378
rect 1104 4335 1133 4369
rect 1167 4335 1225 4369
rect 1259 4335 1317 4369
rect 1351 4335 1409 4369
rect 1443 4335 1501 4369
rect 1535 4335 1593 4369
rect 1627 4335 1685 4369
rect 1719 4335 1777 4369
rect 1811 4335 1869 4369
rect 1903 4335 1961 4369
rect 1995 4335 2053 4369
rect 2087 4335 2145 4369
rect 2179 4335 2237 4369
rect 2271 4335 2329 4369
rect 2363 4335 2421 4369
rect 2455 4335 2513 4369
rect 2547 4335 2605 4369
rect 2639 4335 2697 4369
rect 2731 4335 2789 4369
rect 2823 4335 2881 4369
rect 2915 4335 2973 4369
rect 3007 4335 3065 4369
rect 3099 4335 3157 4369
rect 3191 4335 3249 4369
rect 3283 4335 3341 4369
rect 3375 4335 3433 4369
rect 3467 4335 3525 4369
rect 3559 4335 3617 4369
rect 3651 4335 3709 4369
rect 3743 4335 3801 4369
rect 3835 4335 3893 4369
rect 3927 4335 3985 4369
rect 4019 4335 4077 4369
rect 4111 4335 4169 4369
rect 4203 4335 4261 4369
rect 4295 4335 4353 4369
rect 4387 4335 4445 4369
rect 4479 4335 4537 4369
rect 4571 4335 4629 4369
rect 4663 4335 4721 4369
rect 4755 4335 4813 4369
rect 4847 4335 4905 4369
rect 4939 4335 4997 4369
rect 5031 4335 5089 4369
rect 5123 4335 5181 4369
rect 5215 4335 5273 4369
rect 5307 4335 5365 4369
rect 1104 4326 5388 4335
rect 5440 4326 5452 4378
rect 5504 4326 5516 4378
rect 5568 4369 5580 4378
rect 5632 4369 5644 4378
rect 5696 4369 9827 4378
rect 9879 4369 9891 4378
rect 5632 4335 5641 4369
rect 5696 4335 5733 4369
rect 5767 4335 5825 4369
rect 5859 4335 5917 4369
rect 5951 4335 6009 4369
rect 6043 4335 6101 4369
rect 6135 4335 6193 4369
rect 6227 4335 6285 4369
rect 6319 4335 6377 4369
rect 6411 4335 6469 4369
rect 6503 4335 6561 4369
rect 6595 4335 6653 4369
rect 6687 4335 6745 4369
rect 6779 4335 6837 4369
rect 6871 4335 6929 4369
rect 6963 4335 7021 4369
rect 7055 4335 7113 4369
rect 7147 4335 7205 4369
rect 7239 4335 7297 4369
rect 7331 4335 7389 4369
rect 7423 4335 7481 4369
rect 7515 4335 7573 4369
rect 7607 4335 7665 4369
rect 7699 4335 7757 4369
rect 7791 4335 7849 4369
rect 7883 4335 7941 4369
rect 7975 4335 8033 4369
rect 8067 4335 8125 4369
rect 8159 4335 8217 4369
rect 8251 4335 8309 4369
rect 8343 4335 8401 4369
rect 8435 4335 8493 4369
rect 8527 4335 8585 4369
rect 8619 4335 8677 4369
rect 8711 4335 8769 4369
rect 8803 4335 8861 4369
rect 8895 4335 8953 4369
rect 8987 4335 9045 4369
rect 9079 4335 9137 4369
rect 9171 4335 9229 4369
rect 9263 4335 9321 4369
rect 9355 4335 9413 4369
rect 9447 4335 9505 4369
rect 9539 4335 9597 4369
rect 9631 4335 9689 4369
rect 9723 4335 9781 4369
rect 9815 4335 9827 4369
rect 5568 4326 5580 4335
rect 5632 4326 5644 4335
rect 5696 4326 9827 4335
rect 9879 4326 9891 4335
rect 9943 4326 9955 4378
rect 10007 4326 10019 4378
rect 10071 4369 10083 4378
rect 10135 4369 14266 4378
rect 14318 4369 14330 4378
rect 14382 4369 14394 4378
rect 10135 4335 10149 4369
rect 10183 4335 10241 4369
rect 10275 4335 10333 4369
rect 10367 4335 10425 4369
rect 10459 4335 10517 4369
rect 10551 4335 10609 4369
rect 10643 4335 10701 4369
rect 10735 4335 10793 4369
rect 10827 4335 10885 4369
rect 10919 4335 10977 4369
rect 11011 4335 11069 4369
rect 11103 4335 11161 4369
rect 11195 4335 11253 4369
rect 11287 4335 11345 4369
rect 11379 4335 11437 4369
rect 11471 4335 11529 4369
rect 11563 4335 11621 4369
rect 11655 4335 11713 4369
rect 11747 4335 11805 4369
rect 11839 4335 11897 4369
rect 11931 4335 11989 4369
rect 12023 4335 12081 4369
rect 12115 4335 12173 4369
rect 12207 4335 12265 4369
rect 12299 4335 12357 4369
rect 12391 4335 12449 4369
rect 12483 4335 12541 4369
rect 12575 4335 12633 4369
rect 12667 4335 12725 4369
rect 12759 4335 12817 4369
rect 12851 4335 12909 4369
rect 12943 4335 13001 4369
rect 13035 4335 13093 4369
rect 13127 4335 13185 4369
rect 13219 4335 13277 4369
rect 13311 4335 13369 4369
rect 13403 4335 13461 4369
rect 13495 4335 13553 4369
rect 13587 4335 13645 4369
rect 13679 4335 13737 4369
rect 13771 4335 13829 4369
rect 13863 4335 13921 4369
rect 13955 4335 14013 4369
rect 14047 4335 14105 4369
rect 14139 4335 14197 4369
rect 14231 4335 14266 4369
rect 14323 4335 14330 4369
rect 10071 4326 10083 4335
rect 10135 4326 14266 4335
rect 14318 4326 14330 4335
rect 14382 4326 14394 4335
rect 14446 4326 14458 4378
rect 14510 4326 14522 4378
rect 14574 4369 18705 4378
rect 14599 4335 14657 4369
rect 14691 4335 14749 4369
rect 14783 4335 14841 4369
rect 14875 4335 14933 4369
rect 14967 4335 15025 4369
rect 15059 4335 15117 4369
rect 15151 4335 15209 4369
rect 15243 4335 15301 4369
rect 15335 4335 15393 4369
rect 15427 4335 15485 4369
rect 15519 4335 15577 4369
rect 15611 4335 15669 4369
rect 15703 4335 15761 4369
rect 15795 4335 15853 4369
rect 15887 4335 15945 4369
rect 15979 4335 16037 4369
rect 16071 4335 16129 4369
rect 16163 4335 16221 4369
rect 16255 4335 16313 4369
rect 16347 4335 16405 4369
rect 16439 4335 16497 4369
rect 16531 4335 16589 4369
rect 16623 4335 16681 4369
rect 16715 4335 16773 4369
rect 16807 4335 16865 4369
rect 16899 4335 16957 4369
rect 16991 4335 17049 4369
rect 17083 4335 17141 4369
rect 17175 4335 17233 4369
rect 17267 4335 17325 4369
rect 17359 4335 17417 4369
rect 17451 4335 17509 4369
rect 17543 4335 17601 4369
rect 17635 4335 17693 4369
rect 17727 4335 17785 4369
rect 17819 4335 17877 4369
rect 17911 4335 17969 4369
rect 18003 4335 18061 4369
rect 18095 4335 18153 4369
rect 18187 4335 18245 4369
rect 18279 4335 18337 4369
rect 18371 4335 18429 4369
rect 18463 4335 18521 4369
rect 18555 4335 18613 4369
rect 18647 4335 18705 4369
rect 14574 4326 18705 4335
rect 18757 4326 18769 4378
rect 18821 4369 18833 4378
rect 18831 4335 18833 4369
rect 18821 4326 18833 4335
rect 18885 4326 18897 4378
rect 18949 4326 18961 4378
rect 19013 4326 19019 4378
rect 1104 4304 19019 4326
rect 2409 4267 2467 4273
rect 2409 4233 2421 4267
rect 2455 4264 2467 4267
rect 4982 4264 4988 4276
rect 2455 4236 4988 4264
rect 2455 4233 2467 4236
rect 2409 4227 2467 4233
rect 4982 4224 4988 4236
rect 5040 4224 5046 4276
rect 6178 4224 6184 4276
rect 6236 4264 6242 4276
rect 6236 4236 7880 4264
rect 6236 4224 6242 4236
rect 3601 4199 3731 4205
rect 3601 4165 3613 4199
rect 3647 4165 3685 4199
rect 3719 4196 3731 4199
rect 4321 4199 4379 4205
rect 4321 4196 4333 4199
rect 3719 4168 4333 4196
rect 3719 4165 3731 4168
rect 3601 4159 3731 4165
rect 4261 4165 4333 4168
rect 4367 4196 4379 4199
rect 4430 4196 4436 4208
rect 4367 4168 4436 4196
rect 4367 4165 4379 4168
rect 4261 4159 4379 4165
rect 2222 4128 2228 4140
rect 2183 4100 2228 4128
rect 2222 4088 2228 4100
rect 2280 4088 2286 4140
rect 2962 4131 3020 4137
rect 2962 4097 2974 4131
rect 3008 4128 3020 4131
rect 3329 4131 3387 4137
rect 3329 4128 3341 4131
rect 3008 4100 3341 4128
rect 3008 4097 3020 4100
rect 2962 4091 3020 4097
rect 3329 4097 3341 4100
rect 3375 4128 3387 4131
rect 4045 4131 4103 4137
rect 4045 4128 4057 4131
rect 3375 4100 4057 4128
rect 3375 4097 3387 4100
rect 3329 4091 3387 4097
rect 4045 4097 4057 4100
rect 4091 4097 4103 4131
rect 4045 4091 4103 4097
rect 4261 4136 4319 4159
rect 4430 4156 4436 4168
rect 4488 4196 4494 4208
rect 5258 4196 5264 4208
rect 4488 4168 5264 4196
rect 4488 4156 4494 4168
rect 5258 4156 5264 4168
rect 5316 4156 5322 4208
rect 7282 4196 7288 4208
rect 6656 4168 7288 4196
rect 4261 4102 4273 4136
rect 4307 4102 4319 4136
rect 4261 4096 4319 4102
rect 4706 4088 4712 4140
rect 4764 4128 4770 4140
rect 6656 4128 6684 4168
rect 7282 4156 7288 4168
rect 7340 4156 7346 4208
rect 7852 4196 7880 4236
rect 7926 4224 7932 4276
rect 7984 4264 7990 4276
rect 8021 4267 8079 4273
rect 8021 4264 8033 4267
rect 7984 4236 8033 4264
rect 7984 4224 7990 4236
rect 8021 4233 8033 4236
rect 8067 4233 8079 4267
rect 8386 4264 8392 4276
rect 8347 4236 8392 4264
rect 8021 4227 8079 4233
rect 8386 4224 8392 4236
rect 8444 4224 8450 4276
rect 9030 4264 9036 4276
rect 8956 4236 9036 4264
rect 8846 4196 8852 4208
rect 7852 4168 8852 4196
rect 8846 4156 8852 4168
rect 8904 4156 8910 4208
rect 8956 4205 8984 4236
rect 9030 4224 9036 4236
rect 9088 4224 9094 4276
rect 11146 4224 11152 4276
rect 11204 4264 11210 4276
rect 11701 4267 11759 4273
rect 11701 4264 11713 4267
rect 11204 4236 11713 4264
rect 11204 4224 11210 4236
rect 11701 4233 11713 4236
rect 11747 4233 11759 4267
rect 11701 4227 11759 4233
rect 11882 4224 11888 4276
rect 11940 4264 11946 4276
rect 11940 4236 12848 4264
rect 11940 4224 11946 4236
rect 8943 4199 9001 4205
rect 8943 4165 8955 4199
rect 8989 4165 9001 4199
rect 8943 4159 9001 4165
rect 9398 4156 9404 4208
rect 9456 4196 9462 4208
rect 11790 4196 11796 4208
rect 9456 4168 11796 4196
rect 9456 4156 9462 4168
rect 11790 4156 11796 4168
rect 11848 4156 11854 4208
rect 11997 4199 12055 4205
rect 11997 4165 12009 4199
rect 12043 4196 12055 4199
rect 12645 4199 12775 4205
rect 12645 4196 12657 4199
rect 12043 4168 12657 4196
rect 12043 4165 12115 4168
rect 11997 4159 12115 4165
rect 12645 4165 12657 4168
rect 12691 4165 12729 4199
rect 12763 4196 12775 4199
rect 12820 4196 12848 4236
rect 14641 4199 14771 4205
rect 14641 4196 14653 4199
rect 12763 4168 14653 4196
rect 12763 4165 12775 4168
rect 12645 4159 12775 4165
rect 14641 4165 14653 4168
rect 14687 4165 14725 4199
rect 14759 4196 14771 4199
rect 15361 4199 15419 4205
rect 15361 4196 15373 4199
rect 14759 4168 15373 4196
rect 14759 4165 14771 4168
rect 14641 4159 14771 4165
rect 15301 4165 15373 4168
rect 15407 4165 15419 4199
rect 15301 4159 15419 4165
rect 6822 4128 6828 4140
rect 4764 4100 6684 4128
rect 6783 4100 6828 4128
rect 4764 4088 4770 4100
rect 6822 4088 6828 4100
rect 6880 4088 6886 4140
rect 7466 4088 7472 4140
rect 7524 4128 7530 4140
rect 11882 4128 11888 4140
rect 7524 4100 11888 4128
rect 7524 4088 7530 4100
rect 11882 4088 11888 4100
rect 11940 4088 11946 4140
rect 12057 4136 12115 4159
rect 12057 4102 12069 4136
rect 12103 4102 12115 4136
rect 12057 4096 12115 4102
rect 12273 4131 12331 4137
rect 12273 4097 12285 4131
rect 12319 4128 12331 4131
rect 12989 4131 13047 4137
rect 12989 4128 13001 4131
rect 12319 4100 13001 4128
rect 12319 4097 12331 4100
rect 12273 4091 12331 4097
rect 12989 4097 13001 4100
rect 13035 4128 13047 4131
rect 13356 4131 13414 4137
rect 13356 4128 13368 4131
rect 13035 4100 13368 4128
rect 13035 4097 13047 4100
rect 12989 4091 13047 4097
rect 13356 4097 13368 4100
rect 13402 4097 13414 4131
rect 13356 4091 13414 4097
rect 14002 4131 14060 4137
rect 14002 4097 14014 4131
rect 14048 4128 14060 4131
rect 14369 4131 14427 4137
rect 14369 4128 14381 4131
rect 14048 4100 14381 4128
rect 14048 4097 14060 4100
rect 14002 4091 14060 4097
rect 14369 4097 14381 4100
rect 14415 4128 14427 4131
rect 15085 4131 15143 4137
rect 15085 4128 15097 4131
rect 14415 4100 15097 4128
rect 14415 4097 14427 4100
rect 14369 4091 14427 4097
rect 15085 4097 15097 4100
rect 15131 4097 15143 4131
rect 15085 4091 15143 4097
rect 15301 4136 15359 4159
rect 15301 4102 15313 4136
rect 15347 4102 15359 4136
rect 15301 4096 15359 4102
rect 2869 4063 2927 4069
rect 2869 4029 2881 4063
rect 2915 4029 2927 4063
rect 2869 4023 2927 4029
rect 3145 4063 3203 4069
rect 3145 4029 3157 4063
rect 3191 4060 3203 4063
rect 3191 4032 6684 4060
rect 3191 4029 3203 4032
rect 3145 4023 3203 4029
rect 2498 3884 2504 3936
rect 2556 3924 2562 3936
rect 2884 3924 2912 4023
rect 3043 3995 3101 4001
rect 3043 3961 3055 3995
rect 3089 3992 3101 3995
rect 3421 3995 3479 4001
rect 3421 3992 3433 3995
rect 3089 3964 3433 3992
rect 3089 3961 3101 3964
rect 3043 3955 3101 3961
rect 3421 3961 3433 3964
rect 3467 3992 3479 3995
rect 4045 3995 4103 4001
rect 4045 3992 4057 3995
rect 3467 3964 4057 3992
rect 3467 3961 3479 3964
rect 3421 3955 3479 3961
rect 4045 3961 4057 3964
rect 4091 3961 4103 3995
rect 4045 3955 4103 3961
rect 4522 3952 4528 4004
rect 4580 3992 4586 4004
rect 6656 4001 6684 4032
rect 7098 4020 7104 4072
rect 7156 4060 7162 4072
rect 7745 4063 7803 4069
rect 7745 4060 7757 4063
rect 7156 4032 7757 4060
rect 7156 4020 7162 4032
rect 7745 4029 7757 4032
rect 7791 4029 7803 4063
rect 7745 4023 7803 4029
rect 7834 4020 7840 4072
rect 7892 4060 7898 4072
rect 7929 4063 7987 4069
rect 7929 4060 7941 4063
rect 7892 4032 7941 4060
rect 7892 4020 7898 4032
rect 7929 4029 7941 4032
rect 7975 4029 7987 4063
rect 11054 4060 11060 4072
rect 7929 4023 7987 4029
rect 8404 4032 11060 4060
rect 5077 3995 5135 4001
rect 5077 3992 5089 3995
rect 4580 3964 5089 3992
rect 4580 3952 4586 3964
rect 5077 3961 5089 3964
rect 5123 3961 5135 3995
rect 5077 3955 5135 3961
rect 6641 3995 6699 4001
rect 6641 3961 6653 3995
rect 6687 3961 6699 3995
rect 6641 3955 6699 3961
rect 6914 3952 6920 4004
rect 6972 3992 6978 4004
rect 8404 3992 8432 4032
rect 11054 4020 11060 4032
rect 11112 4020 11118 4072
rect 11146 4020 11152 4072
rect 11204 4060 11210 4072
rect 13173 4063 13231 4069
rect 13173 4060 13185 4063
rect 11204 4032 13185 4060
rect 11204 4020 11210 4032
rect 13173 4029 13185 4032
rect 13219 4029 13231 4063
rect 13173 4023 13231 4029
rect 13449 4063 13507 4069
rect 13449 4029 13461 4063
rect 13495 4060 13507 4063
rect 13630 4060 13636 4072
rect 13495 4032 13636 4060
rect 13495 4029 13507 4032
rect 13449 4023 13507 4029
rect 13630 4020 13636 4032
rect 13688 4060 13694 4072
rect 13909 4063 13967 4069
rect 13909 4060 13921 4063
rect 13688 4032 13921 4060
rect 13688 4020 13694 4032
rect 13909 4029 13921 4032
rect 13955 4029 13967 4063
rect 14185 4063 14243 4069
rect 14185 4060 14197 4063
rect 13909 4023 13967 4029
rect 14016 4032 14197 4060
rect 6972 3964 8432 3992
rect 6972 3952 6978 3964
rect 8478 3952 8484 4004
rect 8536 3992 8542 4004
rect 12273 3995 12331 4001
rect 8536 3964 11836 3992
rect 8536 3952 8542 3964
rect 4154 3924 4160 3936
rect 2556 3896 4160 3924
rect 2556 3884 2562 3896
rect 4154 3884 4160 3896
rect 4212 3884 4218 3936
rect 4617 3927 4675 3933
rect 4617 3893 4629 3927
rect 4663 3924 4675 3927
rect 4706 3924 4712 3936
rect 4663 3896 4712 3924
rect 4663 3893 4675 3896
rect 4617 3887 4675 3893
rect 4706 3884 4712 3896
rect 4764 3884 4770 3936
rect 4982 3884 4988 3936
rect 5040 3924 5046 3936
rect 9122 3924 9128 3936
rect 5040 3896 9128 3924
rect 5040 3884 5046 3896
rect 9122 3884 9128 3896
rect 9180 3884 9186 3936
rect 9398 3884 9404 3936
rect 9456 3924 9462 3936
rect 10229 3927 10287 3933
rect 10229 3924 10241 3927
rect 9456 3896 10241 3924
rect 9456 3884 9462 3896
rect 10229 3893 10241 3896
rect 10275 3893 10287 3927
rect 11808 3924 11836 3964
rect 12273 3961 12285 3995
rect 12319 3992 12331 3995
rect 12897 3995 12955 4001
rect 12897 3992 12909 3995
rect 12319 3964 12909 3992
rect 12319 3961 12331 3964
rect 12273 3955 12331 3961
rect 12897 3961 12909 3964
rect 12943 3992 12955 3995
rect 13275 3995 13333 4001
rect 13275 3992 13287 3995
rect 12943 3964 13287 3992
rect 12943 3961 12955 3964
rect 12897 3955 12955 3961
rect 13275 3961 13287 3964
rect 13321 3961 13333 3995
rect 13275 3955 13333 3961
rect 13722 3952 13728 4004
rect 13780 3992 13786 4004
rect 14016 3992 14044 4032
rect 14185 4029 14197 4032
rect 14231 4029 14243 4063
rect 14185 4023 14243 4029
rect 13780 3964 14044 3992
rect 14083 3995 14141 4001
rect 13780 3952 13786 3964
rect 14083 3961 14095 3995
rect 14129 3992 14141 3995
rect 14461 3995 14519 4001
rect 14461 3992 14473 3995
rect 14129 3964 14473 3992
rect 14129 3961 14141 3964
rect 14083 3955 14141 3961
rect 14461 3961 14473 3964
rect 14507 3992 14519 3995
rect 15085 3995 15143 4001
rect 15085 3992 15097 3995
rect 14507 3964 15097 3992
rect 14507 3961 14519 3964
rect 14461 3955 14519 3961
rect 15085 3961 15097 3964
rect 15131 3961 15143 3995
rect 15085 3955 15143 3961
rect 12986 3924 12992 3936
rect 11808 3896 12992 3924
rect 10229 3887 10287 3893
rect 12986 3884 12992 3896
rect 13044 3884 13050 3936
rect 13078 3884 13084 3936
rect 13136 3924 13142 3936
rect 15657 3927 15715 3933
rect 15657 3924 15669 3927
rect 13136 3896 15669 3924
rect 13136 3884 13142 3896
rect 15657 3893 15669 3896
rect 15703 3893 15715 3927
rect 15657 3887 15715 3893
rect 1104 3834 18860 3856
rect 1104 3825 3169 3834
rect 1104 3791 1133 3825
rect 1167 3791 1225 3825
rect 1259 3791 1317 3825
rect 1351 3791 1409 3825
rect 1443 3791 1501 3825
rect 1535 3791 1593 3825
rect 1627 3791 1685 3825
rect 1719 3791 1777 3825
rect 1811 3791 1869 3825
rect 1903 3791 1961 3825
rect 1995 3791 2053 3825
rect 2087 3791 2145 3825
rect 2179 3791 2237 3825
rect 2271 3791 2329 3825
rect 2363 3791 2421 3825
rect 2455 3791 2513 3825
rect 2547 3791 2605 3825
rect 2639 3791 2697 3825
rect 2731 3791 2789 3825
rect 2823 3791 2881 3825
rect 2915 3791 2973 3825
rect 3007 3791 3065 3825
rect 3099 3791 3157 3825
rect 1104 3782 3169 3791
rect 3221 3782 3233 3834
rect 3285 3782 3297 3834
rect 3349 3825 3361 3834
rect 3349 3782 3361 3791
rect 3413 3782 3425 3834
rect 3477 3825 7608 3834
rect 3477 3791 3525 3825
rect 3559 3791 3617 3825
rect 3651 3791 3709 3825
rect 3743 3791 3801 3825
rect 3835 3791 3893 3825
rect 3927 3791 3985 3825
rect 4019 3791 4077 3825
rect 4111 3791 4169 3825
rect 4203 3791 4261 3825
rect 4295 3791 4353 3825
rect 4387 3791 4445 3825
rect 4479 3791 4537 3825
rect 4571 3791 4629 3825
rect 4663 3791 4721 3825
rect 4755 3791 4813 3825
rect 4847 3791 4905 3825
rect 4939 3791 4997 3825
rect 5031 3791 5089 3825
rect 5123 3791 5181 3825
rect 5215 3791 5273 3825
rect 5307 3791 5365 3825
rect 5399 3791 5457 3825
rect 5491 3791 5549 3825
rect 5583 3791 5641 3825
rect 5675 3791 5733 3825
rect 5767 3791 5825 3825
rect 5859 3791 5917 3825
rect 5951 3791 6009 3825
rect 6043 3791 6101 3825
rect 6135 3791 6193 3825
rect 6227 3791 6285 3825
rect 6319 3791 6377 3825
rect 6411 3791 6469 3825
rect 6503 3791 6561 3825
rect 6595 3791 6653 3825
rect 6687 3791 6745 3825
rect 6779 3791 6837 3825
rect 6871 3791 6929 3825
rect 6963 3791 7021 3825
rect 7055 3791 7113 3825
rect 7147 3791 7205 3825
rect 7239 3791 7297 3825
rect 7331 3791 7389 3825
rect 7423 3791 7481 3825
rect 7515 3791 7573 3825
rect 7607 3791 7608 3825
rect 3477 3782 7608 3791
rect 7660 3825 7672 3834
rect 7660 3791 7665 3825
rect 7660 3782 7672 3791
rect 7724 3782 7736 3834
rect 7788 3825 7800 3834
rect 7852 3825 7864 3834
rect 7916 3825 12047 3834
rect 12099 3825 12111 3834
rect 12163 3825 12175 3834
rect 7791 3791 7800 3825
rect 7916 3791 7941 3825
rect 7975 3791 8033 3825
rect 8067 3791 8125 3825
rect 8159 3791 8217 3825
rect 8251 3791 8309 3825
rect 8343 3791 8401 3825
rect 8435 3791 8493 3825
rect 8527 3791 8585 3825
rect 8619 3791 8677 3825
rect 8711 3791 8769 3825
rect 8803 3791 8861 3825
rect 8895 3791 8953 3825
rect 8987 3791 9045 3825
rect 9079 3791 9137 3825
rect 9171 3791 9229 3825
rect 9263 3791 9321 3825
rect 9355 3791 9413 3825
rect 9447 3791 9505 3825
rect 9539 3791 9597 3825
rect 9631 3791 9689 3825
rect 9723 3791 9781 3825
rect 9815 3791 9873 3825
rect 9907 3791 9965 3825
rect 9999 3791 10057 3825
rect 10091 3791 10149 3825
rect 10183 3791 10241 3825
rect 10275 3791 10333 3825
rect 10367 3791 10425 3825
rect 10459 3791 10517 3825
rect 10551 3791 10609 3825
rect 10643 3791 10701 3825
rect 10735 3791 10793 3825
rect 10827 3791 10885 3825
rect 10919 3791 10977 3825
rect 11011 3791 11069 3825
rect 11103 3791 11161 3825
rect 11195 3791 11253 3825
rect 11287 3791 11345 3825
rect 11379 3791 11437 3825
rect 11471 3791 11529 3825
rect 11563 3791 11621 3825
rect 11655 3791 11713 3825
rect 11747 3791 11805 3825
rect 11839 3791 11897 3825
rect 11931 3791 11989 3825
rect 12023 3791 12047 3825
rect 12163 3791 12173 3825
rect 7788 3782 7800 3791
rect 7852 3782 7864 3791
rect 7916 3782 12047 3791
rect 12099 3782 12111 3791
rect 12163 3782 12175 3791
rect 12227 3782 12239 3834
rect 12291 3825 12303 3834
rect 12299 3791 12303 3825
rect 12291 3782 12303 3791
rect 12355 3825 16486 3834
rect 12355 3791 12357 3825
rect 12391 3791 12449 3825
rect 12483 3791 12541 3825
rect 12575 3791 12633 3825
rect 12667 3791 12725 3825
rect 12759 3791 12817 3825
rect 12851 3791 12909 3825
rect 12943 3791 13001 3825
rect 13035 3791 13093 3825
rect 13127 3791 13185 3825
rect 13219 3791 13277 3825
rect 13311 3791 13369 3825
rect 13403 3791 13461 3825
rect 13495 3791 13553 3825
rect 13587 3791 13645 3825
rect 13679 3791 13737 3825
rect 13771 3791 13829 3825
rect 13863 3791 13921 3825
rect 13955 3791 14013 3825
rect 14047 3791 14105 3825
rect 14139 3791 14197 3825
rect 14231 3791 14289 3825
rect 14323 3791 14381 3825
rect 14415 3791 14473 3825
rect 14507 3791 14565 3825
rect 14599 3791 14657 3825
rect 14691 3791 14749 3825
rect 14783 3791 14841 3825
rect 14875 3791 14933 3825
rect 14967 3791 15025 3825
rect 15059 3791 15117 3825
rect 15151 3791 15209 3825
rect 15243 3791 15301 3825
rect 15335 3791 15393 3825
rect 15427 3791 15485 3825
rect 15519 3791 15577 3825
rect 15611 3791 15669 3825
rect 15703 3791 15761 3825
rect 15795 3791 15853 3825
rect 15887 3791 15945 3825
rect 15979 3791 16037 3825
rect 16071 3791 16129 3825
rect 16163 3791 16221 3825
rect 16255 3791 16313 3825
rect 16347 3791 16405 3825
rect 16439 3791 16486 3825
rect 12355 3782 16486 3791
rect 16538 3782 16550 3834
rect 16602 3825 16614 3834
rect 16602 3782 16614 3791
rect 16666 3782 16678 3834
rect 16730 3782 16742 3834
rect 16794 3825 18860 3834
rect 16807 3791 16865 3825
rect 16899 3791 16957 3825
rect 16991 3791 17049 3825
rect 17083 3791 17141 3825
rect 17175 3791 17233 3825
rect 17267 3791 17325 3825
rect 17359 3791 17417 3825
rect 17451 3791 17509 3825
rect 17543 3791 17601 3825
rect 17635 3791 17693 3825
rect 17727 3791 17785 3825
rect 17819 3791 17877 3825
rect 17911 3791 17969 3825
rect 18003 3791 18061 3825
rect 18095 3791 18153 3825
rect 18187 3791 18245 3825
rect 18279 3791 18337 3825
rect 18371 3791 18429 3825
rect 18463 3791 18521 3825
rect 18555 3791 18613 3825
rect 18647 3791 18705 3825
rect 18739 3791 18797 3825
rect 18831 3791 18860 3825
rect 16794 3782 18860 3791
rect 1104 3760 18860 3782
rect 1936 3723 1994 3729
rect 1936 3689 1948 3723
rect 1982 3720 1994 3723
rect 1982 3692 4108 3720
rect 1982 3689 1994 3692
rect 1936 3683 1994 3689
rect 1847 3655 1905 3661
rect 1847 3621 1859 3655
rect 1893 3652 1905 3655
rect 2225 3655 2283 3661
rect 2225 3652 2237 3655
rect 1893 3624 2237 3652
rect 1893 3621 1905 3624
rect 1847 3615 1905 3621
rect 2225 3621 2237 3624
rect 2271 3652 2283 3655
rect 2849 3655 2907 3661
rect 2849 3652 2861 3655
rect 2271 3624 2861 3652
rect 2271 3621 2283 3624
rect 2225 3615 2283 3621
rect 2849 3621 2861 3624
rect 2895 3621 2907 3655
rect 4080 3652 4108 3692
rect 4154 3680 4160 3732
rect 4212 3720 4218 3732
rect 4985 3723 5043 3729
rect 4985 3720 4997 3723
rect 4212 3692 4997 3720
rect 4212 3680 4218 3692
rect 4985 3689 4997 3692
rect 5031 3720 5043 3723
rect 6730 3720 6736 3732
rect 5031 3692 6736 3720
rect 5031 3689 5043 3692
rect 4985 3683 5043 3689
rect 6730 3680 6736 3692
rect 6788 3680 6794 3732
rect 16022 3720 16028 3732
rect 6840 3692 16028 3720
rect 6840 3652 6868 3692
rect 16022 3680 16028 3692
rect 16080 3680 16086 3732
rect 4080 3624 6868 3652
rect 6907 3655 6965 3661
rect 2849 3615 2907 3621
rect 6907 3621 6919 3655
rect 6953 3652 6965 3655
rect 7285 3655 7343 3661
rect 7285 3652 7297 3655
rect 6953 3624 7297 3652
rect 6953 3621 6965 3624
rect 6907 3615 6965 3621
rect 7285 3621 7297 3624
rect 7331 3652 7343 3655
rect 7909 3655 7967 3661
rect 7909 3652 7921 3655
rect 7331 3624 7921 3652
rect 7331 3621 7343 3624
rect 7285 3615 7343 3621
rect 7909 3621 7921 3624
rect 7955 3621 7967 3655
rect 8478 3652 8484 3664
rect 8439 3624 8484 3652
rect 7909 3615 7967 3621
rect 8478 3612 8484 3624
rect 8536 3612 8542 3664
rect 9214 3612 9220 3664
rect 9272 3652 9278 3664
rect 9309 3655 9367 3661
rect 9309 3652 9321 3655
rect 9272 3624 9321 3652
rect 9272 3612 9278 3624
rect 9309 3621 9321 3624
rect 9355 3621 9367 3655
rect 11146 3652 11152 3664
rect 11107 3624 11152 3652
rect 9309 3615 9367 3621
rect 11146 3612 11152 3624
rect 11204 3612 11210 3664
rect 11790 3612 11796 3664
rect 11848 3652 11854 3664
rect 11977 3655 12035 3661
rect 11977 3652 11989 3655
rect 11848 3624 11989 3652
rect 11848 3612 11854 3624
rect 11977 3621 11989 3624
rect 12023 3621 12035 3655
rect 11977 3615 12035 3621
rect 12549 3655 12607 3661
rect 12549 3621 12561 3655
rect 12595 3652 12607 3655
rect 13173 3655 13231 3661
rect 13173 3652 13185 3655
rect 12595 3624 13185 3652
rect 12595 3621 12607 3624
rect 12549 3615 12607 3621
rect 13173 3621 13185 3624
rect 13219 3652 13231 3655
rect 13551 3655 13609 3661
rect 13551 3652 13563 3655
rect 13219 3624 13563 3652
rect 13219 3621 13231 3624
rect 13173 3615 13231 3621
rect 13551 3621 13563 3624
rect 13597 3621 13609 3655
rect 13551 3615 13609 3621
rect 1673 3587 1731 3593
rect 1673 3553 1685 3587
rect 1719 3584 1731 3587
rect 2498 3584 2504 3596
rect 1719 3556 2504 3584
rect 1719 3553 1731 3556
rect 1673 3547 1731 3553
rect 2498 3544 2504 3556
rect 2556 3544 2562 3596
rect 9398 3584 9404 3596
rect 6288 3556 9404 3584
rect 6288 3525 6316 3556
rect 9398 3544 9404 3556
rect 9456 3544 9462 3596
rect 13446 3584 13452 3596
rect 9692 3556 13452 3584
rect 1766 3519 1824 3525
rect 1766 3485 1778 3519
rect 1812 3516 1824 3519
rect 2133 3519 2191 3525
rect 2133 3516 2145 3519
rect 1812 3488 2145 3516
rect 1812 3485 1824 3488
rect 1766 3479 1824 3485
rect 2133 3485 2145 3488
rect 2179 3516 2191 3519
rect 2849 3519 2907 3525
rect 2849 3516 2861 3519
rect 2179 3488 2861 3516
rect 2179 3485 2191 3488
rect 2133 3479 2191 3485
rect 2849 3485 2861 3488
rect 2895 3485 2907 3519
rect 2849 3479 2907 3485
rect 3065 3514 3123 3520
rect 3065 3480 3077 3514
rect 3111 3480 3123 3514
rect 3065 3457 3123 3480
rect 6273 3519 6331 3525
rect 6273 3485 6285 3519
rect 6319 3485 6331 3519
rect 6730 3516 6736 3528
rect 6691 3488 6736 3516
rect 6273 3479 6331 3485
rect 6730 3476 6736 3488
rect 6788 3476 6794 3528
rect 6826 3519 6884 3525
rect 6826 3485 6838 3519
rect 6872 3516 6884 3519
rect 7193 3519 7251 3525
rect 7193 3516 7205 3519
rect 6872 3488 7205 3516
rect 6872 3485 6884 3488
rect 6826 3479 6884 3485
rect 7193 3485 7205 3488
rect 7239 3516 7251 3519
rect 7909 3519 7967 3525
rect 7909 3516 7921 3519
rect 7239 3488 7921 3516
rect 7239 3485 7251 3488
rect 7193 3479 7251 3485
rect 7909 3485 7921 3488
rect 7955 3485 7967 3519
rect 7909 3479 7967 3485
rect 8125 3516 8183 3520
rect 8294 3516 8300 3528
rect 8125 3514 8300 3516
rect 8125 3480 8137 3514
rect 8171 3488 8300 3514
rect 8171 3480 8183 3488
rect 2405 3451 2535 3457
rect 2405 3417 2417 3451
rect 2451 3417 2489 3451
rect 2523 3448 2535 3451
rect 3065 3451 3183 3457
rect 3065 3448 3137 3451
rect 2523 3420 3137 3448
rect 2523 3417 2535 3420
rect 2405 3411 2535 3417
rect 3125 3417 3137 3420
rect 3171 3448 3183 3451
rect 4430 3448 4436 3460
rect 3171 3420 4436 3448
rect 3171 3417 3183 3420
rect 3125 3411 3183 3417
rect 2958 3340 2964 3392
rect 3016 3380 3022 3392
rect 3252 3380 3280 3420
rect 4430 3408 4436 3420
rect 4488 3408 4494 3460
rect 8125 3457 8183 3480
rect 8294 3476 8300 3488
rect 8352 3476 8358 3528
rect 9122 3516 9128 3528
rect 9083 3488 9128 3516
rect 9122 3476 9128 3488
rect 9180 3476 9186 3528
rect 7009 3451 7067 3457
rect 7009 3417 7021 3451
rect 7055 3417 7067 3451
rect 7009 3411 7067 3417
rect 7465 3451 7595 3457
rect 7465 3417 7477 3451
rect 7511 3417 7549 3451
rect 7583 3448 7595 3451
rect 8125 3451 8243 3457
rect 8125 3448 8197 3451
rect 7583 3420 8197 3448
rect 7583 3417 7595 3420
rect 7465 3411 7595 3417
rect 8185 3417 8197 3420
rect 8231 3417 8243 3451
rect 9692 3448 9720 3556
rect 13446 3544 13452 3556
rect 13504 3544 13510 3596
rect 13722 3584 13728 3596
rect 13683 3556 13728 3584
rect 13722 3544 13728 3556
rect 13780 3544 13786 3596
rect 10226 3516 10232 3528
rect 10187 3488 10232 3516
rect 10226 3476 10232 3488
rect 10284 3476 10290 3528
rect 10962 3516 10968 3528
rect 10923 3488 10968 3516
rect 10962 3476 10968 3488
rect 11020 3476 11026 3528
rect 12333 3514 12391 3520
rect 12333 3480 12345 3514
rect 12379 3480 12391 3514
rect 8185 3411 8243 3417
rect 8404 3420 9720 3448
rect 3016 3352 3280 3380
rect 3421 3383 3479 3389
rect 3016 3340 3022 3352
rect 3421 3349 3433 3383
rect 3467 3380 3479 3383
rect 6914 3380 6920 3392
rect 3467 3352 6920 3380
rect 3467 3349 3479 3352
rect 3421 3343 3479 3349
rect 6914 3340 6920 3352
rect 6972 3340 6978 3392
rect 7024 3380 7052 3411
rect 8404 3380 8432 3420
rect 11698 3408 11704 3460
rect 11756 3448 11762 3460
rect 12333 3457 12391 3480
rect 12549 3519 12607 3525
rect 12549 3485 12561 3519
rect 12595 3516 12607 3519
rect 13265 3519 13323 3525
rect 13265 3516 13277 3519
rect 12595 3488 13277 3516
rect 12595 3485 12607 3488
rect 12549 3479 12607 3485
rect 13265 3485 13277 3488
rect 13311 3516 13323 3519
rect 13632 3519 13690 3525
rect 13632 3516 13644 3519
rect 13311 3488 13644 3516
rect 13311 3485 13323 3488
rect 13265 3479 13323 3485
rect 13632 3485 13644 3488
rect 13678 3485 13690 3519
rect 13632 3479 13690 3485
rect 12273 3451 12391 3457
rect 11756 3420 12112 3448
rect 11756 3408 11762 3420
rect 7024 3352 8432 3380
rect 8662 3340 8668 3392
rect 8720 3380 8726 3392
rect 10045 3383 10103 3389
rect 10045 3380 10057 3383
rect 8720 3352 10057 3380
rect 8720 3340 8726 3352
rect 10045 3349 10057 3352
rect 10091 3349 10103 3383
rect 12084 3380 12112 3420
rect 12273 3417 12285 3451
rect 12319 3448 12391 3451
rect 12710 3448 12716 3460
rect 12319 3420 12716 3448
rect 12319 3417 12331 3420
rect 12273 3411 12331 3417
rect 12710 3408 12716 3420
rect 12768 3448 12774 3460
rect 12921 3451 13051 3457
rect 12921 3448 12933 3451
rect 12768 3420 12933 3448
rect 12768 3408 12774 3420
rect 12921 3417 12933 3420
rect 12967 3417 13005 3451
rect 13039 3417 13051 3451
rect 12921 3411 13051 3417
rect 13449 3451 13507 3457
rect 13449 3417 13461 3451
rect 13495 3417 13507 3451
rect 13449 3411 13507 3417
rect 13464 3380 13492 3411
rect 12084 3352 13492 3380
rect 10045 3343 10103 3349
rect 1104 3290 19019 3312
rect 1104 3281 5388 3290
rect 1104 3247 1133 3281
rect 1167 3247 1225 3281
rect 1259 3247 1317 3281
rect 1351 3247 1409 3281
rect 1443 3247 1501 3281
rect 1535 3247 1593 3281
rect 1627 3247 1685 3281
rect 1719 3247 1777 3281
rect 1811 3247 1869 3281
rect 1903 3247 1961 3281
rect 1995 3247 2053 3281
rect 2087 3247 2145 3281
rect 2179 3247 2237 3281
rect 2271 3247 2329 3281
rect 2363 3247 2421 3281
rect 2455 3247 2513 3281
rect 2547 3247 2605 3281
rect 2639 3247 2697 3281
rect 2731 3247 2789 3281
rect 2823 3247 2881 3281
rect 2915 3247 2973 3281
rect 3007 3247 3065 3281
rect 3099 3247 3157 3281
rect 3191 3247 3249 3281
rect 3283 3247 3341 3281
rect 3375 3247 3433 3281
rect 3467 3247 3525 3281
rect 3559 3247 3617 3281
rect 3651 3247 3709 3281
rect 3743 3247 3801 3281
rect 3835 3247 3893 3281
rect 3927 3247 3985 3281
rect 4019 3247 4077 3281
rect 4111 3247 4169 3281
rect 4203 3247 4261 3281
rect 4295 3247 4353 3281
rect 4387 3247 4445 3281
rect 4479 3247 4537 3281
rect 4571 3247 4629 3281
rect 4663 3247 4721 3281
rect 4755 3247 4813 3281
rect 4847 3247 4905 3281
rect 4939 3247 4997 3281
rect 5031 3247 5089 3281
rect 5123 3247 5181 3281
rect 5215 3247 5273 3281
rect 5307 3247 5365 3281
rect 1104 3238 5388 3247
rect 5440 3238 5452 3290
rect 5504 3238 5516 3290
rect 5568 3281 5580 3290
rect 5632 3281 5644 3290
rect 5696 3281 9827 3290
rect 9879 3281 9891 3290
rect 5632 3247 5641 3281
rect 5696 3247 5733 3281
rect 5767 3247 5825 3281
rect 5859 3247 5917 3281
rect 5951 3247 6009 3281
rect 6043 3247 6101 3281
rect 6135 3247 6193 3281
rect 6227 3247 6285 3281
rect 6319 3247 6377 3281
rect 6411 3247 6469 3281
rect 6503 3247 6561 3281
rect 6595 3247 6653 3281
rect 6687 3247 6745 3281
rect 6779 3247 6837 3281
rect 6871 3247 6929 3281
rect 6963 3247 7021 3281
rect 7055 3247 7113 3281
rect 7147 3247 7205 3281
rect 7239 3247 7297 3281
rect 7331 3247 7389 3281
rect 7423 3247 7481 3281
rect 7515 3247 7573 3281
rect 7607 3247 7665 3281
rect 7699 3247 7757 3281
rect 7791 3247 7849 3281
rect 7883 3247 7941 3281
rect 7975 3247 8033 3281
rect 8067 3247 8125 3281
rect 8159 3247 8217 3281
rect 8251 3247 8309 3281
rect 8343 3247 8401 3281
rect 8435 3247 8493 3281
rect 8527 3247 8585 3281
rect 8619 3247 8677 3281
rect 8711 3247 8769 3281
rect 8803 3247 8861 3281
rect 8895 3247 8953 3281
rect 8987 3247 9045 3281
rect 9079 3247 9137 3281
rect 9171 3247 9229 3281
rect 9263 3247 9321 3281
rect 9355 3247 9413 3281
rect 9447 3247 9505 3281
rect 9539 3247 9597 3281
rect 9631 3247 9689 3281
rect 9723 3247 9781 3281
rect 9815 3247 9827 3281
rect 5568 3238 5580 3247
rect 5632 3238 5644 3247
rect 5696 3238 9827 3247
rect 9879 3238 9891 3247
rect 9943 3238 9955 3290
rect 10007 3238 10019 3290
rect 10071 3281 10083 3290
rect 10135 3281 14266 3290
rect 14318 3281 14330 3290
rect 14382 3281 14394 3290
rect 10135 3247 10149 3281
rect 10183 3247 10241 3281
rect 10275 3247 10333 3281
rect 10367 3247 10425 3281
rect 10459 3247 10517 3281
rect 10551 3247 10609 3281
rect 10643 3247 10701 3281
rect 10735 3247 10793 3281
rect 10827 3247 10885 3281
rect 10919 3247 10977 3281
rect 11011 3247 11069 3281
rect 11103 3247 11161 3281
rect 11195 3247 11253 3281
rect 11287 3247 11345 3281
rect 11379 3247 11437 3281
rect 11471 3247 11529 3281
rect 11563 3247 11621 3281
rect 11655 3247 11713 3281
rect 11747 3247 11805 3281
rect 11839 3247 11897 3281
rect 11931 3247 11989 3281
rect 12023 3247 12081 3281
rect 12115 3247 12173 3281
rect 12207 3247 12265 3281
rect 12299 3247 12357 3281
rect 12391 3247 12449 3281
rect 12483 3247 12541 3281
rect 12575 3247 12633 3281
rect 12667 3247 12725 3281
rect 12759 3247 12817 3281
rect 12851 3247 12909 3281
rect 12943 3247 13001 3281
rect 13035 3247 13093 3281
rect 13127 3247 13185 3281
rect 13219 3247 13277 3281
rect 13311 3247 13369 3281
rect 13403 3247 13461 3281
rect 13495 3247 13553 3281
rect 13587 3247 13645 3281
rect 13679 3247 13737 3281
rect 13771 3247 13829 3281
rect 13863 3247 13921 3281
rect 13955 3247 14013 3281
rect 14047 3247 14105 3281
rect 14139 3247 14197 3281
rect 14231 3247 14266 3281
rect 14323 3247 14330 3281
rect 10071 3238 10083 3247
rect 10135 3238 14266 3247
rect 14318 3238 14330 3247
rect 14382 3238 14394 3247
rect 14446 3238 14458 3290
rect 14510 3238 14522 3290
rect 14574 3281 18705 3290
rect 14599 3247 14657 3281
rect 14691 3247 14749 3281
rect 14783 3247 14841 3281
rect 14875 3247 14933 3281
rect 14967 3247 15025 3281
rect 15059 3247 15117 3281
rect 15151 3247 15209 3281
rect 15243 3247 15301 3281
rect 15335 3247 15393 3281
rect 15427 3247 15485 3281
rect 15519 3247 15577 3281
rect 15611 3247 15669 3281
rect 15703 3247 15761 3281
rect 15795 3247 15853 3281
rect 15887 3247 15945 3281
rect 15979 3247 16037 3281
rect 16071 3247 16129 3281
rect 16163 3247 16221 3281
rect 16255 3247 16313 3281
rect 16347 3247 16405 3281
rect 16439 3247 16497 3281
rect 16531 3247 16589 3281
rect 16623 3247 16681 3281
rect 16715 3247 16773 3281
rect 16807 3247 16865 3281
rect 16899 3247 16957 3281
rect 16991 3247 17049 3281
rect 17083 3247 17141 3281
rect 17175 3247 17233 3281
rect 17267 3247 17325 3281
rect 17359 3247 17417 3281
rect 17451 3247 17509 3281
rect 17543 3247 17601 3281
rect 17635 3247 17693 3281
rect 17727 3247 17785 3281
rect 17819 3247 17877 3281
rect 17911 3247 17969 3281
rect 18003 3247 18061 3281
rect 18095 3247 18153 3281
rect 18187 3247 18245 3281
rect 18279 3247 18337 3281
rect 18371 3247 18429 3281
rect 18463 3247 18521 3281
rect 18555 3247 18613 3281
rect 18647 3247 18705 3281
rect 14574 3238 18705 3247
rect 18757 3238 18769 3290
rect 18821 3281 18833 3290
rect 18831 3247 18833 3281
rect 18821 3238 18833 3247
rect 18885 3238 18897 3290
rect 18949 3238 18961 3290
rect 19013 3238 19019 3290
rect 1104 3216 19019 3238
rect 1946 3176 1952 3188
rect 1859 3148 1952 3176
rect 1946 3136 1952 3148
rect 2004 3176 2010 3188
rect 7098 3176 7104 3188
rect 2004 3148 7104 3176
rect 2004 3136 2010 3148
rect 7098 3136 7104 3148
rect 7156 3136 7162 3188
rect 7193 3179 7251 3185
rect 7193 3145 7205 3179
rect 7239 3176 7251 3179
rect 7926 3176 7932 3188
rect 7239 3148 7932 3176
rect 7239 3145 7251 3148
rect 7193 3139 7251 3145
rect 7926 3136 7932 3148
rect 7984 3136 7990 3188
rect 9214 3176 9220 3188
rect 8588 3148 9220 3176
rect 2958 3117 2964 3120
rect 2245 3111 2303 3117
rect 2245 3077 2257 3111
rect 2291 3108 2303 3111
rect 2893 3111 2964 3117
rect 3016 3117 3022 3120
rect 2893 3108 2905 3111
rect 2291 3080 2905 3108
rect 2291 3077 2363 3080
rect 2245 3071 2363 3077
rect 2893 3077 2905 3080
rect 2939 3077 2964 3111
rect 2893 3071 2964 3077
rect 2305 3048 2363 3071
rect 2958 3068 2964 3071
rect 3016 3071 3023 3117
rect 3421 3111 3479 3117
rect 3421 3077 3433 3111
rect 3467 3108 3479 3111
rect 4246 3108 4252 3120
rect 3467 3080 4252 3108
rect 3467 3077 3479 3080
rect 3421 3071 3479 3077
rect 3016 3068 3022 3071
rect 4246 3068 4252 3080
rect 4304 3068 4310 3120
rect 4342 3111 4400 3117
rect 4342 3077 4354 3111
rect 4388 3108 4400 3111
rect 4714 3111 4772 3117
rect 4714 3108 4726 3111
rect 4388 3080 4726 3108
rect 4388 3077 4400 3080
rect 4342 3071 4400 3077
rect 4714 3077 4726 3080
rect 4760 3077 4772 3111
rect 4714 3071 4772 3077
rect 4898 3111 4956 3117
rect 4898 3077 4910 3111
rect 4944 3108 4956 3111
rect 5550 3111 5608 3117
rect 5550 3108 5562 3111
rect 4944 3080 5562 3108
rect 4944 3077 4956 3080
rect 4898 3071 4956 3077
rect 5550 3077 5562 3080
rect 5596 3108 5608 3111
rect 7374 3108 7380 3120
rect 5596 3080 7380 3108
rect 5596 3077 5608 3080
rect 5550 3071 5608 3077
rect 2305 3014 2317 3048
rect 2351 3014 2363 3048
rect 2305 3008 2363 3014
rect 2521 3043 2579 3049
rect 2521 3009 2533 3043
rect 2567 3040 2579 3043
rect 3237 3043 3295 3049
rect 3237 3040 3249 3043
rect 2567 3012 3249 3040
rect 2567 3009 2579 3012
rect 2521 3003 2579 3009
rect 3237 3009 3249 3012
rect 3283 3040 3295 3043
rect 3604 3043 3662 3049
rect 3604 3040 3616 3043
rect 3283 3012 3616 3040
rect 3283 3009 3295 3012
rect 3237 3003 3295 3009
rect 3604 3009 3616 3012
rect 3650 3009 3662 3043
rect 3604 3003 3662 3009
rect 3697 3043 3755 3049
rect 3697 3009 3709 3043
rect 3743 3040 3755 3043
rect 4154 3040 4160 3052
rect 3743 3012 4160 3040
rect 3743 3009 3755 3012
rect 3697 3003 3755 3009
rect 4154 3000 4160 3012
rect 4212 3000 4218 3052
rect 4522 3040 4528 3052
rect 4483 3012 4528 3040
rect 4522 3000 4528 3012
rect 4580 3000 4586 3052
rect 4729 3040 4772 3071
rect 5178 3043 5236 3049
rect 5178 3040 5190 3043
rect 4729 3012 5190 3040
rect 5178 3009 5190 3012
rect 5224 3009 5236 3043
rect 5178 3003 5236 3009
rect 5258 2932 5264 2984
rect 5316 2972 5322 2984
rect 5552 2972 5580 3071
rect 7374 3068 7380 3080
rect 7432 3068 7438 3120
rect 7489 3111 7547 3117
rect 7489 3077 7501 3111
rect 7535 3108 7547 3111
rect 8137 3111 8267 3117
rect 8137 3108 8149 3111
rect 7535 3080 8149 3108
rect 7535 3077 7607 3080
rect 7489 3071 7607 3077
rect 8137 3077 8149 3080
rect 8183 3077 8221 3111
rect 8255 3108 8267 3111
rect 8588 3108 8616 3148
rect 9214 3136 9220 3148
rect 9272 3136 9278 3188
rect 10870 3136 10876 3188
rect 10928 3176 10934 3188
rect 13722 3176 13728 3188
rect 10928 3148 13728 3176
rect 10928 3136 10934 3148
rect 13722 3136 13728 3148
rect 13780 3136 13786 3188
rect 8255 3080 8616 3108
rect 8255 3077 8267 3080
rect 8137 3071 8267 3077
rect 7549 3048 7607 3071
rect 8662 3068 8668 3120
rect 8720 3117 8726 3120
rect 8720 3111 8735 3117
rect 8723 3077 8735 3111
rect 9398 3108 9404 3120
rect 9359 3080 9404 3108
rect 8720 3071 8735 3077
rect 8720 3068 8726 3071
rect 9398 3068 9404 3080
rect 9456 3068 9462 3120
rect 12710 3117 12716 3120
rect 11997 3111 12055 3117
rect 11997 3077 12009 3111
rect 12043 3108 12055 3111
rect 12645 3111 12716 3117
rect 12768 3117 12774 3120
rect 12645 3108 12657 3111
rect 12043 3080 12657 3108
rect 12043 3077 12115 3080
rect 11997 3071 12115 3077
rect 12645 3077 12657 3080
rect 12691 3077 12716 3111
rect 12645 3071 12716 3077
rect 7549 3014 7561 3048
rect 7595 3014 7607 3048
rect 7549 3008 7607 3014
rect 7765 3043 7823 3049
rect 7765 3009 7777 3043
rect 7811 3040 7823 3043
rect 8481 3043 8539 3049
rect 8481 3040 8493 3043
rect 7811 3012 8493 3040
rect 7811 3009 7823 3012
rect 7765 3003 7823 3009
rect 8481 3009 8493 3012
rect 8527 3040 8539 3043
rect 8848 3043 8906 3049
rect 8848 3040 8860 3043
rect 8527 3012 8860 3040
rect 8527 3009 8539 3012
rect 8481 3003 8539 3009
rect 8848 3009 8860 3012
rect 8894 3009 8906 3043
rect 8848 3003 8906 3009
rect 9030 3000 9036 3052
rect 9088 3040 9094 3052
rect 10686 3040 10692 3052
rect 9088 3012 10692 3040
rect 9088 3000 9094 3012
rect 10686 3000 10692 3012
rect 10744 3000 10750 3052
rect 12057 3048 12115 3071
rect 12710 3068 12716 3071
rect 12768 3071 12775 3117
rect 12768 3068 12774 3071
rect 12894 3068 12900 3120
rect 12952 3108 12958 3120
rect 13173 3111 13231 3117
rect 13173 3108 13185 3111
rect 12952 3080 13185 3108
rect 12952 3068 12958 3080
rect 13173 3077 13185 3080
rect 13219 3077 13231 3111
rect 13173 3071 13231 3077
rect 13446 3068 13452 3120
rect 13504 3108 13510 3120
rect 13504 3080 16574 3108
rect 13504 3068 13510 3080
rect 12057 3014 12069 3048
rect 12103 3014 12115 3048
rect 12057 3008 12115 3014
rect 12273 3043 12331 3049
rect 12273 3009 12285 3043
rect 12319 3040 12331 3043
rect 12989 3043 13047 3049
rect 12989 3040 13001 3043
rect 12319 3012 13001 3040
rect 12319 3009 12331 3012
rect 12273 3003 12331 3009
rect 12989 3009 13001 3012
rect 13035 3040 13047 3043
rect 13356 3043 13414 3049
rect 13356 3040 13368 3043
rect 13035 3012 13368 3040
rect 13035 3009 13047 3012
rect 12989 3003 13047 3009
rect 13356 3009 13368 3012
rect 13402 3009 13414 3043
rect 13906 3040 13912 3052
rect 13867 3012 13912 3040
rect 13356 3003 13414 3009
rect 13906 3000 13912 3012
rect 13964 3000 13970 3052
rect 5316 2944 5580 2972
rect 5951 2975 6009 2981
rect 5316 2932 5322 2944
rect 5951 2941 5963 2975
rect 5997 2972 6009 2975
rect 8941 2975 8999 2981
rect 5997 2944 8892 2972
rect 5997 2941 6009 2944
rect 5951 2935 6009 2941
rect 2521 2907 2579 2913
rect 2521 2873 2533 2907
rect 2567 2904 2579 2907
rect 3145 2907 3203 2913
rect 3145 2904 3157 2907
rect 2567 2876 3157 2904
rect 2567 2873 2579 2876
rect 2521 2867 2579 2873
rect 3145 2873 3157 2876
rect 3191 2904 3203 2907
rect 3523 2907 3581 2913
rect 3523 2904 3535 2907
rect 3191 2876 3535 2904
rect 3191 2873 3203 2876
rect 3145 2867 3203 2873
rect 3523 2873 3535 2876
rect 3569 2873 3581 2907
rect 3523 2867 3581 2873
rect 4250 2907 4308 2913
rect 4250 2873 4262 2907
rect 4296 2904 4308 2907
rect 4622 2907 4680 2913
rect 4622 2904 4634 2907
rect 4296 2876 4634 2904
rect 4296 2873 4308 2876
rect 4250 2867 4308 2873
rect 4622 2873 4634 2876
rect 4668 2904 4680 2907
rect 5178 2907 5236 2913
rect 5178 2904 5190 2907
rect 4668 2876 5190 2904
rect 4668 2873 4680 2876
rect 4622 2867 4680 2873
rect 5178 2873 5190 2876
rect 5224 2873 5236 2907
rect 5178 2867 5236 2873
rect 7765 2907 7823 2913
rect 7765 2873 7777 2907
rect 7811 2904 7823 2907
rect 8389 2907 8447 2913
rect 8389 2904 8401 2907
rect 7811 2876 8401 2904
rect 7811 2873 7823 2876
rect 7765 2867 7823 2873
rect 8389 2873 8401 2876
rect 8435 2904 8447 2907
rect 8767 2907 8825 2913
rect 8767 2904 8779 2907
rect 8435 2876 8779 2904
rect 8435 2873 8447 2876
rect 8389 2867 8447 2873
rect 8767 2873 8779 2876
rect 8813 2873 8825 2907
rect 8864 2904 8892 2944
rect 8941 2941 8953 2975
rect 8987 2972 8999 2975
rect 13449 2975 13507 2981
rect 8987 2944 10732 2972
rect 8987 2941 8999 2944
rect 8941 2935 8999 2941
rect 10704 2913 10732 2944
rect 10980 2944 13400 2972
rect 10689 2907 10747 2913
rect 8864 2876 10640 2904
rect 8767 2867 8825 2873
rect 7466 2796 7472 2848
rect 7524 2836 7530 2848
rect 9582 2836 9588 2848
rect 7524 2808 9588 2836
rect 7524 2796 7530 2808
rect 9582 2796 9588 2808
rect 9640 2796 9646 2848
rect 10612 2836 10640 2876
rect 10689 2873 10701 2907
rect 10735 2904 10747 2907
rect 10870 2904 10876 2916
rect 10735 2876 10876 2904
rect 10735 2873 10747 2876
rect 10689 2867 10747 2873
rect 10870 2864 10876 2876
rect 10928 2864 10934 2916
rect 10980 2836 11008 2944
rect 11698 2904 11704 2916
rect 11659 2876 11704 2904
rect 11698 2864 11704 2876
rect 11756 2864 11762 2916
rect 12273 2907 12331 2913
rect 12273 2873 12285 2907
rect 12319 2904 12331 2907
rect 12897 2907 12955 2913
rect 12897 2904 12909 2907
rect 12319 2876 12909 2904
rect 12319 2873 12331 2876
rect 12273 2867 12331 2873
rect 12897 2873 12909 2876
rect 12943 2904 12955 2907
rect 13275 2907 13333 2913
rect 13275 2904 13287 2907
rect 12943 2876 13287 2904
rect 12943 2873 12955 2876
rect 12897 2867 12955 2873
rect 13275 2873 13287 2876
rect 13321 2873 13333 2907
rect 13372 2904 13400 2944
rect 13449 2941 13461 2975
rect 13495 2972 13507 2975
rect 13722 2972 13728 2984
rect 13495 2944 13728 2972
rect 13495 2941 13507 2944
rect 13449 2935 13507 2941
rect 13722 2932 13728 2944
rect 13780 2932 13786 2984
rect 15378 2904 15384 2916
rect 13372 2876 15384 2904
rect 13275 2867 13333 2873
rect 15378 2864 15384 2876
rect 15436 2904 15442 2916
rect 15746 2904 15752 2916
rect 15436 2876 15752 2904
rect 15436 2864 15442 2876
rect 15746 2864 15752 2876
rect 15804 2864 15810 2916
rect 16546 2904 16574 3080
rect 16850 2904 16856 2916
rect 16546 2876 16856 2904
rect 16850 2864 16856 2876
rect 16908 2864 16914 2916
rect 10612 2808 11008 2836
rect 12434 2796 12440 2848
rect 12492 2836 12498 2848
rect 14093 2839 14151 2845
rect 14093 2836 14105 2839
rect 12492 2808 14105 2836
rect 12492 2796 12498 2808
rect 14093 2805 14105 2808
rect 14139 2805 14151 2839
rect 14093 2799 14151 2805
rect 1104 2746 18860 2768
rect 1104 2737 3169 2746
rect 1104 2703 1133 2737
rect 1167 2703 1225 2737
rect 1259 2703 1317 2737
rect 1351 2703 1409 2737
rect 1443 2703 1501 2737
rect 1535 2703 1593 2737
rect 1627 2703 1685 2737
rect 1719 2703 1777 2737
rect 1811 2703 1869 2737
rect 1903 2703 1961 2737
rect 1995 2703 2053 2737
rect 2087 2703 2145 2737
rect 2179 2703 2237 2737
rect 2271 2703 2329 2737
rect 2363 2703 2421 2737
rect 2455 2703 2513 2737
rect 2547 2703 2605 2737
rect 2639 2703 2697 2737
rect 2731 2703 2789 2737
rect 2823 2703 2881 2737
rect 2915 2703 2973 2737
rect 3007 2703 3065 2737
rect 3099 2703 3157 2737
rect 1104 2694 3169 2703
rect 3221 2694 3233 2746
rect 3285 2694 3297 2746
rect 3349 2737 3361 2746
rect 3349 2694 3361 2703
rect 3413 2694 3425 2746
rect 3477 2737 7608 2746
rect 3477 2703 3525 2737
rect 3559 2703 3617 2737
rect 3651 2703 3709 2737
rect 3743 2703 3801 2737
rect 3835 2703 3893 2737
rect 3927 2703 3985 2737
rect 4019 2703 4077 2737
rect 4111 2703 4169 2737
rect 4203 2703 4261 2737
rect 4295 2703 4353 2737
rect 4387 2703 4445 2737
rect 4479 2703 4537 2737
rect 4571 2703 4629 2737
rect 4663 2703 4721 2737
rect 4755 2703 4813 2737
rect 4847 2703 4905 2737
rect 4939 2703 4997 2737
rect 5031 2703 5089 2737
rect 5123 2703 5181 2737
rect 5215 2703 5273 2737
rect 5307 2703 5365 2737
rect 5399 2703 5457 2737
rect 5491 2703 5549 2737
rect 5583 2703 5641 2737
rect 5675 2703 5733 2737
rect 5767 2703 5825 2737
rect 5859 2703 5917 2737
rect 5951 2703 6009 2737
rect 6043 2703 6101 2737
rect 6135 2703 6193 2737
rect 6227 2703 6285 2737
rect 6319 2703 6377 2737
rect 6411 2703 6469 2737
rect 6503 2703 6561 2737
rect 6595 2703 6653 2737
rect 6687 2703 6745 2737
rect 6779 2703 6837 2737
rect 6871 2703 6929 2737
rect 6963 2703 7021 2737
rect 7055 2703 7113 2737
rect 7147 2703 7205 2737
rect 7239 2703 7297 2737
rect 7331 2703 7389 2737
rect 7423 2703 7481 2737
rect 7515 2703 7573 2737
rect 7607 2703 7608 2737
rect 3477 2694 7608 2703
rect 7660 2737 7672 2746
rect 7660 2703 7665 2737
rect 7660 2694 7672 2703
rect 7724 2694 7736 2746
rect 7788 2737 7800 2746
rect 7852 2737 7864 2746
rect 7916 2737 12047 2746
rect 12099 2737 12111 2746
rect 12163 2737 12175 2746
rect 7791 2703 7800 2737
rect 7916 2703 7941 2737
rect 7975 2703 8033 2737
rect 8067 2703 8125 2737
rect 8159 2703 8217 2737
rect 8251 2703 8309 2737
rect 8343 2703 8401 2737
rect 8435 2703 8493 2737
rect 8527 2703 8585 2737
rect 8619 2703 8677 2737
rect 8711 2703 8769 2737
rect 8803 2703 8861 2737
rect 8895 2703 8953 2737
rect 8987 2703 9045 2737
rect 9079 2703 9137 2737
rect 9171 2703 9229 2737
rect 9263 2703 9321 2737
rect 9355 2703 9413 2737
rect 9447 2703 9505 2737
rect 9539 2703 9597 2737
rect 9631 2703 9689 2737
rect 9723 2703 9781 2737
rect 9815 2703 9873 2737
rect 9907 2703 9965 2737
rect 9999 2703 10057 2737
rect 10091 2703 10149 2737
rect 10183 2703 10241 2737
rect 10275 2703 10333 2737
rect 10367 2703 10425 2737
rect 10459 2703 10517 2737
rect 10551 2703 10609 2737
rect 10643 2703 10701 2737
rect 10735 2703 10793 2737
rect 10827 2703 10885 2737
rect 10919 2703 10977 2737
rect 11011 2703 11069 2737
rect 11103 2703 11161 2737
rect 11195 2703 11253 2737
rect 11287 2703 11345 2737
rect 11379 2703 11437 2737
rect 11471 2703 11529 2737
rect 11563 2703 11621 2737
rect 11655 2703 11713 2737
rect 11747 2703 11805 2737
rect 11839 2703 11897 2737
rect 11931 2703 11989 2737
rect 12023 2703 12047 2737
rect 12163 2703 12173 2737
rect 7788 2694 7800 2703
rect 7852 2694 7864 2703
rect 7916 2694 12047 2703
rect 12099 2694 12111 2703
rect 12163 2694 12175 2703
rect 12227 2694 12239 2746
rect 12291 2737 12303 2746
rect 12299 2703 12303 2737
rect 12291 2694 12303 2703
rect 12355 2737 16486 2746
rect 12355 2703 12357 2737
rect 12391 2703 12449 2737
rect 12483 2703 12541 2737
rect 12575 2703 12633 2737
rect 12667 2703 12725 2737
rect 12759 2703 12817 2737
rect 12851 2703 12909 2737
rect 12943 2703 13001 2737
rect 13035 2703 13093 2737
rect 13127 2703 13185 2737
rect 13219 2703 13277 2737
rect 13311 2703 13369 2737
rect 13403 2703 13461 2737
rect 13495 2703 13553 2737
rect 13587 2703 13645 2737
rect 13679 2703 13737 2737
rect 13771 2703 13829 2737
rect 13863 2703 13921 2737
rect 13955 2703 14013 2737
rect 14047 2703 14105 2737
rect 14139 2703 14197 2737
rect 14231 2703 14289 2737
rect 14323 2703 14381 2737
rect 14415 2703 14473 2737
rect 14507 2703 14565 2737
rect 14599 2703 14657 2737
rect 14691 2703 14749 2737
rect 14783 2703 14841 2737
rect 14875 2703 14933 2737
rect 14967 2703 15025 2737
rect 15059 2703 15117 2737
rect 15151 2703 15209 2737
rect 15243 2703 15301 2737
rect 15335 2703 15393 2737
rect 15427 2703 15485 2737
rect 15519 2703 15577 2737
rect 15611 2703 15669 2737
rect 15703 2703 15761 2737
rect 15795 2703 15853 2737
rect 15887 2703 15945 2737
rect 15979 2703 16037 2737
rect 16071 2703 16129 2737
rect 16163 2703 16221 2737
rect 16255 2703 16313 2737
rect 16347 2703 16405 2737
rect 16439 2703 16486 2737
rect 12355 2694 16486 2703
rect 16538 2694 16550 2746
rect 16602 2737 16614 2746
rect 16602 2694 16614 2703
rect 16666 2694 16678 2746
rect 16730 2694 16742 2746
rect 16794 2737 18860 2746
rect 16807 2703 16865 2737
rect 16899 2703 16957 2737
rect 16991 2703 17049 2737
rect 17083 2703 17141 2737
rect 17175 2703 17233 2737
rect 17267 2703 17325 2737
rect 17359 2703 17417 2737
rect 17451 2703 17509 2737
rect 17543 2703 17601 2737
rect 17635 2703 17693 2737
rect 17727 2703 17785 2737
rect 17819 2703 17877 2737
rect 17911 2703 17969 2737
rect 18003 2703 18061 2737
rect 18095 2703 18153 2737
rect 18187 2703 18245 2737
rect 18279 2703 18337 2737
rect 18371 2703 18429 2737
rect 18463 2703 18521 2737
rect 18555 2703 18613 2737
rect 18647 2703 18705 2737
rect 18739 2703 18797 2737
rect 18831 2703 18860 2737
rect 16794 2694 18860 2703
rect 1104 2672 18860 2694
rect 3421 2635 3479 2641
rect 3421 2601 3433 2635
rect 3467 2632 3479 2635
rect 5997 2635 6055 2641
rect 3467 2604 5948 2632
rect 3467 2601 3479 2604
rect 3421 2595 3479 2601
rect 1847 2567 1905 2573
rect 1847 2533 1859 2567
rect 1893 2564 1905 2567
rect 2225 2567 2283 2573
rect 2225 2564 2237 2567
rect 1893 2536 2237 2564
rect 1893 2533 1905 2536
rect 1847 2527 1905 2533
rect 2225 2533 2237 2536
rect 2271 2564 2283 2567
rect 2849 2567 2907 2573
rect 2849 2564 2861 2567
rect 2271 2536 2861 2564
rect 2271 2533 2283 2536
rect 2225 2527 2283 2533
rect 2849 2533 2861 2536
rect 2895 2533 2907 2567
rect 2849 2527 2907 2533
rect 4423 2567 4481 2573
rect 4423 2533 4435 2567
rect 4469 2564 4481 2567
rect 4801 2567 4859 2573
rect 4801 2564 4813 2567
rect 4469 2536 4813 2564
rect 4469 2533 4481 2536
rect 4423 2527 4481 2533
rect 4801 2533 4813 2536
rect 4847 2564 4859 2567
rect 5425 2567 5483 2573
rect 5425 2564 5437 2567
rect 4847 2536 5437 2564
rect 4847 2533 4859 2536
rect 4801 2527 4859 2533
rect 5425 2533 5437 2536
rect 5471 2533 5483 2567
rect 5920 2564 5948 2604
rect 5997 2601 6009 2635
rect 6043 2632 6055 2635
rect 7006 2632 7012 2644
rect 6043 2604 7012 2632
rect 6043 2601 6055 2604
rect 5997 2595 6055 2601
rect 7006 2592 7012 2604
rect 7064 2592 7070 2644
rect 8202 2592 8208 2644
rect 8260 2632 8266 2644
rect 9125 2635 9183 2641
rect 9125 2632 9137 2635
rect 8260 2604 9137 2632
rect 8260 2592 8266 2604
rect 9125 2601 9137 2604
rect 9171 2601 9183 2635
rect 9125 2595 9183 2601
rect 12894 2592 12900 2644
rect 12952 2632 12958 2644
rect 14277 2635 14335 2641
rect 14277 2632 14289 2635
rect 12952 2604 14289 2632
rect 12952 2592 12958 2604
rect 14277 2601 14289 2604
rect 14323 2601 14335 2635
rect 14277 2595 14335 2601
rect 9582 2564 9588 2576
rect 5920 2536 9588 2564
rect 5425 2527 5483 2533
rect 9582 2524 9588 2536
rect 9640 2524 9646 2576
rect 9697 2567 9755 2573
rect 9697 2533 9709 2567
rect 9743 2564 9755 2567
rect 10321 2567 10379 2573
rect 10321 2564 10333 2567
rect 9743 2536 10333 2564
rect 9743 2533 9755 2536
rect 9697 2527 9755 2533
rect 10321 2533 10333 2536
rect 10367 2564 10379 2567
rect 10699 2567 10757 2573
rect 10699 2564 10711 2567
rect 10367 2536 10711 2564
rect 10367 2533 10379 2536
rect 10321 2527 10379 2533
rect 10699 2533 10711 2536
rect 10745 2533 10757 2567
rect 11977 2567 12035 2573
rect 11977 2564 11989 2567
rect 10699 2527 10757 2533
rect 10796 2536 11989 2564
rect 1673 2499 1731 2505
rect 1673 2465 1685 2499
rect 1719 2496 1731 2499
rect 2498 2496 2504 2508
rect 1719 2468 2504 2496
rect 1719 2465 1731 2468
rect 1673 2459 1731 2465
rect 2498 2456 2504 2468
rect 2556 2456 2562 2508
rect 4154 2456 4160 2508
rect 4212 2496 4218 2508
rect 4249 2499 4307 2505
rect 4249 2496 4261 2499
rect 4212 2468 4261 2496
rect 4212 2456 4218 2468
rect 4249 2465 4261 2468
rect 4295 2465 4307 2499
rect 4249 2459 4307 2465
rect 4525 2499 4583 2505
rect 4525 2465 4537 2499
rect 4571 2496 4583 2499
rect 4614 2496 4620 2508
rect 4571 2468 4620 2496
rect 4571 2465 4583 2468
rect 4525 2459 4583 2465
rect 4614 2456 4620 2468
rect 4672 2456 4678 2508
rect 8018 2456 8024 2508
rect 8076 2496 8082 2508
rect 10597 2499 10655 2505
rect 10597 2496 10609 2499
rect 8076 2468 10609 2496
rect 8076 2456 8082 2468
rect 10597 2465 10609 2468
rect 10643 2496 10655 2499
rect 10796 2496 10824 2536
rect 11977 2533 11989 2536
rect 12023 2533 12035 2567
rect 11977 2527 12035 2533
rect 12549 2567 12607 2573
rect 12549 2533 12561 2567
rect 12595 2564 12607 2567
rect 13173 2567 13231 2573
rect 13173 2564 13185 2567
rect 12595 2536 13185 2564
rect 12595 2533 12607 2536
rect 12549 2527 12607 2533
rect 13173 2533 13185 2536
rect 13219 2564 13231 2567
rect 13551 2567 13609 2573
rect 13551 2564 13563 2567
rect 13219 2536 13563 2564
rect 13219 2533 13231 2536
rect 13173 2527 13231 2533
rect 13551 2533 13563 2536
rect 13597 2533 13609 2567
rect 13551 2527 13609 2533
rect 14849 2567 14907 2573
rect 14849 2533 14861 2567
rect 14895 2564 14907 2567
rect 15473 2567 15531 2573
rect 15473 2564 15485 2567
rect 14895 2536 15485 2564
rect 14895 2533 14907 2536
rect 14849 2527 14907 2533
rect 15473 2533 15485 2536
rect 15519 2564 15531 2567
rect 15851 2567 15909 2573
rect 15851 2564 15863 2567
rect 15519 2536 15863 2564
rect 15519 2533 15531 2536
rect 15473 2527 15531 2533
rect 15851 2533 15863 2536
rect 15897 2533 15909 2567
rect 15851 2527 15909 2533
rect 10643 2468 10824 2496
rect 10643 2465 10655 2468
rect 10597 2459 10655 2465
rect 11698 2456 11704 2508
rect 11756 2496 11762 2508
rect 13449 2499 13507 2505
rect 13449 2496 13461 2499
rect 11756 2468 13461 2496
rect 11756 2456 11762 2468
rect 13449 2465 13461 2468
rect 13495 2465 13507 2499
rect 13722 2496 13728 2508
rect 13635 2468 13728 2496
rect 13449 2459 13507 2465
rect 13722 2456 13728 2468
rect 13780 2496 13786 2508
rect 16025 2499 16083 2505
rect 16025 2496 16037 2499
rect 13780 2468 16037 2496
rect 13780 2456 13786 2468
rect 16025 2465 16037 2468
rect 16071 2465 16083 2499
rect 16025 2459 16083 2465
rect 1766 2431 1824 2437
rect 1766 2397 1778 2431
rect 1812 2428 1824 2431
rect 2133 2431 2191 2437
rect 2133 2428 2145 2431
rect 1812 2400 2145 2428
rect 1812 2397 1824 2400
rect 1766 2391 1824 2397
rect 2133 2397 2145 2400
rect 2179 2428 2191 2431
rect 2849 2431 2907 2437
rect 2849 2428 2861 2431
rect 2179 2400 2861 2428
rect 2179 2397 2191 2400
rect 2133 2391 2191 2397
rect 2849 2397 2861 2400
rect 2895 2397 2907 2431
rect 2849 2391 2907 2397
rect 3065 2426 3123 2432
rect 3065 2392 3077 2426
rect 3111 2392 3123 2426
rect 1946 2360 1952 2372
rect 1907 2332 1952 2360
rect 1946 2320 1952 2332
rect 2004 2320 2010 2372
rect 3065 2369 3123 2392
rect 4342 2431 4400 2437
rect 4342 2397 4354 2431
rect 4388 2428 4400 2431
rect 4709 2431 4767 2437
rect 4709 2428 4721 2431
rect 4388 2400 4721 2428
rect 4388 2397 4400 2400
rect 4342 2391 4400 2397
rect 4709 2397 4721 2400
rect 4755 2428 4767 2431
rect 5425 2431 5483 2437
rect 5425 2428 5437 2431
rect 4755 2400 5437 2428
rect 4755 2397 4767 2400
rect 4709 2391 4767 2397
rect 5425 2397 5437 2400
rect 5471 2397 5483 2431
rect 5425 2391 5483 2397
rect 5641 2426 5699 2432
rect 5641 2392 5653 2426
rect 5687 2392 5699 2426
rect 5641 2369 5699 2392
rect 9481 2426 9539 2432
rect 9481 2392 9493 2426
rect 9527 2392 9539 2426
rect 9481 2369 9539 2392
rect 9697 2431 9755 2437
rect 9697 2397 9709 2431
rect 9743 2428 9755 2431
rect 10413 2431 10471 2437
rect 10413 2428 10425 2431
rect 9743 2400 10425 2428
rect 9743 2397 9755 2400
rect 9697 2391 9755 2397
rect 10413 2397 10425 2400
rect 10459 2428 10471 2431
rect 10780 2431 10838 2437
rect 10780 2428 10792 2431
rect 10459 2400 10792 2428
rect 10459 2397 10471 2400
rect 10413 2391 10471 2397
rect 10780 2397 10792 2400
rect 10826 2397 10838 2431
rect 10780 2391 10838 2397
rect 10870 2388 10876 2440
rect 10928 2428 10934 2440
rect 10928 2400 10973 2428
rect 12333 2426 12391 2432
rect 10928 2388 10934 2400
rect 12333 2392 12345 2426
rect 12379 2392 12391 2426
rect 12333 2369 12391 2392
rect 12549 2431 12607 2437
rect 12549 2397 12561 2431
rect 12595 2428 12607 2431
rect 13265 2431 13323 2437
rect 13265 2428 13277 2431
rect 12595 2400 13277 2428
rect 12595 2397 12607 2400
rect 12549 2391 12607 2397
rect 13265 2397 13277 2400
rect 13311 2428 13323 2431
rect 13632 2431 13690 2437
rect 13632 2428 13644 2431
rect 13311 2400 13644 2428
rect 13311 2397 13323 2400
rect 13265 2391 13323 2397
rect 13632 2397 13644 2400
rect 13678 2397 13690 2431
rect 13632 2391 13690 2397
rect 14633 2426 14691 2432
rect 14633 2392 14645 2426
rect 14679 2392 14691 2426
rect 14633 2369 14691 2392
rect 14849 2431 14907 2437
rect 14849 2397 14861 2431
rect 14895 2428 14907 2431
rect 15565 2431 15623 2437
rect 15565 2428 15577 2431
rect 14895 2400 15577 2428
rect 14895 2397 14907 2400
rect 14849 2391 14907 2397
rect 15565 2397 15577 2400
rect 15611 2428 15623 2431
rect 15932 2431 15990 2437
rect 15932 2428 15944 2431
rect 15611 2400 15944 2428
rect 15611 2397 15623 2400
rect 15565 2391 15623 2397
rect 15932 2397 15944 2400
rect 15978 2397 15990 2431
rect 17494 2428 17500 2440
rect 17455 2400 17500 2428
rect 15932 2391 15990 2397
rect 17494 2388 17500 2400
rect 17552 2388 17558 2440
rect 2405 2363 2535 2369
rect 2405 2329 2417 2363
rect 2451 2329 2489 2363
rect 2523 2360 2535 2363
rect 3065 2363 3183 2369
rect 3065 2360 3137 2363
rect 2523 2332 3137 2360
rect 2523 2329 2535 2332
rect 2405 2323 2535 2329
rect 3125 2329 3137 2332
rect 3171 2360 3183 2363
rect 4981 2363 5111 2369
rect 4981 2360 4993 2363
rect 3171 2332 4993 2360
rect 3171 2329 3183 2332
rect 3125 2323 3183 2329
rect 4908 2292 4936 2332
rect 4981 2329 4993 2332
rect 5027 2329 5065 2363
rect 5099 2360 5111 2363
rect 5641 2363 5759 2369
rect 5641 2360 5713 2363
rect 5099 2332 5713 2360
rect 5099 2329 5111 2332
rect 4981 2323 5111 2329
rect 5701 2329 5713 2332
rect 5747 2329 5759 2363
rect 5701 2323 5759 2329
rect 9421 2363 9539 2369
rect 9421 2329 9433 2363
rect 9467 2360 9539 2363
rect 10069 2363 10199 2369
rect 10069 2360 10081 2363
rect 9467 2332 10081 2360
rect 9467 2329 9479 2332
rect 9421 2323 9479 2329
rect 10069 2329 10081 2332
rect 10115 2329 10153 2363
rect 10187 2360 10199 2363
rect 12273 2363 12391 2369
rect 10187 2332 11836 2360
rect 10187 2329 10199 2332
rect 10069 2323 10199 2329
rect 5258 2292 5264 2304
rect 4908 2264 5264 2292
rect 5258 2252 5264 2264
rect 5316 2252 5322 2304
rect 9306 2252 9312 2304
rect 9364 2292 9370 2304
rect 10244 2292 10272 2332
rect 9364 2264 10272 2292
rect 11808 2292 11836 2332
rect 12273 2329 12285 2363
rect 12319 2360 12391 2363
rect 12921 2363 13051 2369
rect 12921 2360 12933 2363
rect 12319 2332 12933 2360
rect 12319 2329 12331 2332
rect 12273 2323 12331 2329
rect 12921 2329 12933 2332
rect 12967 2329 13005 2363
rect 13039 2360 13051 2363
rect 14573 2363 14691 2369
rect 14573 2360 14585 2363
rect 13039 2332 14585 2360
rect 13039 2329 13051 2332
rect 12921 2323 13051 2329
rect 12710 2292 12716 2304
rect 11808 2264 12716 2292
rect 9364 2252 9370 2264
rect 12710 2252 12716 2264
rect 12768 2292 12774 2304
rect 13096 2292 13124 2332
rect 14573 2329 14585 2332
rect 14619 2360 14691 2363
rect 15221 2363 15351 2369
rect 15221 2360 15233 2363
rect 14619 2332 15233 2360
rect 14619 2329 14631 2332
rect 14573 2323 14631 2329
rect 15221 2329 15233 2332
rect 15267 2329 15305 2363
rect 15339 2329 15351 2363
rect 15746 2360 15752 2372
rect 15707 2332 15752 2360
rect 15221 2323 15351 2329
rect 15746 2320 15752 2332
rect 15804 2320 15810 2372
rect 12768 2264 13124 2292
rect 12768 2252 12774 2264
rect 17402 2252 17408 2304
rect 17460 2292 17466 2304
rect 17681 2295 17739 2301
rect 17681 2292 17693 2295
rect 17460 2264 17693 2292
rect 17460 2252 17466 2264
rect 17681 2261 17693 2264
rect 17727 2261 17739 2295
rect 17681 2255 17739 2261
rect 1104 2202 19019 2224
rect 1104 2193 5388 2202
rect 1104 2159 1133 2193
rect 1167 2159 1225 2193
rect 1259 2159 1317 2193
rect 1351 2159 1409 2193
rect 1443 2159 1501 2193
rect 1535 2159 1593 2193
rect 1627 2159 1685 2193
rect 1719 2159 1777 2193
rect 1811 2159 1869 2193
rect 1903 2159 1961 2193
rect 1995 2159 2053 2193
rect 2087 2159 2145 2193
rect 2179 2159 2237 2193
rect 2271 2159 2329 2193
rect 2363 2159 2421 2193
rect 2455 2159 2513 2193
rect 2547 2159 2605 2193
rect 2639 2159 2697 2193
rect 2731 2159 2789 2193
rect 2823 2159 2881 2193
rect 2915 2159 2973 2193
rect 3007 2159 3065 2193
rect 3099 2159 3157 2193
rect 3191 2159 3249 2193
rect 3283 2159 3341 2193
rect 3375 2159 3433 2193
rect 3467 2159 3525 2193
rect 3559 2159 3617 2193
rect 3651 2159 3709 2193
rect 3743 2159 3801 2193
rect 3835 2159 3893 2193
rect 3927 2159 3985 2193
rect 4019 2159 4077 2193
rect 4111 2159 4169 2193
rect 4203 2159 4261 2193
rect 4295 2159 4353 2193
rect 4387 2159 4445 2193
rect 4479 2159 4537 2193
rect 4571 2159 4629 2193
rect 4663 2159 4721 2193
rect 4755 2159 4813 2193
rect 4847 2159 4905 2193
rect 4939 2159 4997 2193
rect 5031 2159 5089 2193
rect 5123 2159 5181 2193
rect 5215 2159 5273 2193
rect 5307 2159 5365 2193
rect 1104 2150 5388 2159
rect 5440 2150 5452 2202
rect 5504 2150 5516 2202
rect 5568 2193 5580 2202
rect 5632 2193 5644 2202
rect 5696 2193 9827 2202
rect 9879 2193 9891 2202
rect 5632 2159 5641 2193
rect 5696 2159 5733 2193
rect 5767 2159 5825 2193
rect 5859 2159 5917 2193
rect 5951 2159 6009 2193
rect 6043 2159 6101 2193
rect 6135 2159 6193 2193
rect 6227 2159 6285 2193
rect 6319 2159 6377 2193
rect 6411 2159 6469 2193
rect 6503 2159 6561 2193
rect 6595 2159 6653 2193
rect 6687 2159 6745 2193
rect 6779 2159 6837 2193
rect 6871 2159 6929 2193
rect 6963 2159 7021 2193
rect 7055 2159 7113 2193
rect 7147 2159 7205 2193
rect 7239 2159 7297 2193
rect 7331 2159 7389 2193
rect 7423 2159 7481 2193
rect 7515 2159 7573 2193
rect 7607 2159 7665 2193
rect 7699 2159 7757 2193
rect 7791 2159 7849 2193
rect 7883 2159 7941 2193
rect 7975 2159 8033 2193
rect 8067 2159 8125 2193
rect 8159 2159 8217 2193
rect 8251 2159 8309 2193
rect 8343 2159 8401 2193
rect 8435 2159 8493 2193
rect 8527 2159 8585 2193
rect 8619 2159 8677 2193
rect 8711 2159 8769 2193
rect 8803 2159 8861 2193
rect 8895 2159 8953 2193
rect 8987 2159 9045 2193
rect 9079 2159 9137 2193
rect 9171 2159 9229 2193
rect 9263 2159 9321 2193
rect 9355 2159 9413 2193
rect 9447 2159 9505 2193
rect 9539 2159 9597 2193
rect 9631 2159 9689 2193
rect 9723 2159 9781 2193
rect 9815 2159 9827 2193
rect 5568 2150 5580 2159
rect 5632 2150 5644 2159
rect 5696 2150 9827 2159
rect 9879 2150 9891 2159
rect 9943 2150 9955 2202
rect 10007 2150 10019 2202
rect 10071 2193 10083 2202
rect 10135 2193 14266 2202
rect 14318 2193 14330 2202
rect 14382 2193 14394 2202
rect 10135 2159 10149 2193
rect 10183 2159 10241 2193
rect 10275 2159 10333 2193
rect 10367 2159 10425 2193
rect 10459 2159 10517 2193
rect 10551 2159 10609 2193
rect 10643 2159 10701 2193
rect 10735 2159 10793 2193
rect 10827 2159 10885 2193
rect 10919 2159 10977 2193
rect 11011 2159 11069 2193
rect 11103 2159 11161 2193
rect 11195 2159 11253 2193
rect 11287 2159 11345 2193
rect 11379 2159 11437 2193
rect 11471 2159 11529 2193
rect 11563 2159 11621 2193
rect 11655 2159 11713 2193
rect 11747 2159 11805 2193
rect 11839 2159 11897 2193
rect 11931 2159 11989 2193
rect 12023 2159 12081 2193
rect 12115 2159 12173 2193
rect 12207 2159 12265 2193
rect 12299 2159 12357 2193
rect 12391 2159 12449 2193
rect 12483 2159 12541 2193
rect 12575 2159 12633 2193
rect 12667 2159 12725 2193
rect 12759 2159 12817 2193
rect 12851 2159 12909 2193
rect 12943 2159 13001 2193
rect 13035 2159 13093 2193
rect 13127 2159 13185 2193
rect 13219 2159 13277 2193
rect 13311 2159 13369 2193
rect 13403 2159 13461 2193
rect 13495 2159 13553 2193
rect 13587 2159 13645 2193
rect 13679 2159 13737 2193
rect 13771 2159 13829 2193
rect 13863 2159 13921 2193
rect 13955 2159 14013 2193
rect 14047 2159 14105 2193
rect 14139 2159 14197 2193
rect 14231 2159 14266 2193
rect 14323 2159 14330 2193
rect 10071 2150 10083 2159
rect 10135 2150 14266 2159
rect 14318 2150 14330 2159
rect 14382 2150 14394 2159
rect 14446 2150 14458 2202
rect 14510 2150 14522 2202
rect 14574 2193 18705 2202
rect 14599 2159 14657 2193
rect 14691 2159 14749 2193
rect 14783 2159 14841 2193
rect 14875 2159 14933 2193
rect 14967 2159 15025 2193
rect 15059 2159 15117 2193
rect 15151 2159 15209 2193
rect 15243 2159 15301 2193
rect 15335 2159 15393 2193
rect 15427 2159 15485 2193
rect 15519 2159 15577 2193
rect 15611 2159 15669 2193
rect 15703 2159 15761 2193
rect 15795 2159 15853 2193
rect 15887 2159 15945 2193
rect 15979 2159 16037 2193
rect 16071 2159 16129 2193
rect 16163 2159 16221 2193
rect 16255 2159 16313 2193
rect 16347 2159 16405 2193
rect 16439 2159 16497 2193
rect 16531 2159 16589 2193
rect 16623 2159 16681 2193
rect 16715 2159 16773 2193
rect 16807 2159 16865 2193
rect 16899 2159 16957 2193
rect 16991 2159 17049 2193
rect 17083 2159 17141 2193
rect 17175 2159 17233 2193
rect 17267 2159 17325 2193
rect 17359 2159 17417 2193
rect 17451 2159 17509 2193
rect 17543 2159 17601 2193
rect 17635 2159 17693 2193
rect 17727 2159 17785 2193
rect 17819 2159 17877 2193
rect 17911 2159 17969 2193
rect 18003 2159 18061 2193
rect 18095 2159 18153 2193
rect 18187 2159 18245 2193
rect 18279 2159 18337 2193
rect 18371 2159 18429 2193
rect 18463 2159 18521 2193
rect 18555 2159 18613 2193
rect 18647 2159 18705 2193
rect 14574 2150 18705 2159
rect 18757 2150 18769 2202
rect 18821 2193 18833 2202
rect 18831 2159 18833 2193
rect 18821 2150 18833 2159
rect 18885 2150 18897 2202
rect 18949 2150 18961 2202
rect 19013 2150 19019 2202
rect 1104 2128 19019 2150
rect 10686 2048 10692 2100
rect 10744 2088 10750 2100
rect 17494 2088 17500 2100
rect 10744 2060 17500 2088
rect 10744 2048 10750 2060
rect 17494 2048 17500 2060
rect 17552 2048 17558 2100
<< via1 >>
rect 5388 7633 5440 7642
rect 5388 7599 5399 7633
rect 5399 7599 5440 7633
rect 5388 7590 5440 7599
rect 5452 7633 5504 7642
rect 5452 7599 5457 7633
rect 5457 7599 5491 7633
rect 5491 7599 5504 7633
rect 5452 7590 5504 7599
rect 5516 7633 5568 7642
rect 5580 7633 5632 7642
rect 5644 7633 5696 7642
rect 9827 7633 9879 7642
rect 9891 7633 9943 7642
rect 5516 7599 5549 7633
rect 5549 7599 5568 7633
rect 5580 7599 5583 7633
rect 5583 7599 5632 7633
rect 5644 7599 5675 7633
rect 5675 7599 5696 7633
rect 9827 7599 9873 7633
rect 9873 7599 9879 7633
rect 9891 7599 9907 7633
rect 9907 7599 9943 7633
rect 5516 7590 5568 7599
rect 5580 7590 5632 7599
rect 5644 7590 5696 7599
rect 9827 7590 9879 7599
rect 9891 7590 9943 7599
rect 9955 7633 10007 7642
rect 9955 7599 9965 7633
rect 9965 7599 9999 7633
rect 9999 7599 10007 7633
rect 9955 7590 10007 7599
rect 10019 7633 10071 7642
rect 10083 7633 10135 7642
rect 14266 7633 14318 7642
rect 14330 7633 14382 7642
rect 14394 7633 14446 7642
rect 10019 7599 10057 7633
rect 10057 7599 10071 7633
rect 10083 7599 10091 7633
rect 10091 7599 10135 7633
rect 14266 7599 14289 7633
rect 14289 7599 14318 7633
rect 14330 7599 14381 7633
rect 14381 7599 14382 7633
rect 14394 7599 14415 7633
rect 14415 7599 14446 7633
rect 10019 7590 10071 7599
rect 10083 7590 10135 7599
rect 14266 7590 14318 7599
rect 14330 7590 14382 7599
rect 14394 7590 14446 7599
rect 14458 7633 14510 7642
rect 14458 7599 14473 7633
rect 14473 7599 14507 7633
rect 14507 7599 14510 7633
rect 14458 7590 14510 7599
rect 14522 7633 14574 7642
rect 18705 7633 18757 7642
rect 14522 7599 14565 7633
rect 14565 7599 14574 7633
rect 18705 7599 18739 7633
rect 18739 7599 18757 7633
rect 14522 7590 14574 7599
rect 18705 7590 18757 7599
rect 18769 7633 18821 7642
rect 18769 7599 18797 7633
rect 18797 7599 18821 7633
rect 18769 7590 18821 7599
rect 18833 7590 18885 7642
rect 18897 7590 18949 7642
rect 18961 7590 19013 7642
rect 1124 7488 1176 7540
rect 3332 7488 3384 7540
rect 5724 7531 5776 7540
rect 5724 7497 5733 7531
rect 5733 7497 5767 7531
rect 5767 7497 5776 7531
rect 5724 7488 5776 7497
rect 7932 7531 7984 7540
rect 7932 7497 7941 7531
rect 7941 7497 7975 7531
rect 7975 7497 7984 7531
rect 7932 7488 7984 7497
rect 12440 7531 12492 7540
rect 12440 7497 12449 7531
rect 12449 7497 12483 7531
rect 12483 7497 12492 7531
rect 12440 7488 12492 7497
rect 14648 7531 14700 7540
rect 14648 7497 14657 7531
rect 14657 7497 14691 7531
rect 14691 7497 14700 7531
rect 14648 7488 14700 7497
rect 16580 7488 16632 7540
rect 18420 7488 18472 7540
rect 7288 7420 7340 7472
rect 7012 7352 7064 7404
rect 7472 7352 7524 7404
rect 10232 7420 10284 7472
rect 13820 7352 13872 7404
rect 16856 7395 16908 7404
rect 16856 7361 16865 7395
rect 16865 7361 16899 7395
rect 16899 7361 16908 7395
rect 16856 7352 16908 7361
rect 7932 7284 7984 7336
rect 13360 7284 13412 7336
rect 10324 7259 10376 7268
rect 10324 7225 10333 7259
rect 10333 7225 10367 7259
rect 10367 7225 10376 7259
rect 10324 7216 10376 7225
rect 11060 7148 11112 7200
rect 3169 7089 3221 7098
rect 3169 7055 3191 7089
rect 3191 7055 3221 7089
rect 3169 7046 3221 7055
rect 3233 7089 3285 7098
rect 3233 7055 3249 7089
rect 3249 7055 3283 7089
rect 3283 7055 3285 7089
rect 3233 7046 3285 7055
rect 3297 7089 3349 7098
rect 3361 7089 3413 7098
rect 3297 7055 3341 7089
rect 3341 7055 3349 7089
rect 3361 7055 3375 7089
rect 3375 7055 3413 7089
rect 3297 7046 3349 7055
rect 3361 7046 3413 7055
rect 3425 7089 3477 7098
rect 3425 7055 3433 7089
rect 3433 7055 3467 7089
rect 3467 7055 3477 7089
rect 3425 7046 3477 7055
rect 7608 7046 7660 7098
rect 7672 7089 7724 7098
rect 7672 7055 7699 7089
rect 7699 7055 7724 7089
rect 7672 7046 7724 7055
rect 7736 7089 7788 7098
rect 7800 7089 7852 7098
rect 7864 7089 7916 7098
rect 12047 7089 12099 7098
rect 12111 7089 12163 7098
rect 12175 7089 12227 7098
rect 7736 7055 7757 7089
rect 7757 7055 7788 7089
rect 7800 7055 7849 7089
rect 7849 7055 7852 7089
rect 7864 7055 7883 7089
rect 7883 7055 7916 7089
rect 12047 7055 12081 7089
rect 12081 7055 12099 7089
rect 12111 7055 12115 7089
rect 12115 7055 12163 7089
rect 12175 7055 12207 7089
rect 12207 7055 12227 7089
rect 7736 7046 7788 7055
rect 7800 7046 7852 7055
rect 7864 7046 7916 7055
rect 12047 7046 12099 7055
rect 12111 7046 12163 7055
rect 12175 7046 12227 7055
rect 12239 7089 12291 7098
rect 12239 7055 12265 7089
rect 12265 7055 12291 7089
rect 12239 7046 12291 7055
rect 12303 7046 12355 7098
rect 16486 7089 16538 7098
rect 16486 7055 16497 7089
rect 16497 7055 16531 7089
rect 16531 7055 16538 7089
rect 16486 7046 16538 7055
rect 16550 7089 16602 7098
rect 16614 7089 16666 7098
rect 16550 7055 16589 7089
rect 16589 7055 16602 7089
rect 16614 7055 16623 7089
rect 16623 7055 16666 7089
rect 16550 7046 16602 7055
rect 16614 7046 16666 7055
rect 16678 7089 16730 7098
rect 16678 7055 16681 7089
rect 16681 7055 16715 7089
rect 16715 7055 16730 7089
rect 16678 7046 16730 7055
rect 16742 7089 16794 7098
rect 16742 7055 16773 7089
rect 16773 7055 16794 7089
rect 16742 7046 16794 7055
rect 5388 6545 5440 6554
rect 5388 6511 5399 6545
rect 5399 6511 5440 6545
rect 5388 6502 5440 6511
rect 5452 6545 5504 6554
rect 5452 6511 5457 6545
rect 5457 6511 5491 6545
rect 5491 6511 5504 6545
rect 5452 6502 5504 6511
rect 5516 6545 5568 6554
rect 5580 6545 5632 6554
rect 5644 6545 5696 6554
rect 9827 6545 9879 6554
rect 9891 6545 9943 6554
rect 5516 6511 5549 6545
rect 5549 6511 5568 6545
rect 5580 6511 5583 6545
rect 5583 6511 5632 6545
rect 5644 6511 5675 6545
rect 5675 6511 5696 6545
rect 9827 6511 9873 6545
rect 9873 6511 9879 6545
rect 9891 6511 9907 6545
rect 9907 6511 9943 6545
rect 5516 6502 5568 6511
rect 5580 6502 5632 6511
rect 5644 6502 5696 6511
rect 9827 6502 9879 6511
rect 9891 6502 9943 6511
rect 9955 6545 10007 6554
rect 9955 6511 9965 6545
rect 9965 6511 9999 6545
rect 9999 6511 10007 6545
rect 9955 6502 10007 6511
rect 10019 6545 10071 6554
rect 10083 6545 10135 6554
rect 14266 6545 14318 6554
rect 14330 6545 14382 6554
rect 14394 6545 14446 6554
rect 10019 6511 10057 6545
rect 10057 6511 10071 6545
rect 10083 6511 10091 6545
rect 10091 6511 10135 6545
rect 14266 6511 14289 6545
rect 14289 6511 14318 6545
rect 14330 6511 14381 6545
rect 14381 6511 14382 6545
rect 14394 6511 14415 6545
rect 14415 6511 14446 6545
rect 10019 6502 10071 6511
rect 10083 6502 10135 6511
rect 14266 6502 14318 6511
rect 14330 6502 14382 6511
rect 14394 6502 14446 6511
rect 14458 6545 14510 6554
rect 14458 6511 14473 6545
rect 14473 6511 14507 6545
rect 14507 6511 14510 6545
rect 14458 6502 14510 6511
rect 14522 6545 14574 6554
rect 18705 6545 18757 6554
rect 14522 6511 14565 6545
rect 14565 6511 14574 6545
rect 18705 6511 18739 6545
rect 18739 6511 18757 6545
rect 14522 6502 14574 6511
rect 18705 6502 18757 6511
rect 18769 6545 18821 6554
rect 18769 6511 18797 6545
rect 18797 6511 18821 6545
rect 18769 6502 18821 6511
rect 18833 6502 18885 6554
rect 18897 6502 18949 6554
rect 18961 6502 19013 6554
rect 8024 6307 8076 6316
rect 8024 6273 8033 6307
rect 8033 6273 8067 6307
rect 8067 6273 8076 6307
rect 8024 6264 8076 6273
rect 8208 6307 8260 6316
rect 8208 6273 8217 6307
rect 8217 6273 8251 6307
rect 8251 6273 8260 6307
rect 8208 6264 8260 6273
rect 10968 6060 11020 6112
rect 3169 6001 3221 6010
rect 3169 5967 3191 6001
rect 3191 5967 3221 6001
rect 3169 5958 3221 5967
rect 3233 6001 3285 6010
rect 3233 5967 3249 6001
rect 3249 5967 3283 6001
rect 3283 5967 3285 6001
rect 3233 5958 3285 5967
rect 3297 6001 3349 6010
rect 3361 6001 3413 6010
rect 3297 5967 3341 6001
rect 3341 5967 3349 6001
rect 3361 5967 3375 6001
rect 3375 5967 3413 6001
rect 3297 5958 3349 5967
rect 3361 5958 3413 5967
rect 3425 6001 3477 6010
rect 3425 5967 3433 6001
rect 3433 5967 3467 6001
rect 3467 5967 3477 6001
rect 3425 5958 3477 5967
rect 7608 5958 7660 6010
rect 7672 6001 7724 6010
rect 7672 5967 7699 6001
rect 7699 5967 7724 6001
rect 7672 5958 7724 5967
rect 7736 6001 7788 6010
rect 7800 6001 7852 6010
rect 7864 6001 7916 6010
rect 12047 6001 12099 6010
rect 12111 6001 12163 6010
rect 12175 6001 12227 6010
rect 7736 5967 7757 6001
rect 7757 5967 7788 6001
rect 7800 5967 7849 6001
rect 7849 5967 7852 6001
rect 7864 5967 7883 6001
rect 7883 5967 7916 6001
rect 12047 5967 12081 6001
rect 12081 5967 12099 6001
rect 12111 5967 12115 6001
rect 12115 5967 12163 6001
rect 12175 5967 12207 6001
rect 12207 5967 12227 6001
rect 7736 5958 7788 5967
rect 7800 5958 7852 5967
rect 7864 5958 7916 5967
rect 12047 5958 12099 5967
rect 12111 5958 12163 5967
rect 12175 5958 12227 5967
rect 12239 6001 12291 6010
rect 12239 5967 12265 6001
rect 12265 5967 12291 6001
rect 12239 5958 12291 5967
rect 12303 5958 12355 6010
rect 16486 6001 16538 6010
rect 16486 5967 16497 6001
rect 16497 5967 16531 6001
rect 16531 5967 16538 6001
rect 16486 5958 16538 5967
rect 16550 6001 16602 6010
rect 16614 6001 16666 6010
rect 16550 5967 16589 6001
rect 16589 5967 16602 6001
rect 16614 5967 16623 6001
rect 16623 5967 16666 6001
rect 16550 5958 16602 5967
rect 16614 5958 16666 5967
rect 16678 6001 16730 6010
rect 16678 5967 16681 6001
rect 16681 5967 16715 6001
rect 16715 5967 16730 6001
rect 16678 5958 16730 5967
rect 16742 6001 16794 6010
rect 16742 5967 16773 6001
rect 16773 5967 16794 6001
rect 16742 5958 16794 5967
rect 8024 5856 8076 5908
rect 8116 5720 8168 5772
rect 6920 5695 6972 5704
rect 6920 5661 6929 5695
rect 6929 5661 6963 5695
rect 6963 5661 6972 5695
rect 6920 5652 6972 5661
rect 7472 5584 7524 5636
rect 11520 5627 11572 5636
rect 11520 5593 11529 5627
rect 11529 5593 11563 5627
rect 11563 5593 11572 5627
rect 11520 5584 11572 5593
rect 11704 5627 11756 5636
rect 11704 5593 11713 5627
rect 11713 5593 11747 5627
rect 11747 5593 11756 5627
rect 11704 5584 11756 5593
rect 12808 5627 12860 5636
rect 12808 5593 12817 5627
rect 12817 5593 12851 5627
rect 12851 5593 12860 5627
rect 12808 5584 12860 5593
rect 12900 5584 12952 5636
rect 4620 5516 4672 5568
rect 7380 5516 7432 5568
rect 13084 5516 13136 5568
rect 15108 5516 15160 5568
rect 5388 5457 5440 5466
rect 5388 5423 5399 5457
rect 5399 5423 5440 5457
rect 5388 5414 5440 5423
rect 5452 5457 5504 5466
rect 5452 5423 5457 5457
rect 5457 5423 5491 5457
rect 5491 5423 5504 5457
rect 5452 5414 5504 5423
rect 5516 5457 5568 5466
rect 5580 5457 5632 5466
rect 5644 5457 5696 5466
rect 9827 5457 9879 5466
rect 9891 5457 9943 5466
rect 5516 5423 5549 5457
rect 5549 5423 5568 5457
rect 5580 5423 5583 5457
rect 5583 5423 5632 5457
rect 5644 5423 5675 5457
rect 5675 5423 5696 5457
rect 9827 5423 9873 5457
rect 9873 5423 9879 5457
rect 9891 5423 9907 5457
rect 9907 5423 9943 5457
rect 5516 5414 5568 5423
rect 5580 5414 5632 5423
rect 5644 5414 5696 5423
rect 9827 5414 9879 5423
rect 9891 5414 9943 5423
rect 9955 5457 10007 5466
rect 9955 5423 9965 5457
rect 9965 5423 9999 5457
rect 9999 5423 10007 5457
rect 9955 5414 10007 5423
rect 10019 5457 10071 5466
rect 10083 5457 10135 5466
rect 14266 5457 14318 5466
rect 14330 5457 14382 5466
rect 14394 5457 14446 5466
rect 10019 5423 10057 5457
rect 10057 5423 10071 5457
rect 10083 5423 10091 5457
rect 10091 5423 10135 5457
rect 14266 5423 14289 5457
rect 14289 5423 14318 5457
rect 14330 5423 14381 5457
rect 14381 5423 14382 5457
rect 14394 5423 14415 5457
rect 14415 5423 14446 5457
rect 10019 5414 10071 5423
rect 10083 5414 10135 5423
rect 14266 5414 14318 5423
rect 14330 5414 14382 5423
rect 14394 5414 14446 5423
rect 14458 5457 14510 5466
rect 14458 5423 14473 5457
rect 14473 5423 14507 5457
rect 14507 5423 14510 5457
rect 14458 5414 14510 5423
rect 14522 5457 14574 5466
rect 18705 5457 18757 5466
rect 14522 5423 14565 5457
rect 14565 5423 14574 5457
rect 18705 5423 18739 5457
rect 18739 5423 18757 5457
rect 14522 5414 14574 5423
rect 18705 5414 18757 5423
rect 18769 5457 18821 5466
rect 18769 5423 18797 5457
rect 18797 5423 18821 5457
rect 18769 5414 18821 5423
rect 18833 5414 18885 5466
rect 18897 5414 18949 5466
rect 18961 5414 19013 5466
rect 7012 5355 7064 5364
rect 4436 5244 4488 5296
rect 7012 5321 7021 5355
rect 7021 5321 7055 5355
rect 7055 5321 7064 5355
rect 7012 5312 7064 5321
rect 7380 5312 7432 5364
rect 6736 5176 6788 5228
rect 3056 5151 3108 5160
rect 3056 5117 3065 5151
rect 3065 5117 3099 5151
rect 3099 5117 3108 5151
rect 3056 5108 3108 5117
rect 9220 5224 9272 5228
rect 9220 5190 9241 5224
rect 9241 5190 9272 5224
rect 9220 5176 9272 5190
rect 11060 5312 11112 5364
rect 11520 5312 11572 5364
rect 10324 5287 10376 5296
rect 10324 5253 10333 5287
rect 10333 5253 10367 5287
rect 10367 5253 10376 5287
rect 12440 5312 12492 5364
rect 10324 5244 10376 5253
rect 13820 5244 13872 5296
rect 12992 5176 13044 5228
rect 13360 5176 13412 5228
rect 8116 5151 8168 5160
rect 4252 5040 4304 5092
rect 8116 5117 8125 5151
rect 8125 5117 8159 5151
rect 8159 5117 8168 5151
rect 8116 5108 8168 5117
rect 9680 5108 9732 5160
rect 4160 4972 4212 5024
rect 6828 4972 6880 5024
rect 11888 5108 11940 5160
rect 12900 5108 12952 5160
rect 13912 5040 13964 5092
rect 9312 4972 9364 5024
rect 10508 4972 10560 5024
rect 15200 4972 15252 5024
rect 3169 4913 3221 4922
rect 3169 4879 3191 4913
rect 3191 4879 3221 4913
rect 3169 4870 3221 4879
rect 3233 4913 3285 4922
rect 3233 4879 3249 4913
rect 3249 4879 3283 4913
rect 3283 4879 3285 4913
rect 3233 4870 3285 4879
rect 3297 4913 3349 4922
rect 3361 4913 3413 4922
rect 3297 4879 3341 4913
rect 3341 4879 3349 4913
rect 3361 4879 3375 4913
rect 3375 4879 3413 4913
rect 3297 4870 3349 4879
rect 3361 4870 3413 4879
rect 3425 4913 3477 4922
rect 3425 4879 3433 4913
rect 3433 4879 3467 4913
rect 3467 4879 3477 4913
rect 3425 4870 3477 4879
rect 7608 4870 7660 4922
rect 7672 4913 7724 4922
rect 7672 4879 7699 4913
rect 7699 4879 7724 4913
rect 7672 4870 7724 4879
rect 7736 4913 7788 4922
rect 7800 4913 7852 4922
rect 7864 4913 7916 4922
rect 12047 4913 12099 4922
rect 12111 4913 12163 4922
rect 12175 4913 12227 4922
rect 7736 4879 7757 4913
rect 7757 4879 7788 4913
rect 7800 4879 7849 4913
rect 7849 4879 7852 4913
rect 7864 4879 7883 4913
rect 7883 4879 7916 4913
rect 12047 4879 12081 4913
rect 12081 4879 12099 4913
rect 12111 4879 12115 4913
rect 12115 4879 12163 4913
rect 12175 4879 12207 4913
rect 12207 4879 12227 4913
rect 7736 4870 7788 4879
rect 7800 4870 7852 4879
rect 7864 4870 7916 4879
rect 12047 4870 12099 4879
rect 12111 4870 12163 4879
rect 12175 4870 12227 4879
rect 12239 4913 12291 4922
rect 12239 4879 12265 4913
rect 12265 4879 12291 4913
rect 12239 4870 12291 4879
rect 12303 4870 12355 4922
rect 16486 4913 16538 4922
rect 16486 4879 16497 4913
rect 16497 4879 16531 4913
rect 16531 4879 16538 4913
rect 16486 4870 16538 4879
rect 16550 4913 16602 4922
rect 16614 4913 16666 4922
rect 16550 4879 16589 4913
rect 16589 4879 16602 4913
rect 16614 4879 16623 4913
rect 16623 4879 16666 4913
rect 16550 4870 16602 4879
rect 16614 4870 16666 4879
rect 16678 4913 16730 4922
rect 16678 4879 16681 4913
rect 16681 4879 16715 4913
rect 16715 4879 16730 4913
rect 16678 4870 16730 4879
rect 16742 4913 16794 4922
rect 16742 4879 16773 4913
rect 16773 4879 16794 4913
rect 16742 4870 16794 4879
rect 6920 4768 6972 4820
rect 3056 4700 3108 4752
rect 8300 4700 8352 4752
rect 2780 4564 2832 4616
rect 8024 4632 8076 4684
rect 8208 4632 8260 4684
rect 6828 4607 6880 4616
rect 6828 4573 6837 4607
rect 6837 4573 6871 4607
rect 6871 4573 6880 4607
rect 6828 4564 6880 4573
rect 7380 4564 7432 4616
rect 7840 4564 7892 4616
rect 10324 4632 10376 4684
rect 9036 4564 9088 4616
rect 9588 4564 9640 4616
rect 10508 4607 10560 4616
rect 10508 4573 10517 4607
rect 10517 4573 10551 4607
rect 10551 4573 10560 4607
rect 10508 4564 10560 4573
rect 4988 4496 5040 4548
rect 6184 4539 6236 4548
rect 6184 4505 6193 4539
rect 6193 4505 6227 4539
rect 6227 4505 6236 4539
rect 6184 4496 6236 4505
rect 8116 4496 8168 4548
rect 8392 4496 8444 4548
rect 9312 4539 9364 4548
rect 9312 4505 9321 4539
rect 9321 4505 9355 4539
rect 9355 4505 9364 4539
rect 9312 4496 9364 4505
rect 10692 4539 10744 4548
rect 10692 4505 10701 4539
rect 10701 4505 10735 4539
rect 10735 4505 10744 4539
rect 10692 4496 10744 4505
rect 11980 4700 12032 4752
rect 11704 4632 11756 4684
rect 10968 4564 11020 4616
rect 11888 4496 11940 4548
rect 12808 4768 12860 4820
rect 12348 4700 12400 4752
rect 13728 4700 13780 4752
rect 12440 4632 12492 4684
rect 16856 4700 16908 4752
rect 12348 4564 12400 4616
rect 15108 4632 15160 4684
rect 13084 4564 13136 4616
rect 15200 4607 15252 4616
rect 15200 4573 15209 4607
rect 15209 4573 15243 4607
rect 15243 4573 15252 4607
rect 15200 4564 15252 4573
rect 15384 4539 15436 4548
rect 2228 4428 2280 4480
rect 4436 4428 4488 4480
rect 6828 4428 6880 4480
rect 7288 4428 7340 4480
rect 8852 4428 8904 4480
rect 9404 4428 9456 4480
rect 10232 4428 10284 4480
rect 10968 4428 11020 4480
rect 11060 4428 11112 4480
rect 12348 4471 12400 4480
rect 12348 4437 12357 4471
rect 12357 4437 12391 4471
rect 12391 4437 12400 4471
rect 12348 4428 12400 4437
rect 15384 4505 15393 4539
rect 15393 4505 15427 4539
rect 15427 4505 15436 4539
rect 15384 4496 15436 4505
rect 16028 4471 16080 4480
rect 16028 4437 16037 4471
rect 16037 4437 16071 4471
rect 16071 4437 16080 4471
rect 16028 4428 16080 4437
rect 16856 4428 16908 4480
rect 5388 4369 5440 4378
rect 5388 4335 5399 4369
rect 5399 4335 5440 4369
rect 5388 4326 5440 4335
rect 5452 4369 5504 4378
rect 5452 4335 5457 4369
rect 5457 4335 5491 4369
rect 5491 4335 5504 4369
rect 5452 4326 5504 4335
rect 5516 4369 5568 4378
rect 5580 4369 5632 4378
rect 5644 4369 5696 4378
rect 9827 4369 9879 4378
rect 9891 4369 9943 4378
rect 5516 4335 5549 4369
rect 5549 4335 5568 4369
rect 5580 4335 5583 4369
rect 5583 4335 5632 4369
rect 5644 4335 5675 4369
rect 5675 4335 5696 4369
rect 9827 4335 9873 4369
rect 9873 4335 9879 4369
rect 9891 4335 9907 4369
rect 9907 4335 9943 4369
rect 5516 4326 5568 4335
rect 5580 4326 5632 4335
rect 5644 4326 5696 4335
rect 9827 4326 9879 4335
rect 9891 4326 9943 4335
rect 9955 4369 10007 4378
rect 9955 4335 9965 4369
rect 9965 4335 9999 4369
rect 9999 4335 10007 4369
rect 9955 4326 10007 4335
rect 10019 4369 10071 4378
rect 10083 4369 10135 4378
rect 14266 4369 14318 4378
rect 14330 4369 14382 4378
rect 14394 4369 14446 4378
rect 10019 4335 10057 4369
rect 10057 4335 10071 4369
rect 10083 4335 10091 4369
rect 10091 4335 10135 4369
rect 14266 4335 14289 4369
rect 14289 4335 14318 4369
rect 14330 4335 14381 4369
rect 14381 4335 14382 4369
rect 14394 4335 14415 4369
rect 14415 4335 14446 4369
rect 10019 4326 10071 4335
rect 10083 4326 10135 4335
rect 14266 4326 14318 4335
rect 14330 4326 14382 4335
rect 14394 4326 14446 4335
rect 14458 4369 14510 4378
rect 14458 4335 14473 4369
rect 14473 4335 14507 4369
rect 14507 4335 14510 4369
rect 14458 4326 14510 4335
rect 14522 4369 14574 4378
rect 18705 4369 18757 4378
rect 14522 4335 14565 4369
rect 14565 4335 14574 4369
rect 18705 4335 18739 4369
rect 18739 4335 18757 4369
rect 14522 4326 14574 4335
rect 18705 4326 18757 4335
rect 18769 4369 18821 4378
rect 18769 4335 18797 4369
rect 18797 4335 18821 4369
rect 18769 4326 18821 4335
rect 18833 4326 18885 4378
rect 18897 4326 18949 4378
rect 18961 4326 19013 4378
rect 4988 4224 5040 4276
rect 6184 4224 6236 4276
rect 2228 4131 2280 4140
rect 2228 4097 2237 4131
rect 2237 4097 2271 4131
rect 2271 4097 2280 4131
rect 2228 4088 2280 4097
rect 4436 4156 4488 4208
rect 5264 4156 5316 4208
rect 4712 4088 4764 4140
rect 7288 4156 7340 4208
rect 7932 4224 7984 4276
rect 8392 4267 8444 4276
rect 8392 4233 8401 4267
rect 8401 4233 8435 4267
rect 8435 4233 8444 4267
rect 8392 4224 8444 4233
rect 8852 4156 8904 4208
rect 9036 4224 9088 4276
rect 11152 4224 11204 4276
rect 11888 4224 11940 4276
rect 9404 4156 9456 4208
rect 11796 4156 11848 4208
rect 6828 4131 6880 4140
rect 6828 4097 6837 4131
rect 6837 4097 6871 4131
rect 6871 4097 6880 4131
rect 6828 4088 6880 4097
rect 7472 4088 7524 4140
rect 11888 4088 11940 4140
rect 2504 3884 2556 3936
rect 4528 3952 4580 4004
rect 7104 4020 7156 4072
rect 7840 4020 7892 4072
rect 6920 3952 6972 4004
rect 11060 4020 11112 4072
rect 11152 4020 11204 4072
rect 13636 4020 13688 4072
rect 8484 3952 8536 4004
rect 4160 3884 4212 3936
rect 4712 3884 4764 3936
rect 4988 3884 5040 3936
rect 9128 3884 9180 3936
rect 9404 3884 9456 3936
rect 13728 3952 13780 4004
rect 12992 3884 13044 3936
rect 13084 3884 13136 3936
rect 3169 3825 3221 3834
rect 3169 3791 3191 3825
rect 3191 3791 3221 3825
rect 3169 3782 3221 3791
rect 3233 3825 3285 3834
rect 3233 3791 3249 3825
rect 3249 3791 3283 3825
rect 3283 3791 3285 3825
rect 3233 3782 3285 3791
rect 3297 3825 3349 3834
rect 3361 3825 3413 3834
rect 3297 3791 3341 3825
rect 3341 3791 3349 3825
rect 3361 3791 3375 3825
rect 3375 3791 3413 3825
rect 3297 3782 3349 3791
rect 3361 3782 3413 3791
rect 3425 3825 3477 3834
rect 3425 3791 3433 3825
rect 3433 3791 3467 3825
rect 3467 3791 3477 3825
rect 3425 3782 3477 3791
rect 7608 3782 7660 3834
rect 7672 3825 7724 3834
rect 7672 3791 7699 3825
rect 7699 3791 7724 3825
rect 7672 3782 7724 3791
rect 7736 3825 7788 3834
rect 7800 3825 7852 3834
rect 7864 3825 7916 3834
rect 12047 3825 12099 3834
rect 12111 3825 12163 3834
rect 12175 3825 12227 3834
rect 7736 3791 7757 3825
rect 7757 3791 7788 3825
rect 7800 3791 7849 3825
rect 7849 3791 7852 3825
rect 7864 3791 7883 3825
rect 7883 3791 7916 3825
rect 12047 3791 12081 3825
rect 12081 3791 12099 3825
rect 12111 3791 12115 3825
rect 12115 3791 12163 3825
rect 12175 3791 12207 3825
rect 12207 3791 12227 3825
rect 7736 3782 7788 3791
rect 7800 3782 7852 3791
rect 7864 3782 7916 3791
rect 12047 3782 12099 3791
rect 12111 3782 12163 3791
rect 12175 3782 12227 3791
rect 12239 3825 12291 3834
rect 12239 3791 12265 3825
rect 12265 3791 12291 3825
rect 12239 3782 12291 3791
rect 12303 3782 12355 3834
rect 16486 3825 16538 3834
rect 16486 3791 16497 3825
rect 16497 3791 16531 3825
rect 16531 3791 16538 3825
rect 16486 3782 16538 3791
rect 16550 3825 16602 3834
rect 16614 3825 16666 3834
rect 16550 3791 16589 3825
rect 16589 3791 16602 3825
rect 16614 3791 16623 3825
rect 16623 3791 16666 3825
rect 16550 3782 16602 3791
rect 16614 3782 16666 3791
rect 16678 3825 16730 3834
rect 16678 3791 16681 3825
rect 16681 3791 16715 3825
rect 16715 3791 16730 3825
rect 16678 3782 16730 3791
rect 16742 3825 16794 3834
rect 16742 3791 16773 3825
rect 16773 3791 16794 3825
rect 16742 3782 16794 3791
rect 4160 3680 4212 3732
rect 6736 3680 6788 3732
rect 16028 3680 16080 3732
rect 8484 3655 8536 3664
rect 8484 3621 8493 3655
rect 8493 3621 8527 3655
rect 8527 3621 8536 3655
rect 8484 3612 8536 3621
rect 9220 3612 9272 3664
rect 11152 3655 11204 3664
rect 11152 3621 11161 3655
rect 11161 3621 11195 3655
rect 11195 3621 11204 3655
rect 11152 3612 11204 3621
rect 11796 3612 11848 3664
rect 2504 3544 2556 3596
rect 9404 3544 9456 3596
rect 6736 3519 6788 3528
rect 6736 3485 6745 3519
rect 6745 3485 6779 3519
rect 6779 3485 6788 3519
rect 6736 3476 6788 3485
rect 2964 3340 3016 3392
rect 4436 3408 4488 3460
rect 8300 3476 8352 3528
rect 9128 3519 9180 3528
rect 9128 3485 9137 3519
rect 9137 3485 9171 3519
rect 9171 3485 9180 3519
rect 9128 3476 9180 3485
rect 13452 3544 13504 3596
rect 13728 3587 13780 3596
rect 13728 3553 13737 3587
rect 13737 3553 13771 3587
rect 13771 3553 13780 3587
rect 13728 3544 13780 3553
rect 10232 3519 10284 3528
rect 10232 3485 10241 3519
rect 10241 3485 10275 3519
rect 10275 3485 10284 3519
rect 10232 3476 10284 3485
rect 10968 3519 11020 3528
rect 10968 3485 10977 3519
rect 10977 3485 11011 3519
rect 11011 3485 11020 3519
rect 10968 3476 11020 3485
rect 6920 3340 6972 3392
rect 11704 3408 11756 3460
rect 8668 3340 8720 3392
rect 12716 3408 12768 3460
rect 5388 3281 5440 3290
rect 5388 3247 5399 3281
rect 5399 3247 5440 3281
rect 5388 3238 5440 3247
rect 5452 3281 5504 3290
rect 5452 3247 5457 3281
rect 5457 3247 5491 3281
rect 5491 3247 5504 3281
rect 5452 3238 5504 3247
rect 5516 3281 5568 3290
rect 5580 3281 5632 3290
rect 5644 3281 5696 3290
rect 9827 3281 9879 3290
rect 9891 3281 9943 3290
rect 5516 3247 5549 3281
rect 5549 3247 5568 3281
rect 5580 3247 5583 3281
rect 5583 3247 5632 3281
rect 5644 3247 5675 3281
rect 5675 3247 5696 3281
rect 9827 3247 9873 3281
rect 9873 3247 9879 3281
rect 9891 3247 9907 3281
rect 9907 3247 9943 3281
rect 5516 3238 5568 3247
rect 5580 3238 5632 3247
rect 5644 3238 5696 3247
rect 9827 3238 9879 3247
rect 9891 3238 9943 3247
rect 9955 3281 10007 3290
rect 9955 3247 9965 3281
rect 9965 3247 9999 3281
rect 9999 3247 10007 3281
rect 9955 3238 10007 3247
rect 10019 3281 10071 3290
rect 10083 3281 10135 3290
rect 14266 3281 14318 3290
rect 14330 3281 14382 3290
rect 14394 3281 14446 3290
rect 10019 3247 10057 3281
rect 10057 3247 10071 3281
rect 10083 3247 10091 3281
rect 10091 3247 10135 3281
rect 14266 3247 14289 3281
rect 14289 3247 14318 3281
rect 14330 3247 14381 3281
rect 14381 3247 14382 3281
rect 14394 3247 14415 3281
rect 14415 3247 14446 3281
rect 10019 3238 10071 3247
rect 10083 3238 10135 3247
rect 14266 3238 14318 3247
rect 14330 3238 14382 3247
rect 14394 3238 14446 3247
rect 14458 3281 14510 3290
rect 14458 3247 14473 3281
rect 14473 3247 14507 3281
rect 14507 3247 14510 3281
rect 14458 3238 14510 3247
rect 14522 3281 14574 3290
rect 18705 3281 18757 3290
rect 14522 3247 14565 3281
rect 14565 3247 14574 3281
rect 18705 3247 18739 3281
rect 18739 3247 18757 3281
rect 14522 3238 14574 3247
rect 18705 3238 18757 3247
rect 18769 3281 18821 3290
rect 18769 3247 18797 3281
rect 18797 3247 18821 3281
rect 18769 3238 18821 3247
rect 18833 3238 18885 3290
rect 18897 3238 18949 3290
rect 18961 3238 19013 3290
rect 1952 3179 2004 3188
rect 1952 3145 1961 3179
rect 1961 3145 1995 3179
rect 1995 3145 2004 3179
rect 1952 3136 2004 3145
rect 7104 3136 7156 3188
rect 7932 3136 7984 3188
rect 2964 3111 3016 3120
rect 2964 3077 2977 3111
rect 2977 3077 3011 3111
rect 3011 3077 3016 3111
rect 2964 3068 3016 3077
rect 4252 3068 4304 3120
rect 4160 3043 4212 3052
rect 4160 3009 4169 3043
rect 4169 3009 4203 3043
rect 4203 3009 4212 3043
rect 4160 3000 4212 3009
rect 4528 3043 4580 3052
rect 4528 3009 4537 3043
rect 4537 3009 4571 3043
rect 4571 3009 4580 3043
rect 4528 3000 4580 3009
rect 5264 2932 5316 2984
rect 7380 3068 7432 3120
rect 9220 3136 9272 3188
rect 10876 3136 10928 3188
rect 13728 3136 13780 3188
rect 8668 3111 8720 3120
rect 8668 3077 8689 3111
rect 8689 3077 8720 3111
rect 9404 3111 9456 3120
rect 8668 3068 8720 3077
rect 9404 3077 9413 3111
rect 9413 3077 9447 3111
rect 9447 3077 9456 3111
rect 9404 3068 9456 3077
rect 12716 3111 12768 3120
rect 12716 3077 12729 3111
rect 12729 3077 12763 3111
rect 12763 3077 12768 3111
rect 9036 3000 9088 3052
rect 10692 3000 10744 3052
rect 12716 3068 12768 3077
rect 12900 3068 12952 3120
rect 13452 3068 13504 3120
rect 13912 3043 13964 3052
rect 13912 3009 13921 3043
rect 13921 3009 13955 3043
rect 13955 3009 13964 3043
rect 13912 3000 13964 3009
rect 7472 2796 7524 2848
rect 9588 2796 9640 2848
rect 10876 2864 10928 2916
rect 11704 2907 11756 2916
rect 11704 2873 11713 2907
rect 11713 2873 11747 2907
rect 11747 2873 11756 2907
rect 11704 2864 11756 2873
rect 13728 2932 13780 2984
rect 15384 2864 15436 2916
rect 15752 2864 15804 2916
rect 16856 2864 16908 2916
rect 12440 2796 12492 2848
rect 3169 2737 3221 2746
rect 3169 2703 3191 2737
rect 3191 2703 3221 2737
rect 3169 2694 3221 2703
rect 3233 2737 3285 2746
rect 3233 2703 3249 2737
rect 3249 2703 3283 2737
rect 3283 2703 3285 2737
rect 3233 2694 3285 2703
rect 3297 2737 3349 2746
rect 3361 2737 3413 2746
rect 3297 2703 3341 2737
rect 3341 2703 3349 2737
rect 3361 2703 3375 2737
rect 3375 2703 3413 2737
rect 3297 2694 3349 2703
rect 3361 2694 3413 2703
rect 3425 2737 3477 2746
rect 3425 2703 3433 2737
rect 3433 2703 3467 2737
rect 3467 2703 3477 2737
rect 3425 2694 3477 2703
rect 7608 2694 7660 2746
rect 7672 2737 7724 2746
rect 7672 2703 7699 2737
rect 7699 2703 7724 2737
rect 7672 2694 7724 2703
rect 7736 2737 7788 2746
rect 7800 2737 7852 2746
rect 7864 2737 7916 2746
rect 12047 2737 12099 2746
rect 12111 2737 12163 2746
rect 12175 2737 12227 2746
rect 7736 2703 7757 2737
rect 7757 2703 7788 2737
rect 7800 2703 7849 2737
rect 7849 2703 7852 2737
rect 7864 2703 7883 2737
rect 7883 2703 7916 2737
rect 12047 2703 12081 2737
rect 12081 2703 12099 2737
rect 12111 2703 12115 2737
rect 12115 2703 12163 2737
rect 12175 2703 12207 2737
rect 12207 2703 12227 2737
rect 7736 2694 7788 2703
rect 7800 2694 7852 2703
rect 7864 2694 7916 2703
rect 12047 2694 12099 2703
rect 12111 2694 12163 2703
rect 12175 2694 12227 2703
rect 12239 2737 12291 2746
rect 12239 2703 12265 2737
rect 12265 2703 12291 2737
rect 12239 2694 12291 2703
rect 12303 2694 12355 2746
rect 16486 2737 16538 2746
rect 16486 2703 16497 2737
rect 16497 2703 16531 2737
rect 16531 2703 16538 2737
rect 16486 2694 16538 2703
rect 16550 2737 16602 2746
rect 16614 2737 16666 2746
rect 16550 2703 16589 2737
rect 16589 2703 16602 2737
rect 16614 2703 16623 2737
rect 16623 2703 16666 2737
rect 16550 2694 16602 2703
rect 16614 2694 16666 2703
rect 16678 2737 16730 2746
rect 16678 2703 16681 2737
rect 16681 2703 16715 2737
rect 16715 2703 16730 2737
rect 16678 2694 16730 2703
rect 16742 2737 16794 2746
rect 16742 2703 16773 2737
rect 16773 2703 16794 2737
rect 16742 2694 16794 2703
rect 7012 2592 7064 2644
rect 8208 2592 8260 2644
rect 12900 2592 12952 2644
rect 9588 2524 9640 2576
rect 2504 2456 2556 2508
rect 4160 2456 4212 2508
rect 4620 2456 4672 2508
rect 8024 2456 8076 2508
rect 11704 2456 11756 2508
rect 13728 2499 13780 2508
rect 13728 2465 13737 2499
rect 13737 2465 13771 2499
rect 13771 2465 13780 2499
rect 13728 2456 13780 2465
rect 1952 2363 2004 2372
rect 1952 2329 1961 2363
rect 1961 2329 1995 2363
rect 1995 2329 2004 2363
rect 1952 2320 2004 2329
rect 10876 2431 10928 2440
rect 10876 2397 10885 2431
rect 10885 2397 10919 2431
rect 10919 2397 10928 2431
rect 10876 2388 10928 2397
rect 17500 2431 17552 2440
rect 17500 2397 17509 2431
rect 17509 2397 17543 2431
rect 17543 2397 17552 2431
rect 17500 2388 17552 2397
rect 5264 2252 5316 2304
rect 9312 2252 9364 2304
rect 12716 2252 12768 2304
rect 15752 2363 15804 2372
rect 15752 2329 15761 2363
rect 15761 2329 15795 2363
rect 15795 2329 15804 2363
rect 15752 2320 15804 2329
rect 17408 2252 17460 2304
rect 5388 2193 5440 2202
rect 5388 2159 5399 2193
rect 5399 2159 5440 2193
rect 5388 2150 5440 2159
rect 5452 2193 5504 2202
rect 5452 2159 5457 2193
rect 5457 2159 5491 2193
rect 5491 2159 5504 2193
rect 5452 2150 5504 2159
rect 5516 2193 5568 2202
rect 5580 2193 5632 2202
rect 5644 2193 5696 2202
rect 9827 2193 9879 2202
rect 9891 2193 9943 2202
rect 5516 2159 5549 2193
rect 5549 2159 5568 2193
rect 5580 2159 5583 2193
rect 5583 2159 5632 2193
rect 5644 2159 5675 2193
rect 5675 2159 5696 2193
rect 9827 2159 9873 2193
rect 9873 2159 9879 2193
rect 9891 2159 9907 2193
rect 9907 2159 9943 2193
rect 5516 2150 5568 2159
rect 5580 2150 5632 2159
rect 5644 2150 5696 2159
rect 9827 2150 9879 2159
rect 9891 2150 9943 2159
rect 9955 2193 10007 2202
rect 9955 2159 9965 2193
rect 9965 2159 9999 2193
rect 9999 2159 10007 2193
rect 9955 2150 10007 2159
rect 10019 2193 10071 2202
rect 10083 2193 10135 2202
rect 14266 2193 14318 2202
rect 14330 2193 14382 2202
rect 14394 2193 14446 2202
rect 10019 2159 10057 2193
rect 10057 2159 10071 2193
rect 10083 2159 10091 2193
rect 10091 2159 10135 2193
rect 14266 2159 14289 2193
rect 14289 2159 14318 2193
rect 14330 2159 14381 2193
rect 14381 2159 14382 2193
rect 14394 2159 14415 2193
rect 14415 2159 14446 2193
rect 10019 2150 10071 2159
rect 10083 2150 10135 2159
rect 14266 2150 14318 2159
rect 14330 2150 14382 2159
rect 14394 2150 14446 2159
rect 14458 2193 14510 2202
rect 14458 2159 14473 2193
rect 14473 2159 14507 2193
rect 14507 2159 14510 2193
rect 14458 2150 14510 2159
rect 14522 2193 14574 2202
rect 18705 2193 18757 2202
rect 14522 2159 14565 2193
rect 14565 2159 14574 2193
rect 18705 2159 18739 2193
rect 18739 2159 18757 2193
rect 14522 2150 14574 2159
rect 18705 2150 18757 2159
rect 18769 2193 18821 2202
rect 18769 2159 18797 2193
rect 18797 2159 18821 2193
rect 18769 2150 18821 2159
rect 18833 2150 18885 2202
rect 18897 2150 18949 2202
rect 18961 2150 19013 2202
rect 10692 2048 10744 2100
rect 17500 2048 17552 2100
<< metal2 >>
rect 1122 9200 1178 10000
rect 3330 9200 3386 10000
rect 5538 9330 5594 10000
rect 7746 9330 7802 10000
rect 9954 9330 10010 10000
rect 12162 9330 12218 10000
rect 14370 9330 14426 10000
rect 5538 9302 5764 9330
rect 5538 9200 5594 9302
rect 1136 7546 1164 9200
rect 3344 7546 3372 9200
rect 5388 7644 5696 7653
rect 5388 7642 5394 7644
rect 5450 7642 5474 7644
rect 5530 7642 5554 7644
rect 5610 7642 5634 7644
rect 5690 7642 5696 7644
rect 5450 7590 5452 7642
rect 5632 7590 5634 7642
rect 5388 7588 5394 7590
rect 5450 7588 5474 7590
rect 5530 7588 5554 7590
rect 5610 7588 5634 7590
rect 5690 7588 5696 7590
rect 5388 7579 5696 7588
rect 5736 7546 5764 9302
rect 7746 9302 7972 9330
rect 7746 9200 7802 9302
rect 7944 7546 7972 9302
rect 9954 9302 10272 9330
rect 9954 9200 10010 9302
rect 9827 7644 10135 7653
rect 9827 7642 9833 7644
rect 9889 7642 9913 7644
rect 9969 7642 9993 7644
rect 10049 7642 10073 7644
rect 10129 7642 10135 7644
rect 9889 7590 9891 7642
rect 10071 7590 10073 7642
rect 9827 7588 9833 7590
rect 9889 7588 9913 7590
rect 9969 7588 9993 7590
rect 10049 7588 10073 7590
rect 10129 7588 10135 7590
rect 9827 7579 10135 7588
rect 1124 7540 1176 7546
rect 1124 7482 1176 7488
rect 3332 7540 3384 7546
rect 3332 7482 3384 7488
rect 5724 7540 5776 7546
rect 5724 7482 5776 7488
rect 7932 7540 7984 7546
rect 7932 7482 7984 7488
rect 10244 7478 10272 9302
rect 12162 9302 12388 9330
rect 12162 9200 12218 9302
rect 12360 7528 12388 9302
rect 14370 9302 14688 9330
rect 14370 9200 14426 9302
rect 14266 7644 14574 7653
rect 14266 7642 14272 7644
rect 14328 7642 14352 7644
rect 14408 7642 14432 7644
rect 14488 7642 14512 7644
rect 14568 7642 14574 7644
rect 14328 7590 14330 7642
rect 14510 7590 14512 7642
rect 14266 7588 14272 7590
rect 14328 7588 14352 7590
rect 14408 7588 14432 7590
rect 14488 7588 14512 7590
rect 14568 7588 14574 7590
rect 14266 7579 14574 7588
rect 14660 7546 14688 9302
rect 16578 9200 16634 10000
rect 18786 9330 18842 10000
rect 18432 9302 18842 9330
rect 16592 7546 16620 9200
rect 18432 7546 18460 9302
rect 18786 9200 18842 9302
rect 18705 7644 19013 7653
rect 18705 7642 18711 7644
rect 18767 7642 18791 7644
rect 18847 7642 18871 7644
rect 18927 7642 18951 7644
rect 19007 7642 19013 7644
rect 18767 7590 18769 7642
rect 18949 7590 18951 7642
rect 18705 7588 18711 7590
rect 18767 7588 18791 7590
rect 18847 7588 18871 7590
rect 18927 7588 18951 7590
rect 19007 7588 19013 7590
rect 18705 7579 19013 7588
rect 12440 7540 12492 7546
rect 12360 7500 12440 7528
rect 12440 7482 12492 7488
rect 14648 7540 14700 7546
rect 14648 7482 14700 7488
rect 16580 7540 16632 7546
rect 16580 7482 16632 7488
rect 18420 7540 18472 7546
rect 18420 7482 18472 7488
rect 7288 7472 7340 7478
rect 7288 7414 7340 7420
rect 10232 7472 10284 7478
rect 10232 7414 10284 7420
rect 7012 7404 7064 7410
rect 7012 7346 7064 7352
rect 3169 7100 3477 7109
rect 3169 7098 3175 7100
rect 3231 7098 3255 7100
rect 3311 7098 3335 7100
rect 3391 7098 3415 7100
rect 3471 7098 3477 7100
rect 3231 7046 3233 7098
rect 3413 7046 3415 7098
rect 3169 7044 3175 7046
rect 3231 7044 3255 7046
rect 3311 7044 3335 7046
rect 3391 7044 3415 7046
rect 3471 7044 3477 7046
rect 3169 7035 3477 7044
rect 5388 6556 5696 6565
rect 5388 6554 5394 6556
rect 5450 6554 5474 6556
rect 5530 6554 5554 6556
rect 5610 6554 5634 6556
rect 5690 6554 5696 6556
rect 5450 6502 5452 6554
rect 5632 6502 5634 6554
rect 5388 6500 5394 6502
rect 5450 6500 5474 6502
rect 5530 6500 5554 6502
rect 5610 6500 5634 6502
rect 5690 6500 5696 6502
rect 5388 6491 5696 6500
rect 3169 6012 3477 6021
rect 3169 6010 3175 6012
rect 3231 6010 3255 6012
rect 3311 6010 3335 6012
rect 3391 6010 3415 6012
rect 3471 6010 3477 6012
rect 3231 5958 3233 6010
rect 3413 5958 3415 6010
rect 3169 5956 3175 5958
rect 3231 5956 3255 5958
rect 3311 5956 3335 5958
rect 3391 5956 3415 5958
rect 3471 5956 3477 5958
rect 3169 5947 3477 5956
rect 6920 5704 6972 5710
rect 6920 5646 6972 5652
rect 4620 5568 4672 5574
rect 4620 5510 4672 5516
rect 4436 5296 4488 5302
rect 4436 5238 4488 5244
rect 3056 5160 3108 5166
rect 3056 5102 3108 5108
rect 3068 4758 3096 5102
rect 4252 5092 4304 5098
rect 4252 5034 4304 5040
rect 4160 5024 4212 5030
rect 4160 4966 4212 4972
rect 3169 4924 3477 4933
rect 3169 4922 3175 4924
rect 3231 4922 3255 4924
rect 3311 4922 3335 4924
rect 3391 4922 3415 4924
rect 3471 4922 3477 4924
rect 3231 4870 3233 4922
rect 3413 4870 3415 4922
rect 3169 4868 3175 4870
rect 3231 4868 3255 4870
rect 3311 4868 3335 4870
rect 3391 4868 3415 4870
rect 3471 4868 3477 4870
rect 3169 4859 3477 4868
rect 3056 4752 3108 4758
rect 3056 4694 3108 4700
rect 2780 4616 2832 4622
rect 2780 4558 2832 4564
rect 2228 4480 2280 4486
rect 2228 4422 2280 4428
rect 2240 4146 2268 4422
rect 2228 4140 2280 4146
rect 2228 4082 2280 4088
rect 2792 4060 2820 4558
rect 2700 4032 2820 4060
rect 2504 3936 2556 3942
rect 2504 3878 2556 3884
rect 2516 3602 2544 3878
rect 2504 3596 2556 3602
rect 2504 3538 2556 3544
rect 1952 3188 2004 3194
rect 1952 3130 2004 3136
rect 1964 2378 1992 3130
rect 2516 2514 2544 3538
rect 2504 2508 2556 2514
rect 2504 2450 2556 2456
rect 2700 2394 2728 4032
rect 4172 3942 4200 4966
rect 4160 3936 4212 3942
rect 4160 3878 4212 3884
rect 3169 3836 3477 3845
rect 3169 3834 3175 3836
rect 3231 3834 3255 3836
rect 3311 3834 3335 3836
rect 3391 3834 3415 3836
rect 3471 3834 3477 3836
rect 3231 3782 3233 3834
rect 3413 3782 3415 3834
rect 3169 3780 3175 3782
rect 3231 3780 3255 3782
rect 3311 3780 3335 3782
rect 3391 3780 3415 3782
rect 3471 3780 3477 3782
rect 3169 3771 3477 3780
rect 4172 3738 4200 3878
rect 4160 3732 4212 3738
rect 4160 3674 4212 3680
rect 2964 3392 3016 3398
rect 2964 3334 3016 3340
rect 2976 3126 3004 3334
rect 2964 3120 3016 3126
rect 2964 3062 3016 3068
rect 4172 3058 4200 3674
rect 4264 3126 4292 5034
rect 4448 4486 4476 5238
rect 4436 4480 4488 4486
rect 4436 4422 4488 4428
rect 4448 4214 4476 4422
rect 4436 4208 4488 4214
rect 4436 4150 4488 4156
rect 4448 3466 4476 4150
rect 4528 4004 4580 4010
rect 4528 3946 4580 3952
rect 4436 3460 4488 3466
rect 4436 3402 4488 3408
rect 4252 3120 4304 3126
rect 4252 3062 4304 3068
rect 4540 3058 4568 3946
rect 4160 3052 4212 3058
rect 4160 2994 4212 3000
rect 4528 3052 4580 3058
rect 4528 2994 4580 3000
rect 3169 2748 3477 2757
rect 3169 2746 3175 2748
rect 3231 2746 3255 2748
rect 3311 2746 3335 2748
rect 3391 2746 3415 2748
rect 3471 2746 3477 2748
rect 3231 2694 3233 2746
rect 3413 2694 3415 2746
rect 3169 2692 3175 2694
rect 3231 2692 3255 2694
rect 3311 2692 3335 2694
rect 3391 2692 3415 2694
rect 3471 2692 3477 2694
rect 3169 2683 3477 2692
rect 4172 2514 4200 2994
rect 4632 2514 4660 5510
rect 5388 5468 5696 5477
rect 5388 5466 5394 5468
rect 5450 5466 5474 5468
rect 5530 5466 5554 5468
rect 5610 5466 5634 5468
rect 5690 5466 5696 5468
rect 5450 5414 5452 5466
rect 5632 5414 5634 5466
rect 5388 5412 5394 5414
rect 5450 5412 5474 5414
rect 5530 5412 5554 5414
rect 5610 5412 5634 5414
rect 5690 5412 5696 5414
rect 5388 5403 5696 5412
rect 6736 5228 6788 5234
rect 6736 5170 6788 5176
rect 4988 4548 5040 4554
rect 4988 4490 5040 4496
rect 6184 4548 6236 4554
rect 6184 4490 6236 4496
rect 5000 4282 5028 4490
rect 5388 4380 5696 4389
rect 5388 4378 5394 4380
rect 5450 4378 5474 4380
rect 5530 4378 5554 4380
rect 5610 4378 5634 4380
rect 5690 4378 5696 4380
rect 5450 4326 5452 4378
rect 5632 4326 5634 4378
rect 5388 4324 5394 4326
rect 5450 4324 5474 4326
rect 5530 4324 5554 4326
rect 5610 4324 5634 4326
rect 5690 4324 5696 4326
rect 5388 4315 5696 4324
rect 6196 4282 6224 4490
rect 4988 4276 5040 4282
rect 4988 4218 5040 4224
rect 6184 4276 6236 4282
rect 6184 4218 6236 4224
rect 4712 4140 4764 4146
rect 4712 4082 4764 4088
rect 4724 3942 4752 4082
rect 5000 3942 5028 4218
rect 5264 4208 5316 4214
rect 5264 4150 5316 4156
rect 4712 3936 4764 3942
rect 4712 3878 4764 3884
rect 4988 3936 5040 3942
rect 4988 3878 5040 3884
rect 5276 2990 5304 4150
rect 6748 3738 6776 5170
rect 6828 5024 6880 5030
rect 6828 4966 6880 4972
rect 6840 4622 6868 4966
rect 6932 4826 6960 5646
rect 7024 5370 7052 7346
rect 7012 5364 7064 5370
rect 7012 5306 7064 5312
rect 6920 4820 6972 4826
rect 6920 4762 6972 4768
rect 6828 4616 6880 4622
rect 6828 4558 6880 4564
rect 6828 4480 6880 4486
rect 6828 4422 6880 4428
rect 6840 4146 6868 4422
rect 6828 4140 6880 4146
rect 6828 4082 6880 4088
rect 6920 4004 6972 4010
rect 6920 3946 6972 3952
rect 6736 3732 6788 3738
rect 6736 3674 6788 3680
rect 6748 3534 6776 3674
rect 6736 3528 6788 3534
rect 6736 3470 6788 3476
rect 6932 3398 6960 3946
rect 6920 3392 6972 3398
rect 6920 3334 6972 3340
rect 5388 3292 5696 3301
rect 5388 3290 5394 3292
rect 5450 3290 5474 3292
rect 5530 3290 5554 3292
rect 5610 3290 5634 3292
rect 5690 3290 5696 3292
rect 5450 3238 5452 3290
rect 5632 3238 5634 3290
rect 5388 3236 5394 3238
rect 5450 3236 5474 3238
rect 5530 3236 5554 3238
rect 5610 3236 5634 3238
rect 5690 3236 5696 3238
rect 5388 3227 5696 3236
rect 5264 2984 5316 2990
rect 5264 2926 5316 2932
rect 4160 2508 4212 2514
rect 4160 2450 4212 2456
rect 4620 2508 4672 2514
rect 4620 2450 4672 2456
rect 1952 2372 2004 2378
rect 1952 2314 2004 2320
rect 2516 2366 2728 2394
rect 2516 800 2544 2366
rect 5276 2310 5304 2926
rect 7024 2650 7052 5306
rect 7300 4486 7328 7414
rect 7472 7404 7524 7410
rect 7472 7346 7524 7352
rect 13820 7404 13872 7410
rect 13820 7346 13872 7352
rect 16856 7404 16908 7410
rect 16856 7346 16908 7352
rect 7484 5642 7512 7346
rect 7932 7336 7984 7342
rect 7932 7278 7984 7284
rect 13360 7336 13412 7342
rect 13360 7278 13412 7284
rect 7608 7100 7916 7109
rect 7608 7098 7614 7100
rect 7670 7098 7694 7100
rect 7750 7098 7774 7100
rect 7830 7098 7854 7100
rect 7910 7098 7916 7100
rect 7670 7046 7672 7098
rect 7852 7046 7854 7098
rect 7608 7044 7614 7046
rect 7670 7044 7694 7046
rect 7750 7044 7774 7046
rect 7830 7044 7854 7046
rect 7910 7044 7916 7046
rect 7608 7035 7916 7044
rect 7608 6012 7916 6021
rect 7608 6010 7614 6012
rect 7670 6010 7694 6012
rect 7750 6010 7774 6012
rect 7830 6010 7854 6012
rect 7910 6010 7916 6012
rect 7670 5958 7672 6010
rect 7852 5958 7854 6010
rect 7608 5956 7614 5958
rect 7670 5956 7694 5958
rect 7750 5956 7774 5958
rect 7830 5956 7854 5958
rect 7910 5956 7916 5958
rect 7608 5947 7916 5956
rect 7472 5636 7524 5642
rect 7472 5578 7524 5584
rect 7380 5568 7432 5574
rect 7380 5510 7432 5516
rect 7392 5370 7420 5510
rect 7380 5364 7432 5370
rect 7380 5306 7432 5312
rect 7392 4622 7420 5306
rect 7380 4616 7432 4622
rect 7380 4558 7432 4564
rect 7288 4480 7340 4486
rect 7288 4422 7340 4428
rect 7300 4214 7328 4422
rect 7288 4208 7340 4214
rect 7288 4150 7340 4156
rect 7484 4146 7512 5578
rect 7608 4924 7916 4933
rect 7608 4922 7614 4924
rect 7670 4922 7694 4924
rect 7750 4922 7774 4924
rect 7830 4922 7854 4924
rect 7910 4922 7916 4924
rect 7670 4870 7672 4922
rect 7852 4870 7854 4922
rect 7608 4868 7614 4870
rect 7670 4868 7694 4870
rect 7750 4868 7774 4870
rect 7830 4868 7854 4870
rect 7910 4868 7916 4870
rect 7608 4859 7916 4868
rect 7840 4616 7892 4622
rect 7840 4558 7892 4564
rect 7472 4140 7524 4146
rect 7472 4082 7524 4088
rect 7852 4078 7880 4558
rect 7944 4282 7972 7278
rect 10324 7268 10376 7274
rect 10324 7210 10376 7216
rect 9827 6556 10135 6565
rect 9827 6554 9833 6556
rect 9889 6554 9913 6556
rect 9969 6554 9993 6556
rect 10049 6554 10073 6556
rect 10129 6554 10135 6556
rect 9889 6502 9891 6554
rect 10071 6502 10073 6554
rect 9827 6500 9833 6502
rect 9889 6500 9913 6502
rect 9969 6500 9993 6502
rect 10049 6500 10073 6502
rect 10129 6500 10135 6502
rect 9827 6491 10135 6500
rect 8024 6316 8076 6322
rect 8024 6258 8076 6264
rect 8208 6316 8260 6322
rect 8208 6258 8260 6264
rect 8036 5914 8064 6258
rect 8024 5908 8076 5914
rect 8024 5850 8076 5856
rect 8116 5772 8168 5778
rect 8116 5714 8168 5720
rect 8128 5166 8156 5714
rect 8116 5160 8168 5166
rect 8116 5102 8168 5108
rect 8024 4684 8076 4690
rect 8024 4626 8076 4632
rect 7932 4276 7984 4282
rect 7932 4218 7984 4224
rect 7104 4072 7156 4078
rect 7104 4014 7156 4020
rect 7840 4072 7892 4078
rect 7840 4014 7892 4020
rect 7116 3194 7144 4014
rect 7608 3836 7916 3845
rect 7608 3834 7614 3836
rect 7670 3834 7694 3836
rect 7750 3834 7774 3836
rect 7830 3834 7854 3836
rect 7910 3834 7916 3836
rect 7670 3782 7672 3834
rect 7852 3782 7854 3834
rect 7608 3780 7614 3782
rect 7670 3780 7694 3782
rect 7750 3780 7774 3782
rect 7830 3780 7854 3782
rect 7910 3780 7916 3782
rect 7608 3771 7916 3780
rect 7378 3360 7434 3369
rect 7378 3295 7434 3304
rect 7104 3188 7156 3194
rect 7104 3130 7156 3136
rect 7116 3097 7144 3130
rect 7392 3126 7420 3295
rect 7944 3194 7972 4218
rect 7932 3188 7984 3194
rect 7932 3130 7984 3136
rect 7380 3120 7432 3126
rect 7102 3088 7158 3097
rect 7380 3062 7432 3068
rect 7102 3023 7158 3032
rect 7472 2848 7524 2854
rect 7472 2790 7524 2796
rect 7012 2644 7064 2650
rect 7012 2586 7064 2592
rect 5264 2304 5316 2310
rect 5264 2246 5316 2252
rect 5388 2204 5696 2213
rect 5388 2202 5394 2204
rect 5450 2202 5474 2204
rect 5530 2202 5554 2204
rect 5610 2202 5634 2204
rect 5690 2202 5696 2204
rect 5450 2150 5452 2202
rect 5632 2150 5634 2202
rect 5388 2148 5394 2150
rect 5450 2148 5474 2150
rect 5530 2148 5554 2150
rect 5610 2148 5634 2150
rect 5690 2148 5696 2150
rect 5388 2139 5696 2148
rect 7484 800 7512 2790
rect 7608 2748 7916 2757
rect 7608 2746 7614 2748
rect 7670 2746 7694 2748
rect 7750 2746 7774 2748
rect 7830 2746 7854 2748
rect 7910 2746 7916 2748
rect 7670 2694 7672 2746
rect 7852 2694 7854 2746
rect 7608 2692 7614 2694
rect 7670 2692 7694 2694
rect 7750 2692 7774 2694
rect 7830 2692 7854 2694
rect 7910 2692 7916 2694
rect 7608 2683 7916 2692
rect 8036 2514 8064 4626
rect 8128 4554 8156 5102
rect 8220 4690 8248 6258
rect 9827 5468 10135 5477
rect 9827 5466 9833 5468
rect 9889 5466 9913 5468
rect 9969 5466 9993 5468
rect 10049 5466 10073 5468
rect 10129 5466 10135 5468
rect 9889 5414 9891 5466
rect 10071 5414 10073 5466
rect 9827 5412 9833 5414
rect 9889 5412 9913 5414
rect 9969 5412 9993 5414
rect 10049 5412 10073 5414
rect 10129 5412 10135 5414
rect 9827 5403 10135 5412
rect 10336 5302 10364 7210
rect 11060 7200 11112 7206
rect 11060 7142 11112 7148
rect 10968 6112 11020 6118
rect 10968 6054 11020 6060
rect 10324 5296 10376 5302
rect 10324 5238 10376 5244
rect 9220 5228 9272 5234
rect 9220 5170 9272 5176
rect 8300 4752 8352 4758
rect 8300 4694 8352 4700
rect 8208 4684 8260 4690
rect 8208 4626 8260 4632
rect 8116 4548 8168 4554
rect 8116 4490 8168 4496
rect 8128 2774 8156 4490
rect 8312 3534 8340 4694
rect 9036 4616 9088 4622
rect 9036 4558 9088 4564
rect 8392 4548 8444 4554
rect 8392 4490 8444 4496
rect 8404 4282 8432 4490
rect 8852 4480 8904 4486
rect 8852 4422 8904 4428
rect 8392 4276 8444 4282
rect 8392 4218 8444 4224
rect 8864 4214 8892 4422
rect 9048 4282 9076 4558
rect 9036 4276 9088 4282
rect 9036 4218 9088 4224
rect 8852 4208 8904 4214
rect 8852 4150 8904 4156
rect 8484 4004 8536 4010
rect 8484 3946 8536 3952
rect 8496 3670 8524 3946
rect 9128 3936 9180 3942
rect 9128 3878 9180 3884
rect 8484 3664 8536 3670
rect 8484 3606 8536 3612
rect 9140 3534 9168 3878
rect 9232 3670 9260 5170
rect 9680 5160 9732 5166
rect 9680 5102 9732 5108
rect 9312 5024 9364 5030
rect 9312 4966 9364 4972
rect 9324 4554 9352 4966
rect 9588 4616 9640 4622
rect 9588 4558 9640 4564
rect 9312 4548 9364 4554
rect 9312 4490 9364 4496
rect 9404 4480 9456 4486
rect 9404 4422 9456 4428
rect 9416 4214 9444 4422
rect 9404 4208 9456 4214
rect 9404 4150 9456 4156
rect 9404 3936 9456 3942
rect 9404 3878 9456 3884
rect 9220 3664 9272 3670
rect 9220 3606 9272 3612
rect 8300 3528 8352 3534
rect 8300 3470 8352 3476
rect 9128 3528 9180 3534
rect 9128 3470 9180 3476
rect 8312 3369 8340 3470
rect 8668 3392 8720 3398
rect 8298 3360 8354 3369
rect 8668 3334 8720 3340
rect 8298 3295 8354 3304
rect 8680 3126 8708 3334
rect 9232 3194 9260 3606
rect 9416 3602 9444 3878
rect 9404 3596 9456 3602
rect 9404 3538 9456 3544
rect 9220 3188 9272 3194
rect 9220 3130 9272 3136
rect 8668 3120 8720 3126
rect 8668 3062 8720 3068
rect 9034 3088 9090 3097
rect 9034 3023 9036 3032
rect 9088 3023 9090 3032
rect 9036 2994 9088 3000
rect 9232 2774 9260 3130
rect 9416 3126 9444 3538
rect 9404 3120 9456 3126
rect 9404 3062 9456 3068
rect 9600 2854 9628 4558
rect 9588 2848 9640 2854
rect 9588 2790 9640 2796
rect 8128 2746 8248 2774
rect 9232 2746 9352 2774
rect 8220 2650 8248 2746
rect 8208 2644 8260 2650
rect 8208 2586 8260 2592
rect 8024 2508 8076 2514
rect 8024 2450 8076 2456
rect 9324 2310 9352 2746
rect 9692 2666 9720 5102
rect 10336 4690 10364 5238
rect 10508 5024 10560 5030
rect 10508 4966 10560 4972
rect 10324 4684 10376 4690
rect 10324 4626 10376 4632
rect 10520 4622 10548 4966
rect 10980 4622 11008 6054
rect 11072 5370 11100 7142
rect 12047 7100 12355 7109
rect 12047 7098 12053 7100
rect 12109 7098 12133 7100
rect 12189 7098 12213 7100
rect 12269 7098 12293 7100
rect 12349 7098 12355 7100
rect 12109 7046 12111 7098
rect 12291 7046 12293 7098
rect 12047 7044 12053 7046
rect 12109 7044 12133 7046
rect 12189 7044 12213 7046
rect 12269 7044 12293 7046
rect 12349 7044 12355 7046
rect 12047 7035 12355 7044
rect 12047 6012 12355 6021
rect 12047 6010 12053 6012
rect 12109 6010 12133 6012
rect 12189 6010 12213 6012
rect 12269 6010 12293 6012
rect 12349 6010 12355 6012
rect 12109 5958 12111 6010
rect 12291 5958 12293 6010
rect 12047 5956 12053 5958
rect 12109 5956 12133 5958
rect 12189 5956 12213 5958
rect 12269 5956 12293 5958
rect 12349 5956 12355 5958
rect 12047 5947 12355 5956
rect 11520 5636 11572 5642
rect 11520 5578 11572 5584
rect 11704 5636 11756 5642
rect 11704 5578 11756 5584
rect 12808 5636 12860 5642
rect 12808 5578 12860 5584
rect 12900 5636 12952 5642
rect 12900 5578 12952 5584
rect 11532 5370 11560 5578
rect 11060 5364 11112 5370
rect 11520 5364 11572 5370
rect 11112 5324 11192 5352
rect 11060 5306 11112 5312
rect 10508 4616 10560 4622
rect 10508 4558 10560 4564
rect 10968 4616 11020 4622
rect 10968 4558 11020 4564
rect 10692 4548 10744 4554
rect 10692 4490 10744 4496
rect 10232 4480 10284 4486
rect 10232 4422 10284 4428
rect 9827 4380 10135 4389
rect 9827 4378 9833 4380
rect 9889 4378 9913 4380
rect 9969 4378 9993 4380
rect 10049 4378 10073 4380
rect 10129 4378 10135 4380
rect 9889 4326 9891 4378
rect 10071 4326 10073 4378
rect 9827 4324 9833 4326
rect 9889 4324 9913 4326
rect 9969 4324 9993 4326
rect 10049 4324 10073 4326
rect 10129 4324 10135 4326
rect 9827 4315 10135 4324
rect 10244 3534 10272 4422
rect 10232 3528 10284 3534
rect 10232 3470 10284 3476
rect 9827 3292 10135 3301
rect 9827 3290 9833 3292
rect 9889 3290 9913 3292
rect 9969 3290 9993 3292
rect 10049 3290 10073 3292
rect 10129 3290 10135 3292
rect 9889 3238 9891 3290
rect 10071 3238 10073 3290
rect 9827 3236 9833 3238
rect 9889 3236 9913 3238
rect 9969 3236 9993 3238
rect 10049 3236 10073 3238
rect 10129 3236 10135 3238
rect 9827 3227 10135 3236
rect 10704 3058 10732 4490
rect 10968 4480 11020 4486
rect 10968 4422 11020 4428
rect 11060 4480 11112 4486
rect 11060 4422 11112 4428
rect 10980 3534 11008 4422
rect 11072 4078 11100 4422
rect 11164 4282 11192 5324
rect 11520 5306 11572 5312
rect 11716 4690 11744 5578
rect 12440 5364 12492 5370
rect 12440 5306 12492 5312
rect 11888 5160 11940 5166
rect 11808 5108 11888 5114
rect 11808 5102 11940 5108
rect 11808 5086 11928 5102
rect 11704 4684 11756 4690
rect 11704 4626 11756 4632
rect 11152 4276 11204 4282
rect 11152 4218 11204 4224
rect 11060 4072 11112 4078
rect 11060 4014 11112 4020
rect 11152 4072 11204 4078
rect 11152 4014 11204 4020
rect 11164 3670 11192 4014
rect 11152 3664 11204 3670
rect 11152 3606 11204 3612
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 11716 3466 11744 4626
rect 11808 4214 11836 5086
rect 12047 4924 12355 4933
rect 12047 4922 12053 4924
rect 12109 4922 12133 4924
rect 12189 4922 12213 4924
rect 12269 4922 12293 4924
rect 12349 4922 12355 4924
rect 12109 4870 12111 4922
rect 12291 4870 12293 4922
rect 12047 4868 12053 4870
rect 12109 4868 12133 4870
rect 12189 4868 12213 4870
rect 12269 4868 12293 4870
rect 12349 4868 12355 4870
rect 12047 4859 12355 4868
rect 11980 4752 12032 4758
rect 12348 4752 12400 4758
rect 12032 4700 12348 4706
rect 11980 4694 12400 4700
rect 11992 4678 12388 4694
rect 12452 4690 12480 5306
rect 12820 4826 12848 5578
rect 12912 5166 12940 5578
rect 13084 5568 13136 5574
rect 13084 5510 13136 5516
rect 12992 5228 13044 5234
rect 12992 5170 13044 5176
rect 12900 5160 12952 5166
rect 12900 5102 12952 5108
rect 12808 4820 12860 4826
rect 12808 4762 12860 4768
rect 12440 4684 12492 4690
rect 12440 4626 12492 4632
rect 12348 4616 12400 4622
rect 12348 4558 12400 4564
rect 11888 4548 11940 4554
rect 11888 4490 11940 4496
rect 11900 4282 11928 4490
rect 12360 4486 12388 4558
rect 12348 4480 12400 4486
rect 12348 4422 12400 4428
rect 11888 4276 11940 4282
rect 11888 4218 11940 4224
rect 11796 4208 11848 4214
rect 11796 4150 11848 4156
rect 11808 3670 11836 4150
rect 11888 4140 11940 4146
rect 11888 4082 11940 4088
rect 11900 4049 11928 4082
rect 11886 4040 11942 4049
rect 11886 3975 11942 3984
rect 12047 3836 12355 3845
rect 12047 3834 12053 3836
rect 12109 3834 12133 3836
rect 12189 3834 12213 3836
rect 12269 3834 12293 3836
rect 12349 3834 12355 3836
rect 12109 3782 12111 3834
rect 12291 3782 12293 3834
rect 12047 3780 12053 3782
rect 12109 3780 12133 3782
rect 12189 3780 12213 3782
rect 12269 3780 12293 3782
rect 12349 3780 12355 3782
rect 12047 3771 12355 3780
rect 11796 3664 11848 3670
rect 11796 3606 11848 3612
rect 11704 3460 11756 3466
rect 11704 3402 11756 3408
rect 10876 3188 10928 3194
rect 10876 3130 10928 3136
rect 10692 3052 10744 3058
rect 10692 2994 10744 3000
rect 9600 2638 9720 2666
rect 9600 2582 9628 2638
rect 9588 2576 9640 2582
rect 9588 2518 9640 2524
rect 9312 2304 9364 2310
rect 9312 2246 9364 2252
rect 9827 2204 10135 2213
rect 9827 2202 9833 2204
rect 9889 2202 9913 2204
rect 9969 2202 9993 2204
rect 10049 2202 10073 2204
rect 10129 2202 10135 2204
rect 9889 2150 9891 2202
rect 10071 2150 10073 2202
rect 9827 2148 9833 2150
rect 9889 2148 9913 2150
rect 9969 2148 9993 2150
rect 10049 2148 10073 2150
rect 10129 2148 10135 2150
rect 9827 2139 10135 2148
rect 10704 2106 10732 2994
rect 10888 2922 10916 3130
rect 11716 2922 11744 3402
rect 10876 2916 10928 2922
rect 10876 2858 10928 2864
rect 11704 2916 11756 2922
rect 11704 2858 11756 2864
rect 10888 2446 10916 2858
rect 11808 2774 11836 3606
rect 12716 3460 12768 3466
rect 12716 3402 12768 3408
rect 12728 3126 12756 3402
rect 12912 3126 12940 5102
rect 13004 3942 13032 5170
rect 13096 4622 13124 5510
rect 13372 5234 13400 7278
rect 13832 5302 13860 7346
rect 16486 7100 16794 7109
rect 16486 7098 16492 7100
rect 16548 7098 16572 7100
rect 16628 7098 16652 7100
rect 16708 7098 16732 7100
rect 16788 7098 16794 7100
rect 16548 7046 16550 7098
rect 16730 7046 16732 7098
rect 16486 7044 16492 7046
rect 16548 7044 16572 7046
rect 16628 7044 16652 7046
rect 16708 7044 16732 7046
rect 16788 7044 16794 7046
rect 16486 7035 16794 7044
rect 14266 6556 14574 6565
rect 14266 6554 14272 6556
rect 14328 6554 14352 6556
rect 14408 6554 14432 6556
rect 14488 6554 14512 6556
rect 14568 6554 14574 6556
rect 14328 6502 14330 6554
rect 14510 6502 14512 6554
rect 14266 6500 14272 6502
rect 14328 6500 14352 6502
rect 14408 6500 14432 6502
rect 14488 6500 14512 6502
rect 14568 6500 14574 6502
rect 14266 6491 14574 6500
rect 16486 6012 16794 6021
rect 16486 6010 16492 6012
rect 16548 6010 16572 6012
rect 16628 6010 16652 6012
rect 16708 6010 16732 6012
rect 16788 6010 16794 6012
rect 16548 5958 16550 6010
rect 16730 5958 16732 6010
rect 16486 5956 16492 5958
rect 16548 5956 16572 5958
rect 16628 5956 16652 5958
rect 16708 5956 16732 5958
rect 16788 5956 16794 5958
rect 16486 5947 16794 5956
rect 15108 5568 15160 5574
rect 15108 5510 15160 5516
rect 14266 5468 14574 5477
rect 14266 5466 14272 5468
rect 14328 5466 14352 5468
rect 14408 5466 14432 5468
rect 14488 5466 14512 5468
rect 14568 5466 14574 5468
rect 14328 5414 14330 5466
rect 14510 5414 14512 5466
rect 14266 5412 14272 5414
rect 14328 5412 14352 5414
rect 14408 5412 14432 5414
rect 14488 5412 14512 5414
rect 14568 5412 14574 5414
rect 14266 5403 14574 5412
rect 13820 5296 13872 5302
rect 13820 5238 13872 5244
rect 13360 5228 13412 5234
rect 13360 5170 13412 5176
rect 13912 5092 13964 5098
rect 13912 5034 13964 5040
rect 13728 4752 13780 4758
rect 13728 4694 13780 4700
rect 13084 4616 13136 4622
rect 13084 4558 13136 4564
rect 13636 4072 13688 4078
rect 13082 4040 13138 4049
rect 13636 4014 13688 4020
rect 13082 3975 13138 3984
rect 13096 3942 13124 3975
rect 12992 3936 13044 3942
rect 12992 3878 13044 3884
rect 13084 3936 13136 3942
rect 13084 3878 13136 3884
rect 13452 3596 13504 3602
rect 13648 3584 13676 4014
rect 13740 4010 13768 4694
rect 13728 4004 13780 4010
rect 13728 3946 13780 3952
rect 13728 3596 13780 3602
rect 13648 3556 13728 3584
rect 13452 3538 13504 3544
rect 13728 3538 13780 3544
rect 13464 3126 13492 3538
rect 13740 3194 13768 3538
rect 13728 3188 13780 3194
rect 13728 3130 13780 3136
rect 12716 3120 12768 3126
rect 12716 3062 12768 3068
rect 12900 3120 12952 3126
rect 12900 3062 12952 3068
rect 13452 3120 13504 3126
rect 13452 3062 13504 3068
rect 12440 2848 12492 2854
rect 12440 2790 12492 2796
rect 11716 2746 11836 2774
rect 12047 2748 12355 2757
rect 12047 2746 12053 2748
rect 12109 2746 12133 2748
rect 12189 2746 12213 2748
rect 12269 2746 12293 2748
rect 12349 2746 12355 2748
rect 11716 2514 11744 2746
rect 12109 2694 12111 2746
rect 12291 2694 12293 2746
rect 12047 2692 12053 2694
rect 12109 2692 12133 2694
rect 12189 2692 12213 2694
rect 12269 2692 12293 2694
rect 12349 2692 12355 2694
rect 12047 2683 12355 2692
rect 11704 2508 11756 2514
rect 11704 2450 11756 2456
rect 10876 2440 10928 2446
rect 10876 2382 10928 2388
rect 10692 2100 10744 2106
rect 10692 2042 10744 2048
rect 12452 800 12480 2790
rect 12728 2310 12756 3062
rect 12912 2650 12940 3062
rect 13740 2990 13768 3130
rect 13924 3058 13952 5034
rect 15120 4690 15148 5510
rect 15200 5024 15252 5030
rect 15200 4966 15252 4972
rect 15108 4684 15160 4690
rect 15108 4626 15160 4632
rect 15212 4622 15240 4966
rect 16486 4924 16794 4933
rect 16486 4922 16492 4924
rect 16548 4922 16572 4924
rect 16628 4922 16652 4924
rect 16708 4922 16732 4924
rect 16788 4922 16794 4924
rect 16548 4870 16550 4922
rect 16730 4870 16732 4922
rect 16486 4868 16492 4870
rect 16548 4868 16572 4870
rect 16628 4868 16652 4870
rect 16708 4868 16732 4870
rect 16788 4868 16794 4870
rect 16486 4859 16794 4868
rect 16868 4758 16896 7346
rect 18705 6556 19013 6565
rect 18705 6554 18711 6556
rect 18767 6554 18791 6556
rect 18847 6554 18871 6556
rect 18927 6554 18951 6556
rect 19007 6554 19013 6556
rect 18767 6502 18769 6554
rect 18949 6502 18951 6554
rect 18705 6500 18711 6502
rect 18767 6500 18791 6502
rect 18847 6500 18871 6502
rect 18927 6500 18951 6502
rect 19007 6500 19013 6502
rect 18705 6491 19013 6500
rect 18705 5468 19013 5477
rect 18705 5466 18711 5468
rect 18767 5466 18791 5468
rect 18847 5466 18871 5468
rect 18927 5466 18951 5468
rect 19007 5466 19013 5468
rect 18767 5414 18769 5466
rect 18949 5414 18951 5466
rect 18705 5412 18711 5414
rect 18767 5412 18791 5414
rect 18847 5412 18871 5414
rect 18927 5412 18951 5414
rect 19007 5412 19013 5414
rect 18705 5403 19013 5412
rect 16856 4752 16908 4758
rect 16856 4694 16908 4700
rect 15200 4616 15252 4622
rect 15200 4558 15252 4564
rect 15384 4548 15436 4554
rect 15384 4490 15436 4496
rect 14266 4380 14574 4389
rect 14266 4378 14272 4380
rect 14328 4378 14352 4380
rect 14408 4378 14432 4380
rect 14488 4378 14512 4380
rect 14568 4378 14574 4380
rect 14328 4326 14330 4378
rect 14510 4326 14512 4378
rect 14266 4324 14272 4326
rect 14328 4324 14352 4326
rect 14408 4324 14432 4326
rect 14488 4324 14512 4326
rect 14568 4324 14574 4326
rect 14266 4315 14574 4324
rect 14266 3292 14574 3301
rect 14266 3290 14272 3292
rect 14328 3290 14352 3292
rect 14408 3290 14432 3292
rect 14488 3290 14512 3292
rect 14568 3290 14574 3292
rect 14328 3238 14330 3290
rect 14510 3238 14512 3290
rect 14266 3236 14272 3238
rect 14328 3236 14352 3238
rect 14408 3236 14432 3238
rect 14488 3236 14512 3238
rect 14568 3236 14574 3238
rect 14266 3227 14574 3236
rect 13912 3052 13964 3058
rect 13912 2994 13964 3000
rect 13728 2984 13780 2990
rect 13728 2926 13780 2932
rect 12900 2644 12952 2650
rect 12900 2586 12952 2592
rect 13740 2514 13768 2926
rect 15396 2922 15424 4490
rect 16028 4480 16080 4486
rect 16028 4422 16080 4428
rect 16856 4480 16908 4486
rect 16856 4422 16908 4428
rect 16040 3738 16068 4422
rect 16486 3836 16794 3845
rect 16486 3834 16492 3836
rect 16548 3834 16572 3836
rect 16628 3834 16652 3836
rect 16708 3834 16732 3836
rect 16788 3834 16794 3836
rect 16548 3782 16550 3834
rect 16730 3782 16732 3834
rect 16486 3780 16492 3782
rect 16548 3780 16572 3782
rect 16628 3780 16652 3782
rect 16708 3780 16732 3782
rect 16788 3780 16794 3782
rect 16486 3771 16794 3780
rect 16028 3732 16080 3738
rect 16028 3674 16080 3680
rect 16868 2922 16896 4422
rect 18705 4380 19013 4389
rect 18705 4378 18711 4380
rect 18767 4378 18791 4380
rect 18847 4378 18871 4380
rect 18927 4378 18951 4380
rect 19007 4378 19013 4380
rect 18767 4326 18769 4378
rect 18949 4326 18951 4378
rect 18705 4324 18711 4326
rect 18767 4324 18791 4326
rect 18847 4324 18871 4326
rect 18927 4324 18951 4326
rect 19007 4324 19013 4326
rect 18705 4315 19013 4324
rect 18705 3292 19013 3301
rect 18705 3290 18711 3292
rect 18767 3290 18791 3292
rect 18847 3290 18871 3292
rect 18927 3290 18951 3292
rect 19007 3290 19013 3292
rect 18767 3238 18769 3290
rect 18949 3238 18951 3290
rect 18705 3236 18711 3238
rect 18767 3236 18791 3238
rect 18847 3236 18871 3238
rect 18927 3236 18951 3238
rect 19007 3236 19013 3238
rect 18705 3227 19013 3236
rect 15384 2916 15436 2922
rect 15384 2858 15436 2864
rect 15752 2916 15804 2922
rect 15752 2858 15804 2864
rect 16856 2916 16908 2922
rect 16856 2858 16908 2864
rect 13728 2508 13780 2514
rect 13728 2450 13780 2456
rect 15764 2378 15792 2858
rect 16486 2748 16794 2757
rect 16486 2746 16492 2748
rect 16548 2746 16572 2748
rect 16628 2746 16652 2748
rect 16708 2746 16732 2748
rect 16788 2746 16794 2748
rect 16548 2694 16550 2746
rect 16730 2694 16732 2746
rect 16486 2692 16492 2694
rect 16548 2692 16572 2694
rect 16628 2692 16652 2694
rect 16708 2692 16732 2694
rect 16788 2692 16794 2694
rect 16486 2683 16794 2692
rect 17500 2440 17552 2446
rect 17500 2382 17552 2388
rect 15752 2372 15804 2378
rect 15752 2314 15804 2320
rect 12716 2304 12768 2310
rect 12716 2246 12768 2252
rect 17408 2304 17460 2310
rect 17408 2246 17460 2252
rect 14266 2204 14574 2213
rect 14266 2202 14272 2204
rect 14328 2202 14352 2204
rect 14408 2202 14432 2204
rect 14488 2202 14512 2204
rect 14568 2202 14574 2204
rect 14328 2150 14330 2202
rect 14510 2150 14512 2202
rect 14266 2148 14272 2150
rect 14328 2148 14352 2150
rect 14408 2148 14432 2150
rect 14488 2148 14512 2150
rect 14568 2148 14574 2150
rect 14266 2139 14574 2148
rect 17420 800 17448 2246
rect 17512 2106 17540 2382
rect 18705 2204 19013 2213
rect 18705 2202 18711 2204
rect 18767 2202 18791 2204
rect 18847 2202 18871 2204
rect 18927 2202 18951 2204
rect 19007 2202 19013 2204
rect 18767 2150 18769 2202
rect 18949 2150 18951 2202
rect 18705 2148 18711 2150
rect 18767 2148 18791 2150
rect 18847 2148 18871 2150
rect 18927 2148 18951 2150
rect 19007 2148 19013 2150
rect 18705 2139 19013 2148
rect 17500 2100 17552 2106
rect 17500 2042 17552 2048
rect 2502 0 2558 800
rect 7470 0 7526 800
rect 12438 0 12494 800
rect 17406 0 17462 800
<< via2 >>
rect 5394 7642 5450 7644
rect 5474 7642 5530 7644
rect 5554 7642 5610 7644
rect 5634 7642 5690 7644
rect 5394 7590 5440 7642
rect 5440 7590 5450 7642
rect 5474 7590 5504 7642
rect 5504 7590 5516 7642
rect 5516 7590 5530 7642
rect 5554 7590 5568 7642
rect 5568 7590 5580 7642
rect 5580 7590 5610 7642
rect 5634 7590 5644 7642
rect 5644 7590 5690 7642
rect 5394 7588 5450 7590
rect 5474 7588 5530 7590
rect 5554 7588 5610 7590
rect 5634 7588 5690 7590
rect 9833 7642 9889 7644
rect 9913 7642 9969 7644
rect 9993 7642 10049 7644
rect 10073 7642 10129 7644
rect 9833 7590 9879 7642
rect 9879 7590 9889 7642
rect 9913 7590 9943 7642
rect 9943 7590 9955 7642
rect 9955 7590 9969 7642
rect 9993 7590 10007 7642
rect 10007 7590 10019 7642
rect 10019 7590 10049 7642
rect 10073 7590 10083 7642
rect 10083 7590 10129 7642
rect 9833 7588 9889 7590
rect 9913 7588 9969 7590
rect 9993 7588 10049 7590
rect 10073 7588 10129 7590
rect 14272 7642 14328 7644
rect 14352 7642 14408 7644
rect 14432 7642 14488 7644
rect 14512 7642 14568 7644
rect 14272 7590 14318 7642
rect 14318 7590 14328 7642
rect 14352 7590 14382 7642
rect 14382 7590 14394 7642
rect 14394 7590 14408 7642
rect 14432 7590 14446 7642
rect 14446 7590 14458 7642
rect 14458 7590 14488 7642
rect 14512 7590 14522 7642
rect 14522 7590 14568 7642
rect 14272 7588 14328 7590
rect 14352 7588 14408 7590
rect 14432 7588 14488 7590
rect 14512 7588 14568 7590
rect 18711 7642 18767 7644
rect 18791 7642 18847 7644
rect 18871 7642 18927 7644
rect 18951 7642 19007 7644
rect 18711 7590 18757 7642
rect 18757 7590 18767 7642
rect 18791 7590 18821 7642
rect 18821 7590 18833 7642
rect 18833 7590 18847 7642
rect 18871 7590 18885 7642
rect 18885 7590 18897 7642
rect 18897 7590 18927 7642
rect 18951 7590 18961 7642
rect 18961 7590 19007 7642
rect 18711 7588 18767 7590
rect 18791 7588 18847 7590
rect 18871 7588 18927 7590
rect 18951 7588 19007 7590
rect 3175 7098 3231 7100
rect 3255 7098 3311 7100
rect 3335 7098 3391 7100
rect 3415 7098 3471 7100
rect 3175 7046 3221 7098
rect 3221 7046 3231 7098
rect 3255 7046 3285 7098
rect 3285 7046 3297 7098
rect 3297 7046 3311 7098
rect 3335 7046 3349 7098
rect 3349 7046 3361 7098
rect 3361 7046 3391 7098
rect 3415 7046 3425 7098
rect 3425 7046 3471 7098
rect 3175 7044 3231 7046
rect 3255 7044 3311 7046
rect 3335 7044 3391 7046
rect 3415 7044 3471 7046
rect 5394 6554 5450 6556
rect 5474 6554 5530 6556
rect 5554 6554 5610 6556
rect 5634 6554 5690 6556
rect 5394 6502 5440 6554
rect 5440 6502 5450 6554
rect 5474 6502 5504 6554
rect 5504 6502 5516 6554
rect 5516 6502 5530 6554
rect 5554 6502 5568 6554
rect 5568 6502 5580 6554
rect 5580 6502 5610 6554
rect 5634 6502 5644 6554
rect 5644 6502 5690 6554
rect 5394 6500 5450 6502
rect 5474 6500 5530 6502
rect 5554 6500 5610 6502
rect 5634 6500 5690 6502
rect 3175 6010 3231 6012
rect 3255 6010 3311 6012
rect 3335 6010 3391 6012
rect 3415 6010 3471 6012
rect 3175 5958 3221 6010
rect 3221 5958 3231 6010
rect 3255 5958 3285 6010
rect 3285 5958 3297 6010
rect 3297 5958 3311 6010
rect 3335 5958 3349 6010
rect 3349 5958 3361 6010
rect 3361 5958 3391 6010
rect 3415 5958 3425 6010
rect 3425 5958 3471 6010
rect 3175 5956 3231 5958
rect 3255 5956 3311 5958
rect 3335 5956 3391 5958
rect 3415 5956 3471 5958
rect 3175 4922 3231 4924
rect 3255 4922 3311 4924
rect 3335 4922 3391 4924
rect 3415 4922 3471 4924
rect 3175 4870 3221 4922
rect 3221 4870 3231 4922
rect 3255 4870 3285 4922
rect 3285 4870 3297 4922
rect 3297 4870 3311 4922
rect 3335 4870 3349 4922
rect 3349 4870 3361 4922
rect 3361 4870 3391 4922
rect 3415 4870 3425 4922
rect 3425 4870 3471 4922
rect 3175 4868 3231 4870
rect 3255 4868 3311 4870
rect 3335 4868 3391 4870
rect 3415 4868 3471 4870
rect 3175 3834 3231 3836
rect 3255 3834 3311 3836
rect 3335 3834 3391 3836
rect 3415 3834 3471 3836
rect 3175 3782 3221 3834
rect 3221 3782 3231 3834
rect 3255 3782 3285 3834
rect 3285 3782 3297 3834
rect 3297 3782 3311 3834
rect 3335 3782 3349 3834
rect 3349 3782 3361 3834
rect 3361 3782 3391 3834
rect 3415 3782 3425 3834
rect 3425 3782 3471 3834
rect 3175 3780 3231 3782
rect 3255 3780 3311 3782
rect 3335 3780 3391 3782
rect 3415 3780 3471 3782
rect 3175 2746 3231 2748
rect 3255 2746 3311 2748
rect 3335 2746 3391 2748
rect 3415 2746 3471 2748
rect 3175 2694 3221 2746
rect 3221 2694 3231 2746
rect 3255 2694 3285 2746
rect 3285 2694 3297 2746
rect 3297 2694 3311 2746
rect 3335 2694 3349 2746
rect 3349 2694 3361 2746
rect 3361 2694 3391 2746
rect 3415 2694 3425 2746
rect 3425 2694 3471 2746
rect 3175 2692 3231 2694
rect 3255 2692 3311 2694
rect 3335 2692 3391 2694
rect 3415 2692 3471 2694
rect 5394 5466 5450 5468
rect 5474 5466 5530 5468
rect 5554 5466 5610 5468
rect 5634 5466 5690 5468
rect 5394 5414 5440 5466
rect 5440 5414 5450 5466
rect 5474 5414 5504 5466
rect 5504 5414 5516 5466
rect 5516 5414 5530 5466
rect 5554 5414 5568 5466
rect 5568 5414 5580 5466
rect 5580 5414 5610 5466
rect 5634 5414 5644 5466
rect 5644 5414 5690 5466
rect 5394 5412 5450 5414
rect 5474 5412 5530 5414
rect 5554 5412 5610 5414
rect 5634 5412 5690 5414
rect 5394 4378 5450 4380
rect 5474 4378 5530 4380
rect 5554 4378 5610 4380
rect 5634 4378 5690 4380
rect 5394 4326 5440 4378
rect 5440 4326 5450 4378
rect 5474 4326 5504 4378
rect 5504 4326 5516 4378
rect 5516 4326 5530 4378
rect 5554 4326 5568 4378
rect 5568 4326 5580 4378
rect 5580 4326 5610 4378
rect 5634 4326 5644 4378
rect 5644 4326 5690 4378
rect 5394 4324 5450 4326
rect 5474 4324 5530 4326
rect 5554 4324 5610 4326
rect 5634 4324 5690 4326
rect 5394 3290 5450 3292
rect 5474 3290 5530 3292
rect 5554 3290 5610 3292
rect 5634 3290 5690 3292
rect 5394 3238 5440 3290
rect 5440 3238 5450 3290
rect 5474 3238 5504 3290
rect 5504 3238 5516 3290
rect 5516 3238 5530 3290
rect 5554 3238 5568 3290
rect 5568 3238 5580 3290
rect 5580 3238 5610 3290
rect 5634 3238 5644 3290
rect 5644 3238 5690 3290
rect 5394 3236 5450 3238
rect 5474 3236 5530 3238
rect 5554 3236 5610 3238
rect 5634 3236 5690 3238
rect 7614 7098 7670 7100
rect 7694 7098 7750 7100
rect 7774 7098 7830 7100
rect 7854 7098 7910 7100
rect 7614 7046 7660 7098
rect 7660 7046 7670 7098
rect 7694 7046 7724 7098
rect 7724 7046 7736 7098
rect 7736 7046 7750 7098
rect 7774 7046 7788 7098
rect 7788 7046 7800 7098
rect 7800 7046 7830 7098
rect 7854 7046 7864 7098
rect 7864 7046 7910 7098
rect 7614 7044 7670 7046
rect 7694 7044 7750 7046
rect 7774 7044 7830 7046
rect 7854 7044 7910 7046
rect 7614 6010 7670 6012
rect 7694 6010 7750 6012
rect 7774 6010 7830 6012
rect 7854 6010 7910 6012
rect 7614 5958 7660 6010
rect 7660 5958 7670 6010
rect 7694 5958 7724 6010
rect 7724 5958 7736 6010
rect 7736 5958 7750 6010
rect 7774 5958 7788 6010
rect 7788 5958 7800 6010
rect 7800 5958 7830 6010
rect 7854 5958 7864 6010
rect 7864 5958 7910 6010
rect 7614 5956 7670 5958
rect 7694 5956 7750 5958
rect 7774 5956 7830 5958
rect 7854 5956 7910 5958
rect 7614 4922 7670 4924
rect 7694 4922 7750 4924
rect 7774 4922 7830 4924
rect 7854 4922 7910 4924
rect 7614 4870 7660 4922
rect 7660 4870 7670 4922
rect 7694 4870 7724 4922
rect 7724 4870 7736 4922
rect 7736 4870 7750 4922
rect 7774 4870 7788 4922
rect 7788 4870 7800 4922
rect 7800 4870 7830 4922
rect 7854 4870 7864 4922
rect 7864 4870 7910 4922
rect 7614 4868 7670 4870
rect 7694 4868 7750 4870
rect 7774 4868 7830 4870
rect 7854 4868 7910 4870
rect 9833 6554 9889 6556
rect 9913 6554 9969 6556
rect 9993 6554 10049 6556
rect 10073 6554 10129 6556
rect 9833 6502 9879 6554
rect 9879 6502 9889 6554
rect 9913 6502 9943 6554
rect 9943 6502 9955 6554
rect 9955 6502 9969 6554
rect 9993 6502 10007 6554
rect 10007 6502 10019 6554
rect 10019 6502 10049 6554
rect 10073 6502 10083 6554
rect 10083 6502 10129 6554
rect 9833 6500 9889 6502
rect 9913 6500 9969 6502
rect 9993 6500 10049 6502
rect 10073 6500 10129 6502
rect 7614 3834 7670 3836
rect 7694 3834 7750 3836
rect 7774 3834 7830 3836
rect 7854 3834 7910 3836
rect 7614 3782 7660 3834
rect 7660 3782 7670 3834
rect 7694 3782 7724 3834
rect 7724 3782 7736 3834
rect 7736 3782 7750 3834
rect 7774 3782 7788 3834
rect 7788 3782 7800 3834
rect 7800 3782 7830 3834
rect 7854 3782 7864 3834
rect 7864 3782 7910 3834
rect 7614 3780 7670 3782
rect 7694 3780 7750 3782
rect 7774 3780 7830 3782
rect 7854 3780 7910 3782
rect 7378 3304 7434 3360
rect 7102 3032 7158 3088
rect 5394 2202 5450 2204
rect 5474 2202 5530 2204
rect 5554 2202 5610 2204
rect 5634 2202 5690 2204
rect 5394 2150 5440 2202
rect 5440 2150 5450 2202
rect 5474 2150 5504 2202
rect 5504 2150 5516 2202
rect 5516 2150 5530 2202
rect 5554 2150 5568 2202
rect 5568 2150 5580 2202
rect 5580 2150 5610 2202
rect 5634 2150 5644 2202
rect 5644 2150 5690 2202
rect 5394 2148 5450 2150
rect 5474 2148 5530 2150
rect 5554 2148 5610 2150
rect 5634 2148 5690 2150
rect 7614 2746 7670 2748
rect 7694 2746 7750 2748
rect 7774 2746 7830 2748
rect 7854 2746 7910 2748
rect 7614 2694 7660 2746
rect 7660 2694 7670 2746
rect 7694 2694 7724 2746
rect 7724 2694 7736 2746
rect 7736 2694 7750 2746
rect 7774 2694 7788 2746
rect 7788 2694 7800 2746
rect 7800 2694 7830 2746
rect 7854 2694 7864 2746
rect 7864 2694 7910 2746
rect 7614 2692 7670 2694
rect 7694 2692 7750 2694
rect 7774 2692 7830 2694
rect 7854 2692 7910 2694
rect 9833 5466 9889 5468
rect 9913 5466 9969 5468
rect 9993 5466 10049 5468
rect 10073 5466 10129 5468
rect 9833 5414 9879 5466
rect 9879 5414 9889 5466
rect 9913 5414 9943 5466
rect 9943 5414 9955 5466
rect 9955 5414 9969 5466
rect 9993 5414 10007 5466
rect 10007 5414 10019 5466
rect 10019 5414 10049 5466
rect 10073 5414 10083 5466
rect 10083 5414 10129 5466
rect 9833 5412 9889 5414
rect 9913 5412 9969 5414
rect 9993 5412 10049 5414
rect 10073 5412 10129 5414
rect 8298 3304 8354 3360
rect 9034 3052 9090 3088
rect 9034 3032 9036 3052
rect 9036 3032 9088 3052
rect 9088 3032 9090 3052
rect 12053 7098 12109 7100
rect 12133 7098 12189 7100
rect 12213 7098 12269 7100
rect 12293 7098 12349 7100
rect 12053 7046 12099 7098
rect 12099 7046 12109 7098
rect 12133 7046 12163 7098
rect 12163 7046 12175 7098
rect 12175 7046 12189 7098
rect 12213 7046 12227 7098
rect 12227 7046 12239 7098
rect 12239 7046 12269 7098
rect 12293 7046 12303 7098
rect 12303 7046 12349 7098
rect 12053 7044 12109 7046
rect 12133 7044 12189 7046
rect 12213 7044 12269 7046
rect 12293 7044 12349 7046
rect 12053 6010 12109 6012
rect 12133 6010 12189 6012
rect 12213 6010 12269 6012
rect 12293 6010 12349 6012
rect 12053 5958 12099 6010
rect 12099 5958 12109 6010
rect 12133 5958 12163 6010
rect 12163 5958 12175 6010
rect 12175 5958 12189 6010
rect 12213 5958 12227 6010
rect 12227 5958 12239 6010
rect 12239 5958 12269 6010
rect 12293 5958 12303 6010
rect 12303 5958 12349 6010
rect 12053 5956 12109 5958
rect 12133 5956 12189 5958
rect 12213 5956 12269 5958
rect 12293 5956 12349 5958
rect 9833 4378 9889 4380
rect 9913 4378 9969 4380
rect 9993 4378 10049 4380
rect 10073 4378 10129 4380
rect 9833 4326 9879 4378
rect 9879 4326 9889 4378
rect 9913 4326 9943 4378
rect 9943 4326 9955 4378
rect 9955 4326 9969 4378
rect 9993 4326 10007 4378
rect 10007 4326 10019 4378
rect 10019 4326 10049 4378
rect 10073 4326 10083 4378
rect 10083 4326 10129 4378
rect 9833 4324 9889 4326
rect 9913 4324 9969 4326
rect 9993 4324 10049 4326
rect 10073 4324 10129 4326
rect 9833 3290 9889 3292
rect 9913 3290 9969 3292
rect 9993 3290 10049 3292
rect 10073 3290 10129 3292
rect 9833 3238 9879 3290
rect 9879 3238 9889 3290
rect 9913 3238 9943 3290
rect 9943 3238 9955 3290
rect 9955 3238 9969 3290
rect 9993 3238 10007 3290
rect 10007 3238 10019 3290
rect 10019 3238 10049 3290
rect 10073 3238 10083 3290
rect 10083 3238 10129 3290
rect 9833 3236 9889 3238
rect 9913 3236 9969 3238
rect 9993 3236 10049 3238
rect 10073 3236 10129 3238
rect 12053 4922 12109 4924
rect 12133 4922 12189 4924
rect 12213 4922 12269 4924
rect 12293 4922 12349 4924
rect 12053 4870 12099 4922
rect 12099 4870 12109 4922
rect 12133 4870 12163 4922
rect 12163 4870 12175 4922
rect 12175 4870 12189 4922
rect 12213 4870 12227 4922
rect 12227 4870 12239 4922
rect 12239 4870 12269 4922
rect 12293 4870 12303 4922
rect 12303 4870 12349 4922
rect 12053 4868 12109 4870
rect 12133 4868 12189 4870
rect 12213 4868 12269 4870
rect 12293 4868 12349 4870
rect 11886 3984 11942 4040
rect 12053 3834 12109 3836
rect 12133 3834 12189 3836
rect 12213 3834 12269 3836
rect 12293 3834 12349 3836
rect 12053 3782 12099 3834
rect 12099 3782 12109 3834
rect 12133 3782 12163 3834
rect 12163 3782 12175 3834
rect 12175 3782 12189 3834
rect 12213 3782 12227 3834
rect 12227 3782 12239 3834
rect 12239 3782 12269 3834
rect 12293 3782 12303 3834
rect 12303 3782 12349 3834
rect 12053 3780 12109 3782
rect 12133 3780 12189 3782
rect 12213 3780 12269 3782
rect 12293 3780 12349 3782
rect 9833 2202 9889 2204
rect 9913 2202 9969 2204
rect 9993 2202 10049 2204
rect 10073 2202 10129 2204
rect 9833 2150 9879 2202
rect 9879 2150 9889 2202
rect 9913 2150 9943 2202
rect 9943 2150 9955 2202
rect 9955 2150 9969 2202
rect 9993 2150 10007 2202
rect 10007 2150 10019 2202
rect 10019 2150 10049 2202
rect 10073 2150 10083 2202
rect 10083 2150 10129 2202
rect 9833 2148 9889 2150
rect 9913 2148 9969 2150
rect 9993 2148 10049 2150
rect 10073 2148 10129 2150
rect 16492 7098 16548 7100
rect 16572 7098 16628 7100
rect 16652 7098 16708 7100
rect 16732 7098 16788 7100
rect 16492 7046 16538 7098
rect 16538 7046 16548 7098
rect 16572 7046 16602 7098
rect 16602 7046 16614 7098
rect 16614 7046 16628 7098
rect 16652 7046 16666 7098
rect 16666 7046 16678 7098
rect 16678 7046 16708 7098
rect 16732 7046 16742 7098
rect 16742 7046 16788 7098
rect 16492 7044 16548 7046
rect 16572 7044 16628 7046
rect 16652 7044 16708 7046
rect 16732 7044 16788 7046
rect 14272 6554 14328 6556
rect 14352 6554 14408 6556
rect 14432 6554 14488 6556
rect 14512 6554 14568 6556
rect 14272 6502 14318 6554
rect 14318 6502 14328 6554
rect 14352 6502 14382 6554
rect 14382 6502 14394 6554
rect 14394 6502 14408 6554
rect 14432 6502 14446 6554
rect 14446 6502 14458 6554
rect 14458 6502 14488 6554
rect 14512 6502 14522 6554
rect 14522 6502 14568 6554
rect 14272 6500 14328 6502
rect 14352 6500 14408 6502
rect 14432 6500 14488 6502
rect 14512 6500 14568 6502
rect 16492 6010 16548 6012
rect 16572 6010 16628 6012
rect 16652 6010 16708 6012
rect 16732 6010 16788 6012
rect 16492 5958 16538 6010
rect 16538 5958 16548 6010
rect 16572 5958 16602 6010
rect 16602 5958 16614 6010
rect 16614 5958 16628 6010
rect 16652 5958 16666 6010
rect 16666 5958 16678 6010
rect 16678 5958 16708 6010
rect 16732 5958 16742 6010
rect 16742 5958 16788 6010
rect 16492 5956 16548 5958
rect 16572 5956 16628 5958
rect 16652 5956 16708 5958
rect 16732 5956 16788 5958
rect 14272 5466 14328 5468
rect 14352 5466 14408 5468
rect 14432 5466 14488 5468
rect 14512 5466 14568 5468
rect 14272 5414 14318 5466
rect 14318 5414 14328 5466
rect 14352 5414 14382 5466
rect 14382 5414 14394 5466
rect 14394 5414 14408 5466
rect 14432 5414 14446 5466
rect 14446 5414 14458 5466
rect 14458 5414 14488 5466
rect 14512 5414 14522 5466
rect 14522 5414 14568 5466
rect 14272 5412 14328 5414
rect 14352 5412 14408 5414
rect 14432 5412 14488 5414
rect 14512 5412 14568 5414
rect 13082 3984 13138 4040
rect 12053 2746 12109 2748
rect 12133 2746 12189 2748
rect 12213 2746 12269 2748
rect 12293 2746 12349 2748
rect 12053 2694 12099 2746
rect 12099 2694 12109 2746
rect 12133 2694 12163 2746
rect 12163 2694 12175 2746
rect 12175 2694 12189 2746
rect 12213 2694 12227 2746
rect 12227 2694 12239 2746
rect 12239 2694 12269 2746
rect 12293 2694 12303 2746
rect 12303 2694 12349 2746
rect 12053 2692 12109 2694
rect 12133 2692 12189 2694
rect 12213 2692 12269 2694
rect 12293 2692 12349 2694
rect 16492 4922 16548 4924
rect 16572 4922 16628 4924
rect 16652 4922 16708 4924
rect 16732 4922 16788 4924
rect 16492 4870 16538 4922
rect 16538 4870 16548 4922
rect 16572 4870 16602 4922
rect 16602 4870 16614 4922
rect 16614 4870 16628 4922
rect 16652 4870 16666 4922
rect 16666 4870 16678 4922
rect 16678 4870 16708 4922
rect 16732 4870 16742 4922
rect 16742 4870 16788 4922
rect 16492 4868 16548 4870
rect 16572 4868 16628 4870
rect 16652 4868 16708 4870
rect 16732 4868 16788 4870
rect 18711 6554 18767 6556
rect 18791 6554 18847 6556
rect 18871 6554 18927 6556
rect 18951 6554 19007 6556
rect 18711 6502 18757 6554
rect 18757 6502 18767 6554
rect 18791 6502 18821 6554
rect 18821 6502 18833 6554
rect 18833 6502 18847 6554
rect 18871 6502 18885 6554
rect 18885 6502 18897 6554
rect 18897 6502 18927 6554
rect 18951 6502 18961 6554
rect 18961 6502 19007 6554
rect 18711 6500 18767 6502
rect 18791 6500 18847 6502
rect 18871 6500 18927 6502
rect 18951 6500 19007 6502
rect 18711 5466 18767 5468
rect 18791 5466 18847 5468
rect 18871 5466 18927 5468
rect 18951 5466 19007 5468
rect 18711 5414 18757 5466
rect 18757 5414 18767 5466
rect 18791 5414 18821 5466
rect 18821 5414 18833 5466
rect 18833 5414 18847 5466
rect 18871 5414 18885 5466
rect 18885 5414 18897 5466
rect 18897 5414 18927 5466
rect 18951 5414 18961 5466
rect 18961 5414 19007 5466
rect 18711 5412 18767 5414
rect 18791 5412 18847 5414
rect 18871 5412 18927 5414
rect 18951 5412 19007 5414
rect 14272 4378 14328 4380
rect 14352 4378 14408 4380
rect 14432 4378 14488 4380
rect 14512 4378 14568 4380
rect 14272 4326 14318 4378
rect 14318 4326 14328 4378
rect 14352 4326 14382 4378
rect 14382 4326 14394 4378
rect 14394 4326 14408 4378
rect 14432 4326 14446 4378
rect 14446 4326 14458 4378
rect 14458 4326 14488 4378
rect 14512 4326 14522 4378
rect 14522 4326 14568 4378
rect 14272 4324 14328 4326
rect 14352 4324 14408 4326
rect 14432 4324 14488 4326
rect 14512 4324 14568 4326
rect 14272 3290 14328 3292
rect 14352 3290 14408 3292
rect 14432 3290 14488 3292
rect 14512 3290 14568 3292
rect 14272 3238 14318 3290
rect 14318 3238 14328 3290
rect 14352 3238 14382 3290
rect 14382 3238 14394 3290
rect 14394 3238 14408 3290
rect 14432 3238 14446 3290
rect 14446 3238 14458 3290
rect 14458 3238 14488 3290
rect 14512 3238 14522 3290
rect 14522 3238 14568 3290
rect 14272 3236 14328 3238
rect 14352 3236 14408 3238
rect 14432 3236 14488 3238
rect 14512 3236 14568 3238
rect 16492 3834 16548 3836
rect 16572 3834 16628 3836
rect 16652 3834 16708 3836
rect 16732 3834 16788 3836
rect 16492 3782 16538 3834
rect 16538 3782 16548 3834
rect 16572 3782 16602 3834
rect 16602 3782 16614 3834
rect 16614 3782 16628 3834
rect 16652 3782 16666 3834
rect 16666 3782 16678 3834
rect 16678 3782 16708 3834
rect 16732 3782 16742 3834
rect 16742 3782 16788 3834
rect 16492 3780 16548 3782
rect 16572 3780 16628 3782
rect 16652 3780 16708 3782
rect 16732 3780 16788 3782
rect 18711 4378 18767 4380
rect 18791 4378 18847 4380
rect 18871 4378 18927 4380
rect 18951 4378 19007 4380
rect 18711 4326 18757 4378
rect 18757 4326 18767 4378
rect 18791 4326 18821 4378
rect 18821 4326 18833 4378
rect 18833 4326 18847 4378
rect 18871 4326 18885 4378
rect 18885 4326 18897 4378
rect 18897 4326 18927 4378
rect 18951 4326 18961 4378
rect 18961 4326 19007 4378
rect 18711 4324 18767 4326
rect 18791 4324 18847 4326
rect 18871 4324 18927 4326
rect 18951 4324 19007 4326
rect 18711 3290 18767 3292
rect 18791 3290 18847 3292
rect 18871 3290 18927 3292
rect 18951 3290 19007 3292
rect 18711 3238 18757 3290
rect 18757 3238 18767 3290
rect 18791 3238 18821 3290
rect 18821 3238 18833 3290
rect 18833 3238 18847 3290
rect 18871 3238 18885 3290
rect 18885 3238 18897 3290
rect 18897 3238 18927 3290
rect 18951 3238 18961 3290
rect 18961 3238 19007 3290
rect 18711 3236 18767 3238
rect 18791 3236 18847 3238
rect 18871 3236 18927 3238
rect 18951 3236 19007 3238
rect 16492 2746 16548 2748
rect 16572 2746 16628 2748
rect 16652 2746 16708 2748
rect 16732 2746 16788 2748
rect 16492 2694 16538 2746
rect 16538 2694 16548 2746
rect 16572 2694 16602 2746
rect 16602 2694 16614 2746
rect 16614 2694 16628 2746
rect 16652 2694 16666 2746
rect 16666 2694 16678 2746
rect 16678 2694 16708 2746
rect 16732 2694 16742 2746
rect 16742 2694 16788 2746
rect 16492 2692 16548 2694
rect 16572 2692 16628 2694
rect 16652 2692 16708 2694
rect 16732 2692 16788 2694
rect 14272 2202 14328 2204
rect 14352 2202 14408 2204
rect 14432 2202 14488 2204
rect 14512 2202 14568 2204
rect 14272 2150 14318 2202
rect 14318 2150 14328 2202
rect 14352 2150 14382 2202
rect 14382 2150 14394 2202
rect 14394 2150 14408 2202
rect 14432 2150 14446 2202
rect 14446 2150 14458 2202
rect 14458 2150 14488 2202
rect 14512 2150 14522 2202
rect 14522 2150 14568 2202
rect 14272 2148 14328 2150
rect 14352 2148 14408 2150
rect 14432 2148 14488 2150
rect 14512 2148 14568 2150
rect 18711 2202 18767 2204
rect 18791 2202 18847 2204
rect 18871 2202 18927 2204
rect 18951 2202 19007 2204
rect 18711 2150 18757 2202
rect 18757 2150 18767 2202
rect 18791 2150 18821 2202
rect 18821 2150 18833 2202
rect 18833 2150 18847 2202
rect 18871 2150 18885 2202
rect 18885 2150 18897 2202
rect 18897 2150 18927 2202
rect 18951 2150 18961 2202
rect 18961 2150 19007 2202
rect 18711 2148 18767 2150
rect 18791 2148 18847 2150
rect 18871 2148 18927 2150
rect 18951 2148 19007 2150
<< metal3 >>
rect 5384 7648 5700 7649
rect 5384 7584 5390 7648
rect 5454 7584 5470 7648
rect 5534 7584 5550 7648
rect 5614 7584 5630 7648
rect 5694 7584 5700 7648
rect 5384 7583 5700 7584
rect 9823 7648 10139 7649
rect 9823 7584 9829 7648
rect 9893 7584 9909 7648
rect 9973 7584 9989 7648
rect 10053 7584 10069 7648
rect 10133 7584 10139 7648
rect 9823 7583 10139 7584
rect 14262 7648 14578 7649
rect 14262 7584 14268 7648
rect 14332 7584 14348 7648
rect 14412 7584 14428 7648
rect 14492 7584 14508 7648
rect 14572 7584 14578 7648
rect 14262 7583 14578 7584
rect 18701 7648 19017 7649
rect 18701 7584 18707 7648
rect 18771 7584 18787 7648
rect 18851 7584 18867 7648
rect 18931 7584 18947 7648
rect 19011 7584 19017 7648
rect 18701 7583 19017 7584
rect 3165 7104 3481 7105
rect 3165 7040 3171 7104
rect 3235 7040 3251 7104
rect 3315 7040 3331 7104
rect 3395 7040 3411 7104
rect 3475 7040 3481 7104
rect 3165 7039 3481 7040
rect 7604 7104 7920 7105
rect 7604 7040 7610 7104
rect 7674 7040 7690 7104
rect 7754 7040 7770 7104
rect 7834 7040 7850 7104
rect 7914 7040 7920 7104
rect 7604 7039 7920 7040
rect 12043 7104 12359 7105
rect 12043 7040 12049 7104
rect 12113 7040 12129 7104
rect 12193 7040 12209 7104
rect 12273 7040 12289 7104
rect 12353 7040 12359 7104
rect 12043 7039 12359 7040
rect 16482 7104 16798 7105
rect 16482 7040 16488 7104
rect 16552 7040 16568 7104
rect 16632 7040 16648 7104
rect 16712 7040 16728 7104
rect 16792 7040 16798 7104
rect 16482 7039 16798 7040
rect 5384 6560 5700 6561
rect 5384 6496 5390 6560
rect 5454 6496 5470 6560
rect 5534 6496 5550 6560
rect 5614 6496 5630 6560
rect 5694 6496 5700 6560
rect 5384 6495 5700 6496
rect 9823 6560 10139 6561
rect 9823 6496 9829 6560
rect 9893 6496 9909 6560
rect 9973 6496 9989 6560
rect 10053 6496 10069 6560
rect 10133 6496 10139 6560
rect 9823 6495 10139 6496
rect 14262 6560 14578 6561
rect 14262 6496 14268 6560
rect 14332 6496 14348 6560
rect 14412 6496 14428 6560
rect 14492 6496 14508 6560
rect 14572 6496 14578 6560
rect 14262 6495 14578 6496
rect 18701 6560 19017 6561
rect 18701 6496 18707 6560
rect 18771 6496 18787 6560
rect 18851 6496 18867 6560
rect 18931 6496 18947 6560
rect 19011 6496 19017 6560
rect 18701 6495 19017 6496
rect 3165 6016 3481 6017
rect 3165 5952 3171 6016
rect 3235 5952 3251 6016
rect 3315 5952 3331 6016
rect 3395 5952 3411 6016
rect 3475 5952 3481 6016
rect 3165 5951 3481 5952
rect 7604 6016 7920 6017
rect 7604 5952 7610 6016
rect 7674 5952 7690 6016
rect 7754 5952 7770 6016
rect 7834 5952 7850 6016
rect 7914 5952 7920 6016
rect 7604 5951 7920 5952
rect 12043 6016 12359 6017
rect 12043 5952 12049 6016
rect 12113 5952 12129 6016
rect 12193 5952 12209 6016
rect 12273 5952 12289 6016
rect 12353 5952 12359 6016
rect 12043 5951 12359 5952
rect 16482 6016 16798 6017
rect 16482 5952 16488 6016
rect 16552 5952 16568 6016
rect 16632 5952 16648 6016
rect 16712 5952 16728 6016
rect 16792 5952 16798 6016
rect 16482 5951 16798 5952
rect 5384 5472 5700 5473
rect 5384 5408 5390 5472
rect 5454 5408 5470 5472
rect 5534 5408 5550 5472
rect 5614 5408 5630 5472
rect 5694 5408 5700 5472
rect 5384 5407 5700 5408
rect 9823 5472 10139 5473
rect 9823 5408 9829 5472
rect 9893 5408 9909 5472
rect 9973 5408 9989 5472
rect 10053 5408 10069 5472
rect 10133 5408 10139 5472
rect 9823 5407 10139 5408
rect 14262 5472 14578 5473
rect 14262 5408 14268 5472
rect 14332 5408 14348 5472
rect 14412 5408 14428 5472
rect 14492 5408 14508 5472
rect 14572 5408 14578 5472
rect 14262 5407 14578 5408
rect 18701 5472 19017 5473
rect 18701 5408 18707 5472
rect 18771 5408 18787 5472
rect 18851 5408 18867 5472
rect 18931 5408 18947 5472
rect 19011 5408 19017 5472
rect 18701 5407 19017 5408
rect 3165 4928 3481 4929
rect 3165 4864 3171 4928
rect 3235 4864 3251 4928
rect 3315 4864 3331 4928
rect 3395 4864 3411 4928
rect 3475 4864 3481 4928
rect 3165 4863 3481 4864
rect 7604 4928 7920 4929
rect 7604 4864 7610 4928
rect 7674 4864 7690 4928
rect 7754 4864 7770 4928
rect 7834 4864 7850 4928
rect 7914 4864 7920 4928
rect 7604 4863 7920 4864
rect 12043 4928 12359 4929
rect 12043 4864 12049 4928
rect 12113 4864 12129 4928
rect 12193 4864 12209 4928
rect 12273 4864 12289 4928
rect 12353 4864 12359 4928
rect 12043 4863 12359 4864
rect 16482 4928 16798 4929
rect 16482 4864 16488 4928
rect 16552 4864 16568 4928
rect 16632 4864 16648 4928
rect 16712 4864 16728 4928
rect 16792 4864 16798 4928
rect 16482 4863 16798 4864
rect 5384 4384 5700 4385
rect 5384 4320 5390 4384
rect 5454 4320 5470 4384
rect 5534 4320 5550 4384
rect 5614 4320 5630 4384
rect 5694 4320 5700 4384
rect 5384 4319 5700 4320
rect 9823 4384 10139 4385
rect 9823 4320 9829 4384
rect 9893 4320 9909 4384
rect 9973 4320 9989 4384
rect 10053 4320 10069 4384
rect 10133 4320 10139 4384
rect 9823 4319 10139 4320
rect 14262 4384 14578 4385
rect 14262 4320 14268 4384
rect 14332 4320 14348 4384
rect 14412 4320 14428 4384
rect 14492 4320 14508 4384
rect 14572 4320 14578 4384
rect 14262 4319 14578 4320
rect 18701 4384 19017 4385
rect 18701 4320 18707 4384
rect 18771 4320 18787 4384
rect 18851 4320 18867 4384
rect 18931 4320 18947 4384
rect 19011 4320 19017 4384
rect 18701 4319 19017 4320
rect 11881 4042 11947 4045
rect 13077 4042 13143 4045
rect 11881 4040 13143 4042
rect 11881 3984 11886 4040
rect 11942 3984 13082 4040
rect 13138 3984 13143 4040
rect 11881 3982 13143 3984
rect 11881 3979 11947 3982
rect 13077 3979 13143 3982
rect 3165 3840 3481 3841
rect 3165 3776 3171 3840
rect 3235 3776 3251 3840
rect 3315 3776 3331 3840
rect 3395 3776 3411 3840
rect 3475 3776 3481 3840
rect 3165 3775 3481 3776
rect 7604 3840 7920 3841
rect 7604 3776 7610 3840
rect 7674 3776 7690 3840
rect 7754 3776 7770 3840
rect 7834 3776 7850 3840
rect 7914 3776 7920 3840
rect 7604 3775 7920 3776
rect 12043 3840 12359 3841
rect 12043 3776 12049 3840
rect 12113 3776 12129 3840
rect 12193 3776 12209 3840
rect 12273 3776 12289 3840
rect 12353 3776 12359 3840
rect 12043 3775 12359 3776
rect 16482 3840 16798 3841
rect 16482 3776 16488 3840
rect 16552 3776 16568 3840
rect 16632 3776 16648 3840
rect 16712 3776 16728 3840
rect 16792 3776 16798 3840
rect 16482 3775 16798 3776
rect 7373 3362 7439 3365
rect 8293 3362 8359 3365
rect 7373 3360 8359 3362
rect 7373 3304 7378 3360
rect 7434 3304 8298 3360
rect 8354 3304 8359 3360
rect 7373 3302 8359 3304
rect 7373 3299 7439 3302
rect 8293 3299 8359 3302
rect 5384 3296 5700 3297
rect 5384 3232 5390 3296
rect 5454 3232 5470 3296
rect 5534 3232 5550 3296
rect 5614 3232 5630 3296
rect 5694 3232 5700 3296
rect 5384 3231 5700 3232
rect 9823 3296 10139 3297
rect 9823 3232 9829 3296
rect 9893 3232 9909 3296
rect 9973 3232 9989 3296
rect 10053 3232 10069 3296
rect 10133 3232 10139 3296
rect 9823 3231 10139 3232
rect 14262 3296 14578 3297
rect 14262 3232 14268 3296
rect 14332 3232 14348 3296
rect 14412 3232 14428 3296
rect 14492 3232 14508 3296
rect 14572 3232 14578 3296
rect 14262 3231 14578 3232
rect 18701 3296 19017 3297
rect 18701 3232 18707 3296
rect 18771 3232 18787 3296
rect 18851 3232 18867 3296
rect 18931 3232 18947 3296
rect 19011 3232 19017 3296
rect 18701 3231 19017 3232
rect 7097 3090 7163 3093
rect 9029 3090 9095 3093
rect 7097 3088 9095 3090
rect 7097 3032 7102 3088
rect 7158 3032 9034 3088
rect 9090 3032 9095 3088
rect 7097 3030 9095 3032
rect 7097 3027 7163 3030
rect 9029 3027 9095 3030
rect 3165 2752 3481 2753
rect 3165 2688 3171 2752
rect 3235 2688 3251 2752
rect 3315 2688 3331 2752
rect 3395 2688 3411 2752
rect 3475 2688 3481 2752
rect 3165 2687 3481 2688
rect 7604 2752 7920 2753
rect 7604 2688 7610 2752
rect 7674 2688 7690 2752
rect 7754 2688 7770 2752
rect 7834 2688 7850 2752
rect 7914 2688 7920 2752
rect 7604 2687 7920 2688
rect 12043 2752 12359 2753
rect 12043 2688 12049 2752
rect 12113 2688 12129 2752
rect 12193 2688 12209 2752
rect 12273 2688 12289 2752
rect 12353 2688 12359 2752
rect 12043 2687 12359 2688
rect 16482 2752 16798 2753
rect 16482 2688 16488 2752
rect 16552 2688 16568 2752
rect 16632 2688 16648 2752
rect 16712 2688 16728 2752
rect 16792 2688 16798 2752
rect 16482 2687 16798 2688
rect 5384 2208 5700 2209
rect 5384 2144 5390 2208
rect 5454 2144 5470 2208
rect 5534 2144 5550 2208
rect 5614 2144 5630 2208
rect 5694 2144 5700 2208
rect 5384 2143 5700 2144
rect 9823 2208 10139 2209
rect 9823 2144 9829 2208
rect 9893 2144 9909 2208
rect 9973 2144 9989 2208
rect 10053 2144 10069 2208
rect 10133 2144 10139 2208
rect 9823 2143 10139 2144
rect 14262 2208 14578 2209
rect 14262 2144 14268 2208
rect 14332 2144 14348 2208
rect 14412 2144 14428 2208
rect 14492 2144 14508 2208
rect 14572 2144 14578 2208
rect 14262 2143 14578 2144
rect 18701 2208 19017 2209
rect 18701 2144 18707 2208
rect 18771 2144 18787 2208
rect 18851 2144 18867 2208
rect 18931 2144 18947 2208
rect 19011 2144 19017 2208
rect 18701 2143 19017 2144
<< via3 >>
rect 5390 7644 5454 7648
rect 5390 7588 5394 7644
rect 5394 7588 5450 7644
rect 5450 7588 5454 7644
rect 5390 7584 5454 7588
rect 5470 7644 5534 7648
rect 5470 7588 5474 7644
rect 5474 7588 5530 7644
rect 5530 7588 5534 7644
rect 5470 7584 5534 7588
rect 5550 7644 5614 7648
rect 5550 7588 5554 7644
rect 5554 7588 5610 7644
rect 5610 7588 5614 7644
rect 5550 7584 5614 7588
rect 5630 7644 5694 7648
rect 5630 7588 5634 7644
rect 5634 7588 5690 7644
rect 5690 7588 5694 7644
rect 5630 7584 5694 7588
rect 9829 7644 9893 7648
rect 9829 7588 9833 7644
rect 9833 7588 9889 7644
rect 9889 7588 9893 7644
rect 9829 7584 9893 7588
rect 9909 7644 9973 7648
rect 9909 7588 9913 7644
rect 9913 7588 9969 7644
rect 9969 7588 9973 7644
rect 9909 7584 9973 7588
rect 9989 7644 10053 7648
rect 9989 7588 9993 7644
rect 9993 7588 10049 7644
rect 10049 7588 10053 7644
rect 9989 7584 10053 7588
rect 10069 7644 10133 7648
rect 10069 7588 10073 7644
rect 10073 7588 10129 7644
rect 10129 7588 10133 7644
rect 10069 7584 10133 7588
rect 14268 7644 14332 7648
rect 14268 7588 14272 7644
rect 14272 7588 14328 7644
rect 14328 7588 14332 7644
rect 14268 7584 14332 7588
rect 14348 7644 14412 7648
rect 14348 7588 14352 7644
rect 14352 7588 14408 7644
rect 14408 7588 14412 7644
rect 14348 7584 14412 7588
rect 14428 7644 14492 7648
rect 14428 7588 14432 7644
rect 14432 7588 14488 7644
rect 14488 7588 14492 7644
rect 14428 7584 14492 7588
rect 14508 7644 14572 7648
rect 14508 7588 14512 7644
rect 14512 7588 14568 7644
rect 14568 7588 14572 7644
rect 14508 7584 14572 7588
rect 18707 7644 18771 7648
rect 18707 7588 18711 7644
rect 18711 7588 18767 7644
rect 18767 7588 18771 7644
rect 18707 7584 18771 7588
rect 18787 7644 18851 7648
rect 18787 7588 18791 7644
rect 18791 7588 18847 7644
rect 18847 7588 18851 7644
rect 18787 7584 18851 7588
rect 18867 7644 18931 7648
rect 18867 7588 18871 7644
rect 18871 7588 18927 7644
rect 18927 7588 18931 7644
rect 18867 7584 18931 7588
rect 18947 7644 19011 7648
rect 18947 7588 18951 7644
rect 18951 7588 19007 7644
rect 19007 7588 19011 7644
rect 18947 7584 19011 7588
rect 3171 7100 3235 7104
rect 3171 7044 3175 7100
rect 3175 7044 3231 7100
rect 3231 7044 3235 7100
rect 3171 7040 3235 7044
rect 3251 7100 3315 7104
rect 3251 7044 3255 7100
rect 3255 7044 3311 7100
rect 3311 7044 3315 7100
rect 3251 7040 3315 7044
rect 3331 7100 3395 7104
rect 3331 7044 3335 7100
rect 3335 7044 3391 7100
rect 3391 7044 3395 7100
rect 3331 7040 3395 7044
rect 3411 7100 3475 7104
rect 3411 7044 3415 7100
rect 3415 7044 3471 7100
rect 3471 7044 3475 7100
rect 3411 7040 3475 7044
rect 7610 7100 7674 7104
rect 7610 7044 7614 7100
rect 7614 7044 7670 7100
rect 7670 7044 7674 7100
rect 7610 7040 7674 7044
rect 7690 7100 7754 7104
rect 7690 7044 7694 7100
rect 7694 7044 7750 7100
rect 7750 7044 7754 7100
rect 7690 7040 7754 7044
rect 7770 7100 7834 7104
rect 7770 7044 7774 7100
rect 7774 7044 7830 7100
rect 7830 7044 7834 7100
rect 7770 7040 7834 7044
rect 7850 7100 7914 7104
rect 7850 7044 7854 7100
rect 7854 7044 7910 7100
rect 7910 7044 7914 7100
rect 7850 7040 7914 7044
rect 12049 7100 12113 7104
rect 12049 7044 12053 7100
rect 12053 7044 12109 7100
rect 12109 7044 12113 7100
rect 12049 7040 12113 7044
rect 12129 7100 12193 7104
rect 12129 7044 12133 7100
rect 12133 7044 12189 7100
rect 12189 7044 12193 7100
rect 12129 7040 12193 7044
rect 12209 7100 12273 7104
rect 12209 7044 12213 7100
rect 12213 7044 12269 7100
rect 12269 7044 12273 7100
rect 12209 7040 12273 7044
rect 12289 7100 12353 7104
rect 12289 7044 12293 7100
rect 12293 7044 12349 7100
rect 12349 7044 12353 7100
rect 12289 7040 12353 7044
rect 16488 7100 16552 7104
rect 16488 7044 16492 7100
rect 16492 7044 16548 7100
rect 16548 7044 16552 7100
rect 16488 7040 16552 7044
rect 16568 7100 16632 7104
rect 16568 7044 16572 7100
rect 16572 7044 16628 7100
rect 16628 7044 16632 7100
rect 16568 7040 16632 7044
rect 16648 7100 16712 7104
rect 16648 7044 16652 7100
rect 16652 7044 16708 7100
rect 16708 7044 16712 7100
rect 16648 7040 16712 7044
rect 16728 7100 16792 7104
rect 16728 7044 16732 7100
rect 16732 7044 16788 7100
rect 16788 7044 16792 7100
rect 16728 7040 16792 7044
rect 5390 6556 5454 6560
rect 5390 6500 5394 6556
rect 5394 6500 5450 6556
rect 5450 6500 5454 6556
rect 5390 6496 5454 6500
rect 5470 6556 5534 6560
rect 5470 6500 5474 6556
rect 5474 6500 5530 6556
rect 5530 6500 5534 6556
rect 5470 6496 5534 6500
rect 5550 6556 5614 6560
rect 5550 6500 5554 6556
rect 5554 6500 5610 6556
rect 5610 6500 5614 6556
rect 5550 6496 5614 6500
rect 5630 6556 5694 6560
rect 5630 6500 5634 6556
rect 5634 6500 5690 6556
rect 5690 6500 5694 6556
rect 5630 6496 5694 6500
rect 9829 6556 9893 6560
rect 9829 6500 9833 6556
rect 9833 6500 9889 6556
rect 9889 6500 9893 6556
rect 9829 6496 9893 6500
rect 9909 6556 9973 6560
rect 9909 6500 9913 6556
rect 9913 6500 9969 6556
rect 9969 6500 9973 6556
rect 9909 6496 9973 6500
rect 9989 6556 10053 6560
rect 9989 6500 9993 6556
rect 9993 6500 10049 6556
rect 10049 6500 10053 6556
rect 9989 6496 10053 6500
rect 10069 6556 10133 6560
rect 10069 6500 10073 6556
rect 10073 6500 10129 6556
rect 10129 6500 10133 6556
rect 10069 6496 10133 6500
rect 14268 6556 14332 6560
rect 14268 6500 14272 6556
rect 14272 6500 14328 6556
rect 14328 6500 14332 6556
rect 14268 6496 14332 6500
rect 14348 6556 14412 6560
rect 14348 6500 14352 6556
rect 14352 6500 14408 6556
rect 14408 6500 14412 6556
rect 14348 6496 14412 6500
rect 14428 6556 14492 6560
rect 14428 6500 14432 6556
rect 14432 6500 14488 6556
rect 14488 6500 14492 6556
rect 14428 6496 14492 6500
rect 14508 6556 14572 6560
rect 14508 6500 14512 6556
rect 14512 6500 14568 6556
rect 14568 6500 14572 6556
rect 14508 6496 14572 6500
rect 18707 6556 18771 6560
rect 18707 6500 18711 6556
rect 18711 6500 18767 6556
rect 18767 6500 18771 6556
rect 18707 6496 18771 6500
rect 18787 6556 18851 6560
rect 18787 6500 18791 6556
rect 18791 6500 18847 6556
rect 18847 6500 18851 6556
rect 18787 6496 18851 6500
rect 18867 6556 18931 6560
rect 18867 6500 18871 6556
rect 18871 6500 18927 6556
rect 18927 6500 18931 6556
rect 18867 6496 18931 6500
rect 18947 6556 19011 6560
rect 18947 6500 18951 6556
rect 18951 6500 19007 6556
rect 19007 6500 19011 6556
rect 18947 6496 19011 6500
rect 3171 6012 3235 6016
rect 3171 5956 3175 6012
rect 3175 5956 3231 6012
rect 3231 5956 3235 6012
rect 3171 5952 3235 5956
rect 3251 6012 3315 6016
rect 3251 5956 3255 6012
rect 3255 5956 3311 6012
rect 3311 5956 3315 6012
rect 3251 5952 3315 5956
rect 3331 6012 3395 6016
rect 3331 5956 3335 6012
rect 3335 5956 3391 6012
rect 3391 5956 3395 6012
rect 3331 5952 3395 5956
rect 3411 6012 3475 6016
rect 3411 5956 3415 6012
rect 3415 5956 3471 6012
rect 3471 5956 3475 6012
rect 3411 5952 3475 5956
rect 7610 6012 7674 6016
rect 7610 5956 7614 6012
rect 7614 5956 7670 6012
rect 7670 5956 7674 6012
rect 7610 5952 7674 5956
rect 7690 6012 7754 6016
rect 7690 5956 7694 6012
rect 7694 5956 7750 6012
rect 7750 5956 7754 6012
rect 7690 5952 7754 5956
rect 7770 6012 7834 6016
rect 7770 5956 7774 6012
rect 7774 5956 7830 6012
rect 7830 5956 7834 6012
rect 7770 5952 7834 5956
rect 7850 6012 7914 6016
rect 7850 5956 7854 6012
rect 7854 5956 7910 6012
rect 7910 5956 7914 6012
rect 7850 5952 7914 5956
rect 12049 6012 12113 6016
rect 12049 5956 12053 6012
rect 12053 5956 12109 6012
rect 12109 5956 12113 6012
rect 12049 5952 12113 5956
rect 12129 6012 12193 6016
rect 12129 5956 12133 6012
rect 12133 5956 12189 6012
rect 12189 5956 12193 6012
rect 12129 5952 12193 5956
rect 12209 6012 12273 6016
rect 12209 5956 12213 6012
rect 12213 5956 12269 6012
rect 12269 5956 12273 6012
rect 12209 5952 12273 5956
rect 12289 6012 12353 6016
rect 12289 5956 12293 6012
rect 12293 5956 12349 6012
rect 12349 5956 12353 6012
rect 12289 5952 12353 5956
rect 16488 6012 16552 6016
rect 16488 5956 16492 6012
rect 16492 5956 16548 6012
rect 16548 5956 16552 6012
rect 16488 5952 16552 5956
rect 16568 6012 16632 6016
rect 16568 5956 16572 6012
rect 16572 5956 16628 6012
rect 16628 5956 16632 6012
rect 16568 5952 16632 5956
rect 16648 6012 16712 6016
rect 16648 5956 16652 6012
rect 16652 5956 16708 6012
rect 16708 5956 16712 6012
rect 16648 5952 16712 5956
rect 16728 6012 16792 6016
rect 16728 5956 16732 6012
rect 16732 5956 16788 6012
rect 16788 5956 16792 6012
rect 16728 5952 16792 5956
rect 5390 5468 5454 5472
rect 5390 5412 5394 5468
rect 5394 5412 5450 5468
rect 5450 5412 5454 5468
rect 5390 5408 5454 5412
rect 5470 5468 5534 5472
rect 5470 5412 5474 5468
rect 5474 5412 5530 5468
rect 5530 5412 5534 5468
rect 5470 5408 5534 5412
rect 5550 5468 5614 5472
rect 5550 5412 5554 5468
rect 5554 5412 5610 5468
rect 5610 5412 5614 5468
rect 5550 5408 5614 5412
rect 5630 5468 5694 5472
rect 5630 5412 5634 5468
rect 5634 5412 5690 5468
rect 5690 5412 5694 5468
rect 5630 5408 5694 5412
rect 9829 5468 9893 5472
rect 9829 5412 9833 5468
rect 9833 5412 9889 5468
rect 9889 5412 9893 5468
rect 9829 5408 9893 5412
rect 9909 5468 9973 5472
rect 9909 5412 9913 5468
rect 9913 5412 9969 5468
rect 9969 5412 9973 5468
rect 9909 5408 9973 5412
rect 9989 5468 10053 5472
rect 9989 5412 9993 5468
rect 9993 5412 10049 5468
rect 10049 5412 10053 5468
rect 9989 5408 10053 5412
rect 10069 5468 10133 5472
rect 10069 5412 10073 5468
rect 10073 5412 10129 5468
rect 10129 5412 10133 5468
rect 10069 5408 10133 5412
rect 14268 5468 14332 5472
rect 14268 5412 14272 5468
rect 14272 5412 14328 5468
rect 14328 5412 14332 5468
rect 14268 5408 14332 5412
rect 14348 5468 14412 5472
rect 14348 5412 14352 5468
rect 14352 5412 14408 5468
rect 14408 5412 14412 5468
rect 14348 5408 14412 5412
rect 14428 5468 14492 5472
rect 14428 5412 14432 5468
rect 14432 5412 14488 5468
rect 14488 5412 14492 5468
rect 14428 5408 14492 5412
rect 14508 5468 14572 5472
rect 14508 5412 14512 5468
rect 14512 5412 14568 5468
rect 14568 5412 14572 5468
rect 14508 5408 14572 5412
rect 18707 5468 18771 5472
rect 18707 5412 18711 5468
rect 18711 5412 18767 5468
rect 18767 5412 18771 5468
rect 18707 5408 18771 5412
rect 18787 5468 18851 5472
rect 18787 5412 18791 5468
rect 18791 5412 18847 5468
rect 18847 5412 18851 5468
rect 18787 5408 18851 5412
rect 18867 5468 18931 5472
rect 18867 5412 18871 5468
rect 18871 5412 18927 5468
rect 18927 5412 18931 5468
rect 18867 5408 18931 5412
rect 18947 5468 19011 5472
rect 18947 5412 18951 5468
rect 18951 5412 19007 5468
rect 19007 5412 19011 5468
rect 18947 5408 19011 5412
rect 3171 4924 3235 4928
rect 3171 4868 3175 4924
rect 3175 4868 3231 4924
rect 3231 4868 3235 4924
rect 3171 4864 3235 4868
rect 3251 4924 3315 4928
rect 3251 4868 3255 4924
rect 3255 4868 3311 4924
rect 3311 4868 3315 4924
rect 3251 4864 3315 4868
rect 3331 4924 3395 4928
rect 3331 4868 3335 4924
rect 3335 4868 3391 4924
rect 3391 4868 3395 4924
rect 3331 4864 3395 4868
rect 3411 4924 3475 4928
rect 3411 4868 3415 4924
rect 3415 4868 3471 4924
rect 3471 4868 3475 4924
rect 3411 4864 3475 4868
rect 7610 4924 7674 4928
rect 7610 4868 7614 4924
rect 7614 4868 7670 4924
rect 7670 4868 7674 4924
rect 7610 4864 7674 4868
rect 7690 4924 7754 4928
rect 7690 4868 7694 4924
rect 7694 4868 7750 4924
rect 7750 4868 7754 4924
rect 7690 4864 7754 4868
rect 7770 4924 7834 4928
rect 7770 4868 7774 4924
rect 7774 4868 7830 4924
rect 7830 4868 7834 4924
rect 7770 4864 7834 4868
rect 7850 4924 7914 4928
rect 7850 4868 7854 4924
rect 7854 4868 7910 4924
rect 7910 4868 7914 4924
rect 7850 4864 7914 4868
rect 12049 4924 12113 4928
rect 12049 4868 12053 4924
rect 12053 4868 12109 4924
rect 12109 4868 12113 4924
rect 12049 4864 12113 4868
rect 12129 4924 12193 4928
rect 12129 4868 12133 4924
rect 12133 4868 12189 4924
rect 12189 4868 12193 4924
rect 12129 4864 12193 4868
rect 12209 4924 12273 4928
rect 12209 4868 12213 4924
rect 12213 4868 12269 4924
rect 12269 4868 12273 4924
rect 12209 4864 12273 4868
rect 12289 4924 12353 4928
rect 12289 4868 12293 4924
rect 12293 4868 12349 4924
rect 12349 4868 12353 4924
rect 12289 4864 12353 4868
rect 16488 4924 16552 4928
rect 16488 4868 16492 4924
rect 16492 4868 16548 4924
rect 16548 4868 16552 4924
rect 16488 4864 16552 4868
rect 16568 4924 16632 4928
rect 16568 4868 16572 4924
rect 16572 4868 16628 4924
rect 16628 4868 16632 4924
rect 16568 4864 16632 4868
rect 16648 4924 16712 4928
rect 16648 4868 16652 4924
rect 16652 4868 16708 4924
rect 16708 4868 16712 4924
rect 16648 4864 16712 4868
rect 16728 4924 16792 4928
rect 16728 4868 16732 4924
rect 16732 4868 16788 4924
rect 16788 4868 16792 4924
rect 16728 4864 16792 4868
rect 5390 4380 5454 4384
rect 5390 4324 5394 4380
rect 5394 4324 5450 4380
rect 5450 4324 5454 4380
rect 5390 4320 5454 4324
rect 5470 4380 5534 4384
rect 5470 4324 5474 4380
rect 5474 4324 5530 4380
rect 5530 4324 5534 4380
rect 5470 4320 5534 4324
rect 5550 4380 5614 4384
rect 5550 4324 5554 4380
rect 5554 4324 5610 4380
rect 5610 4324 5614 4380
rect 5550 4320 5614 4324
rect 5630 4380 5694 4384
rect 5630 4324 5634 4380
rect 5634 4324 5690 4380
rect 5690 4324 5694 4380
rect 5630 4320 5694 4324
rect 9829 4380 9893 4384
rect 9829 4324 9833 4380
rect 9833 4324 9889 4380
rect 9889 4324 9893 4380
rect 9829 4320 9893 4324
rect 9909 4380 9973 4384
rect 9909 4324 9913 4380
rect 9913 4324 9969 4380
rect 9969 4324 9973 4380
rect 9909 4320 9973 4324
rect 9989 4380 10053 4384
rect 9989 4324 9993 4380
rect 9993 4324 10049 4380
rect 10049 4324 10053 4380
rect 9989 4320 10053 4324
rect 10069 4380 10133 4384
rect 10069 4324 10073 4380
rect 10073 4324 10129 4380
rect 10129 4324 10133 4380
rect 10069 4320 10133 4324
rect 14268 4380 14332 4384
rect 14268 4324 14272 4380
rect 14272 4324 14328 4380
rect 14328 4324 14332 4380
rect 14268 4320 14332 4324
rect 14348 4380 14412 4384
rect 14348 4324 14352 4380
rect 14352 4324 14408 4380
rect 14408 4324 14412 4380
rect 14348 4320 14412 4324
rect 14428 4380 14492 4384
rect 14428 4324 14432 4380
rect 14432 4324 14488 4380
rect 14488 4324 14492 4380
rect 14428 4320 14492 4324
rect 14508 4380 14572 4384
rect 14508 4324 14512 4380
rect 14512 4324 14568 4380
rect 14568 4324 14572 4380
rect 14508 4320 14572 4324
rect 18707 4380 18771 4384
rect 18707 4324 18711 4380
rect 18711 4324 18767 4380
rect 18767 4324 18771 4380
rect 18707 4320 18771 4324
rect 18787 4380 18851 4384
rect 18787 4324 18791 4380
rect 18791 4324 18847 4380
rect 18847 4324 18851 4380
rect 18787 4320 18851 4324
rect 18867 4380 18931 4384
rect 18867 4324 18871 4380
rect 18871 4324 18927 4380
rect 18927 4324 18931 4380
rect 18867 4320 18931 4324
rect 18947 4380 19011 4384
rect 18947 4324 18951 4380
rect 18951 4324 19007 4380
rect 19007 4324 19011 4380
rect 18947 4320 19011 4324
rect 3171 3836 3235 3840
rect 3171 3780 3175 3836
rect 3175 3780 3231 3836
rect 3231 3780 3235 3836
rect 3171 3776 3235 3780
rect 3251 3836 3315 3840
rect 3251 3780 3255 3836
rect 3255 3780 3311 3836
rect 3311 3780 3315 3836
rect 3251 3776 3315 3780
rect 3331 3836 3395 3840
rect 3331 3780 3335 3836
rect 3335 3780 3391 3836
rect 3391 3780 3395 3836
rect 3331 3776 3395 3780
rect 3411 3836 3475 3840
rect 3411 3780 3415 3836
rect 3415 3780 3471 3836
rect 3471 3780 3475 3836
rect 3411 3776 3475 3780
rect 7610 3836 7674 3840
rect 7610 3780 7614 3836
rect 7614 3780 7670 3836
rect 7670 3780 7674 3836
rect 7610 3776 7674 3780
rect 7690 3836 7754 3840
rect 7690 3780 7694 3836
rect 7694 3780 7750 3836
rect 7750 3780 7754 3836
rect 7690 3776 7754 3780
rect 7770 3836 7834 3840
rect 7770 3780 7774 3836
rect 7774 3780 7830 3836
rect 7830 3780 7834 3836
rect 7770 3776 7834 3780
rect 7850 3836 7914 3840
rect 7850 3780 7854 3836
rect 7854 3780 7910 3836
rect 7910 3780 7914 3836
rect 7850 3776 7914 3780
rect 12049 3836 12113 3840
rect 12049 3780 12053 3836
rect 12053 3780 12109 3836
rect 12109 3780 12113 3836
rect 12049 3776 12113 3780
rect 12129 3836 12193 3840
rect 12129 3780 12133 3836
rect 12133 3780 12189 3836
rect 12189 3780 12193 3836
rect 12129 3776 12193 3780
rect 12209 3836 12273 3840
rect 12209 3780 12213 3836
rect 12213 3780 12269 3836
rect 12269 3780 12273 3836
rect 12209 3776 12273 3780
rect 12289 3836 12353 3840
rect 12289 3780 12293 3836
rect 12293 3780 12349 3836
rect 12349 3780 12353 3836
rect 12289 3776 12353 3780
rect 16488 3836 16552 3840
rect 16488 3780 16492 3836
rect 16492 3780 16548 3836
rect 16548 3780 16552 3836
rect 16488 3776 16552 3780
rect 16568 3836 16632 3840
rect 16568 3780 16572 3836
rect 16572 3780 16628 3836
rect 16628 3780 16632 3836
rect 16568 3776 16632 3780
rect 16648 3836 16712 3840
rect 16648 3780 16652 3836
rect 16652 3780 16708 3836
rect 16708 3780 16712 3836
rect 16648 3776 16712 3780
rect 16728 3836 16792 3840
rect 16728 3780 16732 3836
rect 16732 3780 16788 3836
rect 16788 3780 16792 3836
rect 16728 3776 16792 3780
rect 5390 3292 5454 3296
rect 5390 3236 5394 3292
rect 5394 3236 5450 3292
rect 5450 3236 5454 3292
rect 5390 3232 5454 3236
rect 5470 3292 5534 3296
rect 5470 3236 5474 3292
rect 5474 3236 5530 3292
rect 5530 3236 5534 3292
rect 5470 3232 5534 3236
rect 5550 3292 5614 3296
rect 5550 3236 5554 3292
rect 5554 3236 5610 3292
rect 5610 3236 5614 3292
rect 5550 3232 5614 3236
rect 5630 3292 5694 3296
rect 5630 3236 5634 3292
rect 5634 3236 5690 3292
rect 5690 3236 5694 3292
rect 5630 3232 5694 3236
rect 9829 3292 9893 3296
rect 9829 3236 9833 3292
rect 9833 3236 9889 3292
rect 9889 3236 9893 3292
rect 9829 3232 9893 3236
rect 9909 3292 9973 3296
rect 9909 3236 9913 3292
rect 9913 3236 9969 3292
rect 9969 3236 9973 3292
rect 9909 3232 9973 3236
rect 9989 3292 10053 3296
rect 9989 3236 9993 3292
rect 9993 3236 10049 3292
rect 10049 3236 10053 3292
rect 9989 3232 10053 3236
rect 10069 3292 10133 3296
rect 10069 3236 10073 3292
rect 10073 3236 10129 3292
rect 10129 3236 10133 3292
rect 10069 3232 10133 3236
rect 14268 3292 14332 3296
rect 14268 3236 14272 3292
rect 14272 3236 14328 3292
rect 14328 3236 14332 3292
rect 14268 3232 14332 3236
rect 14348 3292 14412 3296
rect 14348 3236 14352 3292
rect 14352 3236 14408 3292
rect 14408 3236 14412 3292
rect 14348 3232 14412 3236
rect 14428 3292 14492 3296
rect 14428 3236 14432 3292
rect 14432 3236 14488 3292
rect 14488 3236 14492 3292
rect 14428 3232 14492 3236
rect 14508 3292 14572 3296
rect 14508 3236 14512 3292
rect 14512 3236 14568 3292
rect 14568 3236 14572 3292
rect 14508 3232 14572 3236
rect 18707 3292 18771 3296
rect 18707 3236 18711 3292
rect 18711 3236 18767 3292
rect 18767 3236 18771 3292
rect 18707 3232 18771 3236
rect 18787 3292 18851 3296
rect 18787 3236 18791 3292
rect 18791 3236 18847 3292
rect 18847 3236 18851 3292
rect 18787 3232 18851 3236
rect 18867 3292 18931 3296
rect 18867 3236 18871 3292
rect 18871 3236 18927 3292
rect 18927 3236 18931 3292
rect 18867 3232 18931 3236
rect 18947 3292 19011 3296
rect 18947 3236 18951 3292
rect 18951 3236 19007 3292
rect 19007 3236 19011 3292
rect 18947 3232 19011 3236
rect 3171 2748 3235 2752
rect 3171 2692 3175 2748
rect 3175 2692 3231 2748
rect 3231 2692 3235 2748
rect 3171 2688 3235 2692
rect 3251 2748 3315 2752
rect 3251 2692 3255 2748
rect 3255 2692 3311 2748
rect 3311 2692 3315 2748
rect 3251 2688 3315 2692
rect 3331 2748 3395 2752
rect 3331 2692 3335 2748
rect 3335 2692 3391 2748
rect 3391 2692 3395 2748
rect 3331 2688 3395 2692
rect 3411 2748 3475 2752
rect 3411 2692 3415 2748
rect 3415 2692 3471 2748
rect 3471 2692 3475 2748
rect 3411 2688 3475 2692
rect 7610 2748 7674 2752
rect 7610 2692 7614 2748
rect 7614 2692 7670 2748
rect 7670 2692 7674 2748
rect 7610 2688 7674 2692
rect 7690 2748 7754 2752
rect 7690 2692 7694 2748
rect 7694 2692 7750 2748
rect 7750 2692 7754 2748
rect 7690 2688 7754 2692
rect 7770 2748 7834 2752
rect 7770 2692 7774 2748
rect 7774 2692 7830 2748
rect 7830 2692 7834 2748
rect 7770 2688 7834 2692
rect 7850 2748 7914 2752
rect 7850 2692 7854 2748
rect 7854 2692 7910 2748
rect 7910 2692 7914 2748
rect 7850 2688 7914 2692
rect 12049 2748 12113 2752
rect 12049 2692 12053 2748
rect 12053 2692 12109 2748
rect 12109 2692 12113 2748
rect 12049 2688 12113 2692
rect 12129 2748 12193 2752
rect 12129 2692 12133 2748
rect 12133 2692 12189 2748
rect 12189 2692 12193 2748
rect 12129 2688 12193 2692
rect 12209 2748 12273 2752
rect 12209 2692 12213 2748
rect 12213 2692 12269 2748
rect 12269 2692 12273 2748
rect 12209 2688 12273 2692
rect 12289 2748 12353 2752
rect 12289 2692 12293 2748
rect 12293 2692 12349 2748
rect 12349 2692 12353 2748
rect 12289 2688 12353 2692
rect 16488 2748 16552 2752
rect 16488 2692 16492 2748
rect 16492 2692 16548 2748
rect 16548 2692 16552 2748
rect 16488 2688 16552 2692
rect 16568 2748 16632 2752
rect 16568 2692 16572 2748
rect 16572 2692 16628 2748
rect 16628 2692 16632 2748
rect 16568 2688 16632 2692
rect 16648 2748 16712 2752
rect 16648 2692 16652 2748
rect 16652 2692 16708 2748
rect 16708 2692 16712 2748
rect 16648 2688 16712 2692
rect 16728 2748 16792 2752
rect 16728 2692 16732 2748
rect 16732 2692 16788 2748
rect 16788 2692 16792 2748
rect 16728 2688 16792 2692
rect 5390 2204 5454 2208
rect 5390 2148 5394 2204
rect 5394 2148 5450 2204
rect 5450 2148 5454 2204
rect 5390 2144 5454 2148
rect 5470 2204 5534 2208
rect 5470 2148 5474 2204
rect 5474 2148 5530 2204
rect 5530 2148 5534 2204
rect 5470 2144 5534 2148
rect 5550 2204 5614 2208
rect 5550 2148 5554 2204
rect 5554 2148 5610 2204
rect 5610 2148 5614 2204
rect 5550 2144 5614 2148
rect 5630 2204 5694 2208
rect 5630 2148 5634 2204
rect 5634 2148 5690 2204
rect 5690 2148 5694 2204
rect 5630 2144 5694 2148
rect 9829 2204 9893 2208
rect 9829 2148 9833 2204
rect 9833 2148 9889 2204
rect 9889 2148 9893 2204
rect 9829 2144 9893 2148
rect 9909 2204 9973 2208
rect 9909 2148 9913 2204
rect 9913 2148 9969 2204
rect 9969 2148 9973 2204
rect 9909 2144 9973 2148
rect 9989 2204 10053 2208
rect 9989 2148 9993 2204
rect 9993 2148 10049 2204
rect 10049 2148 10053 2204
rect 9989 2144 10053 2148
rect 10069 2204 10133 2208
rect 10069 2148 10073 2204
rect 10073 2148 10129 2204
rect 10129 2148 10133 2204
rect 10069 2144 10133 2148
rect 14268 2204 14332 2208
rect 14268 2148 14272 2204
rect 14272 2148 14328 2204
rect 14328 2148 14332 2204
rect 14268 2144 14332 2148
rect 14348 2204 14412 2208
rect 14348 2148 14352 2204
rect 14352 2148 14408 2204
rect 14408 2148 14412 2204
rect 14348 2144 14412 2148
rect 14428 2204 14492 2208
rect 14428 2148 14432 2204
rect 14432 2148 14488 2204
rect 14488 2148 14492 2204
rect 14428 2144 14492 2148
rect 14508 2204 14572 2208
rect 14508 2148 14512 2204
rect 14512 2148 14568 2204
rect 14568 2148 14572 2204
rect 14508 2144 14572 2148
rect 18707 2204 18771 2208
rect 18707 2148 18711 2204
rect 18711 2148 18767 2204
rect 18767 2148 18771 2204
rect 18707 2144 18771 2148
rect 18787 2204 18851 2208
rect 18787 2148 18791 2204
rect 18791 2148 18847 2204
rect 18847 2148 18851 2204
rect 18787 2144 18851 2148
rect 18867 2204 18931 2208
rect 18867 2148 18871 2204
rect 18871 2148 18927 2204
rect 18927 2148 18931 2204
rect 18867 2144 18931 2148
rect 18947 2204 19011 2208
rect 18947 2148 18951 2204
rect 18951 2148 19007 2204
rect 19007 2148 19011 2204
rect 18947 2144 19011 2148
<< metal4 >>
rect 3163 7104 3483 7664
rect 3163 7040 3171 7104
rect 3235 7040 3251 7104
rect 3315 7040 3331 7104
rect 3395 7040 3411 7104
rect 3475 7040 3483 7104
rect 3163 6016 3483 7040
rect 3163 5952 3171 6016
rect 3235 5952 3251 6016
rect 3315 5952 3331 6016
rect 3395 5952 3411 6016
rect 3475 5952 3483 6016
rect 3163 4928 3483 5952
rect 3163 4864 3171 4928
rect 3235 4864 3251 4928
rect 3315 4864 3331 4928
rect 3395 4864 3411 4928
rect 3475 4864 3483 4928
rect 3163 3840 3483 4864
rect 3163 3776 3171 3840
rect 3235 3776 3251 3840
rect 3315 3776 3331 3840
rect 3395 3776 3411 3840
rect 3475 3776 3483 3840
rect 3163 2752 3483 3776
rect 3163 2688 3171 2752
rect 3235 2688 3251 2752
rect 3315 2688 3331 2752
rect 3395 2688 3411 2752
rect 3475 2688 3483 2752
rect 3163 2128 3483 2688
rect 5382 7648 5702 7664
rect 5382 7584 5390 7648
rect 5454 7584 5470 7648
rect 5534 7584 5550 7648
rect 5614 7584 5630 7648
rect 5694 7584 5702 7648
rect 5382 6560 5702 7584
rect 5382 6496 5390 6560
rect 5454 6496 5470 6560
rect 5534 6496 5550 6560
rect 5614 6496 5630 6560
rect 5694 6496 5702 6560
rect 5382 5472 5702 6496
rect 5382 5408 5390 5472
rect 5454 5408 5470 5472
rect 5534 5408 5550 5472
rect 5614 5408 5630 5472
rect 5694 5408 5702 5472
rect 5382 4384 5702 5408
rect 5382 4320 5390 4384
rect 5454 4320 5470 4384
rect 5534 4320 5550 4384
rect 5614 4320 5630 4384
rect 5694 4320 5702 4384
rect 5382 3296 5702 4320
rect 5382 3232 5390 3296
rect 5454 3232 5470 3296
rect 5534 3232 5550 3296
rect 5614 3232 5630 3296
rect 5694 3232 5702 3296
rect 5382 2208 5702 3232
rect 5382 2144 5390 2208
rect 5454 2144 5470 2208
rect 5534 2144 5550 2208
rect 5614 2144 5630 2208
rect 5694 2144 5702 2208
rect 5382 2128 5702 2144
rect 7602 7104 7922 7664
rect 7602 7040 7610 7104
rect 7674 7040 7690 7104
rect 7754 7040 7770 7104
rect 7834 7040 7850 7104
rect 7914 7040 7922 7104
rect 7602 6016 7922 7040
rect 7602 5952 7610 6016
rect 7674 5952 7690 6016
rect 7754 5952 7770 6016
rect 7834 5952 7850 6016
rect 7914 5952 7922 6016
rect 7602 4928 7922 5952
rect 7602 4864 7610 4928
rect 7674 4864 7690 4928
rect 7754 4864 7770 4928
rect 7834 4864 7850 4928
rect 7914 4864 7922 4928
rect 7602 3840 7922 4864
rect 7602 3776 7610 3840
rect 7674 3776 7690 3840
rect 7754 3776 7770 3840
rect 7834 3776 7850 3840
rect 7914 3776 7922 3840
rect 7602 2752 7922 3776
rect 7602 2688 7610 2752
rect 7674 2688 7690 2752
rect 7754 2688 7770 2752
rect 7834 2688 7850 2752
rect 7914 2688 7922 2752
rect 7602 2128 7922 2688
rect 9821 7648 10141 7664
rect 9821 7584 9829 7648
rect 9893 7584 9909 7648
rect 9973 7584 9989 7648
rect 10053 7584 10069 7648
rect 10133 7584 10141 7648
rect 9821 6560 10141 7584
rect 9821 6496 9829 6560
rect 9893 6496 9909 6560
rect 9973 6496 9989 6560
rect 10053 6496 10069 6560
rect 10133 6496 10141 6560
rect 9821 5472 10141 6496
rect 9821 5408 9829 5472
rect 9893 5408 9909 5472
rect 9973 5408 9989 5472
rect 10053 5408 10069 5472
rect 10133 5408 10141 5472
rect 9821 4384 10141 5408
rect 9821 4320 9829 4384
rect 9893 4320 9909 4384
rect 9973 4320 9989 4384
rect 10053 4320 10069 4384
rect 10133 4320 10141 4384
rect 9821 3296 10141 4320
rect 9821 3232 9829 3296
rect 9893 3232 9909 3296
rect 9973 3232 9989 3296
rect 10053 3232 10069 3296
rect 10133 3232 10141 3296
rect 9821 2208 10141 3232
rect 9821 2144 9829 2208
rect 9893 2144 9909 2208
rect 9973 2144 9989 2208
rect 10053 2144 10069 2208
rect 10133 2144 10141 2208
rect 9821 2128 10141 2144
rect 12041 7104 12361 7664
rect 12041 7040 12049 7104
rect 12113 7040 12129 7104
rect 12193 7040 12209 7104
rect 12273 7040 12289 7104
rect 12353 7040 12361 7104
rect 12041 6016 12361 7040
rect 12041 5952 12049 6016
rect 12113 5952 12129 6016
rect 12193 5952 12209 6016
rect 12273 5952 12289 6016
rect 12353 5952 12361 6016
rect 12041 4928 12361 5952
rect 12041 4864 12049 4928
rect 12113 4864 12129 4928
rect 12193 4864 12209 4928
rect 12273 4864 12289 4928
rect 12353 4864 12361 4928
rect 12041 3840 12361 4864
rect 12041 3776 12049 3840
rect 12113 3776 12129 3840
rect 12193 3776 12209 3840
rect 12273 3776 12289 3840
rect 12353 3776 12361 3840
rect 12041 2752 12361 3776
rect 12041 2688 12049 2752
rect 12113 2688 12129 2752
rect 12193 2688 12209 2752
rect 12273 2688 12289 2752
rect 12353 2688 12361 2752
rect 12041 2128 12361 2688
rect 14260 7648 14580 7664
rect 14260 7584 14268 7648
rect 14332 7584 14348 7648
rect 14412 7584 14428 7648
rect 14492 7584 14508 7648
rect 14572 7584 14580 7648
rect 14260 6560 14580 7584
rect 14260 6496 14268 6560
rect 14332 6496 14348 6560
rect 14412 6496 14428 6560
rect 14492 6496 14508 6560
rect 14572 6496 14580 6560
rect 14260 5472 14580 6496
rect 14260 5408 14268 5472
rect 14332 5408 14348 5472
rect 14412 5408 14428 5472
rect 14492 5408 14508 5472
rect 14572 5408 14580 5472
rect 14260 4384 14580 5408
rect 14260 4320 14268 4384
rect 14332 4320 14348 4384
rect 14412 4320 14428 4384
rect 14492 4320 14508 4384
rect 14572 4320 14580 4384
rect 14260 3296 14580 4320
rect 14260 3232 14268 3296
rect 14332 3232 14348 3296
rect 14412 3232 14428 3296
rect 14492 3232 14508 3296
rect 14572 3232 14580 3296
rect 14260 2208 14580 3232
rect 14260 2144 14268 2208
rect 14332 2144 14348 2208
rect 14412 2144 14428 2208
rect 14492 2144 14508 2208
rect 14572 2144 14580 2208
rect 14260 2128 14580 2144
rect 16480 7104 16800 7664
rect 16480 7040 16488 7104
rect 16552 7040 16568 7104
rect 16632 7040 16648 7104
rect 16712 7040 16728 7104
rect 16792 7040 16800 7104
rect 16480 6016 16800 7040
rect 16480 5952 16488 6016
rect 16552 5952 16568 6016
rect 16632 5952 16648 6016
rect 16712 5952 16728 6016
rect 16792 5952 16800 6016
rect 16480 4928 16800 5952
rect 16480 4864 16488 4928
rect 16552 4864 16568 4928
rect 16632 4864 16648 4928
rect 16712 4864 16728 4928
rect 16792 4864 16800 4928
rect 16480 3840 16800 4864
rect 16480 3776 16488 3840
rect 16552 3776 16568 3840
rect 16632 3776 16648 3840
rect 16712 3776 16728 3840
rect 16792 3776 16800 3840
rect 16480 2752 16800 3776
rect 16480 2688 16488 2752
rect 16552 2688 16568 2752
rect 16632 2688 16648 2752
rect 16712 2688 16728 2752
rect 16792 2688 16800 2752
rect 16480 2128 16800 2688
rect 18699 7648 19019 7664
rect 18699 7584 18707 7648
rect 18771 7584 18787 7648
rect 18851 7584 18867 7648
rect 18931 7584 18947 7648
rect 19011 7584 19019 7648
rect 18699 6560 19019 7584
rect 18699 6496 18707 6560
rect 18771 6496 18787 6560
rect 18851 6496 18867 6560
rect 18931 6496 18947 6560
rect 19011 6496 19019 6560
rect 18699 5472 19019 6496
rect 18699 5408 18707 5472
rect 18771 5408 18787 5472
rect 18851 5408 18867 5472
rect 18931 5408 18947 5472
rect 19011 5408 19019 5472
rect 18699 4384 19019 5408
rect 18699 4320 18707 4384
rect 18771 4320 18787 4384
rect 18851 4320 18867 4384
rect 18931 4320 18947 4384
rect 19011 4320 19019 4384
rect 18699 3296 19019 4320
rect 18699 3232 18707 3296
rect 18771 3232 18787 3296
rect 18851 3232 18867 3296
rect 18931 3232 18947 3296
rect 19011 3232 19019 3296
rect 18699 2208 19019 3232
rect 18699 2144 18707 2208
rect 18771 2144 18787 2208
rect 18851 2144 18867 2208
rect 18931 2144 18947 2208
rect 19011 2144 19019 2208
rect 18699 2128 19019 2144
<< labels >>
rlabel metal1 s 9982 7072 9982 7072 4 vccd1
rlabel metal2 s 10061 7616 10061 7616 4 vssd1
rlabel metal2 s 11178 3842 11178 3842 4 _00_
rlabel metal2 s 16882 3672 16882 3672 4 _01_
rlabel metal2 s 16054 4080 16054 4080 4 _02_
rlabel metal1 s 13202 4488 13202 4488 4 _03_
rlabel metal1 s 4922 4046 4922 4046 4 _04_
rlabel metal1 s 14122 4046 14122 4046 4 _05_
rlabel metal1 s 4600 2482 4600 2482 4 _06_
rlabel metal2 s 8700 3094 8700 3094 4 _07_
rlabel metal2 s 10534 4794 10534 4794 4 _08_
rlabel metal2 s 10994 3978 10994 3978 4 _09_
rlabel metal2 s 15226 4794 15226 4794 4 _10_
rlabel metal1 s 16721 4590 16721 4590 4 _11_
rlabel metal1 s 12788 4794 12788 4794 4 _12_
rlabel metal1 s 16238 4624 16238 4624 4 _13_
rlabel metal1 s 11638 5338 11638 5338 4 _14_
rlabel metal1 s 13248 4590 13248 4590 4 _15_
rlabel metal1 s 6394 4624 6394 4624 4 _16_
rlabel metal2 s 6854 4284 6854 4284 4 _17_
rlabel metal1 s 8188 5882 8188 5882 4 _18_
rlabel metal1 s 11178 4590 11178 4590 4 _19_
rlabel metal2 s 6854 4794 6854 4794 4 _20_
rlabel metal1 s 7084 4794 7084 4794 4 _21_
rlabel metal2 s 8418 4386 8418 4386 4 _22_
rlabel metal2 s 10258 3978 10258 3978 4 _23_
rlabel metal1 s 9798 4590 9798 4590 4 clk
rlabel metal2 s 9430 3502 9430 3502 4 clknet_0_clk
rlabel metal1 s 2116 2482 2116 2482 4 clknet_1_0__leaf_clk
rlabel metal1 s 14904 2482 14904 2482 4 clknet_1_1__leaf_clk
rlabel metal1 s 10212 7446 10212 7446 4 comp
rlabel metal1 s 1426 7514 1426 7514 4 dq[0]
rlabel metal1 s 3726 7514 3726 7514 4 dq[1]
rlabel metal2 s 5750 8415 5750 8415 4 dq[2]
rlabel metal2 s 7958 8415 7958 8415 4 dq[3]
rlabel metal2 s 12374 8415 12374 8415 4 dq[4]
rlabel metal2 s 14674 8415 14674 8415 4 dq[5]
rlabel metal1 s 16836 7514 16836 7514 4 dq[6]
rlabel metal1 s 18354 7514 18354 7514 4 dq[7]
rlabel metal2 s 17434 1520 17434 1520 4 last_cycle
rlabel metal2 s 12466 4998 12466 4998 4 net1
rlabel metal1 s 18078 7344 18078 7344 4 net10
rlabel metal2 s 1978 2754 1978 2754 4 net11
rlabel metal2 s 13938 4046 13938 4046 4 net12
rlabel metal1 s 13708 4182 13708 4182 4 net13
rlabel metal2 s 9338 2519 9338 2519 4 net14
rlabel metal2 s 4554 3502 4554 3502 4 net15
rlabel metal2 s 2254 4284 2254 4284 4 net16
rlabel metal1 s 4692 4522 4692 4522 4 net2
rlabel metal1 s 1886 7344 1886 7344 4 net3
rlabel metal1 s 8004 4250 8004 4250 4 net4
rlabel metal1 s 6532 2618 6532 2618 4 net5
rlabel metal2 s 13110 3961 13110 3961 4 net6
rlabel metal1 s 7774 4454 7774 4454 4 net7
rlabel metal1 s 14168 7378 14168 7378 4 net8
rlabel metal2 s 16882 6052 16882 6052 4 net9
rlabel metal2 s 2714 3213 2714 3213 4 rst_n
rlabel metal1 s 7222 5100 7222 5100 4 sr\[1\]
rlabel metal1 s 8694 2618 8694 2618 4 sr\[2\]
rlabel metal1 s 9338 2482 9338 2482 4 sr\[3\]
rlabel metal1 s 12604 2482 12604 2482 4 sr\[4\]
rlabel metal1 s 13478 3400 13478 3400 4 sr\[5\]
rlabel metal1 s 13064 3094 13064 3094 4 sr\[6\]
rlabel metal2 s 15778 2618 15778 2618 4 sr\[7\]
rlabel metal2 s 12466 1792 12466 1792 4 valid
flabel metal2 s 7470 0 7526 800 0 FreeSans 280 90 0 0 clk
port 1 nsew
flabel metal2 s 9954 9200 10010 10000 0 FreeSans 280 90 0 0 comp
port 2 nsew
flabel metal2 s 1122 9200 1178 10000 0 FreeSans 280 90 0 0 dq[0]
port 3 nsew
flabel metal2 s 3330 9200 3386 10000 0 FreeSans 280 90 0 0 dq[1]
port 4 nsew
flabel metal2 s 5538 9200 5594 10000 0 FreeSans 280 90 0 0 dq[2]
port 5 nsew
flabel metal2 s 7746 9200 7802 10000 0 FreeSans 280 90 0 0 dq[3]
port 6 nsew
flabel metal2 s 12162 9200 12218 10000 0 FreeSans 280 90 0 0 dq[4]
port 7 nsew
flabel metal2 s 14370 9200 14426 10000 0 FreeSans 280 90 0 0 dq[5]
port 8 nsew
flabel metal2 s 16578 9200 16634 10000 0 FreeSans 280 90 0 0 dq[6]
port 9 nsew
flabel metal2 s 18786 9200 18842 10000 0 FreeSans 280 90 0 0 dq[7]
port 10 nsew
flabel metal2 s 17406 0 17462 800 0 FreeSans 280 90 0 0 last_cycle
port 11 nsew
flabel metal2 s 2502 0 2558 800 0 FreeSans 280 90 0 0 rst_n
port 12 nsew
flabel metal2 s 12438 0 12494 800 0 FreeSans 280 90 0 0 valid
port 13 nsew
flabel metal4 s 3163 2128 3483 7664 0 FreeSans 2400 90 0 0 vccd1
port 14 nsew
flabel metal4 s 7602 2128 7922 7664 0 FreeSans 2400 90 0 0 vccd1
port 14 nsew
flabel metal4 s 12041 2128 12361 7664 0 FreeSans 2400 90 0 0 vccd1
port 14 nsew
flabel metal4 s 16480 2128 16800 7664 0 FreeSans 2400 90 0 0 vccd1
port 14 nsew
flabel metal4 s 5382 2128 5702 7664 0 FreeSans 2400 90 0 0 vssd1
port 15 nsew
flabel metal4 s 9821 2128 10141 7664 0 FreeSans 2400 90 0 0 vssd1
port 15 nsew
flabel metal4 s 14260 2128 14580 7664 0 FreeSans 2400 90 0 0 vssd1
port 15 nsew
flabel metal4 s 18699 2128 19019 7664 0 FreeSans 2400 90 0 0 vssd1
port 15 nsew
flabel metal1 1409 2703 1443 2737 0 FreeSans 200 0 0 0 FILLER_0_3.VPWR
flabel metal1 1409 2159 1443 2193 0 FreeSans 200 0 0 0 FILLER_0_3.VGND
flabel nwell 1409 2703 1443 2737 0 FreeSans 200 0 0 0 FILLER_0_3.VPB
flabel pwell 1409 2159 1443 2193 0 FreeSans 200 0 0 0 FILLER_0_3.VNB
rlabel comment 1380 2176 1380 2176 4 FILLER_0_3.decap_3
flabel metal1 1409 2703 1443 2737 0 FreeSans 200 0 0 0 FILLER_1_3.VPWR
flabel metal1 1409 3247 1443 3281 0 FreeSans 200 0 0 0 FILLER_1_3.VGND
flabel nwell 1409 2703 1443 2737 0 FreeSans 200 0 0 0 FILLER_1_3.VPB
flabel pwell 1409 3247 1443 3281 0 FreeSans 200 0 0 0 FILLER_1_3.VNB
rlabel comment 1380 3264 1380 3264 2 FILLER_1_3.decap_6
flabel metal1 1133 2703 1167 2737 0 FreeSans 200 0 0 0 PHY_0.VPWR
flabel metal1 1133 2159 1167 2193 0 FreeSans 200 0 0 0 PHY_0.VGND
flabel nwell 1133 2703 1167 2737 0 FreeSans 200 0 0 0 PHY_0.VPB
flabel pwell 1133 2159 1167 2193 0 FreeSans 200 0 0 0 PHY_0.VNB
rlabel comment 1104 2176 1104 2176 4 PHY_0.decap_3
flabel metal1 1133 2703 1167 2737 0 FreeSans 200 0 0 0 PHY_2.VPWR
flabel metal1 1133 3247 1167 3281 0 FreeSans 200 0 0 0 PHY_2.VGND
flabel nwell 1133 2703 1167 2737 0 FreeSans 200 0 0 0 PHY_2.VPB
flabel pwell 1133 3247 1167 3281 0 FreeSans 200 0 0 0 PHY_2.VNB
rlabel comment 1104 3264 1104 3264 2 PHY_2.decap_3
flabel locali 3432 2601 3466 2635 0 FreeSans 400 0 0 0 _61_.Q
flabel locali 3432 2533 3466 2567 0 FreeSans 400 0 0 0 _61_.Q
flabel locali 3432 2465 3466 2499 0 FreeSans 400 0 0 0 _61_.Q
flabel locali 3432 2261 3466 2295 0 FreeSans 400 0 0 0 _61_.Q
flabel locali 3137 2329 3171 2363 0 FreeSans 400 0 0 0 _61_.RESET_B
flabel locali 1961 2465 1995 2499 0 FreeSans 400 0 0 0 _61_.D
flabel locali 1686 2465 1720 2499 0 FreeSans 400 0 0 0 _61_.CLK
flabel locali 1686 2397 1720 2431 0 FreeSans 400 0 0 0 _61_.CLK
flabel locali 3137 2397 3171 2431 0 FreeSans 400 0 0 0 _61_.RESET_B
flabel metal1 1685 2159 1719 2193 0 FreeSans 200 0 0 0 _61_.VGND
flabel metal1 1685 2703 1719 2737 0 FreeSans 200 0 0 0 _61_.VPWR
flabel nwell 1685 2703 1719 2737 0 FreeSans 200 0 0 0 _61_.VPB
flabel pwell 1685 2159 1719 2193 0 FreeSans 200 0 0 0 _61_.VNB
rlabel comment 1656 2176 1656 2176 4 _61_.dfrtp_1
flabel locali 1962 2805 1996 2839 0 FreeSans 400 0 0 0 _62_.Q
flabel locali 1962 2873 1996 2907 0 FreeSans 400 0 0 0 _62_.Q
flabel locali 1962 2941 1996 2975 0 FreeSans 400 0 0 0 _62_.Q
flabel locali 1962 3145 1996 3179 0 FreeSans 400 0 0 0 _62_.Q
flabel locali 2257 3077 2291 3111 0 FreeSans 400 0 0 0 _62_.RESET_B
flabel locali 3433 2941 3467 2975 0 FreeSans 400 0 0 0 _62_.D
flabel locali 3708 2941 3742 2975 0 FreeSans 400 0 0 0 _62_.CLK
flabel locali 3708 3009 3742 3043 0 FreeSans 400 0 0 0 _62_.CLK
flabel locali 2257 3009 2291 3043 0 FreeSans 400 0 0 0 _62_.RESET_B
flabel metal1 3709 3247 3743 3281 0 FreeSans 200 0 0 0 _62_.VGND
flabel metal1 3709 2703 3743 2737 0 FreeSans 200 0 0 0 _62_.VPWR
flabel nwell 3709 2703 3743 2737 0 FreeSans 200 0 0 0 _62_.VPB
flabel pwell 3709 3247 3743 3281 0 FreeSans 200 0 0 0 _62_.VNB
rlabel comment 3772 3264 3772 3264 8 _62_.dfrtp_1
flabel metal1 3516 2162 3569 2194 0 FreeSans 200 0 0 0 FILLER_0_26.VGND
flabel metal1 3517 2706 3569 2737 0 FreeSans 200 0 0 0 FILLER_0_26.VPWR
flabel nwell 3524 2711 3558 2729 0 FreeSans 200 0 0 0 FILLER_0_26.VPB
flabel pwell 3527 2166 3559 2188 0 FreeSans 200 0 0 0 FILLER_0_26.VNB
rlabel comment 3496 2176 3496 2176 4 FILLER_0_26.fill_2
flabel metal1 3801 2159 3835 2193 0 FreeSans 200 0 0 0 FILLER_0_29.VGND
flabel metal1 3801 2703 3835 2737 0 FreeSans 200 0 0 0 FILLER_0_29.VPWR
flabel nwell 3801 2703 3835 2737 0 FreeSans 200 0 0 0 FILLER_0_29.VPB
flabel pwell 3801 2159 3835 2193 0 FreeSans 200 0 0 0 FILLER_0_29.VNB
rlabel comment 3772 2176 3772 2176 4 FILLER_0_29.decap_4
flabel metal1 4162 2703 4198 2733 0 FreeSans 250 0 0 0 FILLER_0_33.VPWR
flabel metal1 4162 2163 4198 2192 0 FreeSans 250 0 0 0 FILLER_0_33.VGND
flabel nwell 4171 2710 4191 2727 0 FreeSans 200 0 0 0 FILLER_0_33.VPB
flabel pwell 4168 2165 4192 2187 0 FreeSans 200 0 0 0 FILLER_0_33.VNB
rlabel comment 4140 2176 4140 2176 4 FILLER_0_33.fill_1
flabel metal1 3801 3247 3835 3281 0 FreeSans 200 0 0 0 FILLER_1_29.VGND
flabel metal1 3801 2703 3835 2737 0 FreeSans 200 0 0 0 FILLER_1_29.VPWR
flabel nwell 3801 2703 3835 2737 0 FreeSans 200 0 0 0 FILLER_1_29.VPB
flabel pwell 3801 3247 3835 3281 0 FreeSans 200 0 0 0 FILLER_1_29.VNB
rlabel comment 3772 3264 3772 3264 2 FILLER_1_29.decap_4
flabel metal1 3702 2700 3755 2729 0 FreeSans 200 0 0 0 TAP_20.VPWR
flabel metal1 3701 2158 3752 2196 0 FreeSans 200 0 0 0 TAP_20.VGND
rlabel comment 3680 2176 3680 2176 4 TAP_20.tapvpwrvgnd_1
flabel locali 6008 2601 6042 2635 0 FreeSans 400 0 0 0 _55_.Q
flabel locali 6008 2533 6042 2567 0 FreeSans 400 0 0 0 _55_.Q
flabel locali 6008 2465 6042 2499 0 FreeSans 400 0 0 0 _55_.Q
flabel locali 6008 2261 6042 2295 0 FreeSans 400 0 0 0 _55_.Q
flabel locali 5713 2329 5747 2363 0 FreeSans 400 0 0 0 _55_.RESET_B
flabel locali 4537 2465 4571 2499 0 FreeSans 400 0 0 0 _55_.D
flabel locali 4262 2465 4296 2499 0 FreeSans 400 0 0 0 _55_.CLK
flabel locali 4262 2397 4296 2431 0 FreeSans 400 0 0 0 _55_.CLK
flabel locali 5713 2397 5747 2431 0 FreeSans 400 0 0 0 _55_.RESET_B
flabel metal1 4261 2159 4295 2193 0 FreeSans 200 0 0 0 _55_.VGND
flabel metal1 4261 2703 4295 2737 0 FreeSans 200 0 0 0 _55_.VPWR
flabel nwell 4261 2703 4295 2737 0 FreeSans 200 0 0 0 _55_.VPB
flabel pwell 4261 2159 4295 2193 0 FreeSans 200 0 0 0 _55_.VNB
rlabel comment 4232 2176 4232 2176 4 _55_.dfrtp_1
flabel locali 4542 2941 4576 2975 0 FreeSans 200 0 0 0 _60_.D
flabel locali 4542 3009 4576 3043 0 FreeSans 200 0 0 0 _60_.D
flabel locali 4169 2703 4203 2737 3 FreeSans 400 0 0 0 _60_.VPWR
flabel locali 5934 2805 5968 2839 0 FreeSans 400 0 0 0 _60_.Q
flabel locali 5934 2873 5968 2907 0 FreeSans 400 0 0 0 _60_.Q
flabel locali 5934 3145 5968 3179 0 FreeSans 400 0 0 0 _60_.Q
flabel locali 4910 3077 4944 3111 0 FreeSans 400 0 0 0 _60_.SET_B
flabel locali 4170 2941 4204 2975 0 FreeSans 400 0 0 0 _60_.CLK
flabel locali 4170 3009 4204 3043 0 FreeSans 400 0 0 0 _60_.CLK
flabel locali 4169 3247 4203 3281 3 FreeSans 400 0 0 0 _60_.VGND
flabel nwell 4169 2703 4203 2737 0 FreeSans 200 0 0 0 _60_.VPB
flabel nwell 4186 2720 4186 2720 3 FreeSans 400 0 0 0 _60_.VPB
flabel pwell 4169 3247 4203 3281 0 FreeSans 200 0 0 0 _60_.VNB
flabel pwell 4186 3264 4186 3264 3 FreeSans 400 0 0 0 _60_.VNB
flabel metal1 4169 2703 4203 2737 0 FreeSans 200 0 0 0 _60_.VPWR
flabel metal1 4169 3247 4203 3281 0 FreeSans 200 0 0 0 _60_.VGND
rlabel comment 4140 3264 4140 3264 2 _60_.dfstp_1
flabel metal1 6092 2162 6145 2194 0 FreeSans 200 0 0 0 FILLER_0_54.VGND
flabel metal1 6093 2706 6145 2737 0 FreeSans 200 0 0 0 FILLER_0_54.VPWR
flabel nwell 6100 2711 6134 2729 0 FreeSans 200 0 0 0 FILLER_0_54.VPB
flabel pwell 6103 2166 6135 2188 0 FreeSans 200 0 0 0 FILLER_0_54.VNB
rlabel comment 6072 2176 6072 2176 4 FILLER_0_54.fill_2
flabel metal1 6377 2159 6411 2193 0 FreeSans 200 0 0 0 FILLER_0_57.VGND
flabel metal1 6377 2703 6411 2737 0 FreeSans 200 0 0 0 FILLER_0_57.VPWR
flabel nwell 6377 2703 6411 2737 0 FreeSans 200 0 0 0 FILLER_0_57.VPB
flabel pwell 6377 2159 6411 2193 0 FreeSans 200 0 0 0 FILLER_0_57.VNB
rlabel comment 6348 2176 6348 2176 4 FILLER_0_57.decap_12
flabel metal1 6092 3246 6145 3278 0 FreeSans 200 0 0 0 FILLER_1_54.VGND
flabel metal1 6093 2703 6145 2734 0 FreeSans 200 0 0 0 FILLER_1_54.VPWR
flabel nwell 6100 2711 6134 2729 0 FreeSans 200 0 0 0 FILLER_1_54.VPB
flabel pwell 6103 3252 6135 3274 0 FreeSans 200 0 0 0 FILLER_1_54.VNB
rlabel comment 6072 3264 6072 3264 2 FILLER_1_54.fill_2
flabel metal1 6377 2703 6411 2737 0 FreeSans 200 0 0 0 FILLER_1_57.VPWR
flabel metal1 6377 3247 6411 3281 0 FreeSans 200 0 0 0 FILLER_1_57.VGND
flabel nwell 6377 2703 6411 2737 0 FreeSans 200 0 0 0 FILLER_1_57.VPB
flabel pwell 6377 3247 6411 3281 0 FreeSans 200 0 0 0 FILLER_1_57.VNB
rlabel comment 6348 3264 6348 3264 2 FILLER_1_57.decap_8
flabel metal1 7106 2707 7142 2737 0 FreeSans 250 0 0 0 FILLER_1_65.VPWR
flabel metal1 7106 3248 7142 3277 0 FreeSans 250 0 0 0 FILLER_1_65.VGND
flabel nwell 7115 2713 7135 2730 0 FreeSans 200 0 0 0 FILLER_1_65.VPB
flabel pwell 7112 3253 7136 3275 0 FreeSans 200 0 0 0 FILLER_1_65.VNB
rlabel comment 7084 3264 7084 3264 2 FILLER_1_65.fill_1
flabel metal1 6278 2700 6331 2729 0 FreeSans 200 0 0 0 TAP_21.VPWR
flabel metal1 6277 2158 6328 2196 0 FreeSans 200 0 0 0 TAP_21.VGND
rlabel comment 6256 2176 6256 2176 4 TAP_21.tapvpwrvgnd_1
flabel metal1 6278 2711 6331 2740 0 FreeSans 200 0 0 0 TAP_26.VPWR
flabel metal1 6277 3244 6328 3282 0 FreeSans 200 0 0 0 TAP_26.VGND
rlabel comment 6256 3264 6256 3264 2 TAP_26.tapvpwrvgnd_1
flabel metal1 7481 2159 7515 2193 0 FreeSans 200 0 0 0 FILLER_0_69.VGND
flabel metal1 7481 2703 7515 2737 0 FreeSans 200 0 0 0 FILLER_0_69.VPWR
flabel nwell 7481 2703 7515 2737 0 FreeSans 200 0 0 0 FILLER_0_69.VPB
flabel pwell 7481 2159 7515 2193 0 FreeSans 200 0 0 0 FILLER_0_69.VNB
rlabel comment 7452 2176 7452 2176 4 FILLER_0_69.decap_12
flabel metal1 8585 2703 8619 2737 0 FreeSans 200 0 0 0 FILLER_0_81.VPWR
flabel metal1 8585 2159 8619 2193 0 FreeSans 200 0 0 0 FILLER_0_81.VGND
flabel nwell 8585 2703 8619 2737 0 FreeSans 200 0 0 0 FILLER_0_81.VPB
flabel pwell 8585 2159 8619 2193 0 FreeSans 200 0 0 0 FILLER_0_81.VNB
rlabel comment 8556 2176 8556 2176 4 FILLER_0_81.decap_3
flabel metal1 8944 2162 8997 2194 0 FreeSans 200 0 0 0 FILLER_0_85.VGND
flabel metal1 8945 2706 8997 2737 0 FreeSans 200 0 0 0 FILLER_0_85.VPWR
flabel nwell 8952 2711 8986 2729 0 FreeSans 200 0 0 0 FILLER_0_85.VPB
flabel pwell 8955 2166 8987 2188 0 FreeSans 200 0 0 0 FILLER_0_85.VNB
rlabel comment 8924 2176 8924 2176 4 FILLER_0_85.fill_2
flabel metal1 9045 3247 9079 3281 0 FreeSans 200 0 0 0 FILLER_1_86.VGND
flabel metal1 9045 2703 9079 2737 0 FreeSans 200 0 0 0 FILLER_1_86.VPWR
flabel nwell 9045 2703 9079 2737 0 FreeSans 200 0 0 0 FILLER_1_86.VPB
flabel pwell 9045 3247 9079 3281 0 FreeSans 200 0 0 0 FILLER_1_86.VNB
rlabel comment 9016 3264 9016 3264 2 FILLER_1_86.decap_4
flabel metal1 8854 2700 8907 2729 0 FreeSans 200 0 0 0 TAP_22.VPWR
flabel metal1 8853 2158 8904 2196 0 FreeSans 200 0 0 0 TAP_22.VGND
rlabel comment 8832 2176 8832 2176 4 TAP_22.tapvpwrvgnd_1
flabel locali 7206 2805 7240 2839 0 FreeSans 400 0 0 0 _56_.Q
flabel locali 7206 2873 7240 2907 0 FreeSans 400 0 0 0 _56_.Q
flabel locali 7206 2941 7240 2975 0 FreeSans 400 0 0 0 _56_.Q
flabel locali 7206 3145 7240 3179 0 FreeSans 400 0 0 0 _56_.Q
flabel locali 7501 3077 7535 3111 0 FreeSans 400 0 0 0 _56_.RESET_B
flabel locali 8677 2941 8711 2975 0 FreeSans 400 0 0 0 _56_.D
flabel locali 8952 2941 8986 2975 0 FreeSans 400 0 0 0 _56_.CLK
flabel locali 8952 3009 8986 3043 0 FreeSans 400 0 0 0 _56_.CLK
flabel locali 7501 3009 7535 3043 0 FreeSans 400 0 0 0 _56_.RESET_B
flabel metal1 8953 3247 8987 3281 0 FreeSans 200 0 0 0 _56_.VGND
flabel metal1 8953 2703 8987 2737 0 FreeSans 200 0 0 0 _56_.VPWR
flabel nwell 8953 2703 8987 2737 0 FreeSans 200 0 0 0 _56_.VPB
flabel pwell 8953 3247 8987 3281 0 FreeSans 200 0 0 0 _56_.VNB
rlabel comment 9016 3264 9016 3264 8 _56_.dfrtp_1
flabel locali 9138 2601 9172 2635 0 FreeSans 400 0 0 0 _57_.Q
flabel locali 9138 2533 9172 2567 0 FreeSans 400 0 0 0 _57_.Q
flabel locali 9138 2465 9172 2499 0 FreeSans 400 0 0 0 _57_.Q
flabel locali 9138 2261 9172 2295 0 FreeSans 400 0 0 0 _57_.Q
flabel locali 9433 2329 9467 2363 0 FreeSans 400 0 0 0 _57_.RESET_B
flabel locali 10609 2465 10643 2499 0 FreeSans 400 0 0 0 _57_.D
flabel locali 10884 2465 10918 2499 0 FreeSans 400 0 0 0 _57_.CLK
flabel locali 10884 2397 10918 2431 0 FreeSans 400 0 0 0 _57_.CLK
flabel locali 9433 2397 9467 2431 0 FreeSans 400 0 0 0 _57_.RESET_B
flabel metal1 10885 2159 10919 2193 0 FreeSans 200 0 0 0 _57_.VGND
flabel metal1 10885 2703 10919 2737 0 FreeSans 200 0 0 0 _57_.VPWR
flabel nwell 10885 2703 10919 2737 0 FreeSans 200 0 0 0 _57_.VPB
flabel pwell 10885 2159 10919 2193 0 FreeSans 200 0 0 0 _57_.VNB
rlabel comment 10948 2176 10948 2176 6 _57_.dfrtp_1
flabel metal1 10977 2159 11011 2193 0 FreeSans 200 0 0 0 FILLER_0_107.VGND
flabel metal1 10977 2703 11011 2737 0 FreeSans 200 0 0 0 FILLER_0_107.VPWR
flabel nwell 10977 2703 11011 2737 0 FreeSans 200 0 0 0 FILLER_0_107.VPB
flabel pwell 10977 2159 11011 2193 0 FreeSans 200 0 0 0 FILLER_0_107.VNB
rlabel comment 10948 2176 10948 2176 4 FILLER_0_107.decap_4
flabel locali 10977 2941 11011 2975 0 FreeSans 200 0 0 0 clkbuf_1_1__f_clk.X
flabel locali 11069 2941 11103 2975 0 FreeSans 200 0 0 0 clkbuf_1_1__f_clk.X
flabel locali 11069 3009 11103 3043 0 FreeSans 200 0 0 0 clkbuf_1_1__f_clk.X
flabel locali 10977 3009 11011 3043 0 FreeSans 200 0 0 0 clkbuf_1_1__f_clk.X
flabel locali 10977 3077 11011 3111 0 FreeSans 200 0 0 0 clkbuf_1_1__f_clk.X
flabel locali 11069 3077 11103 3111 0 FreeSans 200 0 0 0 clkbuf_1_1__f_clk.X
flabel locali 9413 3077 9447 3111 0 FreeSans 200 0 0 0 clkbuf_1_1__f_clk.A
flabel locali 9413 3009 9447 3043 0 FreeSans 200 0 0 0 clkbuf_1_1__f_clk.A
flabel pwell 9413 3247 9447 3281 0 FreeSans 200 0 0 0 clkbuf_1_1__f_clk.VNB
flabel pwell 9430 3264 9430 3264 0 FreeSans 200 0 0 0 clkbuf_1_1__f_clk.VNB
flabel nwell 9413 2703 9447 2737 0 FreeSans 200 0 0 0 clkbuf_1_1__f_clk.VPB
flabel nwell 9430 2720 9430 2720 0 FreeSans 200 0 0 0 clkbuf_1_1__f_clk.VPB
flabel metal1 9413 3247 9447 3281 0 FreeSans 200 0 0 0 clkbuf_1_1__f_clk.VGND
flabel metal1 9413 2703 9447 2737 0 FreeSans 200 0 0 0 clkbuf_1_1__f_clk.VPWR
rlabel comment 9384 3264 9384 3264 2 clkbuf_1_1__f_clk.clkbuf_16
flabel metal1 11338 2703 11374 2733 0 FreeSans 250 0 0 0 FILLER_0_111.VPWR
flabel metal1 11338 2163 11374 2192 0 FreeSans 250 0 0 0 FILLER_0_111.VGND
flabel nwell 11347 2710 11367 2727 0 FreeSans 200 0 0 0 FILLER_0_111.VPB
flabel pwell 11344 2165 11368 2187 0 FreeSans 200 0 0 0 FILLER_0_111.VNB
rlabel comment 11316 2176 11316 2176 4 FILLER_0_111.fill_1
flabel metal1 11529 2159 11563 2193 0 FreeSans 200 0 0 0 FILLER_0_113.VGND
flabel metal1 11529 2703 11563 2737 0 FreeSans 200 0 0 0 FILLER_0_113.VPWR
flabel nwell 11529 2703 11563 2737 0 FreeSans 200 0 0 0 FILLER_0_113.VPB
flabel pwell 11529 2159 11563 2193 0 FreeSans 200 0 0 0 FILLER_0_113.VNB
rlabel comment 11500 2176 11500 2176 4 FILLER_0_113.decap_4
flabel metal1 11890 2703 11926 2733 0 FreeSans 250 0 0 0 FILLER_0_117.VPWR
flabel metal1 11890 2163 11926 2192 0 FreeSans 250 0 0 0 FILLER_0_117.VGND
flabel nwell 11899 2710 11919 2727 0 FreeSans 200 0 0 0 FILLER_0_117.VPB
flabel pwell 11896 2165 11920 2187 0 FreeSans 200 0 0 0 FILLER_0_117.VNB
rlabel comment 11868 2176 11868 2176 4 FILLER_0_117.fill_1
flabel metal1 11244 3246 11297 3278 0 FreeSans 200 0 0 0 FILLER_1_110.VGND
flabel metal1 11245 2703 11297 2734 0 FreeSans 200 0 0 0 FILLER_1_110.VPWR
flabel nwell 11252 2711 11286 2729 0 FreeSans 200 0 0 0 FILLER_1_110.VPB
flabel pwell 11255 3252 11287 3274 0 FreeSans 200 0 0 0 FILLER_1_110.VNB
rlabel comment 11224 3264 11224 3264 2 FILLER_1_110.fill_2
flabel metal1 11520 3246 11573 3278 0 FreeSans 200 0 0 0 FILLER_1_113.VGND
flabel metal1 11521 2703 11573 2734 0 FreeSans 200 0 0 0 FILLER_1_113.VPWR
flabel nwell 11528 2711 11562 2729 0 FreeSans 200 0 0 0 FILLER_1_113.VPB
flabel pwell 11531 3252 11563 3274 0 FreeSans 200 0 0 0 FILLER_1_113.VNB
rlabel comment 11500 3264 11500 3264 2 FILLER_1_113.fill_2
flabel metal1 11430 2700 11483 2729 0 FreeSans 200 0 0 0 TAP_23.VPWR
flabel metal1 11429 2158 11480 2196 0 FreeSans 200 0 0 0 TAP_23.VGND
rlabel comment 11408 2176 11408 2176 4 TAP_23.tapvpwrvgnd_1
flabel metal1 11430 2711 11483 2740 0 FreeSans 200 0 0 0 TAP_27.VPWR
flabel metal1 11429 3244 11480 3282 0 FreeSans 200 0 0 0 TAP_27.VGND
rlabel comment 11408 3264 11408 3264 2 TAP_27.tapvpwrvgnd_1
flabel locali 11990 2601 12024 2635 0 FreeSans 400 0 0 0 _64_.Q
flabel locali 11990 2533 12024 2567 0 FreeSans 400 0 0 0 _64_.Q
flabel locali 11990 2465 12024 2499 0 FreeSans 400 0 0 0 _64_.Q
flabel locali 11990 2261 12024 2295 0 FreeSans 400 0 0 0 _64_.Q
flabel locali 12285 2329 12319 2363 0 FreeSans 400 0 0 0 _64_.RESET_B
flabel locali 13461 2465 13495 2499 0 FreeSans 400 0 0 0 _64_.D
flabel locali 13736 2465 13770 2499 0 FreeSans 400 0 0 0 _64_.CLK
flabel locali 13736 2397 13770 2431 0 FreeSans 400 0 0 0 _64_.CLK
flabel locali 12285 2397 12319 2431 0 FreeSans 400 0 0 0 _64_.RESET_B
flabel metal1 13737 2159 13771 2193 0 FreeSans 200 0 0 0 _64_.VGND
flabel metal1 13737 2703 13771 2737 0 FreeSans 200 0 0 0 _64_.VPWR
flabel nwell 13737 2703 13771 2737 0 FreeSans 200 0 0 0 _64_.VPB
flabel pwell 13737 2159 13771 2193 0 FreeSans 200 0 0 0 _64_.VNB
rlabel comment 13800 2176 13800 2176 6 _64_.dfrtp_1
flabel locali 11714 2805 11748 2839 0 FreeSans 400 0 0 0 _65_.Q
flabel locali 11714 2873 11748 2907 0 FreeSans 400 0 0 0 _65_.Q
flabel locali 11714 2941 11748 2975 0 FreeSans 400 0 0 0 _65_.Q
flabel locali 11714 3145 11748 3179 0 FreeSans 400 0 0 0 _65_.Q
flabel locali 12009 3077 12043 3111 0 FreeSans 400 0 0 0 _65_.RESET_B
flabel locali 13185 2941 13219 2975 0 FreeSans 400 0 0 0 _65_.D
flabel locali 13460 2941 13494 2975 0 FreeSans 400 0 0 0 _65_.CLK
flabel locali 13460 3009 13494 3043 0 FreeSans 400 0 0 0 _65_.CLK
flabel locali 12009 3009 12043 3043 0 FreeSans 400 0 0 0 _65_.RESET_B
flabel metal1 13461 3247 13495 3281 0 FreeSans 200 0 0 0 _65_.VGND
flabel metal1 13461 2703 13495 2737 0 FreeSans 200 0 0 0 _65_.VPWR
flabel nwell 13461 2703 13495 2737 0 FreeSans 200 0 0 0 _65_.VPB
flabel pwell 13461 3247 13495 3281 0 FreeSans 200 0 0 0 _65_.VNB
rlabel comment 13524 3264 13524 3264 8 _65_.dfrtp_1
flabel metal1 13820 2162 13873 2194 0 FreeSans 200 0 0 0 FILLER_0_138.VGND
flabel metal1 13821 2706 13873 2737 0 FreeSans 200 0 0 0 FILLER_0_138.VPWR
flabel nwell 13828 2711 13862 2729 0 FreeSans 200 0 0 0 FILLER_0_138.VPB
flabel pwell 13831 2166 13863 2188 0 FreeSans 200 0 0 0 FILLER_0_138.VNB
rlabel comment 13800 2176 13800 2176 4 FILLER_0_138.fill_2
flabel metal1 14096 2162 14149 2194 0 FreeSans 200 0 0 0 FILLER_0_141.VGND
flabel metal1 14097 2706 14149 2737 0 FreeSans 200 0 0 0 FILLER_0_141.VPWR
flabel nwell 14104 2711 14138 2729 0 FreeSans 200 0 0 0 FILLER_0_141.VPB
flabel pwell 14107 2166 14139 2188 0 FreeSans 200 0 0 0 FILLER_0_141.VNB
rlabel comment 14076 2176 14076 2176 4 FILLER_0_141.fill_2
flabel metal1 13553 3247 13587 3281 0 FreeSans 200 0 0 0 FILLER_1_135.VGND
flabel metal1 13553 2703 13587 2737 0 FreeSans 200 0 0 0 FILLER_1_135.VPWR
flabel nwell 13553 2703 13587 2737 0 FreeSans 200 0 0 0 FILLER_1_135.VPB
flabel pwell 13553 3247 13587 3281 0 FreeSans 200 0 0 0 FILLER_1_135.VNB
rlabel comment 13524 3264 13524 3264 2 FILLER_1_135.decap_4
flabel metal1 14289 3247 14323 3281 0 FreeSans 200 0 0 0 FILLER_1_143.VGND
flabel metal1 14289 2703 14323 2737 0 FreeSans 200 0 0 0 FILLER_1_143.VPWR
flabel nwell 14289 2703 14323 2737 0 FreeSans 200 0 0 0 FILLER_1_143.VPB
flabel pwell 14289 3247 14323 3281 0 FreeSans 200 0 0 0 FILLER_1_143.VNB
rlabel comment 14260 3264 14260 3264 2 FILLER_1_143.decap_12
flabel metal1 14006 2700 14059 2729 0 FreeSans 200 0 0 0 TAP_24.VPWR
flabel metal1 14005 2158 14056 2196 0 FreeSans 200 0 0 0 TAP_24.VGND
rlabel comment 13984 2176 13984 2176 4 TAP_24.tapvpwrvgnd_1
flabel locali 14290 2601 14324 2635 0 FreeSans 400 0 0 0 _59_.Q
flabel locali 14290 2533 14324 2567 0 FreeSans 400 0 0 0 _59_.Q
flabel locali 14290 2465 14324 2499 0 FreeSans 400 0 0 0 _59_.Q
flabel locali 14290 2261 14324 2295 0 FreeSans 400 0 0 0 _59_.Q
flabel locali 14585 2329 14619 2363 0 FreeSans 400 0 0 0 _59_.RESET_B
flabel locali 15761 2465 15795 2499 0 FreeSans 400 0 0 0 _59_.D
flabel locali 16036 2465 16070 2499 0 FreeSans 400 0 0 0 _59_.CLK
flabel locali 16036 2397 16070 2431 0 FreeSans 400 0 0 0 _59_.CLK
flabel locali 14585 2397 14619 2431 0 FreeSans 400 0 0 0 _59_.RESET_B
flabel metal1 16037 2159 16071 2193 0 FreeSans 200 0 0 0 _59_.VGND
flabel metal1 16037 2703 16071 2737 0 FreeSans 200 0 0 0 _59_.VPWR
flabel nwell 16037 2703 16071 2737 0 FreeSans 200 0 0 0 _59_.VPB
flabel pwell 16037 2159 16071 2193 0 FreeSans 200 0 0 0 _59_.VNB
rlabel comment 16100 2176 16100 2176 6 _59_.dfrtp_1
flabel metal1 13921 2703 13955 2737 0 FreeSans 200 0 0 0 output12.VPWR
flabel metal1 13921 3247 13955 3281 0 FreeSans 200 0 0 0 output12.VGND
flabel locali 13921 2703 13955 2737 0 FreeSans 200 0 0 0 output12.VPWR
flabel locali 13921 3247 13955 3281 0 FreeSans 200 0 0 0 output12.VGND
flabel locali 14104 3145 14138 3179 0 FreeSans 200 0 0 0 output12.X
flabel locali 14104 2873 14138 2907 0 FreeSans 200 0 0 0 output12.X
flabel locali 14104 2805 14138 2839 0 FreeSans 200 0 0 0 output12.X
flabel locali 13921 3009 13955 3043 0 FreeSans 200 0 0 0 output12.A
flabel nwell 13921 2703 13955 2737 0 FreeSans 200 0 0 0 output12.VPB
flabel pwell 13921 3247 13955 3281 0 FreeSans 200 0 0 0 output12.VNB
rlabel comment 13892 3264 13892 3264 2 output12.buf_2
flabel metal1 16129 2159 16163 2193 0 FreeSans 200 0 0 0 FILLER_0_163.VGND
flabel metal1 16129 2703 16163 2737 0 FreeSans 200 0 0 0 FILLER_0_163.VPWR
flabel nwell 16129 2703 16163 2737 0 FreeSans 200 0 0 0 FILLER_0_163.VPB
flabel pwell 16129 2159 16163 2193 0 FreeSans 200 0 0 0 FILLER_0_163.VNB
rlabel comment 16100 2176 16100 2176 4 FILLER_0_163.decap_4
flabel metal1 16490 2703 16526 2733 0 FreeSans 250 0 0 0 FILLER_0_167.VPWR
flabel metal1 16490 2163 16526 2192 0 FreeSans 250 0 0 0 FILLER_0_167.VGND
flabel nwell 16499 2710 16519 2727 0 FreeSans 200 0 0 0 FILLER_0_167.VPB
flabel pwell 16496 2165 16520 2187 0 FreeSans 200 0 0 0 FILLER_0_167.VNB
rlabel comment 16468 2176 16468 2176 4 FILLER_0_167.fill_1
flabel metal1 16681 2703 16715 2737 0 FreeSans 200 0 0 0 FILLER_0_169.VPWR
flabel metal1 16681 2159 16715 2193 0 FreeSans 200 0 0 0 FILLER_0_169.VGND
flabel nwell 16681 2703 16715 2737 0 FreeSans 200 0 0 0 FILLER_0_169.VPB
flabel pwell 16681 2159 16715 2193 0 FreeSans 200 0 0 0 FILLER_0_169.VNB
rlabel comment 16652 2176 16652 2176 4 FILLER_0_169.decap_8
flabel metal1 15393 3247 15427 3281 0 FreeSans 200 0 0 0 FILLER_1_155.VGND
flabel metal1 15393 2703 15427 2737 0 FreeSans 200 0 0 0 FILLER_1_155.VPWR
flabel nwell 15393 2703 15427 2737 0 FreeSans 200 0 0 0 FILLER_1_155.VPB
flabel pwell 15393 3247 15427 3281 0 FreeSans 200 0 0 0 FILLER_1_155.VNB
rlabel comment 15364 3264 15364 3264 2 FILLER_1_155.decap_12
flabel metal1 16490 2707 16526 2737 0 FreeSans 250 0 0 0 FILLER_1_167.VPWR
flabel metal1 16490 3248 16526 3277 0 FreeSans 250 0 0 0 FILLER_1_167.VGND
flabel nwell 16499 2713 16519 2730 0 FreeSans 200 0 0 0 FILLER_1_167.VPB
flabel pwell 16496 3253 16520 3275 0 FreeSans 200 0 0 0 FILLER_1_167.VNB
rlabel comment 16468 3264 16468 3264 2 FILLER_1_167.fill_1
flabel metal1 16681 3247 16715 3281 0 FreeSans 200 0 0 0 FILLER_1_169.VGND
flabel metal1 16681 2703 16715 2737 0 FreeSans 200 0 0 0 FILLER_1_169.VPWR
flabel nwell 16681 2703 16715 2737 0 FreeSans 200 0 0 0 FILLER_1_169.VPB
flabel pwell 16681 3247 16715 3281 0 FreeSans 200 0 0 0 FILLER_1_169.VNB
rlabel comment 16652 3264 16652 3264 2 FILLER_1_169.decap_12
flabel metal1 16582 2700 16635 2729 0 FreeSans 200 0 0 0 TAP_25.VPWR
flabel metal1 16581 2158 16632 2196 0 FreeSans 200 0 0 0 TAP_25.VGND
rlabel comment 16560 2176 16560 2176 4 TAP_25.tapvpwrvgnd_1
flabel metal1 16582 2711 16635 2740 0 FreeSans 200 0 0 0 TAP_28.VPWR
flabel metal1 16581 3244 16632 3282 0 FreeSans 200 0 0 0 TAP_28.VGND
rlabel comment 16560 3264 16560 3264 2 TAP_28.tapvpwrvgnd_1
flabel metal1 17410 2703 17446 2733 0 FreeSans 250 0 0 0 FILLER_0_177.VPWR
flabel metal1 17410 2163 17446 2192 0 FreeSans 250 0 0 0 FILLER_0_177.VGND
flabel nwell 17419 2710 17439 2727 0 FreeSans 200 0 0 0 FILLER_0_177.VPB
flabel pwell 17416 2165 17440 2187 0 FreeSans 200 0 0 0 FILLER_0_177.VNB
rlabel comment 17388 2176 17388 2176 4 FILLER_0_177.fill_1
flabel metal1 17877 2703 17911 2737 0 FreeSans 200 0 0 0 FILLER_0_182.VPWR
flabel metal1 17877 2159 17911 2193 0 FreeSans 200 0 0 0 FILLER_0_182.VGND
flabel nwell 17877 2703 17911 2737 0 FreeSans 200 0 0 0 FILLER_0_182.VPB
flabel pwell 17877 2159 17911 2193 0 FreeSans 200 0 0 0 FILLER_0_182.VNB
rlabel comment 17848 2176 17848 2176 4 FILLER_0_182.decap_8
flabel metal1 17785 2703 17819 2737 0 FreeSans 200 0 0 0 FILLER_1_181.VPWR
flabel metal1 17785 3247 17819 3281 0 FreeSans 200 0 0 0 FILLER_1_181.VGND
flabel nwell 17785 2703 17819 2737 0 FreeSans 200 0 0 0 FILLER_1_181.VPB
flabel pwell 17785 3247 17819 3281 0 FreeSans 200 0 0 0 FILLER_1_181.VNB
rlabel comment 17756 3264 17756 3264 2 FILLER_1_181.decap_8
flabel metal1 18514 2707 18550 2737 0 FreeSans 250 0 0 0 FILLER_1_189.VPWR
flabel metal1 18514 3248 18550 3277 0 FreeSans 250 0 0 0 FILLER_1_189.VGND
flabel nwell 18523 2713 18543 2730 0 FreeSans 200 0 0 0 FILLER_1_189.VPB
flabel pwell 18520 3253 18544 3275 0 FreeSans 200 0 0 0 FILLER_1_189.VNB
rlabel comment 18492 3264 18492 3264 2 FILLER_1_189.fill_1
flabel metal1 18797 2703 18831 2737 0 FreeSans 200 0 0 0 PHY_1.VPWR
flabel metal1 18797 2159 18831 2193 0 FreeSans 200 0 0 0 PHY_1.VGND
flabel nwell 18797 2703 18831 2737 0 FreeSans 200 0 0 0 PHY_1.VPB
flabel pwell 18797 2159 18831 2193 0 FreeSans 200 0 0 0 PHY_1.VNB
rlabel comment 18860 2176 18860 2176 6 PHY_1.decap_3
flabel metal1 18797 2703 18831 2737 0 FreeSans 200 0 0 0 PHY_3.VPWR
flabel metal1 18797 3247 18831 3281 0 FreeSans 200 0 0 0 PHY_3.VGND
flabel nwell 18797 2703 18831 2737 0 FreeSans 200 0 0 0 PHY_3.VPB
flabel pwell 18797 3247 18831 3281 0 FreeSans 200 0 0 0 PHY_3.VNB
rlabel comment 18860 3264 18860 3264 8 PHY_3.decap_3
flabel metal1 17509 2703 17543 2737 0 FreeSans 200 0 0 0 output11.VPWR
flabel metal1 17509 2159 17543 2193 0 FreeSans 200 0 0 0 output11.VGND
flabel locali 17509 2703 17543 2737 0 FreeSans 200 0 0 0 output11.VPWR
flabel locali 17509 2159 17543 2193 0 FreeSans 200 0 0 0 output11.VGND
flabel locali 17692 2261 17726 2295 0 FreeSans 200 0 0 0 output11.X
flabel locali 17692 2533 17726 2567 0 FreeSans 200 0 0 0 output11.X
flabel locali 17692 2601 17726 2635 0 FreeSans 200 0 0 0 output11.X
flabel locali 17509 2397 17543 2431 0 FreeSans 200 0 0 0 output11.A
flabel nwell 17509 2703 17543 2737 0 FreeSans 200 0 0 0 output11.VPB
flabel pwell 17509 2159 17543 2193 0 FreeSans 200 0 0 0 output11.VNB
rlabel comment 17480 2176 17480 2176 4 output11.buf_2
flabel metal1 1409 3791 1443 3825 0 FreeSans 200 0 0 0 FILLER_2_3.VPWR
flabel metal1 1409 3247 1443 3281 0 FreeSans 200 0 0 0 FILLER_2_3.VGND
flabel nwell 1409 3791 1443 3825 0 FreeSans 200 0 0 0 FILLER_2_3.VPB
flabel pwell 1409 3247 1443 3281 0 FreeSans 200 0 0 0 FILLER_2_3.VNB
rlabel comment 1380 3264 1380 3264 4 FILLER_2_3.decap_3
flabel metal1 1133 3791 1167 3825 0 FreeSans 200 0 0 0 PHY_4.VPWR
flabel metal1 1133 3247 1167 3281 0 FreeSans 200 0 0 0 PHY_4.VGND
flabel nwell 1133 3791 1167 3825 0 FreeSans 200 0 0 0 PHY_4.VPB
flabel pwell 1133 3247 1167 3281 0 FreeSans 200 0 0 0 PHY_4.VNB
rlabel comment 1104 3264 1104 3264 4 PHY_4.decap_3
flabel locali 3432 3689 3466 3723 0 FreeSans 400 0 0 0 _51_.Q
flabel locali 3432 3621 3466 3655 0 FreeSans 400 0 0 0 _51_.Q
flabel locali 3432 3553 3466 3587 0 FreeSans 400 0 0 0 _51_.Q
flabel locali 3432 3349 3466 3383 0 FreeSans 400 0 0 0 _51_.Q
flabel locali 3137 3417 3171 3451 0 FreeSans 400 0 0 0 _51_.RESET_B
flabel locali 1961 3553 1995 3587 0 FreeSans 400 0 0 0 _51_.D
flabel locali 1686 3553 1720 3587 0 FreeSans 400 0 0 0 _51_.CLK
flabel locali 1686 3485 1720 3519 0 FreeSans 400 0 0 0 _51_.CLK
flabel locali 3137 3485 3171 3519 0 FreeSans 400 0 0 0 _51_.RESET_B
flabel metal1 1685 3247 1719 3281 0 FreeSans 200 0 0 0 _51_.VGND
flabel metal1 1685 3791 1719 3825 0 FreeSans 200 0 0 0 _51_.VPWR
flabel nwell 1685 3791 1719 3825 0 FreeSans 200 0 0 0 _51_.VPB
flabel pwell 1685 3247 1719 3281 0 FreeSans 200 0 0 0 _51_.VNB
rlabel comment 1656 3264 1656 3264 4 _51_.dfrtp_1
flabel metal1 3516 3250 3569 3282 0 FreeSans 200 0 0 0 FILLER_2_26.VGND
flabel metal1 3517 3794 3569 3825 0 FreeSans 200 0 0 0 FILLER_2_26.VPWR
flabel nwell 3524 3799 3558 3817 0 FreeSans 200 0 0 0 FILLER_2_26.VPB
flabel pwell 3527 3254 3559 3276 0 FreeSans 200 0 0 0 FILLER_2_26.VNB
rlabel comment 3496 3264 3496 3264 4 FILLER_2_26.fill_2
flabel metal1 3801 3791 3835 3825 0 FreeSans 200 0 0 0 FILLER_2_29.VPWR
flabel metal1 3801 3247 3835 3281 0 FreeSans 200 0 0 0 FILLER_2_29.VGND
flabel nwell 3801 3791 3835 3825 0 FreeSans 200 0 0 0 FILLER_2_29.VPB
flabel pwell 3801 3247 3835 3281 0 FreeSans 200 0 0 0 FILLER_2_29.VNB
rlabel comment 3772 3264 3772 3264 4 FILLER_2_29.decap_8
flabel metal1 3702 3788 3755 3817 0 FreeSans 200 0 0 0 TAP_29.VPWR
flabel metal1 3701 3246 3752 3284 0 FreeSans 200 0 0 0 TAP_29.VGND
rlabel comment 3680 3264 3680 3264 4 TAP_29.tapvpwrvgnd_1
flabel locali 4721 3553 4755 3587 0 FreeSans 200 0 0 0 clkbuf_1_0__f_clk.X
flabel locali 4629 3553 4663 3587 0 FreeSans 200 0 0 0 clkbuf_1_0__f_clk.X
flabel locali 4629 3485 4663 3519 0 FreeSans 200 0 0 0 clkbuf_1_0__f_clk.X
flabel locali 4721 3485 4755 3519 0 FreeSans 200 0 0 0 clkbuf_1_0__f_clk.X
flabel locali 4721 3417 4755 3451 0 FreeSans 200 0 0 0 clkbuf_1_0__f_clk.X
flabel locali 4629 3417 4663 3451 0 FreeSans 200 0 0 0 clkbuf_1_0__f_clk.X
flabel locali 6285 3417 6319 3451 0 FreeSans 200 0 0 0 clkbuf_1_0__f_clk.A
flabel locali 6285 3485 6319 3519 0 FreeSans 200 0 0 0 clkbuf_1_0__f_clk.A
flabel pwell 6285 3247 6319 3281 0 FreeSans 200 0 0 0 clkbuf_1_0__f_clk.VNB
flabel pwell 6302 3264 6302 3264 0 FreeSans 200 0 0 0 clkbuf_1_0__f_clk.VNB
flabel nwell 6285 3791 6319 3825 0 FreeSans 200 0 0 0 clkbuf_1_0__f_clk.VPB
flabel nwell 6302 3808 6302 3808 0 FreeSans 200 0 0 0 clkbuf_1_0__f_clk.VPB
flabel metal1 6285 3247 6319 3281 0 FreeSans 200 0 0 0 clkbuf_1_0__f_clk.VGND
flabel metal1 6285 3791 6319 3825 0 FreeSans 200 0 0 0 clkbuf_1_0__f_clk.VPWR
rlabel comment 6348 3264 6348 3264 6 clkbuf_1_0__f_clk.clkbuf_16
flabel metal1 6377 3247 6411 3281 0 FreeSans 200 0 0 0 FILLER_2_57.VGND
flabel metal1 6377 3791 6411 3825 0 FreeSans 200 0 0 0 FILLER_2_57.VPWR
flabel nwell 6377 3791 6411 3825 0 FreeSans 200 0 0 0 FILLER_2_57.VPB
flabel pwell 6377 3247 6411 3281 0 FreeSans 200 0 0 0 FILLER_2_57.VNB
rlabel comment 6348 3264 6348 3264 4 FILLER_2_57.decap_4
flabel locali 8492 3689 8526 3723 0 FreeSans 400 0 0 0 _50_.Q
flabel locali 8492 3621 8526 3655 0 FreeSans 400 0 0 0 _50_.Q
flabel locali 8492 3553 8526 3587 0 FreeSans 400 0 0 0 _50_.Q
flabel locali 8492 3349 8526 3383 0 FreeSans 400 0 0 0 _50_.Q
flabel locali 8197 3417 8231 3451 0 FreeSans 400 0 0 0 _50_.RESET_B
flabel locali 7021 3553 7055 3587 0 FreeSans 400 0 0 0 _50_.D
flabel locali 6746 3553 6780 3587 0 FreeSans 400 0 0 0 _50_.CLK
flabel locali 6746 3485 6780 3519 0 FreeSans 400 0 0 0 _50_.CLK
flabel locali 8197 3485 8231 3519 0 FreeSans 400 0 0 0 _50_.RESET_B
flabel metal1 6745 3247 6779 3281 0 FreeSans 200 0 0 0 _50_.VGND
flabel metal1 6745 3791 6779 3825 0 FreeSans 200 0 0 0 _50_.VPWR
flabel nwell 6745 3791 6779 3825 0 FreeSans 200 0 0 0 _50_.VPB
flabel pwell 6745 3247 6779 3281 0 FreeSans 200 0 0 0 _50_.VNB
rlabel comment 6716 3264 6716 3264 4 _50_.dfrtp_1
flabel metal1 8585 3791 8619 3825 0 FreeSans 200 0 0 0 FILLER_2_81.VPWR
flabel metal1 8585 3247 8619 3281 0 FreeSans 200 0 0 0 FILLER_2_81.VGND
flabel nwell 8585 3791 8619 3825 0 FreeSans 200 0 0 0 FILLER_2_81.VPB
flabel pwell 8585 3247 8619 3281 0 FreeSans 200 0 0 0 FILLER_2_81.VNB
rlabel comment 8556 3264 8556 3264 4 FILLER_2_81.decap_3
flabel metal1 8944 3250 8997 3282 0 FreeSans 200 0 0 0 FILLER_2_85.VGND
flabel metal1 8945 3794 8997 3825 0 FreeSans 200 0 0 0 FILLER_2_85.VPWR
flabel nwell 8952 3799 8986 3817 0 FreeSans 200 0 0 0 FILLER_2_85.VPB
flabel pwell 8955 3254 8987 3276 0 FreeSans 200 0 0 0 FILLER_2_85.VNB
rlabel comment 8924 3264 8924 3264 4 FILLER_2_85.fill_2
flabel metal1 8854 3788 8907 3817 0 FreeSans 200 0 0 0 TAP_30.VPWR
flabel metal1 8853 3246 8904 3284 0 FreeSans 200 0 0 0 TAP_30.VGND
rlabel comment 8832 3264 8832 3264 4 TAP_30.tapvpwrvgnd_1
flabel metal1 9137 3791 9171 3825 0 FreeSans 200 0 0 0 fanout14.VPWR
flabel metal1 9137 3247 9171 3281 0 FreeSans 200 0 0 0 fanout14.VGND
flabel locali 9137 3791 9171 3825 0 FreeSans 200 0 0 0 fanout14.VPWR
flabel locali 9137 3247 9171 3281 0 FreeSans 200 0 0 0 fanout14.VGND
flabel locali 9320 3349 9354 3383 0 FreeSans 200 0 0 0 fanout14.X
flabel locali 9320 3621 9354 3655 0 FreeSans 200 0 0 0 fanout14.X
flabel locali 9320 3689 9354 3723 0 FreeSans 200 0 0 0 fanout14.X
flabel locali 9137 3485 9171 3519 0 FreeSans 200 0 0 0 fanout14.A
flabel nwell 9137 3791 9171 3825 0 FreeSans 200 0 0 0 fanout14.VPB
flabel pwell 9137 3247 9171 3281 0 FreeSans 200 0 0 0 fanout14.VNB
rlabel comment 9108 3264 9108 3264 4 fanout14.buf_2
flabel metal1 10333 3791 10367 3825 0 FreeSans 200 0 0 0 FILLER_2_100.VPWR
flabel metal1 10333 3247 10367 3281 0 FreeSans 200 0 0 0 FILLER_2_100.VGND
flabel nwell 10333 3791 10367 3825 0 FreeSans 200 0 0 0 FILLER_2_100.VPB
flabel pwell 10333 3247 10367 3281 0 FreeSans 200 0 0 0 FILLER_2_100.VNB
rlabel comment 10304 3264 10304 3264 4 FILLER_2_100.decap_6
flabel metal1 10878 3791 10914 3821 0 FreeSans 250 0 0 0 FILLER_2_106.VPWR
flabel metal1 10878 3251 10914 3280 0 FreeSans 250 0 0 0 FILLER_2_106.VGND
flabel nwell 10887 3798 10907 3815 0 FreeSans 200 0 0 0 FILLER_2_106.VPB
flabel pwell 10884 3253 10908 3275 0 FreeSans 200 0 0 0 FILLER_2_106.VNB
rlabel comment 10856 3264 10856 3264 4 FILLER_2_106.fill_1
flabel metal1 9505 3791 9539 3825 0 FreeSans 200 0 0 0 FILLER_2_91.VPWR
flabel metal1 9505 3247 9539 3281 0 FreeSans 200 0 0 0 FILLER_2_91.VGND
flabel nwell 9505 3791 9539 3825 0 FreeSans 200 0 0 0 FILLER_2_91.VPB
flabel pwell 9505 3247 9539 3281 0 FreeSans 200 0 0 0 FILLER_2_91.VNB
rlabel comment 9476 3264 9476 3264 4 FILLER_2_91.decap_6
flabel metal1 10977 3247 11011 3281 0 FreeSans 200 180 0 0 _27_.VGND
flabel metal1 10977 3791 11011 3825 0 FreeSans 200 180 0 0 _27_.VPWR
flabel locali 11161 3349 11195 3383 0 FreeSans 200 180 0 0 _27_.X
flabel locali 11161 3621 11195 3655 0 FreeSans 200 180 0 0 _27_.X
flabel locali 11161 3689 11195 3723 0 FreeSans 200 180 0 0 _27_.X
flabel locali 10977 3485 11011 3519 0 FreeSans 200 180 0 0 _27_.A
flabel nwell 10977 3791 11011 3825 0 FreeSans 200 180 0 0 _27_.VPB
flabel pwell 10977 3247 11011 3281 0 FreeSans 200 180 0 0 _27_.VNB
rlabel comment 11224 3264 11224 3264 6 _27_.clkbuf_1
flabel metal1 10241 3247 10275 3281 0 FreeSans 200 180 0 0 _48_.VGND
flabel metal1 10241 3791 10275 3825 0 FreeSans 200 180 0 0 _48_.VPWR
flabel locali 10057 3349 10091 3383 0 FreeSans 200 180 0 0 _48_.X
flabel locali 10057 3621 10091 3655 0 FreeSans 200 180 0 0 _48_.X
flabel locali 10057 3689 10091 3723 0 FreeSans 200 180 0 0 _48_.X
flabel locali 10241 3485 10275 3519 0 FreeSans 200 180 0 0 _48_.A
flabel nwell 10241 3791 10275 3825 0 FreeSans 200 180 0 0 _48_.VPB
flabel pwell 10241 3247 10275 3281 0 FreeSans 200 180 0 0 _48_.VNB
rlabel comment 10028 3264 10028 3264 4 _48_.clkbuf_1
flabel metal1 11253 3791 11287 3825 0 FreeSans 200 0 0 0 FILLER_2_110.VPWR
flabel metal1 11253 3247 11287 3281 0 FreeSans 200 0 0 0 FILLER_2_110.VGND
flabel nwell 11253 3791 11287 3825 0 FreeSans 200 0 0 0 FILLER_2_110.VPB
flabel pwell 11253 3247 11287 3281 0 FreeSans 200 0 0 0 FILLER_2_110.VNB
rlabel comment 11224 3264 11224 3264 4 FILLER_2_110.decap_8
flabel locali 11990 3689 12024 3723 0 FreeSans 400 0 0 0 _58_.Q
flabel locali 11990 3621 12024 3655 0 FreeSans 400 0 0 0 _58_.Q
flabel locali 11990 3553 12024 3587 0 FreeSans 400 0 0 0 _58_.Q
flabel locali 11990 3349 12024 3383 0 FreeSans 400 0 0 0 _58_.Q
flabel locali 12285 3417 12319 3451 0 FreeSans 400 0 0 0 _58_.RESET_B
flabel locali 13461 3553 13495 3587 0 FreeSans 400 0 0 0 _58_.D
flabel locali 13736 3553 13770 3587 0 FreeSans 400 0 0 0 _58_.CLK
flabel locali 13736 3485 13770 3519 0 FreeSans 400 0 0 0 _58_.CLK
flabel locali 12285 3485 12319 3519 0 FreeSans 400 0 0 0 _58_.RESET_B
flabel metal1 13737 3247 13771 3281 0 FreeSans 200 0 0 0 _58_.VGND
flabel metal1 13737 3791 13771 3825 0 FreeSans 200 0 0 0 _58_.VPWR
flabel nwell 13737 3791 13771 3825 0 FreeSans 200 0 0 0 _58_.VPB
flabel pwell 13737 3247 13771 3281 0 FreeSans 200 0 0 0 _58_.VNB
rlabel comment 13800 3264 13800 3264 6 _58_.dfrtp_1
flabel metal1 13820 3250 13873 3282 0 FreeSans 200 0 0 0 FILLER_2_138.VGND
flabel metal1 13821 3794 13873 3825 0 FreeSans 200 0 0 0 FILLER_2_138.VPWR
flabel nwell 13828 3799 13862 3817 0 FreeSans 200 0 0 0 FILLER_2_138.VPB
flabel pwell 13831 3254 13863 3276 0 FreeSans 200 0 0 0 FILLER_2_138.VNB
rlabel comment 13800 3264 13800 3264 4 FILLER_2_138.fill_2
flabel metal1 14105 3247 14139 3281 0 FreeSans 200 0 0 0 FILLER_2_141.VGND
flabel metal1 14105 3791 14139 3825 0 FreeSans 200 0 0 0 FILLER_2_141.VPWR
flabel nwell 14105 3791 14139 3825 0 FreeSans 200 0 0 0 FILLER_2_141.VPB
flabel pwell 14105 3247 14139 3281 0 FreeSans 200 0 0 0 FILLER_2_141.VNB
rlabel comment 14076 3264 14076 3264 4 FILLER_2_141.decap_12
flabel metal1 14006 3788 14059 3817 0 FreeSans 200 0 0 0 TAP_31.VPWR
flabel metal1 14005 3246 14056 3284 0 FreeSans 200 0 0 0 TAP_31.VGND
rlabel comment 13984 3264 13984 3264 4 TAP_31.tapvpwrvgnd_1
flabel metal1 15209 3247 15243 3281 0 FreeSans 200 0 0 0 FILLER_2_153.VGND
flabel metal1 15209 3791 15243 3825 0 FreeSans 200 0 0 0 FILLER_2_153.VPWR
flabel nwell 15209 3791 15243 3825 0 FreeSans 200 0 0 0 FILLER_2_153.VPB
flabel pwell 15209 3247 15243 3281 0 FreeSans 200 0 0 0 FILLER_2_153.VNB
rlabel comment 15180 3264 15180 3264 4 FILLER_2_153.decap_12
flabel metal1 16313 3247 16347 3281 0 FreeSans 200 0 0 0 FILLER_2_165.VGND
flabel metal1 16313 3791 16347 3825 0 FreeSans 200 0 0 0 FILLER_2_165.VPWR
flabel nwell 16313 3791 16347 3825 0 FreeSans 200 0 0 0 FILLER_2_165.VPB
flabel pwell 16313 3247 16347 3281 0 FreeSans 200 0 0 0 FILLER_2_165.VNB
rlabel comment 16284 3264 16284 3264 4 FILLER_2_165.decap_12
flabel metal1 17417 3247 17451 3281 0 FreeSans 200 0 0 0 FILLER_2_177.VGND
flabel metal1 17417 3791 17451 3825 0 FreeSans 200 0 0 0 FILLER_2_177.VPWR
flabel nwell 17417 3791 17451 3825 0 FreeSans 200 0 0 0 FILLER_2_177.VPB
flabel pwell 17417 3247 17451 3281 0 FreeSans 200 0 0 0 FILLER_2_177.VNB
rlabel comment 17388 3264 17388 3264 4 FILLER_2_177.decap_12
flabel metal1 18514 3791 18550 3821 0 FreeSans 250 0 0 0 FILLER_2_189.VPWR
flabel metal1 18514 3251 18550 3280 0 FreeSans 250 0 0 0 FILLER_2_189.VGND
flabel nwell 18523 3798 18543 3815 0 FreeSans 200 0 0 0 FILLER_2_189.VPB
flabel pwell 18520 3253 18544 3275 0 FreeSans 200 0 0 0 FILLER_2_189.VNB
rlabel comment 18492 3264 18492 3264 4 FILLER_2_189.fill_1
flabel metal1 18797 3791 18831 3825 0 FreeSans 200 0 0 0 PHY_5.VPWR
flabel metal1 18797 3247 18831 3281 0 FreeSans 200 0 0 0 PHY_5.VGND
flabel nwell 18797 3791 18831 3825 0 FreeSans 200 0 0 0 PHY_5.VPB
flabel pwell 18797 3247 18831 3281 0 FreeSans 200 0 0 0 PHY_5.VNB
rlabel comment 18860 3264 18860 3264 6 PHY_5.decap_3
flabel metal1 2138 3795 2174 3825 0 FreeSans 250 0 0 0 FILLER_3_11.VPWR
flabel metal1 2138 4336 2174 4365 0 FreeSans 250 0 0 0 FILLER_3_11.VGND
flabel nwell 2147 3801 2167 3818 0 FreeSans 200 0 0 0 FILLER_3_11.VPB
flabel pwell 2144 4341 2168 4363 0 FreeSans 200 0 0 0 FILLER_3_11.VNB
rlabel comment 2116 4352 2116 4352 2 FILLER_3_11.fill_1
flabel metal1 2513 4335 2547 4369 0 FreeSans 200 0 0 0 FILLER_3_15.VGND
flabel metal1 2513 3791 2547 3825 0 FreeSans 200 0 0 0 FILLER_3_15.VPWR
flabel nwell 2513 3791 2547 3825 0 FreeSans 200 0 0 0 FILLER_3_15.VPB
flabel pwell 2513 4335 2547 4369 0 FreeSans 200 0 0 0 FILLER_3_15.VNB
rlabel comment 2484 4352 2484 4352 2 FILLER_3_15.decap_4
flabel metal1 1409 3791 1443 3825 0 FreeSans 200 0 0 0 FILLER_3_3.VPWR
flabel metal1 1409 4335 1443 4369 0 FreeSans 200 0 0 0 FILLER_3_3.VGND
flabel nwell 1409 3791 1443 3825 0 FreeSans 200 0 0 0 FILLER_3_3.VPB
flabel pwell 1409 4335 1443 4369 0 FreeSans 200 0 0 0 FILLER_3_3.VNB
rlabel comment 1380 4352 1380 4352 2 FILLER_3_3.decap_8
flabel metal1 1133 3791 1167 3825 0 FreeSans 200 0 0 0 PHY_6.VPWR
flabel metal1 1133 4335 1167 4369 0 FreeSans 200 0 0 0 PHY_6.VGND
flabel nwell 1133 3791 1167 3825 0 FreeSans 200 0 0 0 PHY_6.VPB
flabel pwell 1133 4335 1167 4369 0 FreeSans 200 0 0 0 PHY_6.VNB
rlabel comment 1104 4352 1104 4352 2 PHY_6.decap_3
flabel locali 4628 3893 4662 3927 0 FreeSans 400 0 0 0 _53_.Q
flabel locali 4628 3961 4662 3995 0 FreeSans 400 0 0 0 _53_.Q
flabel locali 4628 4029 4662 4063 0 FreeSans 400 0 0 0 _53_.Q
flabel locali 4628 4233 4662 4267 0 FreeSans 400 0 0 0 _53_.Q
flabel locali 4333 4165 4367 4199 0 FreeSans 400 0 0 0 _53_.RESET_B
flabel locali 3157 4029 3191 4063 0 FreeSans 400 0 0 0 _53_.D
flabel locali 2882 4029 2916 4063 0 FreeSans 400 0 0 0 _53_.CLK
flabel locali 2882 4097 2916 4131 0 FreeSans 400 0 0 0 _53_.CLK
flabel locali 4333 4097 4367 4131 0 FreeSans 400 0 0 0 _53_.RESET_B
flabel metal1 2881 4335 2915 4369 0 FreeSans 200 0 0 0 _53_.VGND
flabel metal1 2881 3791 2915 3825 0 FreeSans 200 0 0 0 _53_.VPWR
flabel nwell 2881 3791 2915 3825 0 FreeSans 200 0 0 0 _53_.VPB
flabel pwell 2881 4335 2915 4369 0 FreeSans 200 0 0 0 _53_.VNB
rlabel comment 2852 4352 2852 4352 2 _53_.dfrtp_1
flabel metal1 2237 4335 2271 4369 0 FreeSans 200 180 0 0 input2.VGND
flabel metal1 2237 3791 2271 3825 0 FreeSans 200 180 0 0 input2.VPWR
flabel locali 2421 4233 2455 4267 0 FreeSans 200 180 0 0 input2.X
flabel locali 2421 3961 2455 3995 0 FreeSans 200 180 0 0 input2.X
flabel locali 2421 3893 2455 3927 0 FreeSans 200 180 0 0 input2.X
flabel locali 2237 4097 2271 4131 0 FreeSans 200 180 0 0 input2.A
flabel nwell 2237 3791 2271 3825 0 FreeSans 200 180 0 0 input2.VPB
flabel pwell 2237 4335 2271 4369 0 FreeSans 200 180 0 0 input2.VNB
rlabel comment 2484 4352 2484 4352 8 input2.clkbuf_1
flabel metal1 4721 4335 4755 4369 0 FreeSans 200 0 0 0 FILLER_3_39.VGND
flabel metal1 4721 3791 4755 3825 0 FreeSans 200 0 0 0 FILLER_3_39.VPWR
flabel nwell 4721 3791 4755 3825 0 FreeSans 200 0 0 0 FILLER_3_39.VPB
flabel pwell 4721 4335 4755 4369 0 FreeSans 200 0 0 0 FILLER_3_39.VNB
rlabel comment 4692 4352 4692 4352 2 FILLER_3_39.decap_4
flabel locali 5108 4029 5142 4063 0 FreeSans 200 0 0 0 _60__15.LO
flabel locali 5235 4093 5269 4127 0 FreeSans 200 0 0 0 _60__15.HI
flabel nwell 5273 3791 5307 3825 0 FreeSans 200 0 0 0 _60__15.VPB
flabel pwell 5273 4335 5307 4369 0 FreeSans 200 0 0 0 _60__15.VNB
flabel metal1 5273 4335 5307 4369 0 FreeSans 200 0 0 0 _60__15.VGND
flabel metal1 5273 3791 5307 3825 0 FreeSans 200 0 0 0 _60__15.VPWR
rlabel comment 5336 4352 5336 4352 8 _60__15.conb_1
flabel comment 5291 4079 5291 4079 0 FreeSans 200 90 0 0 _60__15.resistive_li1_ok
flabel comment 5103 4079 5103 4079 0 FreeSans 200 90 0 0 _60__15.resistive_li1_ok
flabel comment 5150 4094 5150 4094 0 FreeSans 200 90 0 0 _60__15.no_jumper_check
flabel comment 5253 4094 5253 4094 0 FreeSans 200 90 0 0 _60__15.no_jumper_check
flabel metal1 5365 3791 5399 3825 0 FreeSans 200 0 0 0 FILLER_3_46.VPWR
flabel metal1 5365 4335 5399 4369 0 FreeSans 200 0 0 0 FILLER_3_46.VGND
flabel nwell 5365 3791 5399 3825 0 FreeSans 200 0 0 0 FILLER_3_46.VPB
flabel pwell 5365 4335 5399 4369 0 FreeSans 200 0 0 0 FILLER_3_46.VNB
rlabel comment 5336 4352 5336 4352 2 FILLER_3_46.decap_8
flabel metal1 6092 4334 6145 4366 0 FreeSans 200 0 0 0 FILLER_3_54.VGND
flabel metal1 6093 3791 6145 3822 0 FreeSans 200 0 0 0 FILLER_3_54.VPWR
flabel nwell 6100 3799 6134 3817 0 FreeSans 200 0 0 0 FILLER_3_54.VPB
flabel pwell 6103 4340 6135 4362 0 FreeSans 200 0 0 0 FILLER_3_54.VNB
rlabel comment 6072 4352 6072 4352 2 FILLER_3_54.fill_2
flabel metal1 6377 3791 6411 3825 0 FreeSans 200 0 0 0 FILLER_3_57.VPWR
flabel metal1 6377 4335 6411 4369 0 FreeSans 200 0 0 0 FILLER_3_57.VGND
flabel nwell 6377 3791 6411 3825 0 FreeSans 200 0 0 0 FILLER_3_57.VPB
flabel pwell 6377 4335 6411 4369 0 FreeSans 200 0 0 0 FILLER_3_57.VNB
rlabel comment 6348 4352 6348 4352 2 FILLER_3_57.decap_3
flabel metal1 6929 3791 6963 3825 0 FreeSans 200 0 0 0 FILLER_3_63.VPWR
flabel metal1 6929 4335 6963 4369 0 FreeSans 200 0 0 0 FILLER_3_63.VGND
flabel nwell 6929 3791 6963 3825 0 FreeSans 200 0 0 0 FILLER_3_63.VPB
flabel pwell 6929 4335 6963 4369 0 FreeSans 200 0 0 0 FILLER_3_63.VNB
rlabel comment 6900 4352 6900 4352 2 FILLER_3_63.decap_8
flabel metal1 6278 3799 6331 3828 0 FreeSans 200 0 0 0 TAP_32.VPWR
flabel metal1 6277 4332 6328 4370 0 FreeSans 200 0 0 0 TAP_32.VGND
rlabel comment 6256 4352 6256 4352 2 TAP_32.tapvpwrvgnd_1
flabel metal1 6837 4335 6871 4369 0 FreeSans 200 180 0 0 _39_.VGND
flabel metal1 6837 3791 6871 3825 0 FreeSans 200 180 0 0 _39_.VPWR
flabel locali 6653 4233 6687 4267 0 FreeSans 200 180 0 0 _39_.X
flabel locali 6653 3961 6687 3995 0 FreeSans 200 180 0 0 _39_.X
flabel locali 6653 3893 6687 3927 0 FreeSans 200 180 0 0 _39_.X
flabel locali 6837 4097 6871 4131 0 FreeSans 200 180 0 0 _39_.A
flabel nwell 6837 3791 6871 3825 0 FreeSans 200 180 0 0 _39_.VPB
flabel pwell 6837 4335 6871 4369 0 FreeSans 200 180 0 0 _39_.VNB
rlabel comment 6624 4352 6624 4352 2 _39_.clkbuf_1
flabel metal1 8493 4335 8527 4369 0 FreeSans 200 0 0 0 FILLER_3_80.VGND
flabel metal1 8493 3791 8527 3825 0 FreeSans 200 0 0 0 FILLER_3_80.VPWR
flabel nwell 8493 3791 8527 3825 0 FreeSans 200 0 0 0 FILLER_3_80.VPB
flabel pwell 8493 4335 8527 4369 0 FreeSans 200 0 0 0 FILLER_3_80.VNB
rlabel comment 8464 4352 8464 4352 2 FILLER_3_80.decap_4
flabel metal1 8854 3795 8890 3825 0 FreeSans 250 0 0 0 FILLER_3_84.VPWR
flabel metal1 8854 4336 8890 4365 0 FreeSans 250 0 0 0 FILLER_3_84.VGND
flabel nwell 8863 3801 8883 3818 0 FreeSans 200 0 0 0 FILLER_3_84.VPB
flabel pwell 8860 4341 8884 4363 0 FreeSans 200 0 0 0 FILLER_3_84.VNB
rlabel comment 8832 4352 8832 4352 2 FILLER_3_84.fill_1
flabel metal1 8400 4335 8434 4369 0 FreeSans 200 0 0 0 _46_.VGND
flabel metal1 8400 3791 8434 3825 0 FreeSans 200 0 0 0 _46_.VPWR
flabel locali 7756 4029 7790 4063 0 FreeSans 250 0 0 0 _46_.S
flabel locali 7848 4029 7882 4063 0 FreeSans 250 0 0 0 _46_.S
flabel locali 7940 4165 7974 4199 0 FreeSans 250 0 0 0 _46_.A1
flabel locali 7940 4097 7974 4131 0 FreeSans 250 0 0 0 _46_.A1
flabel locali 8032 4097 8066 4131 0 FreeSans 250 0 0 0 _46_.A0
flabel locali 8400 4233 8434 4267 0 FreeSans 250 0 0 0 _46_.X
flabel locali 8400 3961 8434 3995 0 FreeSans 250 0 0 0 _46_.X
flabel locali 8400 3893 8434 3927 0 FreeSans 250 0 0 0 _46_.X
flabel nwell 8356 3791 8390 3825 0 FreeSans 250 0 0 0 _46_.VPB
flabel pwell 8346 4335 8380 4369 0 FreeSans 250 0 0 0 _46_.VNB
rlabel comment 8464 4352 8464 4352 8 _46_.mux2_1
flabel locali 10517 4029 10551 4063 0 FreeSans 200 0 0 0 clkbuf_0_clk.X
flabel locali 10609 4029 10643 4063 0 FreeSans 200 0 0 0 clkbuf_0_clk.X
flabel locali 10609 4097 10643 4131 0 FreeSans 200 0 0 0 clkbuf_0_clk.X
flabel locali 10517 4097 10551 4131 0 FreeSans 200 0 0 0 clkbuf_0_clk.X
flabel locali 10517 4165 10551 4199 0 FreeSans 200 0 0 0 clkbuf_0_clk.X
flabel locali 10609 4165 10643 4199 0 FreeSans 200 0 0 0 clkbuf_0_clk.X
flabel locali 8953 4165 8987 4199 0 FreeSans 200 0 0 0 clkbuf_0_clk.A
flabel locali 8953 4097 8987 4131 0 FreeSans 200 0 0 0 clkbuf_0_clk.A
flabel pwell 8953 4335 8987 4369 0 FreeSans 200 0 0 0 clkbuf_0_clk.VNB
flabel pwell 8970 4352 8970 4352 0 FreeSans 200 0 0 0 clkbuf_0_clk.VNB
flabel nwell 8953 3791 8987 3825 0 FreeSans 200 0 0 0 clkbuf_0_clk.VPB
flabel nwell 8970 3808 8970 3808 0 FreeSans 200 0 0 0 clkbuf_0_clk.VPB
flabel metal1 8953 4335 8987 4369 0 FreeSans 200 0 0 0 clkbuf_0_clk.VGND
flabel metal1 8953 3791 8987 3825 0 FreeSans 200 0 0 0 clkbuf_0_clk.VPWR
rlabel comment 8924 4352 8924 4352 2 clkbuf_0_clk.clkbuf_16
flabel metal1 10793 3791 10827 3825 0 FreeSans 200 0 0 0 FILLER_3_105.VPWR
flabel metal1 10793 4335 10827 4369 0 FreeSans 200 0 0 0 FILLER_3_105.VGND
flabel nwell 10793 3791 10827 3825 0 FreeSans 200 0 0 0 FILLER_3_105.VPB
flabel pwell 10793 4335 10827 4369 0 FreeSans 200 0 0 0 FILLER_3_105.VNB
rlabel comment 10764 4352 10764 4352 2 FILLER_3_105.decap_6
flabel metal1 11338 3795 11374 3825 0 FreeSans 250 0 0 0 FILLER_3_111.VPWR
flabel metal1 11338 4336 11374 4365 0 FreeSans 250 0 0 0 FILLER_3_111.VGND
flabel nwell 11347 3801 11367 3818 0 FreeSans 200 0 0 0 FILLER_3_111.VPB
flabel pwell 11344 4341 11368 4363 0 FreeSans 200 0 0 0 FILLER_3_111.VNB
rlabel comment 11316 4352 11316 4352 2 FILLER_3_111.fill_1
flabel metal1 11520 4334 11573 4366 0 FreeSans 200 0 0 0 FILLER_3_113.VGND
flabel metal1 11521 3791 11573 3822 0 FreeSans 200 0 0 0 FILLER_3_113.VPWR
flabel nwell 11528 3799 11562 3817 0 FreeSans 200 0 0 0 FILLER_3_113.VPB
flabel pwell 11531 4340 11563 4362 0 FreeSans 200 0 0 0 FILLER_3_113.VNB
rlabel comment 11500 4352 11500 4352 2 FILLER_3_113.fill_2
flabel metal1 11430 3799 11483 3828 0 FreeSans 200 0 0 0 TAP_33.VPWR
flabel metal1 11429 4332 11480 4370 0 FreeSans 200 0 0 0 TAP_33.VGND
rlabel comment 11408 4352 11408 4352 2 TAP_33.tapvpwrvgnd_1
flabel locali 11714 3893 11748 3927 0 FreeSans 400 0 0 0 _49_.Q
flabel locali 11714 3961 11748 3995 0 FreeSans 400 0 0 0 _49_.Q
flabel locali 11714 4029 11748 4063 0 FreeSans 400 0 0 0 _49_.Q
flabel locali 11714 4233 11748 4267 0 FreeSans 400 0 0 0 _49_.Q
flabel locali 12009 4165 12043 4199 0 FreeSans 400 0 0 0 _49_.RESET_B
flabel locali 13185 4029 13219 4063 0 FreeSans 400 0 0 0 _49_.D
flabel locali 13460 4029 13494 4063 0 FreeSans 400 0 0 0 _49_.CLK
flabel locali 13460 4097 13494 4131 0 FreeSans 400 0 0 0 _49_.CLK
flabel locali 12009 4097 12043 4131 0 FreeSans 400 0 0 0 _49_.RESET_B
flabel metal1 13461 4335 13495 4369 0 FreeSans 200 0 0 0 _49_.VGND
flabel metal1 13461 3791 13495 3825 0 FreeSans 200 0 0 0 _49_.VPWR
flabel nwell 13461 3791 13495 3825 0 FreeSans 200 0 0 0 _49_.VPB
flabel pwell 13461 4335 13495 4369 0 FreeSans 200 0 0 0 _49_.VNB
rlabel comment 13524 4352 13524 4352 8 _49_.dfrtp_1
flabel metal1 13553 4335 13587 4369 0 FreeSans 200 0 0 0 FILLER_3_135.VGND
flabel metal1 13553 3791 13587 3825 0 FreeSans 200 0 0 0 FILLER_3_135.VPWR
flabel nwell 13553 3791 13587 3825 0 FreeSans 200 0 0 0 FILLER_3_135.VPB
flabel pwell 13553 4335 13587 4369 0 FreeSans 200 0 0 0 FILLER_3_135.VNB
rlabel comment 13524 4352 13524 4352 2 FILLER_3_135.decap_4
flabel locali 15668 3893 15702 3927 0 FreeSans 400 0 0 0 _54_.Q
flabel locali 15668 3961 15702 3995 0 FreeSans 400 0 0 0 _54_.Q
flabel locali 15668 4029 15702 4063 0 FreeSans 400 0 0 0 _54_.Q
flabel locali 15668 4233 15702 4267 0 FreeSans 400 0 0 0 _54_.Q
flabel locali 15373 4165 15407 4199 0 FreeSans 400 0 0 0 _54_.RESET_B
flabel locali 14197 4029 14231 4063 0 FreeSans 400 0 0 0 _54_.D
flabel locali 13922 4029 13956 4063 0 FreeSans 400 0 0 0 _54_.CLK
flabel locali 13922 4097 13956 4131 0 FreeSans 400 0 0 0 _54_.CLK
flabel locali 15373 4097 15407 4131 0 FreeSans 400 0 0 0 _54_.RESET_B
flabel metal1 13921 4335 13955 4369 0 FreeSans 200 0 0 0 _54_.VGND
flabel metal1 13921 3791 13955 3825 0 FreeSans 200 0 0 0 _54_.VPWR
flabel nwell 13921 3791 13955 3825 0 FreeSans 200 0 0 0 _54_.VPB
flabel pwell 13921 4335 13955 4369 0 FreeSans 200 0 0 0 _54_.VNB
rlabel comment 13892 4352 13892 4352 2 _54_.dfrtp_1
flabel metal1 15761 3791 15795 3825 0 FreeSans 200 0 0 0 FILLER_3_159.VPWR
flabel metal1 15761 4335 15795 4369 0 FreeSans 200 0 0 0 FILLER_3_159.VGND
flabel nwell 15761 3791 15795 3825 0 FreeSans 200 0 0 0 FILLER_3_159.VPB
flabel pwell 15761 4335 15795 4369 0 FreeSans 200 0 0 0 FILLER_3_159.VNB
rlabel comment 15732 4352 15732 4352 2 FILLER_3_159.decap_8
flabel metal1 16490 3795 16526 3825 0 FreeSans 250 0 0 0 FILLER_3_167.VPWR
flabel metal1 16490 4336 16526 4365 0 FreeSans 250 0 0 0 FILLER_3_167.VGND
flabel nwell 16499 3801 16519 3818 0 FreeSans 200 0 0 0 FILLER_3_167.VPB
flabel pwell 16496 4341 16520 4363 0 FreeSans 200 0 0 0 FILLER_3_167.VNB
rlabel comment 16468 4352 16468 4352 2 FILLER_3_167.fill_1
flabel metal1 16681 4335 16715 4369 0 FreeSans 200 0 0 0 FILLER_3_169.VGND
flabel metal1 16681 3791 16715 3825 0 FreeSans 200 0 0 0 FILLER_3_169.VPWR
flabel nwell 16681 3791 16715 3825 0 FreeSans 200 0 0 0 FILLER_3_169.VPB
flabel pwell 16681 4335 16715 4369 0 FreeSans 200 0 0 0 FILLER_3_169.VNB
rlabel comment 16652 4352 16652 4352 2 FILLER_3_169.decap_12
flabel metal1 16582 3799 16635 3828 0 FreeSans 200 0 0 0 TAP_34.VPWR
flabel metal1 16581 4332 16632 4370 0 FreeSans 200 0 0 0 TAP_34.VGND
rlabel comment 16560 4352 16560 4352 2 TAP_34.tapvpwrvgnd_1
flabel metal1 17785 3791 17819 3825 0 FreeSans 200 0 0 0 FILLER_3_181.VPWR
flabel metal1 17785 4335 17819 4369 0 FreeSans 200 0 0 0 FILLER_3_181.VGND
flabel nwell 17785 3791 17819 3825 0 FreeSans 200 0 0 0 FILLER_3_181.VPB
flabel pwell 17785 4335 17819 4369 0 FreeSans 200 0 0 0 FILLER_3_181.VNB
rlabel comment 17756 4352 17756 4352 2 FILLER_3_181.decap_8
flabel metal1 18514 3795 18550 3825 0 FreeSans 250 0 0 0 FILLER_3_189.VPWR
flabel metal1 18514 4336 18550 4365 0 FreeSans 250 0 0 0 FILLER_3_189.VGND
flabel nwell 18523 3801 18543 3818 0 FreeSans 200 0 0 0 FILLER_3_189.VPB
flabel pwell 18520 4341 18544 4363 0 FreeSans 200 0 0 0 FILLER_3_189.VNB
rlabel comment 18492 4352 18492 4352 2 FILLER_3_189.fill_1
flabel metal1 18797 3791 18831 3825 0 FreeSans 200 0 0 0 PHY_7.VPWR
flabel metal1 18797 4335 18831 4369 0 FreeSans 200 0 0 0 PHY_7.VGND
flabel nwell 18797 3791 18831 3825 0 FreeSans 200 0 0 0 PHY_7.VPB
flabel pwell 18797 4335 18831 4369 0 FreeSans 200 0 0 0 PHY_7.VNB
rlabel comment 18860 4352 18860 4352 8 PHY_7.decap_3
flabel metal1 2145 4879 2179 4913 0 FreeSans 200 0 0 0 FILLER_4_11.VPWR
flabel metal1 2145 4335 2179 4369 0 FreeSans 200 0 0 0 FILLER_4_11.VGND
flabel nwell 2145 4879 2179 4913 0 FreeSans 200 0 0 0 FILLER_4_11.VPB
flabel pwell 2145 4335 2179 4369 0 FreeSans 200 0 0 0 FILLER_4_11.VNB
rlabel comment 2116 4352 2116 4352 4 FILLER_4_11.decap_3
flabel metal1 1409 4879 1443 4913 0 FreeSans 200 0 0 0 FILLER_4_3.VPWR
flabel metal1 1409 4335 1443 4369 0 FreeSans 200 0 0 0 FILLER_4_3.VGND
flabel nwell 1409 4879 1443 4913 0 FreeSans 200 0 0 0 FILLER_4_3.VPB
flabel pwell 1409 4335 1443 4369 0 FreeSans 200 0 0 0 FILLER_4_3.VNB
rlabel comment 1380 4352 1380 4352 4 FILLER_4_3.decap_8
flabel metal1 1133 4879 1167 4913 0 FreeSans 200 0 0 0 PHY_8.VPWR
flabel metal1 1133 4335 1167 4369 0 FreeSans 200 0 0 0 PHY_8.VGND
flabel nwell 1133 4879 1167 4913 0 FreeSans 200 0 0 0 PHY_8.VPB
flabel pwell 1133 4335 1167 4369 0 FreeSans 200 0 0 0 PHY_8.VNB
rlabel comment 1104 4352 1104 4352 4 PHY_8.decap_3
flabel locali 3065 4573 3099 4607 0 FreeSans 200 0 0 0 hold1.A
flabel locali 2417 4505 2451 4539 0 FreeSans 200 0 0 0 hold1.X
flabel locali 3065 4641 3099 4675 0 FreeSans 200 0 0 0 hold1.A
flabel locali 2417 4437 2451 4471 0 FreeSans 200 0 0 0 hold1.X
flabel locali 2973 4573 3007 4607 0 FreeSans 200 0 0 0 hold1.A
flabel locali 2973 4641 3007 4675 0 FreeSans 200 0 0 0 hold1.A
flabel locali 2417 4777 2451 4811 0 FreeSans 200 0 0 0 hold1.X
flabel locali 2417 4641 2451 4675 0 FreeSans 200 0 0 0 hold1.X
flabel locali 2417 4709 2451 4743 0 FreeSans 200 0 0 0 hold1.X
flabel locali 2417 4573 2451 4607 0 FreeSans 200 0 0 0 hold1.X
flabel nwell 3065 4879 3099 4913 0 FreeSans 200 0 0 0 hold1.VPB
flabel pwell 3065 4335 3099 4369 0 FreeSans 200 0 0 0 hold1.VNB
flabel metal1 3065 4335 3099 4369 0 FreeSans 200 0 0 0 hold1.VGND
flabel metal1 3065 4879 3099 4913 0 FreeSans 200 0 0 0 hold1.VPWR
rlabel comment 3128 4352 3128 4352 6 hold1.dlygate4sd3_1
flabel locali 4905 4437 4939 4471 0 FreeSans 200 0 0 0 ANTENNA_hold1_A.DIODE
flabel locali 4905 4709 4939 4743 0 FreeSans 200 0 0 0 ANTENNA_hold1_A.DIODE
flabel locali 4997 4709 5031 4743 0 FreeSans 200 0 0 0 ANTENNA_hold1_A.DIODE
flabel locali 4905 4777 4939 4811 0 FreeSans 200 0 0 0 ANTENNA_hold1_A.DIODE
flabel locali 4997 4777 5031 4811 0 FreeSans 200 0 0 0 ANTENNA_hold1_A.DIODE
flabel locali 4997 4641 5031 4675 0 FreeSans 200 0 0 0 ANTENNA_hold1_A.DIODE
flabel locali 4905 4641 4939 4675 0 FreeSans 200 0 0 0 ANTENNA_hold1_A.DIODE
flabel locali 4997 4573 5031 4607 0 FreeSans 200 0 0 0 ANTENNA_hold1_A.DIODE
flabel locali 4905 4573 4939 4607 0 FreeSans 200 0 0 0 ANTENNA_hold1_A.DIODE
flabel locali 4905 4505 4939 4539 0 FreeSans 200 0 0 0 ANTENNA_hold1_A.DIODE
flabel locali 4997 4505 5031 4539 0 FreeSans 200 0 0 0 ANTENNA_hold1_A.DIODE
flabel locali 4997 4437 5031 4471 0 FreeSans 200 0 0 0 ANTENNA_hold1_A.DIODE
flabel metal1 4997 4335 5031 4369 0 FreeSans 200 0 0 0 ANTENNA_hold1_A.VGND
flabel metal1 4997 4879 5031 4913 0 FreeSans 200 0 0 0 ANTENNA_hold1_A.VPWR
flabel nwell 4997 4879 5031 4913 0 FreeSans 200 0 0 0 ANTENNA_hold1_A.VPB
flabel pwell 4997 4335 5031 4369 0 FreeSans 200 0 0 0 ANTENNA_hold1_A.VNB
rlabel comment 5060 4352 5060 4352 6 ANTENNA_hold1_A.diode_2
flabel metal1 3157 4879 3191 4913 0 FreeSans 200 0 0 0 FILLER_4_22.VPWR
flabel metal1 3157 4335 3191 4369 0 FreeSans 200 0 0 0 FILLER_4_22.VGND
flabel nwell 3157 4879 3191 4913 0 FreeSans 200 0 0 0 FILLER_4_22.VPB
flabel pwell 3157 4335 3191 4369 0 FreeSans 200 0 0 0 FILLER_4_22.VNB
rlabel comment 3128 4352 3128 4352 4 FILLER_4_22.decap_6
flabel metal1 3792 4338 3845 4370 0 FreeSans 200 0 0 0 FILLER_4_29.VGND
flabel metal1 3793 4882 3845 4913 0 FreeSans 200 0 0 0 FILLER_4_29.VPWR
flabel nwell 3800 4887 3834 4905 0 FreeSans 200 0 0 0 FILLER_4_29.VPB
flabel pwell 3803 4342 3835 4364 0 FreeSans 200 0 0 0 FILLER_4_29.VNB
rlabel comment 3772 4352 3772 4352 4 FILLER_4_29.fill_2
flabel metal1 4537 4335 4571 4369 0 FreeSans 200 0 0 0 FILLER_4_37.VGND
flabel metal1 4537 4879 4571 4913 0 FreeSans 200 0 0 0 FILLER_4_37.VPWR
flabel nwell 4537 4879 4571 4913 0 FreeSans 200 0 0 0 FILLER_4_37.VPB
flabel pwell 4537 4335 4571 4369 0 FreeSans 200 0 0 0 FILLER_4_37.VNB
rlabel comment 4508 4352 4508 4352 4 FILLER_4_37.decap_4
flabel metal1 5089 4879 5123 4913 0 FreeSans 200 0 0 0 FILLER_4_43.VPWR
flabel metal1 5089 4335 5123 4369 0 FreeSans 200 0 0 0 FILLER_4_43.VGND
flabel nwell 5089 4879 5123 4913 0 FreeSans 200 0 0 0 FILLER_4_43.VPB
flabel pwell 5089 4335 5123 4369 0 FreeSans 200 0 0 0 FILLER_4_43.VNB
rlabel comment 5060 4352 5060 4352 4 FILLER_4_43.decap_8
flabel metal1 3702 4876 3755 4905 0 FreeSans 200 0 0 0 TAP_35.VPWR
flabel metal1 3701 4334 3752 4372 0 FreeSans 200 0 0 0 TAP_35.VGND
rlabel comment 3680 4352 3680 4352 4 TAP_35.tapvpwrvgnd_1
flabel locali 4077 4641 4111 4675 0 FreeSans 200 0 0 0 fanout13.X
flabel locali 4353 4505 4387 4539 0 FreeSans 200 0 0 0 fanout13.A
flabel locali 3985 4505 4019 4539 0 FreeSans 200 0 0 0 fanout13.X
flabel locali 4353 4573 4387 4607 0 FreeSans 200 0 0 0 fanout13.A
flabel locali 3985 4573 4019 4607 0 FreeSans 200 0 0 0 fanout13.X
flabel metal1 4445 4335 4479 4369 0 FreeSans 200 0 0 0 fanout13.VGND
flabel metal1 4445 4879 4479 4913 0 FreeSans 200 0 0 0 fanout13.VPWR
flabel nwell 4445 4879 4479 4913 0 FreeSans 200 0 0 0 fanout13.VPB
flabel pwell 4445 4335 4479 4369 0 FreeSans 200 0 0 0 fanout13.VNB
rlabel comment 4508 4352 4508 4352 6 fanout13.clkbuf_4
flabel metal1 5816 4338 5869 4370 0 FreeSans 200 0 0 0 FILLER_4_51.VGND
flabel metal1 5817 4882 5869 4913 0 FreeSans 200 0 0 0 FILLER_4_51.VPWR
flabel nwell 5824 4887 5858 4905 0 FreeSans 200 0 0 0 FILLER_4_51.VPB
flabel pwell 5827 4342 5859 4364 0 FreeSans 200 0 0 0 FILLER_4_51.VNB
rlabel comment 5796 4352 5796 4352 4 FILLER_4_51.fill_2
flabel metal1 6469 4335 6503 4369 0 FreeSans 200 0 0 0 FILLER_4_58.VGND
flabel metal1 6469 4879 6503 4913 0 FreeSans 200 0 0 0 FILLER_4_58.VPWR
flabel nwell 6469 4879 6503 4913 0 FreeSans 200 0 0 0 FILLER_4_58.VPB
flabel pwell 6469 4335 6503 4369 0 FreeSans 200 0 0 0 FILLER_4_58.VNB
rlabel comment 6440 4352 6440 4352 4 FILLER_4_58.decap_4
flabel locali 6193 4573 6227 4607 0 FreeSans 200 0 0 0 _38_.A
flabel locali 6009 4709 6043 4743 0 FreeSans 200 0 0 0 _38_.X
flabel locali 6377 4573 6411 4607 0 FreeSans 200 0 0 0 _38_.B
flabel nwell 6377 4879 6411 4913 0 FreeSans 200 0 0 0 _38_.VPB
flabel pwell 6377 4335 6411 4369 0 FreeSans 200 0 0 0 _38_.VNB
flabel metal1 6377 4335 6411 4369 0 FreeSans 200 0 0 0 _38_.VGND
flabel metal1 6377 4879 6411 4913 0 FreeSans 200 0 0 0 _38_.VPWR
rlabel comment 6440 4352 6440 4352 6 _38_.or2_1
flabel locali 7021 4573 7055 4607 0 FreeSans 200 0 0 0 _44_.A
flabel locali 7205 4709 7239 4743 0 FreeSans 200 0 0 0 _44_.X
flabel locali 6837 4573 6871 4607 0 FreeSans 200 0 0 0 _44_.B
flabel nwell 6837 4879 6871 4913 0 FreeSans 200 0 0 0 _44_.VPB
flabel pwell 6837 4335 6871 4369 0 FreeSans 200 0 0 0 _44_.VNB
flabel metal1 6837 4335 6871 4369 0 FreeSans 200 0 0 0 _44_.VGND
flabel metal1 6837 4879 6871 4913 0 FreeSans 200 0 0 0 _44_.VPWR
rlabel comment 6808 4352 6808 4352 4 _44_.or2_1
flabel metal1 7297 4879 7331 4913 0 FreeSans 200 0 0 0 FILLER_4_67.VPWR
flabel metal1 7297 4335 7331 4369 0 FreeSans 200 0 0 0 FILLER_4_67.VGND
flabel nwell 7297 4879 7331 4913 0 FreeSans 200 0 0 0 FILLER_4_67.VPB
flabel pwell 7297 4335 7331 4369 0 FreeSans 200 0 0 0 FILLER_4_67.VNB
rlabel comment 7268 4352 7268 4352 4 FILLER_4_67.decap_6
flabel metal1 8668 4338 8721 4370 0 FreeSans 200 0 0 0 FILLER_4_82.VGND
flabel metal1 8669 4882 8721 4913 0 FreeSans 200 0 0 0 FILLER_4_82.VPWR
flabel nwell 8676 4887 8710 4905 0 FreeSans 200 0 0 0 FILLER_4_82.VPB
flabel pwell 8679 4342 8711 4364 0 FreeSans 200 0 0 0 FILLER_4_82.VNB
rlabel comment 8648 4352 8648 4352 4 FILLER_4_82.fill_2
flabel metal1 8944 4338 8997 4370 0 FreeSans 200 0 0 0 FILLER_4_85.VGND
flabel metal1 8945 4882 8997 4913 0 FreeSans 200 0 0 0 FILLER_4_85.VPWR
flabel nwell 8952 4887 8986 4905 0 FreeSans 200 0 0 0 FILLER_4_85.VPB
flabel pwell 8955 4342 8987 4364 0 FreeSans 200 0 0 0 FILLER_4_85.VNB
rlabel comment 8924 4352 8924 4352 4 FILLER_4_85.fill_2
flabel metal1 8854 4876 8907 4905 0 FreeSans 200 0 0 0 TAP_36.VPWR
flabel metal1 8853 4334 8904 4372 0 FreeSans 200 0 0 0 TAP_36.VGND
rlabel comment 8832 4352 8832 4352 4 TAP_36.tapvpwrvgnd_1
flabel metal1 7850 4335 7884 4369 0 FreeSans 200 0 0 0 _37_.VGND
flabel metal1 7850 4879 7884 4913 0 FreeSans 200 0 0 0 _37_.VPWR
flabel locali 8494 4641 8528 4675 0 FreeSans 250 0 0 0 _37_.S
flabel locali 8402 4641 8436 4675 0 FreeSans 250 0 0 0 _37_.S
flabel locali 8310 4505 8344 4539 0 FreeSans 250 0 0 0 _37_.A1
flabel locali 8310 4573 8344 4607 0 FreeSans 250 0 0 0 _37_.A1
flabel locali 8218 4573 8252 4607 0 FreeSans 250 0 0 0 _37_.A0
flabel locali 7850 4437 7884 4471 0 FreeSans 250 0 0 0 _37_.X
flabel locali 7850 4709 7884 4743 0 FreeSans 250 0 0 0 _37_.X
flabel locali 7850 4777 7884 4811 0 FreeSans 250 0 0 0 _37_.X
flabel nwell 7894 4879 7928 4913 0 FreeSans 250 0 0 0 _37_.VPB
flabel pwell 7904 4335 7938 4369 0 FreeSans 250 0 0 0 _37_.VNB
rlabel comment 7820 4352 7820 4352 4 _37_.mux2_1
flabel locali 9321 4573 9355 4607 0 FreeSans 200 0 0 0 _47_.A
flabel locali 9505 4709 9539 4743 0 FreeSans 200 0 0 0 _47_.X
flabel locali 9137 4573 9171 4607 0 FreeSans 200 0 0 0 _47_.B
flabel nwell 9137 4879 9171 4913 0 FreeSans 200 0 0 0 _47_.VPB
flabel pwell 9137 4335 9171 4369 0 FreeSans 200 0 0 0 _47_.VNB
flabel metal1 9137 4335 9171 4369 0 FreeSans 200 0 0 0 _47_.VGND
flabel metal1 9137 4879 9171 4913 0 FreeSans 200 0 0 0 _47_.VPWR
rlabel comment 9108 4352 9108 4352 4 _47_.or2_1
flabel locali 9965 4437 9999 4471 0 FreeSans 200 0 0 0 ANTENNA_clkbuf_0_clk_A.DIODE
flabel locali 9965 4709 9999 4743 0 FreeSans 200 0 0 0 ANTENNA_clkbuf_0_clk_A.DIODE
flabel locali 10057 4709 10091 4743 0 FreeSans 200 0 0 0 ANTENNA_clkbuf_0_clk_A.DIODE
flabel locali 9965 4777 9999 4811 0 FreeSans 200 0 0 0 ANTENNA_clkbuf_0_clk_A.DIODE
flabel locali 10057 4777 10091 4811 0 FreeSans 200 0 0 0 ANTENNA_clkbuf_0_clk_A.DIODE
flabel locali 10057 4641 10091 4675 0 FreeSans 200 0 0 0 ANTENNA_clkbuf_0_clk_A.DIODE
flabel locali 9965 4641 9999 4675 0 FreeSans 200 0 0 0 ANTENNA_clkbuf_0_clk_A.DIODE
flabel locali 10057 4573 10091 4607 0 FreeSans 200 0 0 0 ANTENNA_clkbuf_0_clk_A.DIODE
flabel locali 9965 4573 9999 4607 0 FreeSans 200 0 0 0 ANTENNA_clkbuf_0_clk_A.DIODE
flabel locali 9965 4505 9999 4539 0 FreeSans 200 0 0 0 ANTENNA_clkbuf_0_clk_A.DIODE
flabel locali 10057 4505 10091 4539 0 FreeSans 200 0 0 0 ANTENNA_clkbuf_0_clk_A.DIODE
flabel locali 10057 4437 10091 4471 0 FreeSans 200 0 0 0 ANTENNA_clkbuf_0_clk_A.DIODE
flabel metal1 10057 4335 10091 4369 0 FreeSans 200 0 0 0 ANTENNA_clkbuf_0_clk_A.VGND
flabel metal1 10057 4879 10091 4913 0 FreeSans 200 0 0 0 ANTENNA_clkbuf_0_clk_A.VPWR
flabel nwell 10057 4879 10091 4913 0 FreeSans 200 0 0 0 ANTENNA_clkbuf_0_clk_A.VPB
flabel pwell 10057 4335 10091 4369 0 FreeSans 200 0 0 0 ANTENNA_clkbuf_0_clk_A.VNB
rlabel comment 10120 4352 10120 4352 6 ANTENNA_clkbuf_0_clk_A.diode_2
flabel metal1 10977 4335 11011 4369 0 FreeSans 200 0 0 0 FILLER_4_107.VGND
flabel metal1 10977 4879 11011 4913 0 FreeSans 200 0 0 0 FILLER_4_107.VPWR
flabel nwell 10977 4879 11011 4913 0 FreeSans 200 0 0 0 FILLER_4_107.VPB
flabel pwell 10977 4335 11011 4369 0 FreeSans 200 0 0 0 FILLER_4_107.VNB
rlabel comment 10948 4352 10948 4352 4 FILLER_4_107.decap_4
flabel metal1 9597 4335 9631 4369 0 FreeSans 200 0 0 0 FILLER_4_92.VGND
flabel metal1 9597 4879 9631 4913 0 FreeSans 200 0 0 0 FILLER_4_92.VPWR
flabel nwell 9597 4879 9631 4913 0 FreeSans 200 0 0 0 FILLER_4_92.VPB
flabel pwell 9597 4335 9631 4369 0 FreeSans 200 0 0 0 FILLER_4_92.VNB
rlabel comment 9568 4352 9568 4352 4 FILLER_4_92.decap_4
flabel metal1 10149 4335 10183 4369 0 FreeSans 200 0 0 0 FILLER_4_98.VGND
flabel metal1 10149 4879 10183 4913 0 FreeSans 200 0 0 0 FILLER_4_98.VPWR
flabel nwell 10149 4879 10183 4913 0 FreeSans 200 0 0 0 FILLER_4_98.VPB
flabel pwell 10149 4335 10183 4369 0 FreeSans 200 0 0 0 FILLER_4_98.VNB
rlabel comment 10120 4352 10120 4352 4 FILLER_4_98.decap_4
flabel locali 10701 4573 10735 4607 0 FreeSans 200 0 0 0 _26_.A
flabel locali 10885 4709 10919 4743 0 FreeSans 200 0 0 0 _26_.X
flabel locali 10517 4573 10551 4607 0 FreeSans 200 0 0 0 _26_.B
flabel nwell 10517 4879 10551 4913 0 FreeSans 200 0 0 0 _26_.VPB
flabel pwell 10517 4335 10551 4369 0 FreeSans 200 0 0 0 _26_.VNB
flabel metal1 10517 4335 10551 4369 0 FreeSans 200 0 0 0 _26_.VGND
flabel metal1 10517 4879 10551 4913 0 FreeSans 200 0 0 0 _26_.VPWR
rlabel comment 10488 4352 10488 4352 4 _26_.or2_1
flabel metal1 11621 4335 11655 4369 0 FreeSans 200 0 0 0 FILLER_4_114.VGND
flabel metal1 11621 4879 11655 4913 0 FreeSans 200 0 0 0 FILLER_4_114.VPWR
flabel nwell 11621 4879 11655 4913 0 FreeSans 200 0 0 0 FILLER_4_114.VPB
flabel pwell 11621 4335 11655 4369 0 FreeSans 200 0 0 0 FILLER_4_114.VNB
rlabel comment 11592 4352 11592 4352 4 FILLER_4_114.decap_4
flabel metal1 12817 4335 12851 4369 0 FreeSans 200 0 0 0 FILLER_4_127.VGND
flabel metal1 12817 4879 12851 4913 0 FreeSans 200 0 0 0 FILLER_4_127.VPWR
flabel nwell 12817 4879 12851 4913 0 FreeSans 200 0 0 0 FILLER_4_127.VPB
flabel pwell 12817 4335 12851 4369 0 FreeSans 200 0 0 0 FILLER_4_127.VNB
rlabel comment 12788 4352 12788 4352 4 FILLER_4_127.decap_4
flabel metal1 12724 4335 12758 4369 0 FreeSans 200 0 0 0 _31_.VGND
flabel metal1 12724 4879 12758 4913 0 FreeSans 200 0 0 0 _31_.VPWR
flabel locali 12080 4641 12114 4675 0 FreeSans 250 0 0 0 _31_.S
flabel locali 12172 4641 12206 4675 0 FreeSans 250 0 0 0 _31_.S
flabel locali 12264 4505 12298 4539 0 FreeSans 250 0 0 0 _31_.A1
flabel locali 12264 4573 12298 4607 0 FreeSans 250 0 0 0 _31_.A1
flabel locali 12356 4573 12390 4607 0 FreeSans 250 0 0 0 _31_.A0
flabel locali 12724 4437 12758 4471 0 FreeSans 250 0 0 0 _31_.X
flabel locali 12724 4709 12758 4743 0 FreeSans 250 0 0 0 _31_.X
flabel locali 12724 4777 12758 4811 0 FreeSans 250 0 0 0 _31_.X
flabel nwell 12680 4879 12714 4913 0 FreeSans 250 0 0 0 _31_.VPB
flabel pwell 12670 4335 12704 4369 0 FreeSans 250 0 0 0 _31_.VNB
rlabel comment 12788 4352 12788 4352 6 _31_.mux2_1
flabel metal1 13369 4335 13403 4369 0 FreeSans 200 180 0 0 _36_.VGND
flabel metal1 13369 4879 13403 4913 0 FreeSans 200 180 0 0 _36_.VPWR
flabel locali 13185 4437 13219 4471 0 FreeSans 200 180 0 0 _36_.X
flabel locali 13185 4709 13219 4743 0 FreeSans 200 180 0 0 _36_.X
flabel locali 13185 4777 13219 4811 0 FreeSans 200 180 0 0 _36_.X
flabel locali 13369 4573 13403 4607 0 FreeSans 200 180 0 0 _36_.A
flabel nwell 13369 4879 13403 4913 0 FreeSans 200 180 0 0 _36_.VPB
flabel pwell 13369 4335 13403 4369 0 FreeSans 200 180 0 0 _36_.VNB
rlabel comment 13156 4352 13156 4352 4 _36_.clkbuf_1
flabel metal1 11345 4335 11379 4369 0 FreeSans 200 180 0 0 _42_.VGND
flabel metal1 11345 4879 11379 4913 0 FreeSans 200 180 0 0 _42_.VPWR
flabel locali 11529 4437 11563 4471 0 FreeSans 200 180 0 0 _42_.X
flabel locali 11529 4709 11563 4743 0 FreeSans 200 180 0 0 _42_.X
flabel locali 11529 4777 11563 4811 0 FreeSans 200 180 0 0 _42_.X
flabel locali 11345 4573 11379 4607 0 FreeSans 200 180 0 0 _42_.A
flabel nwell 11345 4879 11379 4913 0 FreeSans 200 180 0 0 _42_.VPB
flabel pwell 11345 4335 11379 4369 0 FreeSans 200 180 0 0 _42_.VNB
rlabel comment 11592 4352 11592 4352 6 _42_.clkbuf_1
flabel metal1 13461 4879 13495 4913 0 FreeSans 200 0 0 0 FILLER_4_134.VPWR
flabel metal1 13461 4335 13495 4369 0 FreeSans 200 0 0 0 FILLER_4_134.VGND
flabel nwell 13461 4879 13495 4913 0 FreeSans 200 0 0 0 FILLER_4_134.VPB
flabel pwell 13461 4335 13495 4369 0 FreeSans 200 0 0 0 FILLER_4_134.VNB
rlabel comment 13432 4352 13432 4352 4 FILLER_4_134.decap_6
flabel metal1 14105 4335 14139 4369 0 FreeSans 200 0 0 0 FILLER_4_141.VGND
flabel metal1 14105 4879 14139 4913 0 FreeSans 200 0 0 0 FILLER_4_141.VPWR
flabel nwell 14105 4879 14139 4913 0 FreeSans 200 0 0 0 FILLER_4_141.VPB
flabel pwell 14105 4335 14139 4369 0 FreeSans 200 0 0 0 FILLER_4_141.VNB
rlabel comment 14076 4352 14076 4352 4 FILLER_4_141.decap_12
flabel metal1 14006 4876 14059 4905 0 FreeSans 200 0 0 0 TAP_37.VPWR
flabel metal1 14005 4334 14056 4372 0 FreeSans 200 0 0 0 TAP_37.VGND
rlabel comment 13984 4352 13984 4352 4 TAP_37.tapvpwrvgnd_1
flabel metal1 15669 4335 15703 4369 0 FreeSans 200 0 0 0 FILLER_4_158.VGND
flabel metal1 15669 4879 15703 4913 0 FreeSans 200 0 0 0 FILLER_4_158.VPWR
flabel nwell 15669 4879 15703 4913 0 FreeSans 200 0 0 0 FILLER_4_158.VPB
flabel pwell 15669 4335 15703 4369 0 FreeSans 200 0 0 0 FILLER_4_158.VNB
rlabel comment 15640 4352 15640 4352 4 FILLER_4_158.decap_4
flabel metal1 16313 4335 16347 4369 0 FreeSans 200 0 0 0 FILLER_4_165.VGND
flabel metal1 16313 4879 16347 4913 0 FreeSans 200 0 0 0 FILLER_4_165.VPWR
flabel nwell 16313 4879 16347 4913 0 FreeSans 200 0 0 0 FILLER_4_165.VPB
flabel pwell 16313 4335 16347 4369 0 FreeSans 200 0 0 0 FILLER_4_165.VNB
rlabel comment 16284 4352 16284 4352 4 FILLER_4_165.decap_4
flabel metal1 16957 4335 16991 4369 0 FreeSans 200 0 0 0 FILLER_4_172.VGND
flabel metal1 16957 4879 16991 4913 0 FreeSans 200 0 0 0 FILLER_4_172.VPWR
flabel nwell 16957 4879 16991 4913 0 FreeSans 200 0 0 0 FILLER_4_172.VPB
flabel pwell 16957 4335 16991 4369 0 FreeSans 200 0 0 0 FILLER_4_172.VNB
rlabel comment 16928 4352 16928 4352 4 FILLER_4_172.decap_12
flabel locali 15393 4573 15427 4607 0 FreeSans 200 0 0 0 _29_.A
flabel locali 15577 4709 15611 4743 0 FreeSans 200 0 0 0 _29_.X
flabel locali 15209 4573 15243 4607 0 FreeSans 200 0 0 0 _29_.B
flabel nwell 15209 4879 15243 4913 0 FreeSans 200 0 0 0 _29_.VPB
flabel pwell 15209 4335 15243 4369 0 FreeSans 200 0 0 0 _29_.VNB
flabel metal1 15209 4335 15243 4369 0 FreeSans 200 0 0 0 _29_.VGND
flabel metal1 15209 4879 15243 4913 0 FreeSans 200 0 0 0 _29_.VPWR
rlabel comment 15180 4352 15180 4352 4 _29_.or2_1
flabel metal1 16865 4335 16899 4369 0 FreeSans 200 180 0 0 _30_.VGND
flabel metal1 16865 4879 16899 4913 0 FreeSans 200 180 0 0 _30_.VPWR
flabel locali 16681 4437 16715 4471 0 FreeSans 200 180 0 0 _30_.X
flabel locali 16681 4709 16715 4743 0 FreeSans 200 180 0 0 _30_.X
flabel locali 16681 4777 16715 4811 0 FreeSans 200 180 0 0 _30_.X
flabel locali 16865 4573 16899 4607 0 FreeSans 200 180 0 0 _30_.A
flabel nwell 16865 4879 16899 4913 0 FreeSans 200 180 0 0 _30_.VPB
flabel pwell 16865 4335 16899 4369 0 FreeSans 200 180 0 0 _30_.VNB
rlabel comment 16652 4352 16652 4352 4 _30_.clkbuf_1
flabel metal1 16221 4335 16255 4369 0 FreeSans 200 180 0 0 _33_.VGND
flabel metal1 16221 4879 16255 4913 0 FreeSans 200 180 0 0 _33_.VPWR
flabel locali 16037 4437 16071 4471 0 FreeSans 200 180 0 0 _33_.X
flabel locali 16037 4709 16071 4743 0 FreeSans 200 180 0 0 _33_.X
flabel locali 16037 4777 16071 4811 0 FreeSans 200 180 0 0 _33_.X
flabel locali 16221 4573 16255 4607 0 FreeSans 200 180 0 0 _33_.A
flabel nwell 16221 4879 16255 4913 0 FreeSans 200 180 0 0 _33_.VPB
flabel pwell 16221 4335 16255 4369 0 FreeSans 200 180 0 0 _33_.VNB
rlabel comment 16008 4352 16008 4352 4 _33_.clkbuf_1
flabel metal1 18061 4879 18095 4913 0 FreeSans 200 0 0 0 FILLER_4_184.VPWR
flabel metal1 18061 4335 18095 4369 0 FreeSans 200 0 0 0 FILLER_4_184.VGND
flabel nwell 18061 4879 18095 4913 0 FreeSans 200 0 0 0 FILLER_4_184.VPB
flabel pwell 18061 4335 18095 4369 0 FreeSans 200 0 0 0 FILLER_4_184.VNB
rlabel comment 18032 4352 18032 4352 4 FILLER_4_184.decap_6
flabel metal1 18797 4879 18831 4913 0 FreeSans 200 0 0 0 PHY_9.VPWR
flabel metal1 18797 4335 18831 4369 0 FreeSans 200 0 0 0 PHY_9.VGND
flabel nwell 18797 4879 18831 4913 0 FreeSans 200 0 0 0 PHY_9.VPB
flabel pwell 18797 4335 18831 4369 0 FreeSans 200 0 0 0 PHY_9.VNB
rlabel comment 18860 4352 18860 4352 6 PHY_9.decap_3
flabel metal1 2513 4879 2547 4913 0 FreeSans 200 0 0 0 FILLER_5_15.VPWR
flabel metal1 2513 5423 2547 5457 0 FreeSans 200 0 0 0 FILLER_5_15.VGND
flabel nwell 2513 4879 2547 4913 0 FreeSans 200 0 0 0 FILLER_5_15.VPB
flabel pwell 2513 5423 2547 5457 0 FreeSans 200 0 0 0 FILLER_5_15.VNB
rlabel comment 2484 5440 2484 5440 2 FILLER_5_15.decap_3
flabel metal1 1409 5423 1443 5457 0 FreeSans 200 0 0 0 FILLER_5_3.VGND
flabel metal1 1409 4879 1443 4913 0 FreeSans 200 0 0 0 FILLER_5_3.VPWR
flabel nwell 1409 4879 1443 4913 0 FreeSans 200 0 0 0 FILLER_5_3.VPB
flabel pwell 1409 5423 1443 5457 0 FreeSans 200 0 0 0 FILLER_5_3.VNB
rlabel comment 1380 5440 1380 5440 2 FILLER_5_3.decap_12
flabel metal1 1133 4879 1167 4913 0 FreeSans 200 0 0 0 PHY_10.VPWR
flabel metal1 1133 5423 1167 5457 0 FreeSans 200 0 0 0 PHY_10.VGND
flabel nwell 1133 4879 1167 4913 0 FreeSans 200 0 0 0 PHY_10.VPB
flabel pwell 1133 5423 1167 5457 0 FreeSans 200 0 0 0 PHY_10.VNB
rlabel comment 1104 5440 1104 5440 2 PHY_10.decap_3
flabel locali 4536 4981 4570 5015 0 FreeSans 400 0 0 0 _52_.Q
flabel locali 4536 5049 4570 5083 0 FreeSans 400 0 0 0 _52_.Q
flabel locali 4536 5117 4570 5151 0 FreeSans 400 0 0 0 _52_.Q
flabel locali 4536 5321 4570 5355 0 FreeSans 400 0 0 0 _52_.Q
flabel locali 4241 5253 4275 5287 0 FreeSans 400 0 0 0 _52_.RESET_B
flabel locali 3065 5117 3099 5151 0 FreeSans 400 0 0 0 _52_.D
flabel locali 2790 5117 2824 5151 0 FreeSans 400 0 0 0 _52_.CLK
flabel locali 2790 5185 2824 5219 0 FreeSans 400 0 0 0 _52_.CLK
flabel locali 4241 5185 4275 5219 0 FreeSans 400 0 0 0 _52_.RESET_B
flabel metal1 2789 5423 2823 5457 0 FreeSans 200 0 0 0 _52_.VGND
flabel metal1 2789 4879 2823 4913 0 FreeSans 200 0 0 0 _52_.VPWR
flabel nwell 2789 4879 2823 4913 0 FreeSans 200 0 0 0 _52_.VPB
flabel pwell 2789 5423 2823 5457 0 FreeSans 200 0 0 0 _52_.VNB
rlabel comment 2760 5440 2760 5440 2 _52_.dfrtp_1
flabel metal1 4629 5423 4663 5457 0 FreeSans 200 0 0 0 FILLER_5_38.VGND
flabel metal1 4629 4879 4663 4913 0 FreeSans 200 0 0 0 FILLER_5_38.VPWR
flabel nwell 4629 4879 4663 4913 0 FreeSans 200 0 0 0 FILLER_5_38.VPB
flabel pwell 4629 5423 4663 5457 0 FreeSans 200 0 0 0 FILLER_5_38.VNB
rlabel comment 4600 5440 4600 5440 2 FILLER_5_38.decap_12
flabel metal1 5733 4879 5767 4913 0 FreeSans 200 0 0 0 FILLER_5_50.VPWR
flabel metal1 5733 5423 5767 5457 0 FreeSans 200 0 0 0 FILLER_5_50.VGND
flabel nwell 5733 4879 5767 4913 0 FreeSans 200 0 0 0 FILLER_5_50.VPB
flabel pwell 5733 5423 5767 5457 0 FreeSans 200 0 0 0 FILLER_5_50.VNB
rlabel comment 5704 5440 5704 5440 2 FILLER_5_50.decap_6
flabel metal1 6377 4879 6411 4913 0 FreeSans 200 0 0 0 FILLER_5_57.VPWR
flabel metal1 6377 5423 6411 5457 0 FreeSans 200 0 0 0 FILLER_5_57.VGND
flabel nwell 6377 4879 6411 4913 0 FreeSans 200 0 0 0 FILLER_5_57.VPB
flabel pwell 6377 5423 6411 5457 0 FreeSans 200 0 0 0 FILLER_5_57.VNB
rlabel comment 6348 5440 6348 5440 2 FILLER_5_57.decap_3
flabel metal1 6278 4887 6331 4916 0 FreeSans 200 0 0 0 TAP_38.VPWR
flabel metal1 6277 5420 6328 5458 0 FreeSans 200 0 0 0 TAP_38.VGND
rlabel comment 6256 5440 6256 5440 2 TAP_38.tapvpwrvgnd_1
flabel metal1 6654 5423 6688 5457 0 FreeSans 200 0 0 0 _43_.VGND
flabel metal1 6654 4879 6688 4913 0 FreeSans 200 0 0 0 _43_.VPWR
flabel locali 7298 5117 7332 5151 0 FreeSans 250 0 0 0 _43_.S
flabel locali 7206 5117 7240 5151 0 FreeSans 250 0 0 0 _43_.S
flabel locali 7114 5253 7148 5287 0 FreeSans 250 0 0 0 _43_.A1
flabel locali 7114 5185 7148 5219 0 FreeSans 250 0 0 0 _43_.A1
flabel locali 7022 5185 7056 5219 0 FreeSans 250 0 0 0 _43_.A0
flabel locali 6654 5321 6688 5355 0 FreeSans 250 0 0 0 _43_.X
flabel locali 6654 5049 6688 5083 0 FreeSans 250 0 0 0 _43_.X
flabel locali 6654 4981 6688 5015 0 FreeSans 250 0 0 0 _43_.X
flabel nwell 6698 4879 6732 4913 0 FreeSans 250 0 0 0 _43_.VPB
flabel pwell 6708 5423 6742 5457 0 FreeSans 250 0 0 0 _43_.VNB
rlabel comment 6624 5440 6624 5440 2 _43_.mux2_1
flabel metal1 7481 5423 7515 5457 0 FreeSans 200 0 0 0 FILLER_5_69.VGND
flabel metal1 7481 4879 7515 4913 0 FreeSans 200 0 0 0 FILLER_5_69.VPWR
flabel nwell 7481 4879 7515 4913 0 FreeSans 200 0 0 0 FILLER_5_69.VPB
flabel pwell 7481 5423 7515 5457 0 FreeSans 200 0 0 0 FILLER_5_69.VNB
rlabel comment 7452 5440 7452 5440 2 FILLER_5_69.decap_4
flabel locali 9596 4981 9630 5015 0 FreeSans 400 0 0 0 _63_.Q
flabel locali 9596 5049 9630 5083 0 FreeSans 400 0 0 0 _63_.Q
flabel locali 9596 5117 9630 5151 0 FreeSans 400 0 0 0 _63_.Q
flabel locali 9596 5321 9630 5355 0 FreeSans 400 0 0 0 _63_.Q
flabel locali 9301 5253 9335 5287 0 FreeSans 400 0 0 0 _63_.RESET_B
flabel locali 8125 5117 8159 5151 0 FreeSans 400 0 0 0 _63_.D
flabel locali 7850 5117 7884 5151 0 FreeSans 400 0 0 0 _63_.CLK
flabel locali 7850 5185 7884 5219 0 FreeSans 400 0 0 0 _63_.CLK
flabel locali 9301 5185 9335 5219 0 FreeSans 400 0 0 0 _63_.RESET_B
flabel metal1 7849 5423 7883 5457 0 FreeSans 200 0 0 0 _63_.VGND
flabel metal1 7849 4879 7883 4913 0 FreeSans 200 0 0 0 _63_.VPWR
flabel nwell 7849 4879 7883 4913 0 FreeSans 200 0 0 0 _63_.VPB
flabel pwell 7849 5423 7883 5457 0 FreeSans 200 0 0 0 _63_.VNB
rlabel comment 7820 5440 7820 5440 2 _63_.dfrtp_1
flabel metal1 10885 4879 10919 4913 0 FreeSans 200 0 0 0 FILLER_5_106.VPWR
flabel metal1 10885 5423 10919 5457 0 FreeSans 200 0 0 0 FILLER_5_106.VGND
flabel nwell 10885 4879 10919 4913 0 FreeSans 200 0 0 0 FILLER_5_106.VPB
flabel pwell 10885 5423 10919 5457 0 FreeSans 200 0 0 0 FILLER_5_106.VNB
rlabel comment 10856 5440 10856 5440 2 FILLER_5_106.decap_6
flabel metal1 9689 5423 9723 5457 0 FreeSans 200 0 0 0 FILLER_5_93.VGND
flabel metal1 9689 4879 9723 4913 0 FreeSans 200 0 0 0 FILLER_5_93.VPWR
flabel nwell 9689 4879 9723 4913 0 FreeSans 200 0 0 0 FILLER_5_93.VPB
flabel pwell 9689 5423 9723 5457 0 FreeSans 200 0 0 0 FILLER_5_93.VNB
rlabel comment 9660 5440 9660 5440 2 FILLER_5_93.decap_4
flabel metal1 10792 5423 10826 5457 0 FreeSans 200 0 0 0 _25_.VGND
flabel metal1 10792 4879 10826 4913 0 FreeSans 200 0 0 0 _25_.VPWR
flabel locali 10148 5117 10182 5151 0 FreeSans 250 0 0 0 _25_.S
flabel locali 10240 5117 10274 5151 0 FreeSans 250 0 0 0 _25_.S
flabel locali 10332 5253 10366 5287 0 FreeSans 250 0 0 0 _25_.A1
flabel locali 10332 5185 10366 5219 0 FreeSans 250 0 0 0 _25_.A1
flabel locali 10424 5185 10458 5219 0 FreeSans 250 0 0 0 _25_.A0
flabel locali 10792 5321 10826 5355 0 FreeSans 250 0 0 0 _25_.X
flabel locali 10792 5049 10826 5083 0 FreeSans 250 0 0 0 _25_.X
flabel locali 10792 4981 10826 5015 0 FreeSans 250 0 0 0 _25_.X
flabel nwell 10748 4879 10782 4913 0 FreeSans 250 0 0 0 _25_.VPB
flabel pwell 10738 5423 10772 5457 0 FreeSans 250 0 0 0 _25_.VNB
rlabel comment 10856 5440 10856 5440 8 _25_.mux2_1
flabel metal1 11520 5422 11573 5454 0 FreeSans 200 0 0 0 FILLER_5_113.VGND
flabel metal1 11521 4879 11573 4910 0 FreeSans 200 0 0 0 FILLER_5_113.VPWR
flabel nwell 11528 4887 11562 4905 0 FreeSans 200 0 0 0 FILLER_5_113.VPB
flabel pwell 11531 5428 11563 5450 0 FreeSans 200 0 0 0 FILLER_5_113.VNB
rlabel comment 11500 5440 11500 5440 2 FILLER_5_113.fill_2
flabel metal1 12541 5423 12575 5457 0 FreeSans 200 0 0 0 FILLER_5_124.VGND
flabel metal1 12541 4879 12575 4913 0 FreeSans 200 0 0 0 FILLER_5_124.VPWR
flabel nwell 12541 4879 12575 4913 0 FreeSans 200 0 0 0 FILLER_5_124.VPB
flabel pwell 12541 5423 12575 5457 0 FreeSans 200 0 0 0 FILLER_5_124.VNB
rlabel comment 12512 5440 12512 5440 2 FILLER_5_124.decap_4
flabel metal1 11430 4887 11483 4916 0 FreeSans 200 0 0 0 TAP_39.VPWR
flabel metal1 11429 5420 11480 5458 0 FreeSans 200 0 0 0 TAP_39.VGND
rlabel comment 11408 5440 11408 5440 2 TAP_39.tapvpwrvgnd_1
flabel metal1 13644 5423 13678 5457 0 FreeSans 200 0 0 0 _28_.VGND
flabel metal1 13644 4879 13678 4913 0 FreeSans 200 0 0 0 _28_.VPWR
flabel locali 13000 5117 13034 5151 0 FreeSans 250 0 0 0 _28_.S
flabel locali 13092 5117 13126 5151 0 FreeSans 250 0 0 0 _28_.S
flabel locali 13184 5253 13218 5287 0 FreeSans 250 0 0 0 _28_.A1
flabel locali 13184 5185 13218 5219 0 FreeSans 250 0 0 0 _28_.A1
flabel locali 13276 5185 13310 5219 0 FreeSans 250 0 0 0 _28_.A0
flabel locali 13644 5321 13678 5355 0 FreeSans 250 0 0 0 _28_.X
flabel locali 13644 5049 13678 5083 0 FreeSans 250 0 0 0 _28_.X
flabel locali 13644 4981 13678 5015 0 FreeSans 250 0 0 0 _28_.X
flabel nwell 13600 4879 13634 4913 0 FreeSans 250 0 0 0 _28_.VPB
flabel pwell 13590 5423 13624 5457 0 FreeSans 250 0 0 0 _28_.VNB
rlabel comment 13708 5440 13708 5440 8 _28_.mux2_1
flabel metal1 11714 5423 11748 5457 0 FreeSans 200 0 0 0 _34_.VGND
flabel metal1 11714 4879 11748 4913 0 FreeSans 200 0 0 0 _34_.VPWR
flabel locali 12358 5117 12392 5151 0 FreeSans 250 0 0 0 _34_.S
flabel locali 12266 5117 12300 5151 0 FreeSans 250 0 0 0 _34_.S
flabel locali 12174 5253 12208 5287 0 FreeSans 250 0 0 0 _34_.A1
flabel locali 12174 5185 12208 5219 0 FreeSans 250 0 0 0 _34_.A1
flabel locali 12082 5185 12116 5219 0 FreeSans 250 0 0 0 _34_.A0
flabel locali 11714 5321 11748 5355 0 FreeSans 250 0 0 0 _34_.X
flabel locali 11714 5049 11748 5083 0 FreeSans 250 0 0 0 _34_.X
flabel locali 11714 4981 11748 5015 0 FreeSans 250 0 0 0 _34_.X
flabel nwell 11758 4879 11792 4913 0 FreeSans 250 0 0 0 _34_.VPB
flabel pwell 11768 5423 11802 5457 0 FreeSans 250 0 0 0 _34_.VNB
rlabel comment 11684 5440 11684 5440 2 _34_.mux2_1
flabel metal1 13737 5423 13771 5457 0 FreeSans 200 0 0 0 FILLER_5_137.VGND
flabel metal1 13737 4879 13771 4913 0 FreeSans 200 0 0 0 FILLER_5_137.VPWR
flabel nwell 13737 4879 13771 4913 0 FreeSans 200 0 0 0 FILLER_5_137.VPB
flabel pwell 13737 5423 13771 5457 0 FreeSans 200 0 0 0 FILLER_5_137.VNB
rlabel comment 13708 5440 13708 5440 2 FILLER_5_137.decap_12
flabel metal1 14841 5423 14875 5457 0 FreeSans 200 0 0 0 FILLER_5_149.VGND
flabel metal1 14841 4879 14875 4913 0 FreeSans 200 0 0 0 FILLER_5_149.VPWR
flabel nwell 14841 4879 14875 4913 0 FreeSans 200 0 0 0 FILLER_5_149.VPB
flabel pwell 14841 5423 14875 5457 0 FreeSans 200 0 0 0 FILLER_5_149.VNB
rlabel comment 14812 5440 14812 5440 2 FILLER_5_149.decap_12
flabel metal1 15945 4879 15979 4913 0 FreeSans 200 0 0 0 FILLER_5_161.VPWR
flabel metal1 15945 5423 15979 5457 0 FreeSans 200 0 0 0 FILLER_5_161.VGND
flabel nwell 15945 4879 15979 4913 0 FreeSans 200 0 0 0 FILLER_5_161.VPB
flabel pwell 15945 5423 15979 5457 0 FreeSans 200 0 0 0 FILLER_5_161.VNB
rlabel comment 15916 5440 15916 5440 2 FILLER_5_161.decap_6
flabel metal1 16490 4883 16526 4913 0 FreeSans 250 0 0 0 FILLER_5_167.VPWR
flabel metal1 16490 5424 16526 5453 0 FreeSans 250 0 0 0 FILLER_5_167.VGND
flabel nwell 16499 4889 16519 4906 0 FreeSans 200 0 0 0 FILLER_5_167.VPB
flabel pwell 16496 5429 16520 5451 0 FreeSans 200 0 0 0 FILLER_5_167.VNB
rlabel comment 16468 5440 16468 5440 2 FILLER_5_167.fill_1
flabel metal1 16681 5423 16715 5457 0 FreeSans 200 0 0 0 FILLER_5_169.VGND
flabel metal1 16681 4879 16715 4913 0 FreeSans 200 0 0 0 FILLER_5_169.VPWR
flabel nwell 16681 4879 16715 4913 0 FreeSans 200 0 0 0 FILLER_5_169.VPB
flabel pwell 16681 5423 16715 5457 0 FreeSans 200 0 0 0 FILLER_5_169.VNB
rlabel comment 16652 5440 16652 5440 2 FILLER_5_169.decap_12
flabel metal1 16582 4887 16635 4916 0 FreeSans 200 0 0 0 TAP_40.VPWR
flabel metal1 16581 5420 16632 5458 0 FreeSans 200 0 0 0 TAP_40.VGND
rlabel comment 16560 5440 16560 5440 2 TAP_40.tapvpwrvgnd_1
flabel metal1 17785 4879 17819 4913 0 FreeSans 200 0 0 0 FILLER_5_181.VPWR
flabel metal1 17785 5423 17819 5457 0 FreeSans 200 0 0 0 FILLER_5_181.VGND
flabel nwell 17785 4879 17819 4913 0 FreeSans 200 0 0 0 FILLER_5_181.VPB
flabel pwell 17785 5423 17819 5457 0 FreeSans 200 0 0 0 FILLER_5_181.VNB
rlabel comment 17756 5440 17756 5440 2 FILLER_5_181.decap_8
flabel metal1 18514 4883 18550 4913 0 FreeSans 250 0 0 0 FILLER_5_189.VPWR
flabel metal1 18514 5424 18550 5453 0 FreeSans 250 0 0 0 FILLER_5_189.VGND
flabel nwell 18523 4889 18543 4906 0 FreeSans 200 0 0 0 FILLER_5_189.VPB
flabel pwell 18520 5429 18544 5451 0 FreeSans 200 0 0 0 FILLER_5_189.VNB
rlabel comment 18492 5440 18492 5440 2 FILLER_5_189.fill_1
flabel metal1 18797 4879 18831 4913 0 FreeSans 200 0 0 0 PHY_11.VPWR
flabel metal1 18797 5423 18831 5457 0 FreeSans 200 0 0 0 PHY_11.VGND
flabel nwell 18797 4879 18831 4913 0 FreeSans 200 0 0 0 PHY_11.VPB
flabel pwell 18797 5423 18831 5457 0 FreeSans 200 0 0 0 PHY_11.VNB
rlabel comment 18860 5440 18860 5440 8 PHY_11.decap_3
flabel metal1 2513 5423 2547 5457 0 FreeSans 200 0 0 0 FILLER_6_15.VGND
flabel metal1 2513 5967 2547 6001 0 FreeSans 200 0 0 0 FILLER_6_15.VPWR
flabel nwell 2513 5967 2547 6001 0 FreeSans 200 0 0 0 FILLER_6_15.VPB
flabel pwell 2513 5423 2547 5457 0 FreeSans 200 0 0 0 FILLER_6_15.VNB
rlabel comment 2484 5440 2484 5440 4 FILLER_6_15.decap_12
flabel metal1 1409 5423 1443 5457 0 FreeSans 200 0 0 0 FILLER_6_3.VGND
flabel metal1 1409 5967 1443 6001 0 FreeSans 200 0 0 0 FILLER_6_3.VPWR
flabel nwell 1409 5967 1443 6001 0 FreeSans 200 0 0 0 FILLER_6_3.VPB
flabel pwell 1409 5423 1443 5457 0 FreeSans 200 0 0 0 FILLER_6_3.VNB
rlabel comment 1380 5440 1380 5440 4 FILLER_6_3.decap_12
flabel metal1 2513 6511 2547 6545 0 FreeSans 200 0 0 0 FILLER_7_15.VGND
flabel metal1 2513 5967 2547 6001 0 FreeSans 200 0 0 0 FILLER_7_15.VPWR
flabel nwell 2513 5967 2547 6001 0 FreeSans 200 0 0 0 FILLER_7_15.VPB
flabel pwell 2513 6511 2547 6545 0 FreeSans 200 0 0 0 FILLER_7_15.VNB
rlabel comment 2484 6528 2484 6528 2 FILLER_7_15.decap_12
flabel metal1 1409 6511 1443 6545 0 FreeSans 200 0 0 0 FILLER_7_3.VGND
flabel metal1 1409 5967 1443 6001 0 FreeSans 200 0 0 0 FILLER_7_3.VPWR
flabel nwell 1409 5967 1443 6001 0 FreeSans 200 0 0 0 FILLER_7_3.VPB
flabel pwell 1409 6511 1443 6545 0 FreeSans 200 0 0 0 FILLER_7_3.VNB
rlabel comment 1380 6528 1380 6528 2 FILLER_7_3.decap_12
flabel metal1 1133 5967 1167 6001 0 FreeSans 200 0 0 0 PHY_12.VPWR
flabel metal1 1133 5423 1167 5457 0 FreeSans 200 0 0 0 PHY_12.VGND
flabel nwell 1133 5967 1167 6001 0 FreeSans 200 0 0 0 PHY_12.VPB
flabel pwell 1133 5423 1167 5457 0 FreeSans 200 0 0 0 PHY_12.VNB
rlabel comment 1104 5440 1104 5440 4 PHY_12.decap_3
flabel metal1 1133 5967 1167 6001 0 FreeSans 200 0 0 0 PHY_14.VPWR
flabel metal1 1133 6511 1167 6545 0 FreeSans 200 0 0 0 PHY_14.VGND
flabel nwell 1133 5967 1167 6001 0 FreeSans 200 0 0 0 PHY_14.VPB
flabel pwell 1133 6511 1167 6545 0 FreeSans 200 0 0 0 PHY_14.VNB
rlabel comment 1104 6528 1104 6528 2 PHY_14.decap_3
flabel metal1 3610 5967 3646 5997 0 FreeSans 250 0 0 0 FILLER_6_27.VPWR
flabel metal1 3610 5427 3646 5456 0 FreeSans 250 0 0 0 FILLER_6_27.VGND
flabel nwell 3619 5974 3639 5991 0 FreeSans 200 0 0 0 FILLER_6_27.VPB
flabel pwell 3616 5429 3640 5451 0 FreeSans 200 0 0 0 FILLER_6_27.VNB
rlabel comment 3588 5440 3588 5440 4 FILLER_6_27.fill_1
flabel metal1 3801 5423 3835 5457 0 FreeSans 200 0 0 0 FILLER_6_29.VGND
flabel metal1 3801 5967 3835 6001 0 FreeSans 200 0 0 0 FILLER_6_29.VPWR
flabel nwell 3801 5967 3835 6001 0 FreeSans 200 0 0 0 FILLER_6_29.VPB
flabel pwell 3801 5423 3835 5457 0 FreeSans 200 0 0 0 FILLER_6_29.VNB
rlabel comment 3772 5440 3772 5440 4 FILLER_6_29.decap_12
flabel metal1 4905 5423 4939 5457 0 FreeSans 200 0 0 0 FILLER_6_41.VGND
flabel metal1 4905 5967 4939 6001 0 FreeSans 200 0 0 0 FILLER_6_41.VPWR
flabel nwell 4905 5967 4939 6001 0 FreeSans 200 0 0 0 FILLER_6_41.VPB
flabel pwell 4905 5423 4939 5457 0 FreeSans 200 0 0 0 FILLER_6_41.VNB
rlabel comment 4876 5440 4876 5440 4 FILLER_6_41.decap_12
flabel metal1 3617 6511 3651 6545 0 FreeSans 200 0 0 0 FILLER_7_27.VGND
flabel metal1 3617 5967 3651 6001 0 FreeSans 200 0 0 0 FILLER_7_27.VPWR
flabel nwell 3617 5967 3651 6001 0 FreeSans 200 0 0 0 FILLER_7_27.VPB
flabel pwell 3617 6511 3651 6545 0 FreeSans 200 0 0 0 FILLER_7_27.VNB
rlabel comment 3588 6528 3588 6528 2 FILLER_7_27.decap_12
flabel metal1 4721 6511 4755 6545 0 FreeSans 200 0 0 0 FILLER_7_39.VGND
flabel metal1 4721 5967 4755 6001 0 FreeSans 200 0 0 0 FILLER_7_39.VPWR
flabel nwell 4721 5967 4755 6001 0 FreeSans 200 0 0 0 FILLER_7_39.VPB
flabel pwell 4721 6511 4755 6545 0 FreeSans 200 0 0 0 FILLER_7_39.VNB
rlabel comment 4692 6528 4692 6528 2 FILLER_7_39.decap_12
flabel metal1 3702 5964 3755 5993 0 FreeSans 200 0 0 0 TAP_41.VPWR
flabel metal1 3701 5422 3752 5460 0 FreeSans 200 0 0 0 TAP_41.VGND
rlabel comment 3680 5440 3680 5440 4 TAP_41.tapvpwrvgnd_1
flabel metal1 6009 5967 6043 6001 0 FreeSans 200 0 0 0 FILLER_6_53.VPWR
flabel metal1 6009 5423 6043 5457 0 FreeSans 200 0 0 0 FILLER_6_53.VGND
flabel nwell 6009 5967 6043 6001 0 FreeSans 200 0 0 0 FILLER_6_53.VPB
flabel pwell 6009 5423 6043 5457 0 FreeSans 200 0 0 0 FILLER_6_53.VNB
rlabel comment 5980 5440 5980 5440 4 FILLER_6_53.decap_8
flabel metal1 7021 5967 7055 6001 0 FreeSans 200 0 0 0 FILLER_6_64.VPWR
flabel metal1 7021 5423 7055 5457 0 FreeSans 200 0 0 0 FILLER_6_64.VGND
flabel nwell 7021 5967 7055 6001 0 FreeSans 200 0 0 0 FILLER_6_64.VPB
flabel pwell 7021 5423 7055 5457 0 FreeSans 200 0 0 0 FILLER_6_64.VNB
rlabel comment 6992 5440 6992 5440 4 FILLER_6_64.decap_6
flabel metal1 5825 6511 5859 6545 0 FreeSans 200 0 0 0 FILLER_7_51.VGND
flabel metal1 5825 5967 5859 6001 0 FreeSans 200 0 0 0 FILLER_7_51.VPWR
flabel nwell 5825 5967 5859 6001 0 FreeSans 200 0 0 0 FILLER_7_51.VPB
flabel pwell 5825 6511 5859 6545 0 FreeSans 200 0 0 0 FILLER_7_51.VNB
rlabel comment 5796 6528 5796 6528 2 FILLER_7_51.decap_4
flabel metal1 6186 5971 6222 6001 0 FreeSans 250 0 0 0 FILLER_7_55.VPWR
flabel metal1 6186 6512 6222 6541 0 FreeSans 250 0 0 0 FILLER_7_55.VGND
flabel nwell 6195 5977 6215 5994 0 FreeSans 200 0 0 0 FILLER_7_55.VPB
flabel pwell 6192 6517 6216 6539 0 FreeSans 200 0 0 0 FILLER_7_55.VNB
rlabel comment 6164 6528 6164 6528 2 FILLER_7_55.fill_1
flabel metal1 6377 6511 6411 6545 0 FreeSans 200 0 0 0 FILLER_7_57.VGND
flabel metal1 6377 5967 6411 6001 0 FreeSans 200 0 0 0 FILLER_7_57.VPWR
flabel nwell 6377 5967 6411 6001 0 FreeSans 200 0 0 0 FILLER_7_57.VPB
flabel pwell 6377 6511 6411 6545 0 FreeSans 200 0 0 0 FILLER_7_57.VNB
rlabel comment 6348 6528 6348 6528 2 FILLER_7_57.decap_12
flabel metal1 6278 5975 6331 6004 0 FreeSans 200 0 0 0 TAP_44.VPWR
flabel metal1 6277 6508 6328 6546 0 FreeSans 200 0 0 0 TAP_44.VGND
rlabel comment 6256 6528 6256 6528 2 TAP_44.tapvpwrvgnd_1
flabel metal1 6929 5423 6963 5457 0 FreeSans 200 180 0 0 _45_.VGND
flabel metal1 6929 5967 6963 6001 0 FreeSans 200 180 0 0 _45_.VPWR
flabel locali 6745 5525 6779 5559 0 FreeSans 200 180 0 0 _45_.X
flabel locali 6745 5797 6779 5831 0 FreeSans 200 180 0 0 _45_.X
flabel locali 6745 5865 6779 5899 0 FreeSans 200 180 0 0 _45_.X
flabel locali 6929 5661 6963 5695 0 FreeSans 200 180 0 0 _45_.A
flabel nwell 6929 5967 6963 6001 0 FreeSans 200 180 0 0 _45_.VPB
flabel pwell 6929 5423 6963 5457 0 FreeSans 200 180 0 0 _45_.VNB
rlabel comment 6716 5440 6716 5440 4 _45_.clkbuf_1
flabel metal1 8401 5423 8435 5457 0 FreeSans 200 0 0 0 FILLER_6_79.VGND
flabel metal1 8401 5967 8435 6001 0 FreeSans 200 0 0 0 FILLER_6_79.VPWR
flabel nwell 8401 5967 8435 6001 0 FreeSans 200 0 0 0 FILLER_6_79.VPB
flabel pwell 8401 5423 8435 5457 0 FreeSans 200 0 0 0 FILLER_6_79.VNB
rlabel comment 8372 5440 8372 5440 4 FILLER_6_79.decap_4
flabel metal1 8762 5967 8798 5997 0 FreeSans 250 0 0 0 FILLER_6_83.VPWR
flabel metal1 8762 5427 8798 5456 0 FreeSans 250 0 0 0 FILLER_6_83.VGND
flabel nwell 8771 5974 8791 5991 0 FreeSans 200 0 0 0 FILLER_6_83.VPB
flabel pwell 8768 5429 8792 5451 0 FreeSans 200 0 0 0 FILLER_6_83.VNB
rlabel comment 8740 5440 8740 5440 4 FILLER_6_83.fill_1
flabel metal1 8953 5423 8987 5457 0 FreeSans 200 0 0 0 FILLER_6_85.VGND
flabel metal1 8953 5967 8987 6001 0 FreeSans 200 0 0 0 FILLER_6_85.VPWR
flabel nwell 8953 5967 8987 6001 0 FreeSans 200 0 0 0 FILLER_6_85.VPB
flabel pwell 8953 5423 8987 5457 0 FreeSans 200 0 0 0 FILLER_6_85.VNB
rlabel comment 8924 5440 8924 5440 4 FILLER_6_85.decap_12
flabel metal1 7481 5967 7515 6001 0 FreeSans 200 0 0 0 FILLER_7_69.VPWR
flabel metal1 7481 6511 7515 6545 0 FreeSans 200 0 0 0 FILLER_7_69.VGND
flabel nwell 7481 5967 7515 6001 0 FreeSans 200 0 0 0 FILLER_7_69.VPB
flabel pwell 7481 6511 7515 6545 0 FreeSans 200 0 0 0 FILLER_7_69.VNB
rlabel comment 7452 6528 7452 6528 2 FILLER_7_69.decap_6
flabel metal1 8493 6511 8527 6545 0 FreeSans 200 0 0 0 FILLER_7_80.VGND
flabel metal1 8493 5967 8527 6001 0 FreeSans 200 0 0 0 FILLER_7_80.VPWR
flabel nwell 8493 5967 8527 6001 0 FreeSans 200 0 0 0 FILLER_7_80.VPB
flabel pwell 8493 6511 8527 6545 0 FreeSans 200 0 0 0 FILLER_7_80.VNB
rlabel comment 8464 6528 8464 6528 2 FILLER_7_80.decap_12
flabel metal1 8854 5964 8907 5993 0 FreeSans 200 0 0 0 TAP_42.VPWR
flabel metal1 8853 5422 8904 5460 0 FreeSans 200 0 0 0 TAP_42.VGND
rlabel comment 8832 5440 8832 5440 4 TAP_42.tapvpwrvgnd_1
flabel metal1 8308 5423 8342 5457 0 FreeSans 200 0 0 0 _40_.VGND
flabel metal1 8308 5967 8342 6001 0 FreeSans 200 0 0 0 _40_.VPWR
flabel locali 7664 5729 7698 5763 0 FreeSans 250 0 0 0 _40_.S
flabel locali 7756 5729 7790 5763 0 FreeSans 250 0 0 0 _40_.S
flabel locali 7848 5593 7882 5627 0 FreeSans 250 0 0 0 _40_.A1
flabel locali 7848 5661 7882 5695 0 FreeSans 250 0 0 0 _40_.A1
flabel locali 7940 5661 7974 5695 0 FreeSans 250 0 0 0 _40_.A0
flabel locali 8308 5525 8342 5559 0 FreeSans 250 0 0 0 _40_.X
flabel locali 8308 5797 8342 5831 0 FreeSans 250 0 0 0 _40_.X
flabel locali 8308 5865 8342 5899 0 FreeSans 250 0 0 0 _40_.X
flabel nwell 8264 5967 8298 6001 0 FreeSans 250 0 0 0 _40_.VPB
flabel pwell 8254 5423 8288 5457 0 FreeSans 250 0 0 0 _40_.VNB
rlabel comment 8372 5440 8372 5440 6 _40_.mux2_1
flabel locali 8217 6273 8251 6307 0 FreeSans 200 0 0 0 _41_.A
flabel locali 8401 6137 8435 6171 0 FreeSans 200 0 0 0 _41_.X
flabel locali 8033 6273 8067 6307 0 FreeSans 200 0 0 0 _41_.B
flabel nwell 8033 5967 8067 6001 0 FreeSans 200 0 0 0 _41_.VPB
flabel pwell 8033 6511 8067 6545 0 FreeSans 200 0 0 0 _41_.VNB
flabel metal1 8033 6511 8067 6545 0 FreeSans 200 0 0 0 _41_.VGND
flabel metal1 8033 5967 8067 6001 0 FreeSans 200 0 0 0 _41_.VPWR
rlabel comment 8004 6528 8004 6528 2 _41_.or2_1
flabel metal1 11161 5423 11195 5457 0 FreeSans 200 0 0 0 FILLER_6_109.VGND
flabel metal1 11161 5967 11195 6001 0 FreeSans 200 0 0 0 FILLER_6_109.VPWR
flabel nwell 11161 5967 11195 6001 0 FreeSans 200 0 0 0 FILLER_6_109.VPB
flabel pwell 11161 5423 11195 5457 0 FreeSans 200 0 0 0 FILLER_6_109.VNB
rlabel comment 11132 5440 11132 5440 4 FILLER_6_109.decap_4
flabel metal1 10057 5423 10091 5457 0 FreeSans 200 0 0 0 FILLER_6_97.VGND
flabel metal1 10057 5967 10091 6001 0 FreeSans 200 0 0 0 FILLER_6_97.VPWR
flabel nwell 10057 5967 10091 6001 0 FreeSans 200 0 0 0 FILLER_6_97.VPB
flabel pwell 10057 5423 10091 5457 0 FreeSans 200 0 0 0 FILLER_6_97.VNB
rlabel comment 10028 5440 10028 5440 4 FILLER_6_97.decap_12
flabel metal1 10701 5967 10735 6001 0 FreeSans 200 0 0 0 FILLER_7_104.VPWR
flabel metal1 10701 6511 10735 6545 0 FreeSans 200 0 0 0 FILLER_7_104.VGND
flabel nwell 10701 5967 10735 6001 0 FreeSans 200 0 0 0 FILLER_7_104.VPB
flabel pwell 10701 6511 10735 6545 0 FreeSans 200 0 0 0 FILLER_7_104.VNB
rlabel comment 10672 6528 10672 6528 2 FILLER_7_104.decap_8
flabel metal1 9597 6511 9631 6545 0 FreeSans 200 0 0 0 FILLER_7_92.VGND
flabel metal1 9597 5967 9631 6001 0 FreeSans 200 0 0 0 FILLER_7_92.VPWR
flabel nwell 9597 5967 9631 6001 0 FreeSans 200 0 0 0 FILLER_7_92.VPB
flabel pwell 9597 6511 9631 6545 0 FreeSans 200 0 0 0 FILLER_7_92.VNB
rlabel comment 9568 6528 9568 6528 2 FILLER_7_92.decap_12
flabel metal1 11989 5967 12023 6001 0 FreeSans 200 0 0 0 FILLER_6_118.VPWR
flabel metal1 11989 5423 12023 5457 0 FreeSans 200 0 0 0 FILLER_6_118.VGND
flabel nwell 11989 5967 12023 6001 0 FreeSans 200 0 0 0 FILLER_6_118.VPB
flabel pwell 11989 5423 12023 5457 0 FreeSans 200 0 0 0 FILLER_6_118.VNB
rlabel comment 11960 5440 11960 5440 4 FILLER_6_118.decap_8
flabel metal1 12718 5967 12754 5997 0 FreeSans 250 0 0 0 FILLER_6_126.VPWR
flabel metal1 12718 5427 12754 5456 0 FreeSans 250 0 0 0 FILLER_6_126.VGND
flabel nwell 12727 5974 12747 5991 0 FreeSans 200 0 0 0 FILLER_6_126.VPB
flabel pwell 12724 5429 12748 5451 0 FreeSans 200 0 0 0 FILLER_6_126.VNB
rlabel comment 12696 5440 12696 5440 4 FILLER_6_126.fill_1
flabel metal1 11529 6511 11563 6545 0 FreeSans 200 0 0 0 FILLER_7_113.VGND
flabel metal1 11529 5967 11563 6001 0 FreeSans 200 0 0 0 FILLER_7_113.VPWR
flabel nwell 11529 5967 11563 6001 0 FreeSans 200 0 0 0 FILLER_7_113.VPB
flabel pwell 11529 6511 11563 6545 0 FreeSans 200 0 0 0 FILLER_7_113.VNB
rlabel comment 11500 6528 11500 6528 2 FILLER_7_113.decap_12
flabel metal1 12633 6511 12667 6545 0 FreeSans 200 0 0 0 FILLER_7_125.VGND
flabel metal1 12633 5967 12667 6001 0 FreeSans 200 0 0 0 FILLER_7_125.VPWR
flabel nwell 12633 5967 12667 6001 0 FreeSans 200 0 0 0 FILLER_7_125.VPB
flabel pwell 12633 6511 12667 6545 0 FreeSans 200 0 0 0 FILLER_7_125.VNB
rlabel comment 12604 6528 12604 6528 2 FILLER_7_125.decap_12
flabel metal1 11430 5975 11483 6004 0 FreeSans 200 0 0 0 TAP_45.VPWR
flabel metal1 11429 6508 11480 6546 0 FreeSans 200 0 0 0 TAP_45.VGND
rlabel comment 11408 6528 11408 6528 2 TAP_45.tapvpwrvgnd_1
flabel locali 13001 5661 13035 5695 0 FreeSans 200 0 0 0 _32_.A
flabel locali 13185 5797 13219 5831 0 FreeSans 200 0 0 0 _32_.X
flabel locali 12817 5661 12851 5695 0 FreeSans 200 0 0 0 _32_.B
flabel nwell 12817 5967 12851 6001 0 FreeSans 200 0 0 0 _32_.VPB
flabel pwell 12817 5423 12851 5457 0 FreeSans 200 0 0 0 _32_.VNB
flabel metal1 12817 5423 12851 5457 0 FreeSans 200 0 0 0 _32_.VGND
flabel metal1 12817 5967 12851 6001 0 FreeSans 200 0 0 0 _32_.VPWR
rlabel comment 12788 5440 12788 5440 4 _32_.or2_1
flabel locali 11713 5661 11747 5695 0 FreeSans 200 0 0 0 _35_.A
flabel locali 11897 5797 11931 5831 0 FreeSans 200 0 0 0 _35_.X
flabel locali 11529 5661 11563 5695 0 FreeSans 200 0 0 0 _35_.B
flabel nwell 11529 5967 11563 6001 0 FreeSans 200 0 0 0 _35_.VPB
flabel pwell 11529 5423 11563 5457 0 FreeSans 200 0 0 0 _35_.VNB
flabel metal1 11529 5423 11563 5457 0 FreeSans 200 0 0 0 _35_.VGND
flabel metal1 11529 5967 11563 6001 0 FreeSans 200 0 0 0 _35_.VPWR
rlabel comment 11500 5440 11500 5440 4 _35_.or2_1
flabel metal1 13277 5967 13311 6001 0 FreeSans 200 0 0 0 FILLER_6_132.VPWR
flabel metal1 13277 5423 13311 5457 0 FreeSans 200 0 0 0 FILLER_6_132.VGND
flabel nwell 13277 5967 13311 6001 0 FreeSans 200 0 0 0 FILLER_6_132.VPB
flabel pwell 13277 5423 13311 5457 0 FreeSans 200 0 0 0 FILLER_6_132.VNB
rlabel comment 13248 5440 13248 5440 4 FILLER_6_132.decap_8
flabel metal1 14105 5423 14139 5457 0 FreeSans 200 0 0 0 FILLER_6_141.VGND
flabel metal1 14105 5967 14139 6001 0 FreeSans 200 0 0 0 FILLER_6_141.VPWR
flabel nwell 14105 5967 14139 6001 0 FreeSans 200 0 0 0 FILLER_6_141.VPB
flabel pwell 14105 5423 14139 5457 0 FreeSans 200 0 0 0 FILLER_6_141.VNB
rlabel comment 14076 5440 14076 5440 4 FILLER_6_141.decap_12
flabel metal1 13737 6511 13771 6545 0 FreeSans 200 0 0 0 FILLER_7_137.VGND
flabel metal1 13737 5967 13771 6001 0 FreeSans 200 0 0 0 FILLER_7_137.VPWR
flabel nwell 13737 5967 13771 6001 0 FreeSans 200 0 0 0 FILLER_7_137.VPB
flabel pwell 13737 6511 13771 6545 0 FreeSans 200 0 0 0 FILLER_7_137.VNB
rlabel comment 13708 6528 13708 6528 2 FILLER_7_137.decap_12
flabel metal1 14841 6511 14875 6545 0 FreeSans 200 0 0 0 FILLER_7_149.VGND
flabel metal1 14841 5967 14875 6001 0 FreeSans 200 0 0 0 FILLER_7_149.VPWR
flabel nwell 14841 5967 14875 6001 0 FreeSans 200 0 0 0 FILLER_7_149.VPB
flabel pwell 14841 6511 14875 6545 0 FreeSans 200 0 0 0 FILLER_7_149.VNB
rlabel comment 14812 6528 14812 6528 2 FILLER_7_149.decap_12
flabel metal1 14006 5964 14059 5993 0 FreeSans 200 0 0 0 TAP_43.VPWR
flabel metal1 14005 5422 14056 5460 0 FreeSans 200 0 0 0 TAP_43.VGND
rlabel comment 13984 5440 13984 5440 4 TAP_43.tapvpwrvgnd_1
flabel metal1 15209 5423 15243 5457 0 FreeSans 200 0 0 0 FILLER_6_153.VGND
flabel metal1 15209 5967 15243 6001 0 FreeSans 200 0 0 0 FILLER_6_153.VPWR
flabel nwell 15209 5967 15243 6001 0 FreeSans 200 0 0 0 FILLER_6_153.VPB
flabel pwell 15209 5423 15243 5457 0 FreeSans 200 0 0 0 FILLER_6_153.VNB
rlabel comment 15180 5440 15180 5440 4 FILLER_6_153.decap_12
flabel metal1 16313 5423 16347 5457 0 FreeSans 200 0 0 0 FILLER_6_165.VGND
flabel metal1 16313 5967 16347 6001 0 FreeSans 200 0 0 0 FILLER_6_165.VPWR
flabel nwell 16313 5967 16347 6001 0 FreeSans 200 0 0 0 FILLER_6_165.VPB
flabel pwell 16313 5423 16347 5457 0 FreeSans 200 0 0 0 FILLER_6_165.VNB
rlabel comment 16284 5440 16284 5440 4 FILLER_6_165.decap_12
flabel metal1 15945 5967 15979 6001 0 FreeSans 200 0 0 0 FILLER_7_161.VPWR
flabel metal1 15945 6511 15979 6545 0 FreeSans 200 0 0 0 FILLER_7_161.VGND
flabel nwell 15945 5967 15979 6001 0 FreeSans 200 0 0 0 FILLER_7_161.VPB
flabel pwell 15945 6511 15979 6545 0 FreeSans 200 0 0 0 FILLER_7_161.VNB
rlabel comment 15916 6528 15916 6528 2 FILLER_7_161.decap_6
flabel metal1 16490 5971 16526 6001 0 FreeSans 250 0 0 0 FILLER_7_167.VPWR
flabel metal1 16490 6512 16526 6541 0 FreeSans 250 0 0 0 FILLER_7_167.VGND
flabel nwell 16499 5977 16519 5994 0 FreeSans 200 0 0 0 FILLER_7_167.VPB
flabel pwell 16496 6517 16520 6539 0 FreeSans 200 0 0 0 FILLER_7_167.VNB
rlabel comment 16468 6528 16468 6528 2 FILLER_7_167.fill_1
flabel metal1 16681 6511 16715 6545 0 FreeSans 200 0 0 0 FILLER_7_169.VGND
flabel metal1 16681 5967 16715 6001 0 FreeSans 200 0 0 0 FILLER_7_169.VPWR
flabel nwell 16681 5967 16715 6001 0 FreeSans 200 0 0 0 FILLER_7_169.VPB
flabel pwell 16681 6511 16715 6545 0 FreeSans 200 0 0 0 FILLER_7_169.VNB
rlabel comment 16652 6528 16652 6528 2 FILLER_7_169.decap_12
flabel metal1 16582 5975 16635 6004 0 FreeSans 200 0 0 0 TAP_46.VPWR
flabel metal1 16581 6508 16632 6546 0 FreeSans 200 0 0 0 TAP_46.VGND
rlabel comment 16560 6528 16560 6528 2 TAP_46.tapvpwrvgnd_1
flabel metal1 17417 5423 17451 5457 0 FreeSans 200 0 0 0 FILLER_6_177.VGND
flabel metal1 17417 5967 17451 6001 0 FreeSans 200 0 0 0 FILLER_6_177.VPWR
flabel nwell 17417 5967 17451 6001 0 FreeSans 200 0 0 0 FILLER_6_177.VPB
flabel pwell 17417 5423 17451 5457 0 FreeSans 200 0 0 0 FILLER_6_177.VNB
rlabel comment 17388 5440 17388 5440 4 FILLER_6_177.decap_12
flabel metal1 18514 5967 18550 5997 0 FreeSans 250 0 0 0 FILLER_6_189.VPWR
flabel metal1 18514 5427 18550 5456 0 FreeSans 250 0 0 0 FILLER_6_189.VGND
flabel nwell 18523 5974 18543 5991 0 FreeSans 200 0 0 0 FILLER_6_189.VPB
flabel pwell 18520 5429 18544 5451 0 FreeSans 200 0 0 0 FILLER_6_189.VNB
rlabel comment 18492 5440 18492 5440 4 FILLER_6_189.fill_1
flabel metal1 17785 5967 17819 6001 0 FreeSans 200 0 0 0 FILLER_7_181.VPWR
flabel metal1 17785 6511 17819 6545 0 FreeSans 200 0 0 0 FILLER_7_181.VGND
flabel nwell 17785 5967 17819 6001 0 FreeSans 200 0 0 0 FILLER_7_181.VPB
flabel pwell 17785 6511 17819 6545 0 FreeSans 200 0 0 0 FILLER_7_181.VNB
rlabel comment 17756 6528 17756 6528 2 FILLER_7_181.decap_8
flabel metal1 18514 5971 18550 6001 0 FreeSans 250 0 0 0 FILLER_7_189.VPWR
flabel metal1 18514 6512 18550 6541 0 FreeSans 250 0 0 0 FILLER_7_189.VGND
flabel nwell 18523 5977 18543 5994 0 FreeSans 200 0 0 0 FILLER_7_189.VPB
flabel pwell 18520 6517 18544 6539 0 FreeSans 200 0 0 0 FILLER_7_189.VNB
rlabel comment 18492 6528 18492 6528 2 FILLER_7_189.fill_1
flabel metal1 18797 5967 18831 6001 0 FreeSans 200 0 0 0 PHY_13.VPWR
flabel metal1 18797 5423 18831 5457 0 FreeSans 200 0 0 0 PHY_13.VGND
flabel nwell 18797 5967 18831 6001 0 FreeSans 200 0 0 0 PHY_13.VPB
flabel pwell 18797 5423 18831 5457 0 FreeSans 200 0 0 0 PHY_13.VNB
rlabel comment 18860 5440 18860 5440 6 PHY_13.decap_3
flabel metal1 18797 5967 18831 6001 0 FreeSans 200 0 0 0 PHY_15.VPWR
flabel metal1 18797 6511 18831 6545 0 FreeSans 200 0 0 0 PHY_15.VGND
flabel nwell 18797 5967 18831 6001 0 FreeSans 200 0 0 0 PHY_15.VPB
flabel pwell 18797 6511 18831 6545 0 FreeSans 200 0 0 0 PHY_15.VNB
rlabel comment 18860 6528 18860 6528 8 PHY_15.decap_3
flabel metal1 2513 6511 2547 6545 0 FreeSans 200 0 0 0 FILLER_8_15.VGND
flabel metal1 2513 7055 2547 7089 0 FreeSans 200 0 0 0 FILLER_8_15.VPWR
flabel nwell 2513 7055 2547 7089 0 FreeSans 200 0 0 0 FILLER_8_15.VPB
flabel pwell 2513 6511 2547 6545 0 FreeSans 200 0 0 0 FILLER_8_15.VNB
rlabel comment 2484 6528 2484 6528 4 FILLER_8_15.decap_12
flabel metal1 1409 6511 1443 6545 0 FreeSans 200 0 0 0 FILLER_8_3.VGND
flabel metal1 1409 7055 1443 7089 0 FreeSans 200 0 0 0 FILLER_8_3.VPWR
flabel nwell 1409 7055 1443 7089 0 FreeSans 200 0 0 0 FILLER_8_3.VPB
flabel pwell 1409 6511 1443 6545 0 FreeSans 200 0 0 0 FILLER_8_3.VNB
rlabel comment 1380 6528 1380 6528 4 FILLER_8_3.decap_12
flabel metal1 1133 7055 1167 7089 0 FreeSans 200 0 0 0 PHY_16.VPWR
flabel metal1 1133 6511 1167 6545 0 FreeSans 200 0 0 0 PHY_16.VGND
flabel nwell 1133 7055 1167 7089 0 FreeSans 200 0 0 0 PHY_16.VPB
flabel pwell 1133 6511 1167 6545 0 FreeSans 200 0 0 0 PHY_16.VNB
rlabel comment 1104 6528 1104 6528 4 PHY_16.decap_3
flabel metal1 3610 7055 3646 7085 0 FreeSans 250 0 0 0 FILLER_8_27.VPWR
flabel metal1 3610 6515 3646 6544 0 FreeSans 250 0 0 0 FILLER_8_27.VGND
flabel nwell 3619 7062 3639 7079 0 FreeSans 200 0 0 0 FILLER_8_27.VPB
flabel pwell 3616 6517 3640 6539 0 FreeSans 200 0 0 0 FILLER_8_27.VNB
rlabel comment 3588 6528 3588 6528 4 FILLER_8_27.fill_1
flabel metal1 3801 6511 3835 6545 0 FreeSans 200 0 0 0 FILLER_8_29.VGND
flabel metal1 3801 7055 3835 7089 0 FreeSans 200 0 0 0 FILLER_8_29.VPWR
flabel nwell 3801 7055 3835 7089 0 FreeSans 200 0 0 0 FILLER_8_29.VPB
flabel pwell 3801 6511 3835 6545 0 FreeSans 200 0 0 0 FILLER_8_29.VNB
rlabel comment 3772 6528 3772 6528 4 FILLER_8_29.decap_12
flabel metal1 4905 6511 4939 6545 0 FreeSans 200 0 0 0 FILLER_8_41.VGND
flabel metal1 4905 7055 4939 7089 0 FreeSans 200 0 0 0 FILLER_8_41.VPWR
flabel nwell 4905 7055 4939 7089 0 FreeSans 200 0 0 0 FILLER_8_41.VPB
flabel pwell 4905 6511 4939 6545 0 FreeSans 200 0 0 0 FILLER_8_41.VNB
rlabel comment 4876 6528 4876 6528 4 FILLER_8_41.decap_12
flabel metal1 3702 7052 3755 7081 0 FreeSans 200 0 0 0 TAP_47.VPWR
flabel metal1 3701 6510 3752 6548 0 FreeSans 200 0 0 0 TAP_47.VGND
rlabel comment 3680 6528 3680 6528 4 TAP_47.tapvpwrvgnd_1
flabel metal1 6009 6511 6043 6545 0 FreeSans 200 0 0 0 FILLER_8_53.VGND
flabel metal1 6009 7055 6043 7089 0 FreeSans 200 0 0 0 FILLER_8_53.VPWR
flabel nwell 6009 7055 6043 7089 0 FreeSans 200 0 0 0 FILLER_8_53.VPB
flabel pwell 6009 6511 6043 6545 0 FreeSans 200 0 0 0 FILLER_8_53.VNB
rlabel comment 5980 6528 5980 6528 4 FILLER_8_53.decap_12
flabel metal1 7113 6511 7147 6545 0 FreeSans 200 0 0 0 FILLER_8_65.VGND
flabel metal1 7113 7055 7147 7089 0 FreeSans 200 0 0 0 FILLER_8_65.VPWR
flabel nwell 7113 7055 7147 7089 0 FreeSans 200 0 0 0 FILLER_8_65.VPB
flabel pwell 7113 6511 7147 6545 0 FreeSans 200 0 0 0 FILLER_8_65.VNB
rlabel comment 7084 6528 7084 6528 4 FILLER_8_65.decap_12
flabel metal1 8217 7055 8251 7089 0 FreeSans 200 0 0 0 FILLER_8_77.VPWR
flabel metal1 8217 6511 8251 6545 0 FreeSans 200 0 0 0 FILLER_8_77.VGND
flabel nwell 8217 7055 8251 7089 0 FreeSans 200 0 0 0 FILLER_8_77.VPB
flabel pwell 8217 6511 8251 6545 0 FreeSans 200 0 0 0 FILLER_8_77.VNB
rlabel comment 8188 6528 8188 6528 4 FILLER_8_77.decap_6
flabel metal1 8762 7055 8798 7085 0 FreeSans 250 0 0 0 FILLER_8_83.VPWR
flabel metal1 8762 6515 8798 6544 0 FreeSans 250 0 0 0 FILLER_8_83.VGND
flabel nwell 8771 7062 8791 7079 0 FreeSans 200 0 0 0 FILLER_8_83.VPB
flabel pwell 8768 6517 8792 6539 0 FreeSans 200 0 0 0 FILLER_8_83.VNB
rlabel comment 8740 6528 8740 6528 4 FILLER_8_83.fill_1
flabel metal1 8953 6511 8987 6545 0 FreeSans 200 0 0 0 FILLER_8_85.VGND
flabel metal1 8953 7055 8987 7089 0 FreeSans 200 0 0 0 FILLER_8_85.VPWR
flabel nwell 8953 7055 8987 7089 0 FreeSans 200 0 0 0 FILLER_8_85.VPB
flabel pwell 8953 6511 8987 6545 0 FreeSans 200 0 0 0 FILLER_8_85.VNB
rlabel comment 8924 6528 8924 6528 4 FILLER_8_85.decap_12
flabel metal1 8854 7052 8907 7081 0 FreeSans 200 0 0 0 TAP_48.VPWR
flabel metal1 8853 6510 8904 6548 0 FreeSans 200 0 0 0 TAP_48.VGND
rlabel comment 8832 6528 8832 6528 4 TAP_48.tapvpwrvgnd_1
flabel metal1 11161 6511 11195 6545 0 FreeSans 200 0 0 0 FILLER_8_109.VGND
flabel metal1 11161 7055 11195 7089 0 FreeSans 200 0 0 0 FILLER_8_109.VPWR
flabel nwell 11161 7055 11195 7089 0 FreeSans 200 0 0 0 FILLER_8_109.VPB
flabel pwell 11161 6511 11195 6545 0 FreeSans 200 0 0 0 FILLER_8_109.VNB
rlabel comment 11132 6528 11132 6528 4 FILLER_8_109.decap_12
flabel metal1 10057 6511 10091 6545 0 FreeSans 200 0 0 0 FILLER_8_97.VGND
flabel metal1 10057 7055 10091 7089 0 FreeSans 200 0 0 0 FILLER_8_97.VPWR
flabel nwell 10057 7055 10091 7089 0 FreeSans 200 0 0 0 FILLER_8_97.VPB
flabel pwell 10057 6511 10091 6545 0 FreeSans 200 0 0 0 FILLER_8_97.VNB
rlabel comment 10028 6528 10028 6528 4 FILLER_8_97.decap_12
flabel metal1 12265 6511 12299 6545 0 FreeSans 200 0 0 0 FILLER_8_121.VGND
flabel metal1 12265 7055 12299 7089 0 FreeSans 200 0 0 0 FILLER_8_121.VPWR
flabel nwell 12265 7055 12299 7089 0 FreeSans 200 0 0 0 FILLER_8_121.VPB
flabel pwell 12265 6511 12299 6545 0 FreeSans 200 0 0 0 FILLER_8_121.VNB
rlabel comment 12236 6528 12236 6528 4 FILLER_8_121.decap_12
flabel metal1 13369 7055 13403 7089 0 FreeSans 200 0 0 0 FILLER_8_133.VPWR
flabel metal1 13369 6511 13403 6545 0 FreeSans 200 0 0 0 FILLER_8_133.VGND
flabel nwell 13369 7055 13403 7089 0 FreeSans 200 0 0 0 FILLER_8_133.VPB
flabel pwell 13369 6511 13403 6545 0 FreeSans 200 0 0 0 FILLER_8_133.VNB
rlabel comment 13340 6528 13340 6528 4 FILLER_8_133.decap_6
flabel metal1 13914 7055 13950 7085 0 FreeSans 250 0 0 0 FILLER_8_139.VPWR
flabel metal1 13914 6515 13950 6544 0 FreeSans 250 0 0 0 FILLER_8_139.VGND
flabel nwell 13923 7062 13943 7079 0 FreeSans 200 0 0 0 FILLER_8_139.VPB
flabel pwell 13920 6517 13944 6539 0 FreeSans 200 0 0 0 FILLER_8_139.VNB
rlabel comment 13892 6528 13892 6528 4 FILLER_8_139.fill_1
flabel metal1 14105 6511 14139 6545 0 FreeSans 200 0 0 0 FILLER_8_141.VGND
flabel metal1 14105 7055 14139 7089 0 FreeSans 200 0 0 0 FILLER_8_141.VPWR
flabel nwell 14105 7055 14139 7089 0 FreeSans 200 0 0 0 FILLER_8_141.VPB
flabel pwell 14105 6511 14139 6545 0 FreeSans 200 0 0 0 FILLER_8_141.VNB
rlabel comment 14076 6528 14076 6528 4 FILLER_8_141.decap_12
flabel metal1 14006 7052 14059 7081 0 FreeSans 200 0 0 0 TAP_49.VPWR
flabel metal1 14005 6510 14056 6548 0 FreeSans 200 0 0 0 TAP_49.VGND
rlabel comment 13984 6528 13984 6528 4 TAP_49.tapvpwrvgnd_1
flabel metal1 15209 6511 15243 6545 0 FreeSans 200 0 0 0 FILLER_8_153.VGND
flabel metal1 15209 7055 15243 7089 0 FreeSans 200 0 0 0 FILLER_8_153.VPWR
flabel nwell 15209 7055 15243 7089 0 FreeSans 200 0 0 0 FILLER_8_153.VPB
flabel pwell 15209 6511 15243 6545 0 FreeSans 200 0 0 0 FILLER_8_153.VNB
rlabel comment 15180 6528 15180 6528 4 FILLER_8_153.decap_12
flabel metal1 16313 6511 16347 6545 0 FreeSans 200 0 0 0 FILLER_8_165.VGND
flabel metal1 16313 7055 16347 7089 0 FreeSans 200 0 0 0 FILLER_8_165.VPWR
flabel nwell 16313 7055 16347 7089 0 FreeSans 200 0 0 0 FILLER_8_165.VPB
flabel pwell 16313 6511 16347 6545 0 FreeSans 200 0 0 0 FILLER_8_165.VNB
rlabel comment 16284 6528 16284 6528 4 FILLER_8_165.decap_12
flabel metal1 17417 6511 17451 6545 0 FreeSans 200 0 0 0 FILLER_8_177.VGND
flabel metal1 17417 7055 17451 7089 0 FreeSans 200 0 0 0 FILLER_8_177.VPWR
flabel nwell 17417 7055 17451 7089 0 FreeSans 200 0 0 0 FILLER_8_177.VPB
flabel pwell 17417 6511 17451 6545 0 FreeSans 200 0 0 0 FILLER_8_177.VNB
rlabel comment 17388 6528 17388 6528 4 FILLER_8_177.decap_12
flabel metal1 18514 7055 18550 7085 0 FreeSans 250 0 0 0 FILLER_8_189.VPWR
flabel metal1 18514 6515 18550 6544 0 FreeSans 250 0 0 0 FILLER_8_189.VGND
flabel nwell 18523 7062 18543 7079 0 FreeSans 200 0 0 0 FILLER_8_189.VPB
flabel pwell 18520 6517 18544 6539 0 FreeSans 200 0 0 0 FILLER_8_189.VNB
rlabel comment 18492 6528 18492 6528 4 FILLER_8_189.fill_1
flabel metal1 18797 7055 18831 7089 0 FreeSans 200 0 0 0 PHY_17.VPWR
flabel metal1 18797 6511 18831 6545 0 FreeSans 200 0 0 0 PHY_17.VGND
flabel nwell 18797 7055 18831 7089 0 FreeSans 200 0 0 0 PHY_17.VPB
flabel pwell 18797 6511 18831 6545 0 FreeSans 200 0 0 0 PHY_17.VNB
rlabel comment 18860 6528 18860 6528 6 PHY_17.decap_3
flabel metal1 3065 7055 3099 7089 0 FreeSans 200 0 0 0 FILLER_9_21.VPWR
flabel metal1 3065 7599 3099 7633 0 FreeSans 200 0 0 0 FILLER_9_21.VGND
flabel nwell 3065 7055 3099 7089 0 FreeSans 200 0 0 0 FILLER_9_21.VPB
flabel pwell 3065 7599 3099 7633 0 FreeSans 200 0 0 0 FILLER_9_21.VNB
rlabel comment 3036 7616 3036 7616 2 FILLER_9_21.decap_6
flabel metal1 1400 7598 1453 7630 0 FreeSans 200 0 0 0 FILLER_9_3.VGND
flabel metal1 1401 7055 1453 7086 0 FreeSans 200 0 0 0 FILLER_9_3.VPWR
flabel nwell 1408 7063 1442 7081 0 FreeSans 200 0 0 0 FILLER_9_3.VPB
flabel pwell 1411 7604 1443 7626 0 FreeSans 200 0 0 0 FILLER_9_3.VNB
rlabel comment 1380 7616 1380 7616 2 FILLER_9_3.fill_2
flabel metal1 1961 7599 1995 7633 0 FreeSans 200 0 0 0 FILLER_9_9.VGND
flabel metal1 1961 7055 1995 7089 0 FreeSans 200 0 0 0 FILLER_9_9.VPWR
flabel nwell 1961 7055 1995 7089 0 FreeSans 200 0 0 0 FILLER_9_9.VPB
flabel pwell 1961 7599 1995 7633 0 FreeSans 200 0 0 0 FILLER_9_9.VNB
rlabel comment 1932 7616 1932 7616 2 FILLER_9_9.decap_12
flabel metal1 1133 7055 1167 7089 0 FreeSans 200 0 0 0 PHY_18.VPWR
flabel metal1 1133 7599 1167 7633 0 FreeSans 200 0 0 0 PHY_18.VGND
flabel nwell 1133 7055 1167 7089 0 FreeSans 200 0 0 0 PHY_18.VPB
flabel pwell 1133 7599 1167 7633 0 FreeSans 200 0 0 0 PHY_18.VNB
rlabel comment 1104 7616 1104 7616 2 PHY_18.decap_3
flabel metal1 1869 7055 1903 7089 0 FreeSans 200 0 0 0 output3.VPWR
flabel metal1 1869 7599 1903 7633 0 FreeSans 200 0 0 0 output3.VGND
flabel locali 1869 7055 1903 7089 0 FreeSans 200 0 0 0 output3.VPWR
flabel locali 1869 7599 1903 7633 0 FreeSans 200 0 0 0 output3.VGND
flabel locali 1686 7497 1720 7531 0 FreeSans 200 0 0 0 output3.X
flabel locali 1686 7225 1720 7259 0 FreeSans 200 0 0 0 output3.X
flabel locali 1686 7157 1720 7191 0 FreeSans 200 0 0 0 output3.X
flabel locali 1869 7361 1903 7395 0 FreeSans 200 0 0 0 output3.A
flabel nwell 1869 7055 1903 7089 0 FreeSans 200 0 0 0 output3.VPB
flabel pwell 1869 7599 1903 7633 0 FreeSans 200 0 0 0 output3.VNB
rlabel comment 1932 7616 1932 7616 8 output3.buf_2
flabel metal1 3610 7059 3646 7089 0 FreeSans 250 0 0 0 FILLER_9_27.VPWR
flabel metal1 3610 7600 3646 7629 0 FreeSans 250 0 0 0 FILLER_9_27.VGND
flabel nwell 3619 7065 3639 7082 0 FreeSans 200 0 0 0 FILLER_9_27.VPB
flabel pwell 3616 7605 3640 7627 0 FreeSans 200 0 0 0 FILLER_9_27.VNB
rlabel comment 3588 7616 3588 7616 2 FILLER_9_27.fill_1
flabel metal1 3792 7598 3845 7630 0 FreeSans 200 0 0 0 FILLER_9_29.VGND
flabel metal1 3793 7055 3845 7086 0 FreeSans 200 0 0 0 FILLER_9_29.VPWR
flabel nwell 3800 7063 3834 7081 0 FreeSans 200 0 0 0 FILLER_9_29.VPB
flabel pwell 3803 7604 3835 7626 0 FreeSans 200 0 0 0 FILLER_9_29.VNB
rlabel comment 3772 7616 3772 7616 2 FILLER_9_29.fill_2
flabel metal1 4353 7599 4387 7633 0 FreeSans 200 0 0 0 FILLER_9_35.VGND
flabel metal1 4353 7055 4387 7089 0 FreeSans 200 0 0 0 FILLER_9_35.VPWR
flabel nwell 4353 7055 4387 7089 0 FreeSans 200 0 0 0 FILLER_9_35.VPB
flabel pwell 4353 7599 4387 7633 0 FreeSans 200 0 0 0 FILLER_9_35.VNB
rlabel comment 4324 7616 4324 7616 2 FILLER_9_35.decap_12
flabel metal1 3702 7063 3755 7092 0 FreeSans 200 0 0 0 TAP_50.VPWR
flabel metal1 3701 7596 3752 7634 0 FreeSans 200 0 0 0 TAP_50.VGND
rlabel comment 3680 7616 3680 7616 2 TAP_50.tapvpwrvgnd_1
flabel metal1 4261 7055 4295 7089 0 FreeSans 200 0 0 0 output4.VPWR
flabel metal1 4261 7599 4295 7633 0 FreeSans 200 0 0 0 output4.VGND
flabel locali 4261 7055 4295 7089 0 FreeSans 200 0 0 0 output4.VPWR
flabel locali 4261 7599 4295 7633 0 FreeSans 200 0 0 0 output4.VGND
flabel locali 4078 7497 4112 7531 0 FreeSans 200 0 0 0 output4.X
flabel locali 4078 7225 4112 7259 0 FreeSans 200 0 0 0 output4.X
flabel locali 4078 7157 4112 7191 0 FreeSans 200 0 0 0 output4.X
flabel locali 4261 7361 4295 7395 0 FreeSans 200 0 0 0 output4.A
flabel nwell 4261 7055 4295 7089 0 FreeSans 200 0 0 0 output4.VPB
flabel pwell 4261 7599 4295 7633 0 FreeSans 200 0 0 0 output4.VNB
rlabel comment 4324 7616 4324 7616 8 output4.buf_2
flabel metal1 5448 7598 5501 7630 0 FreeSans 200 0 0 0 FILLER_9_47.VGND
flabel metal1 5449 7055 5501 7086 0 FreeSans 200 0 0 0 FILLER_9_47.VPWR
flabel nwell 5456 7063 5490 7081 0 FreeSans 200 0 0 0 FILLER_9_47.VPB
flabel pwell 5459 7604 5491 7626 0 FreeSans 200 0 0 0 FILLER_9_47.VNB
rlabel comment 5428 7616 5428 7616 2 FILLER_9_47.fill_2
flabel metal1 6009 7055 6043 7089 0 FreeSans 200 0 0 0 FILLER_9_53.VPWR
flabel metal1 6009 7599 6043 7633 0 FreeSans 200 0 0 0 FILLER_9_53.VGND
flabel nwell 6009 7055 6043 7089 0 FreeSans 200 0 0 0 FILLER_9_53.VPB
flabel pwell 6009 7599 6043 7633 0 FreeSans 200 0 0 0 FILLER_9_53.VNB
rlabel comment 5980 7616 5980 7616 2 FILLER_9_53.decap_3
flabel metal1 6377 7599 6411 7633 0 FreeSans 200 0 0 0 FILLER_9_57.VGND
flabel metal1 6377 7055 6411 7089 0 FreeSans 200 0 0 0 FILLER_9_57.VPWR
flabel nwell 6377 7055 6411 7089 0 FreeSans 200 0 0 0 FILLER_9_57.VPB
flabel pwell 6377 7599 6411 7633 0 FreeSans 200 0 0 0 FILLER_9_57.VNB
rlabel comment 6348 7616 6348 7616 2 FILLER_9_57.decap_12
flabel metal1 6278 7063 6331 7092 0 FreeSans 200 0 0 0 TAP_51.VPWR
flabel metal1 6277 7596 6328 7634 0 FreeSans 200 0 0 0 TAP_51.VGND
rlabel comment 6256 7616 6256 7616 2 TAP_51.tapvpwrvgnd_1
flabel metal1 5917 7055 5951 7089 0 FreeSans 200 0 0 0 output5.VPWR
flabel metal1 5917 7599 5951 7633 0 FreeSans 200 0 0 0 output5.VGND
flabel locali 5917 7055 5951 7089 0 FreeSans 200 0 0 0 output5.VPWR
flabel locali 5917 7599 5951 7633 0 FreeSans 200 0 0 0 output5.VGND
flabel locali 5734 7497 5768 7531 0 FreeSans 200 0 0 0 output5.X
flabel locali 5734 7225 5768 7259 0 FreeSans 200 0 0 0 output5.X
flabel locali 5734 7157 5768 7191 0 FreeSans 200 0 0 0 output5.X
flabel locali 5917 7361 5951 7395 0 FreeSans 200 0 0 0 output5.A
flabel nwell 5917 7055 5951 7089 0 FreeSans 200 0 0 0 output5.VPB
flabel pwell 5917 7599 5951 7633 0 FreeSans 200 0 0 0 output5.VNB
rlabel comment 5980 7616 5980 7616 8 output5.buf_2
flabel metal1 7481 7599 7515 7633 0 FreeSans 200 0 0 0 FILLER_9_69.VGND
flabel metal1 7481 7055 7515 7089 0 FreeSans 200 0 0 0 FILLER_9_69.VPWR
flabel nwell 7481 7055 7515 7089 0 FreeSans 200 0 0 0 FILLER_9_69.VPB
flabel pwell 7481 7599 7515 7633 0 FreeSans 200 0 0 0 FILLER_9_69.VNB
rlabel comment 7452 7616 7452 7616 2 FILLER_9_69.decap_4
flabel metal1 8217 7055 8251 7089 0 FreeSans 200 0 0 0 FILLER_9_77.VPWR
flabel metal1 8217 7599 8251 7633 0 FreeSans 200 0 0 0 FILLER_9_77.VGND
flabel nwell 8217 7055 8251 7089 0 FreeSans 200 0 0 0 FILLER_9_77.VPB
flabel pwell 8217 7599 8251 7633 0 FreeSans 200 0 0 0 FILLER_9_77.VNB
rlabel comment 8188 7616 8188 7616 2 FILLER_9_77.decap_6
flabel metal1 8762 7059 8798 7089 0 FreeSans 250 0 0 0 FILLER_9_83.VPWR
flabel metal1 8762 7600 8798 7629 0 FreeSans 250 0 0 0 FILLER_9_83.VGND
flabel nwell 8771 7065 8791 7082 0 FreeSans 200 0 0 0 FILLER_9_83.VPB
flabel pwell 8768 7605 8792 7627 0 FreeSans 200 0 0 0 FILLER_9_83.VNB
rlabel comment 8740 7616 8740 7616 2 FILLER_9_83.fill_1
flabel metal1 8953 7055 8987 7089 0 FreeSans 200 0 0 0 FILLER_9_85.VPWR
flabel metal1 8953 7599 8987 7633 0 FreeSans 200 0 0 0 FILLER_9_85.VGND
flabel nwell 8953 7055 8987 7089 0 FreeSans 200 0 0 0 FILLER_9_85.VPB
flabel pwell 8953 7599 8987 7633 0 FreeSans 200 0 0 0 FILLER_9_85.VNB
rlabel comment 8924 7616 8924 7616 2 FILLER_9_85.decap_6
flabel metal1 8854 7063 8907 7092 0 FreeSans 200 0 0 0 TAP_52.VPWR
flabel metal1 8853 7596 8904 7634 0 FreeSans 200 0 0 0 TAP_52.VGND
rlabel comment 8832 7616 8832 7616 2 TAP_52.tapvpwrvgnd_1
flabel metal1 8125 7055 8159 7089 0 FreeSans 200 0 0 0 output6.VPWR
flabel metal1 8125 7599 8159 7633 0 FreeSans 200 0 0 0 output6.VGND
flabel locali 8125 7055 8159 7089 0 FreeSans 200 0 0 0 output6.VPWR
flabel locali 8125 7599 8159 7633 0 FreeSans 200 0 0 0 output6.VGND
flabel locali 7942 7497 7976 7531 0 FreeSans 200 0 0 0 output6.X
flabel locali 7942 7225 7976 7259 0 FreeSans 200 0 0 0 output6.X
flabel locali 7942 7157 7976 7191 0 FreeSans 200 0 0 0 output6.X
flabel locali 8125 7361 8159 7395 0 FreeSans 200 0 0 0 output6.A
flabel nwell 8125 7055 8159 7089 0 FreeSans 200 0 0 0 output6.VPB
flabel pwell 8125 7599 8159 7633 0 FreeSans 200 0 0 0 output6.VNB
rlabel comment 8188 7616 8188 7616 8 output6.buf_2
flabel locali 9505 7497 9539 7531 0 FreeSans 200 0 0 0 ANTENNA_input1_A.DIODE
flabel locali 9505 7225 9539 7259 0 FreeSans 200 0 0 0 ANTENNA_input1_A.DIODE
flabel locali 9597 7225 9631 7259 0 FreeSans 200 0 0 0 ANTENNA_input1_A.DIODE
flabel locali 9505 7157 9539 7191 0 FreeSans 200 0 0 0 ANTENNA_input1_A.DIODE
flabel locali 9597 7157 9631 7191 0 FreeSans 200 0 0 0 ANTENNA_input1_A.DIODE
flabel locali 9597 7293 9631 7327 0 FreeSans 200 0 0 0 ANTENNA_input1_A.DIODE
flabel locali 9505 7293 9539 7327 0 FreeSans 200 0 0 0 ANTENNA_input1_A.DIODE
flabel locali 9597 7361 9631 7395 0 FreeSans 200 0 0 0 ANTENNA_input1_A.DIODE
flabel locali 9505 7361 9539 7395 0 FreeSans 200 0 0 0 ANTENNA_input1_A.DIODE
flabel locali 9505 7429 9539 7463 0 FreeSans 200 0 0 0 ANTENNA_input1_A.DIODE
flabel locali 9597 7429 9631 7463 0 FreeSans 200 0 0 0 ANTENNA_input1_A.DIODE
flabel locali 9597 7497 9631 7531 0 FreeSans 200 0 0 0 ANTENNA_input1_A.DIODE
flabel metal1 9597 7599 9631 7633 0 FreeSans 200 0 0 0 ANTENNA_input1_A.VGND
flabel metal1 9597 7055 9631 7089 0 FreeSans 200 0 0 0 ANTENNA_input1_A.VPWR
<< end >>
