magic
tech sky130A
magscale 1 2
timestamp 1671931150
<< pwell >>
rect -201 -4386 201 4386
<< psubdiff >>
rect -165 4316 -69 4350
rect 69 4316 165 4350
rect -165 4254 -131 4316
rect 131 4254 165 4316
rect -165 -4316 -131 -4254
rect 131 -4316 165 -4254
rect -165 -4350 -69 -4316
rect 69 -4350 165 -4316
<< psubdiffcont >>
rect -69 4316 69 4350
rect -165 -4254 -131 4254
rect 131 -4254 165 4254
rect -69 -4350 69 -4316
<< xpolycontact >>
rect -35 3788 35 4220
rect -35 3256 35 3688
rect -35 2720 35 3152
rect -35 2188 35 2620
rect -35 1652 35 2084
rect -35 1120 35 1552
rect -35 584 35 1016
rect -35 52 35 484
rect -35 -484 35 -52
rect -35 -1016 35 -584
rect -35 -1552 35 -1120
rect -35 -2084 35 -1652
rect -35 -2620 35 -2188
rect -35 -3152 35 -2720
rect -35 -3688 35 -3256
rect -35 -4220 35 -3788
<< xpolyres >>
rect -35 3688 35 3788
rect -35 2620 35 2720
rect -35 1552 35 1652
rect -35 484 35 584
rect -35 -584 35 -484
rect -35 -1652 35 -1552
rect -35 -2720 35 -2620
rect -35 -3788 35 -3688
<< locali >>
rect -165 4316 -69 4350
rect 69 4316 165 4350
rect -165 4254 -131 4316
rect 131 4254 165 4316
rect -165 -4316 -131 -4254
rect 131 -4316 165 -4254
rect -165 -4350 -69 -4316
rect 69 -4350 165 -4316
<< viali >>
rect -19 3805 19 4202
rect -19 3274 19 3671
rect -19 2737 19 3134
rect -19 2206 19 2603
rect -19 1669 19 2066
rect -19 1138 19 1535
rect -19 601 19 998
rect -19 70 19 467
rect -19 -467 19 -70
rect -19 -998 19 -601
rect -19 -1535 19 -1138
rect -19 -2066 19 -1669
rect -19 -2603 19 -2206
rect -19 -3134 19 -2737
rect -19 -3671 19 -3274
rect -19 -4202 19 -3805
<< metal1 >>
rect -25 4202 25 4214
rect -25 3805 -19 4202
rect 19 3805 25 4202
rect -25 3793 25 3805
rect -25 3671 25 3683
rect -25 3274 -19 3671
rect 19 3274 25 3671
rect -25 3262 25 3274
rect -25 3134 25 3146
rect -25 2737 -19 3134
rect 19 2737 25 3134
rect -25 2725 25 2737
rect -25 2603 25 2615
rect -25 2206 -19 2603
rect 19 2206 25 2603
rect -25 2194 25 2206
rect -25 2066 25 2078
rect -25 1669 -19 2066
rect 19 1669 25 2066
rect -25 1657 25 1669
rect -25 1535 25 1547
rect -25 1138 -19 1535
rect 19 1138 25 1535
rect -25 1126 25 1138
rect -25 998 25 1010
rect -25 601 -19 998
rect 19 601 25 998
rect -25 589 25 601
rect -25 467 25 479
rect -25 70 -19 467
rect 19 70 25 467
rect -25 58 25 70
rect -25 -70 25 -58
rect -25 -467 -19 -70
rect 19 -467 25 -70
rect -25 -479 25 -467
rect -25 -601 25 -589
rect -25 -998 -19 -601
rect 19 -998 25 -601
rect -25 -1010 25 -998
rect -25 -1138 25 -1126
rect -25 -1535 -19 -1138
rect 19 -1535 25 -1138
rect -25 -1547 25 -1535
rect -25 -1669 25 -1657
rect -25 -2066 -19 -1669
rect 19 -2066 25 -1669
rect -25 -2078 25 -2066
rect -25 -2206 25 -2194
rect -25 -2603 -19 -2206
rect 19 -2603 25 -2206
rect -25 -2615 25 -2603
rect -25 -2737 25 -2725
rect -25 -3134 -19 -2737
rect 19 -3134 25 -2737
rect -25 -3146 25 -3134
rect -25 -3274 25 -3262
rect -25 -3671 -19 -3274
rect 19 -3671 25 -3274
rect -25 -3683 25 -3671
rect -25 -3805 25 -3793
rect -25 -4202 -19 -3805
rect 19 -4202 25 -3805
rect -25 -4214 25 -4202
<< res0p35 >>
rect -37 3686 37 3790
rect -37 2618 37 2722
rect -37 1550 37 1654
rect -37 482 37 586
rect -37 -586 37 -482
rect -37 -1654 37 -1550
rect -37 -2722 37 -2618
rect -37 -3790 37 -3686
<< properties >>
string FIXED_BBOX -148 -4333 148 4333
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 0.50 m 8 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 3.932k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
