magic
tech sky130A
magscale 1 2
timestamp 1671401643
<< nwell >>
rect 716 3220 3972 5658
<< pwell >>
rect 148 3220 716 4488
rect -200 1800 3972 3220
<< nmos >>
rect -4 2010 396 3010
rect 454 2010 854 3010
rect 912 2010 1312 3010
rect 1370 2010 1770 3010
rect 1828 2010 2228 3010
rect 2286 2010 2686 3010
rect 2744 2010 3144 3010
rect 3430 2010 3460 3010
rect 3746 2010 3776 3010
<< pmos >>
rect 912 3439 1312 5439
rect 1370 3439 1770 5439
rect 1828 3439 2228 5439
rect 2286 3439 2686 5439
rect 2744 3439 3144 5439
rect 3430 3439 3460 5439
rect 3746 3439 3776 5439
<< ndiff >>
rect -62 2998 -4 3010
rect -62 2022 -50 2998
rect -16 2022 -4 2998
rect -62 2010 -4 2022
rect 396 2998 454 3010
rect 396 2022 408 2998
rect 442 2022 454 2998
rect 396 2010 454 2022
rect 854 2998 912 3010
rect 854 2022 866 2998
rect 900 2022 912 2998
rect 854 2010 912 2022
rect 1312 2998 1370 3010
rect 1312 2022 1324 2998
rect 1358 2022 1370 2998
rect 1312 2010 1370 2022
rect 1770 2998 1828 3010
rect 1770 2022 1782 2998
rect 1816 2022 1828 2998
rect 1770 2010 1828 2022
rect 2228 2998 2286 3010
rect 2228 2022 2240 2998
rect 2274 2022 2286 2998
rect 2228 2010 2286 2022
rect 2686 2998 2744 3010
rect 2686 2022 2698 2998
rect 2732 2022 2744 2998
rect 2686 2010 2744 2022
rect 3144 2998 3202 3010
rect 3144 2022 3156 2998
rect 3190 2022 3202 2998
rect 3144 2010 3202 2022
rect 3372 2998 3430 3010
rect 3372 2022 3384 2998
rect 3418 2022 3430 2998
rect 3372 2010 3430 2022
rect 3460 2998 3518 3010
rect 3460 2022 3472 2998
rect 3506 2022 3518 2998
rect 3460 2010 3518 2022
rect 3688 2998 3746 3010
rect 3688 2022 3700 2998
rect 3734 2022 3746 2998
rect 3688 2010 3746 2022
rect 3776 2998 3834 3010
rect 3776 2022 3788 2998
rect 3822 2022 3834 2998
rect 3776 2010 3834 2022
<< pdiff >>
rect 854 5427 912 5439
rect 854 3451 866 5427
rect 900 3451 912 5427
rect 854 3439 912 3451
rect 1312 5427 1370 5439
rect 1312 3451 1324 5427
rect 1358 3451 1370 5427
rect 1312 3439 1370 3451
rect 1770 5427 1828 5439
rect 1770 3451 1782 5427
rect 1816 3451 1828 5427
rect 1770 3439 1828 3451
rect 2228 5427 2286 5439
rect 2228 3451 2240 5427
rect 2274 3451 2286 5427
rect 2228 3439 2286 3451
rect 2686 5427 2744 5439
rect 2686 3451 2698 5427
rect 2732 3451 2744 5427
rect 2686 3439 2744 3451
rect 3144 5427 3202 5439
rect 3144 3451 3156 5427
rect 3190 3451 3202 5427
rect 3144 3439 3202 3451
rect 3372 5427 3430 5439
rect 3372 3451 3384 5427
rect 3418 3451 3430 5427
rect 3372 3439 3430 3451
rect 3460 5427 3518 5439
rect 3460 3451 3472 5427
rect 3506 3451 3518 5427
rect 3460 3439 3518 3451
rect 3688 5427 3746 5439
rect 3688 3451 3700 5427
rect 3734 3451 3746 5427
rect 3688 3439 3746 3451
rect 3776 5427 3834 5439
rect 3776 3451 3788 5427
rect 3822 3451 3834 5427
rect 3776 3439 3834 3451
<< ndiffc >>
rect -50 2022 -16 2998
rect 408 2022 442 2998
rect 866 2022 900 2998
rect 1324 2022 1358 2998
rect 1782 2022 1816 2998
rect 2240 2022 2274 2998
rect 2698 2022 2732 2998
rect 3156 2022 3190 2998
rect 3384 2022 3418 2998
rect 3472 2022 3506 2998
rect 3700 2022 3734 2998
rect 3788 2022 3822 2998
<< pdiffc >>
rect 866 3451 900 5427
rect 1324 3451 1358 5427
rect 1782 3451 1816 5427
rect 2240 3451 2274 5427
rect 2698 3451 2732 5427
rect 3156 3451 3190 5427
rect 3384 3451 3418 5427
rect 3472 3451 3506 5427
rect 3700 3451 3734 5427
rect 3788 3451 3822 5427
<< psubdiff >>
rect 184 4418 280 4452
rect 584 4418 680 4452
rect 184 4356 218 4418
rect 646 4356 680 4418
rect 184 3290 218 3352
rect 646 3290 680 3352
rect 184 3256 280 3290
rect 584 3256 680 3290
rect -164 3150 -68 3184
rect 3208 3150 3366 3184
rect 3524 3150 3682 3184
rect 3840 3150 3936 3184
rect -164 3088 -130 3150
rect 3270 3088 3304 3150
rect -164 1870 -130 1932
rect 3586 3088 3620 3150
rect 3270 1870 3304 1932
rect 3902 3088 3936 3150
rect 3586 1870 3620 1932
rect 3902 1870 3936 1932
rect -164 1836 -68 1870
rect 3208 1836 3366 1870
rect 3524 1836 3682 1870
rect 3840 1836 3936 1870
<< nsubdiff >>
rect 752 5588 848 5622
rect 3208 5588 3366 5622
rect 3524 5588 3682 5622
rect 3840 5588 3936 5622
rect 752 5526 786 5588
rect 3270 5526 3304 5588
rect 752 3290 786 3352
rect 3586 5526 3620 5588
rect 3270 3290 3304 3352
rect 3902 5526 3936 5588
rect 3586 3290 3620 3352
rect 3902 3290 3936 3352
rect 752 3256 848 3290
rect 3208 3256 3366 3290
rect 3524 3256 3682 3290
rect 3840 3256 3936 3290
<< psubdiffcont >>
rect 280 4418 584 4452
rect 184 3352 218 4356
rect 646 3352 680 4356
rect 280 3256 584 3290
rect -68 3150 3208 3184
rect 3366 3150 3524 3184
rect 3682 3150 3840 3184
rect -164 1932 -130 3088
rect 3270 1932 3304 3088
rect 3586 1932 3620 3088
rect 3902 1932 3936 3088
rect -68 1836 3208 1870
rect 3366 1836 3524 1870
rect 3682 1836 3840 1870
<< nsubdiffcont >>
rect 848 5588 3208 5622
rect 3366 5588 3524 5622
rect 3682 5588 3840 5622
rect 752 3352 786 5526
rect 3270 3352 3304 5526
rect 3586 3352 3620 5526
rect 3902 3352 3936 5526
rect 848 3256 3208 3290
rect 3366 3256 3524 3290
rect 3682 3256 3840 3290
<< poly >>
rect 912 5520 1312 5536
rect 912 5486 928 5520
rect 1296 5486 1312 5520
rect 912 5439 1312 5486
rect 1370 5520 1770 5536
rect 1370 5486 1386 5520
rect 1754 5486 1770 5520
rect 1370 5439 1770 5486
rect 1828 5520 2228 5536
rect 1828 5486 1844 5520
rect 2212 5486 2228 5520
rect 1828 5439 2228 5486
rect 2286 5520 2686 5536
rect 2286 5486 2302 5520
rect 2670 5486 2686 5520
rect 2286 5439 2686 5486
rect 2744 5520 3144 5536
rect 2744 5486 2760 5520
rect 3128 5486 3144 5520
rect 2744 5439 3144 5486
rect 912 3392 1312 3439
rect 912 3358 928 3392
rect 1296 3358 1312 3392
rect 912 3342 1312 3358
rect 1370 3392 1770 3439
rect 1370 3358 1386 3392
rect 1754 3358 1770 3392
rect 1370 3342 1770 3358
rect 1828 3392 2228 3439
rect 1828 3358 1844 3392
rect 2212 3358 2228 3392
rect 1828 3342 2228 3358
rect 2286 3392 2686 3439
rect 2286 3358 2302 3392
rect 2670 3358 2686 3392
rect 2286 3342 2686 3358
rect 2744 3392 3144 3439
rect 2744 3358 2760 3392
rect 3128 3358 3144 3392
rect 2744 3342 3144 3358
rect 3412 5470 3478 5536
rect 3430 5439 3460 5470
rect 3430 3408 3460 3439
rect 3412 3392 3478 3408
rect 3412 3358 3428 3392
rect 3462 3358 3478 3392
rect 3412 3342 3478 3358
rect 3728 5470 3794 5536
rect 3746 5439 3776 5470
rect 3746 3408 3776 3439
rect 3728 3392 3794 3408
rect 3728 3358 3744 3392
rect 3778 3358 3794 3392
rect 3728 3342 3794 3358
rect -4 3082 396 3098
rect -4 3048 12 3082
rect 380 3048 396 3082
rect -4 3010 396 3048
rect 454 3082 854 3098
rect 454 3048 470 3082
rect 838 3048 854 3082
rect 454 3010 854 3048
rect 912 3082 1312 3098
rect 912 3048 928 3082
rect 1296 3048 1312 3082
rect 912 3010 1312 3048
rect 1370 3082 1770 3098
rect 1370 3048 1386 3082
rect 1754 3048 1770 3082
rect 1370 3010 1770 3048
rect 1828 3082 2228 3098
rect 1828 3048 1844 3082
rect 2212 3048 2228 3082
rect 1828 3010 2228 3048
rect 2286 3082 2686 3098
rect 2286 3048 2302 3082
rect 2670 3048 2686 3082
rect 2286 3010 2686 3048
rect 2744 3082 3144 3098
rect 2744 3048 2760 3082
rect 3128 3048 3144 3082
rect 2744 3010 3144 3048
rect -4 1972 396 2010
rect -4 1938 12 1972
rect 380 1938 396 1972
rect -4 1922 396 1938
rect 454 1972 854 2010
rect 454 1938 470 1972
rect 838 1938 854 1972
rect 454 1922 854 1938
rect 912 1972 1312 2010
rect 912 1938 928 1972
rect 1296 1938 1312 1972
rect 912 1922 1312 1938
rect 1370 1972 1770 2010
rect 1370 1938 1386 1972
rect 1754 1938 1770 1972
rect 1370 1922 1770 1938
rect 1828 1972 2228 2010
rect 1828 1938 1844 1972
rect 2212 1938 2228 1972
rect 1828 1922 2228 1938
rect 2286 1972 2686 2010
rect 2286 1938 2302 1972
rect 2670 1938 2686 1972
rect 2286 1922 2686 1938
rect 2744 1972 3144 2010
rect 2744 1938 2760 1972
rect 3128 1938 3144 1972
rect 2744 1922 3144 1938
rect 3412 3082 3478 3098
rect 3412 3048 3428 3082
rect 3462 3048 3478 3082
rect 3412 3032 3478 3048
rect 3430 3010 3460 3032
rect 3430 1988 3460 2010
rect 3412 1922 3478 1988
rect 3728 3082 3794 3098
rect 3728 3048 3744 3082
rect 3778 3048 3794 3082
rect 3728 3032 3794 3048
rect 3746 3010 3776 3032
rect 3746 1988 3776 2010
rect 3728 1922 3794 1988
<< polycont >>
rect 928 5486 1296 5520
rect 1386 5486 1754 5520
rect 1844 5486 2212 5520
rect 2302 5486 2670 5520
rect 2760 5486 3128 5520
rect 928 3358 1296 3392
rect 1386 3358 1754 3392
rect 1844 3358 2212 3392
rect 2302 3358 2670 3392
rect 2760 3358 3128 3392
rect 3428 3358 3462 3392
rect 3744 3358 3778 3392
rect 12 3048 380 3082
rect 470 3048 838 3082
rect 928 3048 1296 3082
rect 1386 3048 1754 3082
rect 1844 3048 2212 3082
rect 2302 3048 2670 3082
rect 2760 3048 3128 3082
rect 12 1938 380 1972
rect 470 1938 838 1972
rect 928 1938 1296 1972
rect 1386 1938 1754 1972
rect 1844 1938 2212 1972
rect 2302 1938 2670 1972
rect 2760 1938 3128 1972
rect 3428 3048 3462 3082
rect 3744 3048 3778 3082
<< xpolycontact >>
rect 314 3386 384 3818
rect 480 3386 550 3818
<< xpolyres >>
rect 314 4252 550 4322
rect 314 3818 384 4252
rect 480 3818 550 4252
<< locali >>
rect 760 5680 3930 5690
rect 760 5622 770 5680
rect 3920 5622 3930 5680
rect 752 5610 770 5622
rect 3920 5610 3936 5622
rect 752 5588 848 5610
rect 3208 5588 3366 5610
rect 3524 5588 3682 5610
rect 3840 5588 3936 5610
rect 752 5526 786 5588
rect 184 4418 280 4452
rect 584 4418 680 4452
rect 184 4356 218 4418
rect 646 4356 680 4418
rect 310 3386 314 3810
rect 384 3386 390 3810
rect 310 3380 390 3386
rect 184 3290 218 3352
rect 646 3290 680 3352
rect 184 3256 280 3290
rect 584 3256 680 3290
rect 3270 5526 3304 5588
rect 912 5486 928 5520
rect 1296 5486 1312 5520
rect 1370 5486 1386 5520
rect 1754 5486 1770 5520
rect 1828 5486 1844 5520
rect 2212 5486 2228 5520
rect 2286 5486 2302 5520
rect 2670 5486 2686 5520
rect 2744 5486 2760 5520
rect 3128 5486 3144 5520
rect 866 5427 900 5443
rect 866 3435 900 3451
rect 1324 5427 1358 5443
rect 1324 3435 1358 3451
rect 1782 5427 1816 5443
rect 1782 3435 1816 3451
rect 2240 5427 2274 5443
rect 2240 3435 2274 3451
rect 2698 5427 2732 5443
rect 2698 3435 2732 3451
rect 3156 5427 3190 5443
rect 3156 3435 3190 3451
rect 912 3358 928 3392
rect 1296 3358 1312 3392
rect 1370 3358 1386 3392
rect 1754 3358 1770 3392
rect 1828 3358 1844 3392
rect 2212 3358 2228 3392
rect 2286 3358 2302 3392
rect 2670 3358 2686 3392
rect 2744 3358 2760 3392
rect 3128 3358 3144 3392
rect 752 3290 786 3352
rect 3586 5526 3620 5588
rect 3384 5427 3418 5443
rect 3384 3435 3418 3451
rect 3472 5427 3506 5443
rect 3472 3435 3506 3451
rect 3412 3358 3428 3392
rect 3462 3358 3478 3392
rect 3270 3290 3304 3352
rect 3902 5526 3936 5588
rect 3700 5427 3734 5443
rect 3700 3435 3734 3451
rect 3788 5427 3822 5443
rect 3788 3435 3822 3451
rect 3728 3358 3744 3392
rect 3778 3358 3794 3392
rect 3586 3290 3620 3352
rect 3902 3290 3936 3352
rect 752 3256 848 3290
rect 3208 3256 3366 3290
rect 3524 3256 3682 3290
rect 3840 3256 3936 3290
rect 184 3184 680 3256
rect -164 3150 -68 3184
rect 3208 3150 3366 3184
rect 3524 3150 3682 3184
rect 3840 3150 3936 3184
rect -164 3088 -130 3150
rect 3270 3088 3304 3150
rect -4 3048 12 3082
rect 380 3048 396 3082
rect 454 3048 470 3082
rect 838 3048 854 3082
rect 912 3048 928 3082
rect 1296 3048 1312 3082
rect 1370 3048 1386 3082
rect 1754 3048 1770 3082
rect 1828 3048 1844 3082
rect 2212 3048 2228 3082
rect 2286 3048 2302 3082
rect 2670 3048 2686 3082
rect 2744 3048 2760 3082
rect 3128 3048 3144 3082
rect -50 2998 -16 3014
rect -50 2006 -16 2022
rect 408 2998 442 3014
rect 408 2006 442 2022
rect 866 2998 900 3014
rect 866 2006 900 2022
rect 1324 2998 1358 3014
rect 1324 2006 1358 2022
rect 1782 2998 1816 3014
rect 1782 2006 1816 2022
rect 2240 2998 2274 3014
rect 2240 2006 2274 2022
rect 2698 2998 2732 3014
rect 2698 2006 2732 2022
rect 3156 2998 3190 3014
rect 3156 2006 3190 2022
rect -4 1938 12 1972
rect 380 1938 396 1972
rect 454 1938 470 1972
rect 838 1938 854 1972
rect 912 1938 928 1972
rect 1296 1938 1312 1972
rect 1370 1938 1386 1972
rect 1754 1938 1770 1972
rect 1828 1938 1844 1972
rect 2212 1938 2228 1972
rect 2286 1938 2302 1972
rect 2670 1938 2686 1972
rect 2744 1938 2760 1972
rect 3128 1938 3144 1972
rect -164 1870 -130 1932
rect 3586 3088 3620 3150
rect 3412 3048 3428 3082
rect 3462 3048 3478 3082
rect 3384 2998 3418 3014
rect 3384 2006 3418 2022
rect 3472 2998 3506 3014
rect 3472 2006 3506 2022
rect 3270 1870 3304 1932
rect 3902 3088 3936 3150
rect 3728 3048 3744 3082
rect 3778 3048 3794 3082
rect 3700 2998 3734 3014
rect 3700 2006 3734 2022
rect 3788 2998 3822 3014
rect 3788 2006 3822 2022
rect 3586 1870 3620 1932
rect 3902 1870 3936 1932
rect -164 1860 -68 1870
rect 3208 1860 3366 1870
rect 3524 1860 3682 1870
rect 3840 1860 3940 1870
rect -164 1840 -150 1860
rect -170 1780 -150 1840
rect 3920 1780 3940 1860
rect -170 1770 3940 1780
<< viali >>
rect 770 5622 3920 5680
rect 770 5610 848 5622
rect 848 5610 3208 5622
rect 3208 5610 3366 5622
rect 3366 5610 3524 5622
rect 3524 5610 3682 5622
rect 3682 5610 3840 5622
rect 3840 5610 3920 5622
rect 320 3390 380 3800
rect 490 3390 550 3800
rect 928 5486 1296 5520
rect 1386 5486 1754 5520
rect 1844 5486 2212 5520
rect 2302 5486 2670 5520
rect 2760 5486 3128 5520
rect 866 3451 900 5427
rect 1324 3451 1358 5427
rect 1782 3451 1816 5427
rect 2240 3451 2274 5427
rect 2698 3451 2732 5427
rect 3156 3451 3190 5427
rect 928 3358 1296 3392
rect 1386 3358 1754 3392
rect 1844 3358 2212 3392
rect 2302 3358 2670 3392
rect 2760 3358 3128 3392
rect 3384 3451 3418 5427
rect 3472 3451 3506 5427
rect 3428 3358 3462 3392
rect 3700 3451 3734 5427
rect 3788 3451 3822 5427
rect 3744 3358 3778 3392
rect 12 3048 380 3082
rect 470 3048 838 3082
rect 928 3048 1296 3082
rect 1386 3048 1754 3082
rect 1844 3048 2212 3082
rect 2302 3048 2670 3082
rect 2760 3048 3128 3082
rect -50 2022 -16 2998
rect 408 2022 442 2998
rect 866 2022 900 2998
rect 1324 2022 1358 2998
rect 1782 2022 1816 2998
rect 2240 2022 2274 2998
rect 2698 2022 2732 2998
rect 3156 2022 3190 2998
rect 12 1938 380 1972
rect 470 1938 838 1972
rect 928 1938 1296 1972
rect 1386 1938 1754 1972
rect 1844 1938 2212 1972
rect 2302 1938 2670 1972
rect 2760 1938 3128 1972
rect 3428 3048 3462 3082
rect 3384 2022 3418 2998
rect 3472 2022 3506 2998
rect 3744 3048 3778 3082
rect 3700 2022 3734 2998
rect 3788 2022 3822 2998
rect -150 1836 -68 1860
rect -68 1836 3208 1860
rect 3208 1836 3366 1860
rect 3366 1836 3524 1860
rect 3524 1836 3682 1860
rect 3682 1836 3840 1860
rect 3840 1836 3920 1860
rect -150 1780 3920 1836
<< metal1 >>
rect -200 5680 3940 5700
rect -200 5610 770 5680
rect 3920 5610 3940 5680
rect -200 5590 3940 5610
rect 916 5526 956 5590
rect 1268 5526 1308 5590
rect 2184 5526 2224 5590
rect 3100 5526 3140 5590
rect 916 5520 1308 5526
rect 916 5486 928 5520
rect 1296 5486 1308 5520
rect 916 5480 1308 5486
rect 1374 5520 1766 5526
rect 1374 5486 1386 5520
rect 1754 5486 1766 5520
rect 1374 5480 1766 5486
rect 1832 5520 2224 5526
rect 1832 5486 1844 5520
rect 2212 5486 2224 5520
rect 1832 5480 2224 5486
rect 2290 5520 2682 5526
rect 2290 5486 2302 5520
rect 2670 5486 2682 5520
rect 2290 5480 2682 5486
rect 2748 5520 3140 5526
rect 2748 5486 2760 5520
rect 3128 5486 3140 5520
rect 2748 5480 3140 5486
rect 916 5439 956 5480
rect 857 5427 956 5439
rect 310 3810 390 3820
rect 310 3380 320 3810
rect 380 3380 390 3810
rect 310 3370 390 3380
rect 480 3810 560 3820
rect 480 3380 490 3810
rect 550 3380 560 3810
rect 909 5403 956 5427
rect 1268 5439 1308 5480
rect 1720 5450 1760 5480
rect 1720 5439 1800 5450
rect 2184 5439 2224 5480
rect 3100 5439 3140 5480
rect 3820 5439 3900 5590
rect 1268 5427 1367 5439
rect 1268 5403 1315 5427
rect 909 3451 956 3530
rect 857 3439 956 3451
rect 480 3370 560 3380
rect 916 3398 956 3439
rect 1268 3451 1315 3521
rect 1720 5427 1825 5439
rect 1720 5370 1773 5427
rect 1268 3439 1367 3451
rect 1730 3451 1773 3520
rect 2184 5427 2283 5439
rect 2184 5357 2231 5427
rect 1730 3439 1825 3451
rect 2184 3451 2231 3521
rect 2689 5427 2741 5439
rect 2680 3470 2689 3660
rect 2184 3439 2283 3451
rect 3100 5427 3196 5439
rect 3378 5430 3424 5439
rect 3100 5357 3156 5427
rect 2741 3650 2760 3660
rect 2750 3480 2760 3650
rect 3150 3521 3156 5357
rect 2741 3470 2760 3480
rect 2689 3439 2741 3451
rect 3100 3451 3156 3521
rect 3190 3451 3196 5427
rect 3100 3439 3196 3451
rect 3340 5427 3424 5430
rect 3340 3800 3384 5427
rect 3340 3590 3350 3800
rect 3340 3451 3384 3590
rect 3418 3451 3424 5427
rect 3340 3450 3424 3451
rect 3378 3439 3424 3450
rect 3466 5430 3512 5439
rect 3694 5430 3740 5439
rect 3466 5427 3550 5430
rect 3466 3451 3472 5427
rect 3506 4040 3550 5427
rect 3660 5427 3740 5430
rect 3506 4030 3560 4040
rect 3540 3820 3560 4030
rect 3506 3810 3560 3820
rect 3506 3451 3550 3810
rect 3660 3492 3700 5427
rect 3466 3450 3550 3451
rect 3608 3451 3700 3492
rect 3734 3451 3740 5427
rect 3466 3439 3512 3450
rect 3608 3448 3740 3451
rect 1268 3398 1308 3439
rect 1730 3430 1790 3439
rect 1730 3400 1770 3430
rect 916 3392 1308 3398
rect 916 3358 928 3392
rect 1296 3358 1308 3392
rect 916 3352 1308 3358
rect 1370 3392 1770 3400
rect 2184 3398 2224 3439
rect 1370 3358 1386 3392
rect 1754 3358 1770 3392
rect 1370 3340 1770 3358
rect 1832 3392 2224 3398
rect 1832 3358 1844 3392
rect 2212 3358 2224 3392
rect 1832 3352 2224 3358
rect 2290 3392 2690 3400
rect 3100 3398 3140 3439
rect 2290 3358 2302 3392
rect 2670 3358 2690 3392
rect 1370 3280 1600 3340
rect 1700 3320 1770 3340
rect 2290 3320 2690 3358
rect 2748 3392 3140 3398
rect 2748 3358 2760 3392
rect 3128 3358 3140 3392
rect 2748 3352 3140 3358
rect 3400 3400 3480 3410
rect 3400 3340 3410 3400
rect 3470 3340 3480 3400
rect 3400 3330 3480 3340
rect 1700 3280 2690 3320
rect 3608 3250 3652 3448
rect 3694 3439 3740 3448
rect 3782 5427 3900 5439
rect 3782 3451 3788 5427
rect 3822 3451 3900 5427
rect 3782 3450 3900 3451
rect 3782 3439 3828 3450
rect 3730 3400 3810 3410
rect 3730 3340 3740 3400
rect 3800 3340 3810 3400
rect 3730 3330 3810 3340
rect 3320 3200 3652 3250
rect 450 3120 2680 3160
rect -50 3088 10 3090
rect -50 3082 420 3088
rect -50 3048 12 3082
rect 380 3048 420 3082
rect 450 3082 850 3120
rect 450 3080 470 3082
rect -50 3042 420 3048
rect 458 3048 470 3080
rect 838 3048 850 3082
rect 458 3042 850 3048
rect 916 3082 1308 3088
rect 916 3048 928 3082
rect 1296 3048 1308 3082
rect 916 3042 1308 3048
rect -50 3040 10 3042
rect -50 3010 -20 3040
rect 380 3010 420 3042
rect 810 3010 850 3042
rect 1268 3011 1308 3042
rect 1370 3082 1770 3120
rect 2290 3088 2680 3120
rect 1370 3048 1386 3082
rect 1754 3048 1770 3082
rect 1370 3040 1770 3048
rect 1832 3082 2224 3088
rect 1832 3048 1844 3082
rect 2212 3048 2224 3082
rect 1832 3042 2224 3048
rect 1268 3010 1325 3011
rect 2184 3010 2224 3042
rect 2290 3082 2682 3088
rect 2290 3048 2302 3082
rect 2670 3048 2682 3082
rect 2290 3042 2682 3048
rect 2748 3082 3140 3088
rect 2748 3048 2760 3082
rect 3128 3048 3140 3082
rect 2748 3042 3140 3048
rect 2290 3040 2680 3042
rect 3100 3010 3140 3042
rect 3320 3010 3360 3200
rect 3622 3198 3652 3200
rect 3400 3110 3480 3120
rect 3400 3050 3410 3110
rect 3470 3050 3480 3110
rect 3400 3048 3428 3050
rect 3462 3048 3480 3050
rect 3400 3040 3480 3048
rect 3730 3110 3810 3120
rect 3730 3050 3740 3110
rect 3800 3050 3810 3110
rect 3730 3048 3744 3050
rect 3778 3048 3810 3050
rect 3730 3040 3810 3048
rect -59 2998 -7 3010
rect 380 2998 451 3010
rect 380 2980 399 2998
rect -59 2010 -7 2022
rect 352 2022 399 2076
rect 810 2998 909 3010
rect 810 2920 857 2998
rect 352 2010 451 2022
rect 810 2022 857 2100
rect 1268 2998 1367 3010
rect 1268 2920 1315 2998
rect 810 2010 909 2022
rect 1268 2022 1315 2101
rect 1773 2998 1825 3010
rect 1760 2970 1773 2980
rect 1760 2870 1770 2970
rect 1760 2860 1773 2870
rect 1268 2010 1367 2022
rect 2184 2998 2283 3010
rect 1825 2970 1840 2980
rect 1830 2870 1840 2970
rect 2184 2919 2231 2998
rect 1825 2860 1840 2870
rect 1773 2010 1825 2022
rect 2184 2022 2231 2101
rect 2689 2998 2741 3010
rect 2680 2790 2689 2980
rect 2184 2010 2283 2022
rect 3100 2998 3196 3010
rect 2741 2970 2760 2980
rect 2750 2800 2760 2970
rect 3100 2944 3156 2998
rect 2741 2790 2760 2800
rect 3150 2076 3156 2944
rect 2689 2010 2741 2022
rect 3100 2022 3156 2076
rect 3190 2022 3196 2998
rect 3320 2998 3424 3010
rect 3320 2860 3384 2998
rect 3100 2010 3196 2022
rect 3340 2650 3350 2860
rect 3340 2022 3384 2650
rect 3418 2022 3424 2998
rect 3340 2020 3424 2022
rect 3378 2010 3424 2020
rect 3466 2998 3550 3010
rect 3466 2022 3472 2998
rect 3506 2640 3550 2998
rect 3650 3000 3740 3010
rect 3650 2940 3660 3000
rect 3720 2998 3740 3000
rect 3650 2930 3700 2940
rect 3506 2630 3560 2640
rect 3550 2420 3560 2630
rect 3506 2410 3560 2420
rect 3506 2022 3550 2410
rect 3466 2020 3550 2022
rect 3660 2022 3700 2930
rect 3734 2022 3740 2998
rect 3660 2020 3740 2022
rect 3466 2010 3512 2020
rect 3694 2010 3740 2020
rect 3782 3000 3828 3010
rect 3782 2998 3900 3000
rect 3782 2022 3788 2998
rect 3822 2022 3900 2998
rect 3782 2010 3900 2022
rect -50 1980 -20 2010
rect -50 1978 10 1980
rect 352 1978 392 2010
rect 810 1978 850 2010
rect 1268 1978 1308 2010
rect 2184 1978 2224 2010
rect 3100 1978 3140 2010
rect -50 1972 392 1978
rect -50 1938 12 1972
rect 380 1938 392 1972
rect -50 1932 392 1938
rect 458 1972 850 1978
rect 458 1938 470 1972
rect 838 1938 850 1972
rect 458 1932 850 1938
rect 916 1972 1308 1978
rect 916 1938 928 1972
rect 1296 1938 1308 1972
rect 916 1932 1308 1938
rect 1374 1972 1766 1978
rect 1374 1938 1386 1972
rect 1754 1938 1766 1972
rect 1374 1932 1766 1938
rect 1832 1972 2224 1978
rect 1832 1938 1844 1972
rect 2212 1938 2224 1972
rect 1832 1932 2224 1938
rect 2290 1972 2682 1978
rect 2290 1938 2302 1972
rect 2670 1938 2682 1972
rect 2290 1932 2682 1938
rect 2748 1972 3140 1978
rect 2748 1938 2760 1972
rect 3128 1938 3140 1972
rect 2748 1932 3140 1938
rect -50 1930 10 1932
rect -50 1870 -20 1930
rect 352 1870 392 1932
rect 810 1930 850 1932
rect 1268 1870 1308 1932
rect 2184 1870 2224 1932
rect 3100 1870 3140 1932
rect 3820 1870 3900 2010
rect -200 1860 3940 1870
rect -200 1780 -150 1860
rect 3920 1780 3940 1860
rect -200 1760 3940 1780
<< via1 >>
rect 770 5610 3920 5680
rect 320 3800 380 3810
rect 320 3390 380 3800
rect 320 3380 380 3390
rect 490 3800 550 3810
rect 490 3390 550 3800
rect 490 3380 550 3390
rect 857 3451 866 5427
rect 866 3451 900 5427
rect 900 3451 909 5427
rect 1315 3451 1324 5427
rect 1324 3451 1358 5427
rect 1358 3451 1367 5427
rect 1773 3451 1782 5427
rect 1782 3451 1816 5427
rect 1816 3451 1825 5427
rect 2231 3451 2240 5427
rect 2240 3451 2274 5427
rect 2274 3451 2283 5427
rect 2689 3451 2698 5427
rect 2698 3451 2732 5427
rect 2732 3650 2741 5427
rect 2732 3480 2750 3650
rect 2732 3451 2741 3480
rect 3350 3590 3384 3800
rect 3384 3590 3410 3800
rect 3480 3820 3506 4030
rect 3506 3820 3540 4030
rect 1600 3280 1700 3340
rect 3410 3392 3470 3400
rect 3410 3358 3428 3392
rect 3428 3358 3462 3392
rect 3462 3358 3470 3392
rect 3410 3340 3470 3358
rect 3740 3392 3800 3400
rect 3740 3358 3744 3392
rect 3744 3358 3778 3392
rect 3778 3358 3800 3392
rect 3740 3340 3800 3358
rect 3410 3082 3470 3110
rect 3410 3050 3428 3082
rect 3428 3050 3462 3082
rect 3462 3050 3470 3082
rect 3740 3082 3800 3110
rect 3740 3050 3744 3082
rect 3744 3050 3778 3082
rect 3778 3050 3800 3082
rect -59 2022 -50 2998
rect -50 2022 -16 2998
rect -16 2022 -7 2998
rect 399 2022 408 2998
rect 408 2022 442 2998
rect 442 2022 451 2998
rect 857 2022 866 2998
rect 866 2022 900 2998
rect 900 2022 909 2998
rect 1315 2022 1324 2998
rect 1324 2022 1358 2998
rect 1358 2022 1367 2998
rect 1773 2970 1782 2998
rect 1770 2870 1782 2970
rect 1773 2022 1782 2870
rect 1782 2022 1816 2998
rect 1816 2970 1825 2998
rect 1816 2870 1830 2970
rect 1816 2022 1825 2870
rect 2231 2022 2240 2998
rect 2240 2022 2274 2998
rect 2274 2022 2283 2998
rect 2689 2022 2698 2998
rect 2698 2022 2732 2998
rect 2732 2970 2741 2998
rect 2732 2800 2750 2970
rect 2732 2022 2741 2800
rect 3350 2650 3384 2860
rect 3384 2650 3410 2860
rect 3660 2998 3720 3000
rect 3660 2940 3700 2998
rect 3700 2940 3720 2998
rect 3480 2420 3506 2630
rect 3506 2420 3550 2630
rect -150 1780 3920 1860
<< metal2 >>
rect -200 5680 3940 5700
rect -200 5610 770 5680
rect 3920 5610 3940 5680
rect -200 5590 3940 5610
rect 857 5427 909 5439
rect 310 3810 390 3820
rect 310 3380 320 3810
rect 380 3380 390 3810
rect 310 3370 390 3380
rect 480 3810 560 3820
rect 480 3380 490 3810
rect 550 3380 560 3810
rect 857 3439 909 3451
rect 1315 5427 1367 5439
rect 1315 3439 1367 3451
rect 1773 5427 1825 5439
rect 1773 3439 1825 3451
rect 2231 5427 2283 5439
rect 2689 5427 2741 5439
rect 2680 3470 2689 3660
rect 3470 4030 3560 4040
rect 3470 3820 3480 4030
rect 3540 3820 3560 4030
rect 3470 3810 3560 3820
rect 3340 3800 3420 3810
rect 3340 3660 3350 3800
rect 2741 3650 3350 3660
rect 2750 3590 3350 3650
rect 3410 3590 3420 3800
rect 2750 3580 3420 3590
rect 2750 3480 2760 3580
rect 2231 3439 2283 3451
rect 2741 3470 2760 3480
rect 2689 3439 2741 3451
rect 480 3370 560 3380
rect 330 3140 370 3370
rect 500 3240 540 3370
rect 1590 3340 1710 3350
rect 1590 3280 1600 3340
rect 1700 3310 1710 3340
rect 1700 3280 1780 3310
rect 1590 3270 1780 3280
rect 1740 3240 1780 3270
rect 3320 3300 3370 3580
rect 3400 3400 3480 3410
rect 3400 3340 3410 3400
rect 3470 3340 3480 3400
rect 3400 3330 3480 3340
rect 3730 3400 3810 3410
rect 3730 3340 3740 3400
rect 3800 3340 3810 3400
rect 3730 3330 3810 3340
rect 3320 3250 3620 3300
rect 500 3200 1780 3240
rect 330 3100 1820 3140
rect 1780 3010 1820 3100
rect 3400 3110 3480 3120
rect 3400 3050 3410 3110
rect 3470 3050 3480 3110
rect 3400 3040 3480 3050
rect 3580 3010 3620 3250
rect 3730 3110 3810 3120
rect 3730 3050 3740 3110
rect 3800 3050 3810 3110
rect 3730 3040 3810 3050
rect -59 2998 -7 3010
rect -59 2010 -7 2022
rect 399 2998 451 3010
rect 399 2010 451 2022
rect 857 2998 909 3010
rect 857 2010 909 2022
rect 1315 2998 1367 3010
rect 1773 2998 1825 3010
rect 1760 2970 1773 2980
rect 2231 2998 2283 3010
rect 1825 2970 1840 2980
rect 1760 2870 1770 2970
rect 1830 2870 1840 2970
rect 1760 2860 1773 2870
rect 1315 2010 1367 2022
rect 1825 2860 1840 2870
rect 1773 2010 1825 2022
rect 2689 2998 2741 3010
rect 2680 2790 2689 2980
rect 3580 3000 3730 3010
rect 2741 2970 2760 2980
rect 3580 2970 3660 3000
rect 2750 2870 2760 2970
rect 3650 2940 3660 2970
rect 3720 2940 3730 3000
rect 3650 2930 3730 2940
rect 2750 2860 3420 2870
rect 2750 2800 3350 2860
rect 2231 2010 2283 2022
rect 2741 2790 3350 2800
rect 3340 2650 3350 2790
rect 3410 2650 3420 2860
rect 3340 2640 3420 2650
rect 3470 2630 3560 2640
rect 3470 2420 3480 2630
rect 3550 2420 3560 2630
rect 3470 2410 3560 2420
rect 2689 2010 2741 2022
rect -200 1860 3940 1870
rect -200 1780 -150 1860
rect 3920 1780 3940 1860
rect -200 1760 3940 1780
<< via2 >>
rect 3480 3820 3540 4030
rect 3410 3340 3470 3400
rect 3740 3340 3800 3400
rect 3410 3050 3470 3110
rect 3740 3050 3800 3110
rect 3480 2420 3550 2630
<< metal3 >>
rect 3470 4030 3560 4040
rect 3470 3820 3480 4030
rect 3550 3820 3560 4030
rect 3470 3810 3560 3820
rect 3240 3490 3800 3550
rect 3240 3110 3300 3490
rect 3740 3410 3800 3490
rect 3400 3400 3530 3410
rect 3730 3400 3810 3410
rect 3400 3340 3410 3400
rect 3470 3340 3650 3400
rect 3400 3330 3530 3340
rect 3400 3110 3480 3120
rect 3240 3050 3410 3110
rect 3470 3050 3480 3110
rect 3590 3110 3650 3340
rect 3730 3340 3740 3400
rect 3800 3340 3810 3400
rect 3730 3330 3810 3340
rect 3730 3110 3810 3120
rect 3590 3050 3740 3110
rect 3800 3050 3810 3110
rect 3400 3040 3480 3050
rect 3730 3040 3810 3050
rect 3470 2630 3560 2640
rect 3470 2420 3480 2630
rect 3550 2420 3560 2630
rect 3470 2410 3560 2420
<< via3 >>
rect 3480 3820 3540 4030
rect 3540 3820 3550 4030
rect 3480 2420 3550 2630
<< metal4 >>
rect 3470 4030 3560 4040
rect 3470 3820 3480 4030
rect 3550 3930 3560 4030
rect 3550 3820 4090 3930
rect 3470 3810 4090 3820
rect 3950 2640 4090 3810
rect 3470 2630 4090 2640
rect 3470 2420 3480 2630
rect 3550 2520 4090 2630
rect 3550 2420 3560 2520
rect 3470 2410 3560 2420
<< labels >>
rlabel metal4 4010 3760 4090 3930 1 IOUT
rlabel metal3 3240 3210 3300 3250 1 GN
rlabel metal3 3590 3180 3650 3220 1 GP
rlabel metal1 810 2920 850 3020 1 IIN
rlabel metal2 -200 5590 -40 5700 1 VHI
rlabel metal2 -200 1760 -40 1870 1 VLO
rlabel metal2 2950 3580 3030 3660 1 IP
rlabel metal2 2980 2790 3060 2870 1 IN
rlabel metal1 2150 3120 2220 3160 1 VREFN
rlabel metal1 2130 3280 2200 3320 1 VREFP
<< end >>
