magic
tech sky130A
timestamp 1671856587
<< metal1 >>
rect 11600 -3700 11650 -3600
rect 11750 -3700 11800 -3600
rect 11630 -3860 11635 -3820
rect 11705 -3860 11710 -3820
rect 11770 -3860 11775 -3820
rect 11845 -3860 11850 -3820
rect 11600 -4050 11650 -3950
rect 11750 -4050 11800 -3950
rect 8195 -4760 8235 -4755
rect 8195 -4790 8200 -4760
rect 8230 -4790 8235 -4760
rect 8195 -4795 8235 -4790
rect 8250 -4825 8270 -4775
rect 8230 -4830 8270 -4825
rect 8230 -4860 8235 -4830
rect 8265 -4860 8270 -4830
rect 8230 -4865 8270 -4860
rect 8350 -5255 8405 -5250
rect 8350 -5425 8355 -5255
rect 8400 -5425 8405 -5255
rect 8700 -5255 8760 -5250
rect 8510 -5310 8570 -5305
rect 8510 -5370 8515 -5310
rect 8565 -5370 8570 -5310
rect 8510 -5375 8570 -5370
rect 8350 -5430 8405 -5425
rect 8700 -5425 8710 -5255
rect 8755 -5425 8760 -5255
rect 8700 -5430 8760 -5425
rect 3000 -5624 7000 -5500
rect 3000 -5650 3307 -5624
rect 3333 -5650 3467 -5624
rect 3493 -5650 3627 -5624
rect 3653 -5650 3787 -5624
rect 3813 -5650 3947 -5624
rect 3973 -5650 4107 -5624
rect 4133 -5650 4267 -5624
rect 4293 -5650 4427 -5624
rect 4453 -5650 4587 -5624
rect 4613 -5650 4747 -5624
rect 4773 -5650 4907 -5624
rect 4933 -5650 5067 -5624
rect 5093 -5650 5227 -5624
rect 5253 -5650 5387 -5624
rect 5413 -5650 5547 -5624
rect 5573 -5650 5707 -5624
rect 5733 -5650 5867 -5624
rect 5893 -5650 6027 -5624
rect 6053 -5650 6187 -5624
rect 6213 -5650 6347 -5624
rect 6373 -5650 6507 -5624
rect 6533 -5650 6667 -5624
rect 6693 -5650 7000 -5624
rect 3000 -5727 7000 -5650
rect 3000 -5753 3122 -5727
rect 3148 -5753 6855 -5727
rect 6881 -5753 7000 -5727
rect 3000 -5770 7000 -5753
rect 3000 -5887 3270 -5770
rect 3000 -5913 3122 -5887
rect 3148 -5913 3270 -5887
rect 3000 -6047 3270 -5913
rect 3000 -6073 3122 -6047
rect 3148 -6073 3270 -6047
rect 3000 -6207 3270 -6073
rect 3000 -6233 3122 -6207
rect 3148 -6233 3270 -6207
rect 3000 -6367 3270 -6233
rect 3000 -6393 3122 -6367
rect 3148 -6393 3270 -6367
rect 3000 -6527 3270 -6393
rect 3000 -6553 3122 -6527
rect 3148 -6553 3270 -6527
rect 3000 -6687 3270 -6553
rect 3000 -6713 3122 -6687
rect 3148 -6713 3270 -6687
rect 3000 -6847 3270 -6713
rect 3000 -6873 3122 -6847
rect 3148 -6873 3270 -6847
rect 3000 -7007 3270 -6873
rect 3000 -7033 3122 -7007
rect 3148 -7033 3270 -7007
rect 3000 -7167 3270 -7033
rect 3000 -7193 3122 -7167
rect 3148 -7193 3270 -7167
rect 3000 -7327 3270 -7193
rect 3000 -7353 3122 -7327
rect 3148 -7353 3270 -7327
rect 3000 -7487 3270 -7353
rect 3000 -7513 3122 -7487
rect 3148 -7513 3270 -7487
rect 3000 -7647 3270 -7513
rect 3000 -7673 3122 -7647
rect 3148 -7673 3270 -7647
rect 3000 -7807 3270 -7673
rect 3000 -7833 3122 -7807
rect 3148 -7833 3270 -7807
rect 3000 -7967 3270 -7833
rect 3000 -7993 3122 -7967
rect 3148 -7993 3270 -7967
rect 3000 -8127 3270 -7993
rect 3000 -8153 3122 -8127
rect 3148 -8153 3270 -8127
rect 3000 -8287 3270 -8153
rect 3000 -8313 3122 -8287
rect 3148 -8313 3270 -8287
rect 3000 -8447 3270 -8313
rect 3000 -8473 3122 -8447
rect 3148 -8473 3270 -8447
rect 3000 -8607 3270 -8473
rect 3000 -8633 3122 -8607
rect 3148 -8633 3270 -8607
rect 3000 -8767 3270 -8633
rect 3000 -8793 3122 -8767
rect 3148 -8793 3270 -8767
rect 3000 -8927 3270 -8793
rect 3000 -8953 3122 -8927
rect 3148 -8953 3270 -8927
rect 3000 -9087 3270 -8953
rect 3000 -9113 3122 -9087
rect 3148 -9113 3270 -9087
rect 3000 -9230 3270 -9113
rect 6730 -5887 7000 -5770
rect 6730 -5913 6855 -5887
rect 6881 -5913 7000 -5887
rect 6730 -6047 7000 -5913
rect 6730 -6073 6855 -6047
rect 6881 -6073 7000 -6047
rect 6730 -6207 7000 -6073
rect 6730 -6233 6855 -6207
rect 6881 -6233 7000 -6207
rect 6730 -6367 7000 -6233
rect 6730 -6393 6855 -6367
rect 6881 -6393 7000 -6367
rect 6730 -6527 7000 -6393
rect 6730 -6553 6855 -6527
rect 6881 -6553 7000 -6527
rect 6730 -6687 7000 -6553
rect 6730 -6713 6855 -6687
rect 6881 -6713 7000 -6687
rect 6730 -6847 7000 -6713
rect 6730 -6873 6855 -6847
rect 6881 -6873 7000 -6847
rect 6730 -7007 7000 -6873
rect 6730 -7033 6855 -7007
rect 6881 -7033 7000 -7007
rect 6730 -7167 7000 -7033
rect 6730 -7193 6855 -7167
rect 6881 -7193 7000 -7167
rect 6730 -7327 7000 -7193
rect 6730 -7353 6855 -7327
rect 6881 -7353 7000 -7327
rect 6730 -7487 7000 -7353
rect 6730 -7513 6855 -7487
rect 6881 -7513 7000 -7487
rect 6730 -7647 7000 -7513
rect 6730 -7673 6855 -7647
rect 6881 -7673 7000 -7647
rect 6730 -7807 7000 -7673
rect 6730 -7833 6855 -7807
rect 6881 -7833 7000 -7807
rect 6730 -7967 7000 -7833
rect 6730 -7993 6855 -7967
rect 6881 -7993 7000 -7967
rect 6730 -8127 7000 -7993
rect 6730 -8153 6855 -8127
rect 6881 -8153 7000 -8127
rect 6730 -8287 7000 -8153
rect 6730 -8313 6855 -8287
rect 6881 -8313 7000 -8287
rect 6730 -8447 7000 -8313
rect 6730 -8473 6855 -8447
rect 6881 -8473 7000 -8447
rect 6730 -8607 7000 -8473
rect 6730 -8633 6855 -8607
rect 6881 -8633 7000 -8607
rect 6730 -8767 7000 -8633
rect 6730 -8793 6855 -8767
rect 6881 -8793 7000 -8767
rect 6730 -8927 7000 -8793
rect 6730 -8953 6855 -8927
rect 6881 -8953 7000 -8927
rect 6730 -9087 7000 -8953
rect 6730 -9113 6855 -9087
rect 6881 -9113 7000 -9087
rect 6730 -9230 7000 -9113
rect 3000 -9247 7000 -9230
rect 3000 -9273 3122 -9247
rect 3148 -9273 6855 -9247
rect 6881 -9273 7000 -9247
rect 3000 -9352 7000 -9273
rect 3000 -9378 3307 -9352
rect 3333 -9378 3467 -9352
rect 3493 -9378 3627 -9352
rect 3653 -9378 3787 -9352
rect 3813 -9378 3947 -9352
rect 3973 -9378 4107 -9352
rect 4133 -9378 4267 -9352
rect 4293 -9378 4427 -9352
rect 4453 -9378 4587 -9352
rect 4613 -9378 4747 -9352
rect 4773 -9378 4907 -9352
rect 4933 -9378 5067 -9352
rect 5093 -9378 5227 -9352
rect 5253 -9378 5387 -9352
rect 5413 -9378 5547 -9352
rect 5573 -9378 5707 -9352
rect 5733 -9378 5867 -9352
rect 5893 -9378 6027 -9352
rect 6053 -9378 6187 -9352
rect 6213 -9378 6347 -9352
rect 6373 -9378 6507 -9352
rect 6533 -9378 6667 -9352
rect 6693 -9378 7000 -9352
rect 3000 -9500 7000 -9378
rect 9000 -5624 13000 -5500
rect 9000 -5650 9307 -5624
rect 9333 -5650 9467 -5624
rect 9493 -5650 9627 -5624
rect 9653 -5650 9787 -5624
rect 9813 -5650 9947 -5624
rect 9973 -5650 10107 -5624
rect 10133 -5650 10267 -5624
rect 10293 -5650 10427 -5624
rect 10453 -5650 10587 -5624
rect 10613 -5650 10747 -5624
rect 10773 -5650 10907 -5624
rect 10933 -5650 11067 -5624
rect 11093 -5650 11227 -5624
rect 11253 -5650 11387 -5624
rect 11413 -5650 11547 -5624
rect 11573 -5650 11707 -5624
rect 11733 -5650 11867 -5624
rect 11893 -5650 12027 -5624
rect 12053 -5650 12187 -5624
rect 12213 -5650 12347 -5624
rect 12373 -5650 12507 -5624
rect 12533 -5650 12667 -5624
rect 12693 -5650 13000 -5624
rect 9000 -5727 13000 -5650
rect 9000 -5753 9122 -5727
rect 9148 -5753 12855 -5727
rect 12881 -5753 13000 -5727
rect 9000 -5770 13000 -5753
rect 9000 -5887 9270 -5770
rect 9000 -5913 9122 -5887
rect 9148 -5913 9270 -5887
rect 9000 -6047 9270 -5913
rect 9000 -6073 9122 -6047
rect 9148 -6073 9270 -6047
rect 9000 -6207 9270 -6073
rect 9000 -6233 9122 -6207
rect 9148 -6233 9270 -6207
rect 9000 -6367 9270 -6233
rect 9000 -6393 9122 -6367
rect 9148 -6393 9270 -6367
rect 9000 -6527 9270 -6393
rect 9000 -6553 9122 -6527
rect 9148 -6553 9270 -6527
rect 9000 -6687 9270 -6553
rect 9000 -6713 9122 -6687
rect 9148 -6713 9270 -6687
rect 9000 -6847 9270 -6713
rect 9000 -6873 9122 -6847
rect 9148 -6873 9270 -6847
rect 9000 -7007 9270 -6873
rect 9000 -7033 9122 -7007
rect 9148 -7033 9270 -7007
rect 9000 -7167 9270 -7033
rect 9000 -7193 9122 -7167
rect 9148 -7193 9270 -7167
rect 9000 -7327 9270 -7193
rect 9000 -7353 9122 -7327
rect 9148 -7353 9270 -7327
rect 9000 -7487 9270 -7353
rect 9000 -7513 9122 -7487
rect 9148 -7513 9270 -7487
rect 9000 -7647 9270 -7513
rect 9000 -7673 9122 -7647
rect 9148 -7673 9270 -7647
rect 9000 -7807 9270 -7673
rect 9000 -7833 9122 -7807
rect 9148 -7833 9270 -7807
rect 9000 -7967 9270 -7833
rect 9000 -7993 9122 -7967
rect 9148 -7993 9270 -7967
rect 9000 -8127 9270 -7993
rect 9000 -8153 9122 -8127
rect 9148 -8153 9270 -8127
rect 9000 -8287 9270 -8153
rect 9000 -8313 9122 -8287
rect 9148 -8313 9270 -8287
rect 9000 -8447 9270 -8313
rect 9000 -8473 9122 -8447
rect 9148 -8473 9270 -8447
rect 9000 -8607 9270 -8473
rect 9000 -8633 9122 -8607
rect 9148 -8633 9270 -8607
rect 9000 -8767 9270 -8633
rect 9000 -8793 9122 -8767
rect 9148 -8793 9270 -8767
rect 9000 -8927 9270 -8793
rect 9000 -8953 9122 -8927
rect 9148 -8953 9270 -8927
rect 9000 -9087 9270 -8953
rect 9000 -9113 9122 -9087
rect 9148 -9113 9270 -9087
rect 9000 -9230 9270 -9113
rect 12730 -5887 13000 -5770
rect 12730 -5913 12855 -5887
rect 12881 -5913 13000 -5887
rect 12730 -6047 13000 -5913
rect 12730 -6073 12855 -6047
rect 12881 -6073 13000 -6047
rect 12730 -6207 13000 -6073
rect 12730 -6233 12855 -6207
rect 12881 -6233 13000 -6207
rect 12730 -6367 13000 -6233
rect 12730 -6393 12855 -6367
rect 12881 -6393 13000 -6367
rect 12730 -6527 13000 -6393
rect 12730 -6553 12855 -6527
rect 12881 -6553 13000 -6527
rect 12730 -6687 13000 -6553
rect 12730 -6713 12855 -6687
rect 12881 -6713 13000 -6687
rect 12730 -6847 13000 -6713
rect 12730 -6873 12855 -6847
rect 12881 -6873 13000 -6847
rect 12730 -7007 13000 -6873
rect 12730 -7033 12855 -7007
rect 12881 -7033 13000 -7007
rect 12730 -7167 13000 -7033
rect 12730 -7193 12855 -7167
rect 12881 -7193 13000 -7167
rect 12730 -7327 13000 -7193
rect 12730 -7353 12855 -7327
rect 12881 -7353 13000 -7327
rect 12730 -7487 13000 -7353
rect 12730 -7513 12855 -7487
rect 12881 -7513 13000 -7487
rect 12730 -7647 13000 -7513
rect 12730 -7673 12855 -7647
rect 12881 -7673 13000 -7647
rect 12730 -7807 13000 -7673
rect 12730 -7833 12855 -7807
rect 12881 -7833 13000 -7807
rect 12730 -7967 13000 -7833
rect 12730 -7993 12855 -7967
rect 12881 -7993 13000 -7967
rect 12730 -8127 13000 -7993
rect 12730 -8153 12855 -8127
rect 12881 -8153 13000 -8127
rect 12730 -8287 13000 -8153
rect 12730 -8313 12855 -8287
rect 12881 -8313 13000 -8287
rect 12730 -8447 13000 -8313
rect 12730 -8473 12855 -8447
rect 12881 -8473 13000 -8447
rect 12730 -8607 13000 -8473
rect 12730 -8633 12855 -8607
rect 12881 -8633 13000 -8607
rect 12730 -8767 13000 -8633
rect 12730 -8793 12855 -8767
rect 12881 -8793 13000 -8767
rect 12730 -8927 13000 -8793
rect 12730 -8953 12855 -8927
rect 12881 -8953 13000 -8927
rect 12730 -9087 13000 -8953
rect 12730 -9113 12855 -9087
rect 12881 -9113 13000 -9087
rect 12730 -9230 13000 -9113
rect 9000 -9247 13000 -9230
rect 9000 -9273 9122 -9247
rect 9148 -9273 12855 -9247
rect 12881 -9273 13000 -9247
rect 9000 -9352 13000 -9273
rect 9000 -9378 9307 -9352
rect 9333 -9378 9467 -9352
rect 9493 -9378 9627 -9352
rect 9653 -9378 9787 -9352
rect 9813 -9378 9947 -9352
rect 9973 -9378 10107 -9352
rect 10133 -9378 10267 -9352
rect 10293 -9378 10427 -9352
rect 10453 -9378 10587 -9352
rect 10613 -9378 10747 -9352
rect 10773 -9378 10907 -9352
rect 10933 -9378 11067 -9352
rect 11093 -9378 11227 -9352
rect 11253 -9378 11387 -9352
rect 11413 -9378 11547 -9352
rect 11573 -9378 11707 -9352
rect 11733 -9378 11867 -9352
rect 11893 -9378 12027 -9352
rect 12053 -9378 12187 -9352
rect 12213 -9378 12347 -9352
rect 12373 -9378 12507 -9352
rect 12533 -9378 12667 -9352
rect 12693 -9378 13000 -9352
rect 9000 -9500 13000 -9378
rect 15000 -5624 19000 -5500
rect 15000 -5650 15307 -5624
rect 15333 -5650 15467 -5624
rect 15493 -5650 15627 -5624
rect 15653 -5650 15787 -5624
rect 15813 -5650 15947 -5624
rect 15973 -5650 16107 -5624
rect 16133 -5650 16267 -5624
rect 16293 -5650 16427 -5624
rect 16453 -5650 16587 -5624
rect 16613 -5650 16747 -5624
rect 16773 -5650 16907 -5624
rect 16933 -5650 17067 -5624
rect 17093 -5650 17227 -5624
rect 17253 -5650 17387 -5624
rect 17413 -5650 17547 -5624
rect 17573 -5650 17707 -5624
rect 17733 -5650 17867 -5624
rect 17893 -5650 18027 -5624
rect 18053 -5650 18187 -5624
rect 18213 -5650 18347 -5624
rect 18373 -5650 18507 -5624
rect 18533 -5650 18667 -5624
rect 18693 -5650 19000 -5624
rect 15000 -5727 19000 -5650
rect 15000 -5753 15122 -5727
rect 15148 -5753 18855 -5727
rect 18881 -5753 19000 -5727
rect 15000 -5770 19000 -5753
rect 15000 -5887 15270 -5770
rect 15000 -5913 15122 -5887
rect 15148 -5913 15270 -5887
rect 15000 -6047 15270 -5913
rect 15000 -6073 15122 -6047
rect 15148 -6073 15270 -6047
rect 15000 -6207 15270 -6073
rect 15000 -6233 15122 -6207
rect 15148 -6233 15270 -6207
rect 15000 -6367 15270 -6233
rect 15000 -6393 15122 -6367
rect 15148 -6393 15270 -6367
rect 15000 -6527 15270 -6393
rect 15000 -6553 15122 -6527
rect 15148 -6553 15270 -6527
rect 15000 -6687 15270 -6553
rect 15000 -6713 15122 -6687
rect 15148 -6713 15270 -6687
rect 15000 -6847 15270 -6713
rect 15000 -6873 15122 -6847
rect 15148 -6873 15270 -6847
rect 15000 -7007 15270 -6873
rect 15000 -7033 15122 -7007
rect 15148 -7033 15270 -7007
rect 15000 -7167 15270 -7033
rect 15000 -7193 15122 -7167
rect 15148 -7193 15270 -7167
rect 15000 -7327 15270 -7193
rect 15000 -7353 15122 -7327
rect 15148 -7353 15270 -7327
rect 15000 -7487 15270 -7353
rect 15000 -7513 15122 -7487
rect 15148 -7513 15270 -7487
rect 15000 -7647 15270 -7513
rect 15000 -7673 15122 -7647
rect 15148 -7673 15270 -7647
rect 15000 -7807 15270 -7673
rect 15000 -7833 15122 -7807
rect 15148 -7833 15270 -7807
rect 15000 -7967 15270 -7833
rect 15000 -7993 15122 -7967
rect 15148 -7993 15270 -7967
rect 15000 -8127 15270 -7993
rect 15000 -8153 15122 -8127
rect 15148 -8153 15270 -8127
rect 15000 -8287 15270 -8153
rect 15000 -8313 15122 -8287
rect 15148 -8313 15270 -8287
rect 15000 -8447 15270 -8313
rect 15000 -8473 15122 -8447
rect 15148 -8473 15270 -8447
rect 15000 -8607 15270 -8473
rect 15000 -8633 15122 -8607
rect 15148 -8633 15270 -8607
rect 15000 -8767 15270 -8633
rect 15000 -8793 15122 -8767
rect 15148 -8793 15270 -8767
rect 15000 -8927 15270 -8793
rect 15000 -8953 15122 -8927
rect 15148 -8953 15270 -8927
rect 15000 -9087 15270 -8953
rect 15000 -9113 15122 -9087
rect 15148 -9113 15270 -9087
rect 15000 -9230 15270 -9113
rect 18730 -5887 19000 -5770
rect 18730 -5913 18855 -5887
rect 18881 -5913 19000 -5887
rect 18730 -6047 19000 -5913
rect 18730 -6073 18855 -6047
rect 18881 -6073 19000 -6047
rect 18730 -6207 19000 -6073
rect 18730 -6233 18855 -6207
rect 18881 -6233 19000 -6207
rect 18730 -6367 19000 -6233
rect 18730 -6393 18855 -6367
rect 18881 -6393 19000 -6367
rect 18730 -6527 19000 -6393
rect 18730 -6553 18855 -6527
rect 18881 -6553 19000 -6527
rect 18730 -6687 19000 -6553
rect 18730 -6713 18855 -6687
rect 18881 -6713 19000 -6687
rect 18730 -6847 19000 -6713
rect 18730 -6873 18855 -6847
rect 18881 -6873 19000 -6847
rect 18730 -7007 19000 -6873
rect 18730 -7033 18855 -7007
rect 18881 -7033 19000 -7007
rect 18730 -7167 19000 -7033
rect 18730 -7193 18855 -7167
rect 18881 -7193 19000 -7167
rect 18730 -7327 19000 -7193
rect 18730 -7353 18855 -7327
rect 18881 -7353 19000 -7327
rect 18730 -7487 19000 -7353
rect 18730 -7513 18855 -7487
rect 18881 -7513 19000 -7487
rect 18730 -7647 19000 -7513
rect 18730 -7673 18855 -7647
rect 18881 -7673 19000 -7647
rect 18730 -7807 19000 -7673
rect 18730 -7833 18855 -7807
rect 18881 -7833 19000 -7807
rect 18730 -7967 19000 -7833
rect 18730 -7993 18855 -7967
rect 18881 -7993 19000 -7967
rect 18730 -8127 19000 -7993
rect 18730 -8153 18855 -8127
rect 18881 -8153 19000 -8127
rect 18730 -8287 19000 -8153
rect 18730 -8313 18855 -8287
rect 18881 -8313 19000 -8287
rect 18730 -8447 19000 -8313
rect 18730 -8473 18855 -8447
rect 18881 -8473 19000 -8447
rect 18730 -8607 19000 -8473
rect 18730 -8633 18855 -8607
rect 18881 -8633 19000 -8607
rect 18730 -8767 19000 -8633
rect 18730 -8793 18855 -8767
rect 18881 -8793 19000 -8767
rect 18730 -8927 19000 -8793
rect 18730 -8953 18855 -8927
rect 18881 -8953 19000 -8927
rect 18730 -9087 19000 -8953
rect 18730 -9113 18855 -9087
rect 18881 -9113 19000 -9087
rect 18730 -9230 19000 -9113
rect 15000 -9247 19000 -9230
rect 15000 -9273 15122 -9247
rect 15148 -9273 18855 -9247
rect 18881 -9273 19000 -9247
rect 15000 -9352 19000 -9273
rect 15000 -9378 15307 -9352
rect 15333 -9378 15467 -9352
rect 15493 -9378 15627 -9352
rect 15653 -9378 15787 -9352
rect 15813 -9378 15947 -9352
rect 15973 -9378 16107 -9352
rect 16133 -9378 16267 -9352
rect 16293 -9378 16427 -9352
rect 16453 -9378 16587 -9352
rect 16613 -9378 16747 -9352
rect 16773 -9378 16907 -9352
rect 16933 -9378 17067 -9352
rect 17093 -9378 17227 -9352
rect 17253 -9378 17387 -9352
rect 17413 -9378 17547 -9352
rect 17573 -9378 17707 -9352
rect 17733 -9378 17867 -9352
rect 17893 -9378 18027 -9352
rect 18053 -9378 18187 -9352
rect 18213 -9378 18347 -9352
rect 18373 -9378 18507 -9352
rect 18533 -9378 18667 -9352
rect 18693 -9378 19000 -9352
rect 15000 -9500 19000 -9378
rect 21000 -5624 25000 -5500
rect 21000 -5650 21307 -5624
rect 21333 -5650 21467 -5624
rect 21493 -5650 21627 -5624
rect 21653 -5650 21787 -5624
rect 21813 -5650 21947 -5624
rect 21973 -5650 22107 -5624
rect 22133 -5650 22267 -5624
rect 22293 -5650 22427 -5624
rect 22453 -5650 22587 -5624
rect 22613 -5650 22747 -5624
rect 22773 -5650 22907 -5624
rect 22933 -5650 23067 -5624
rect 23093 -5650 23227 -5624
rect 23253 -5650 23387 -5624
rect 23413 -5650 23547 -5624
rect 23573 -5650 23707 -5624
rect 23733 -5650 23867 -5624
rect 23893 -5650 24027 -5624
rect 24053 -5650 24187 -5624
rect 24213 -5650 24347 -5624
rect 24373 -5650 24507 -5624
rect 24533 -5650 24667 -5624
rect 24693 -5650 25000 -5624
rect 21000 -5727 25000 -5650
rect 21000 -5753 21122 -5727
rect 21148 -5753 24855 -5727
rect 24881 -5753 25000 -5727
rect 21000 -5770 25000 -5753
rect 21000 -5887 21270 -5770
rect 21000 -5913 21122 -5887
rect 21148 -5913 21270 -5887
rect 21000 -6047 21270 -5913
rect 21000 -6073 21122 -6047
rect 21148 -6073 21270 -6047
rect 21000 -6207 21270 -6073
rect 21000 -6233 21122 -6207
rect 21148 -6233 21270 -6207
rect 21000 -6367 21270 -6233
rect 21000 -6393 21122 -6367
rect 21148 -6393 21270 -6367
rect 21000 -6527 21270 -6393
rect 21000 -6553 21122 -6527
rect 21148 -6553 21270 -6527
rect 21000 -6687 21270 -6553
rect 21000 -6713 21122 -6687
rect 21148 -6713 21270 -6687
rect 21000 -6847 21270 -6713
rect 21000 -6873 21122 -6847
rect 21148 -6873 21270 -6847
rect 21000 -7007 21270 -6873
rect 21000 -7033 21122 -7007
rect 21148 -7033 21270 -7007
rect 21000 -7167 21270 -7033
rect 21000 -7193 21122 -7167
rect 21148 -7193 21270 -7167
rect 21000 -7327 21270 -7193
rect 21000 -7353 21122 -7327
rect 21148 -7353 21270 -7327
rect 21000 -7487 21270 -7353
rect 21000 -7513 21122 -7487
rect 21148 -7513 21270 -7487
rect 21000 -7647 21270 -7513
rect 21000 -7673 21122 -7647
rect 21148 -7673 21270 -7647
rect 21000 -7807 21270 -7673
rect 21000 -7833 21122 -7807
rect 21148 -7833 21270 -7807
rect 21000 -7967 21270 -7833
rect 21000 -7993 21122 -7967
rect 21148 -7993 21270 -7967
rect 21000 -8127 21270 -7993
rect 21000 -8153 21122 -8127
rect 21148 -8153 21270 -8127
rect 21000 -8287 21270 -8153
rect 21000 -8313 21122 -8287
rect 21148 -8313 21270 -8287
rect 21000 -8447 21270 -8313
rect 21000 -8473 21122 -8447
rect 21148 -8473 21270 -8447
rect 21000 -8607 21270 -8473
rect 21000 -8633 21122 -8607
rect 21148 -8633 21270 -8607
rect 21000 -8767 21270 -8633
rect 21000 -8793 21122 -8767
rect 21148 -8793 21270 -8767
rect 21000 -8927 21270 -8793
rect 21000 -8953 21122 -8927
rect 21148 -8953 21270 -8927
rect 21000 -9087 21270 -8953
rect 21000 -9113 21122 -9087
rect 21148 -9113 21270 -9087
rect 21000 -9230 21270 -9113
rect 24730 -5887 25000 -5770
rect 24730 -5913 24855 -5887
rect 24881 -5913 25000 -5887
rect 24730 -6047 25000 -5913
rect 24730 -6073 24855 -6047
rect 24881 -6073 25000 -6047
rect 24730 -6207 25000 -6073
rect 24730 -6233 24855 -6207
rect 24881 -6233 25000 -6207
rect 24730 -6367 25000 -6233
rect 24730 -6393 24855 -6367
rect 24881 -6393 25000 -6367
rect 24730 -6527 25000 -6393
rect 24730 -6553 24855 -6527
rect 24881 -6553 25000 -6527
rect 24730 -6687 25000 -6553
rect 24730 -6713 24855 -6687
rect 24881 -6713 25000 -6687
rect 24730 -6847 25000 -6713
rect 24730 -6873 24855 -6847
rect 24881 -6873 25000 -6847
rect 24730 -7007 25000 -6873
rect 24730 -7033 24855 -7007
rect 24881 -7033 25000 -7007
rect 24730 -7167 25000 -7033
rect 24730 -7193 24855 -7167
rect 24881 -7193 25000 -7167
rect 24730 -7327 25000 -7193
rect 24730 -7353 24855 -7327
rect 24881 -7353 25000 -7327
rect 24730 -7487 25000 -7353
rect 24730 -7513 24855 -7487
rect 24881 -7513 25000 -7487
rect 24730 -7647 25000 -7513
rect 24730 -7673 24855 -7647
rect 24881 -7673 25000 -7647
rect 24730 -7807 25000 -7673
rect 24730 -7833 24855 -7807
rect 24881 -7833 25000 -7807
rect 24730 -7967 25000 -7833
rect 24730 -7993 24855 -7967
rect 24881 -7993 25000 -7967
rect 24730 -8127 25000 -7993
rect 24730 -8153 24855 -8127
rect 24881 -8153 25000 -8127
rect 24730 -8287 25000 -8153
rect 24730 -8313 24855 -8287
rect 24881 -8313 25000 -8287
rect 24730 -8447 25000 -8313
rect 24730 -8473 24855 -8447
rect 24881 -8473 25000 -8447
rect 24730 -8607 25000 -8473
rect 24730 -8633 24855 -8607
rect 24881 -8633 25000 -8607
rect 24730 -8767 25000 -8633
rect 24730 -8793 24855 -8767
rect 24881 -8793 25000 -8767
rect 24730 -8927 25000 -8793
rect 24730 -8953 24855 -8927
rect 24881 -8953 25000 -8927
rect 24730 -9087 25000 -8953
rect 24730 -9113 24855 -9087
rect 24881 -9113 25000 -9087
rect 24730 -9230 25000 -9113
rect 21000 -9247 25000 -9230
rect 21000 -9273 21122 -9247
rect 21148 -9273 24855 -9247
rect 24881 -9273 25000 -9247
rect 21000 -9352 25000 -9273
rect 21000 -9378 21307 -9352
rect 21333 -9378 21467 -9352
rect 21493 -9378 21627 -9352
rect 21653 -9378 21787 -9352
rect 21813 -9378 21947 -9352
rect 21973 -9378 22107 -9352
rect 22133 -9378 22267 -9352
rect 22293 -9378 22427 -9352
rect 22453 -9378 22587 -9352
rect 22613 -9378 22747 -9352
rect 22773 -9378 22907 -9352
rect 22933 -9378 23067 -9352
rect 23093 -9378 23227 -9352
rect 23253 -9378 23387 -9352
rect 23413 -9378 23547 -9352
rect 23573 -9378 23707 -9352
rect 23733 -9378 23867 -9352
rect 23893 -9378 24027 -9352
rect 24053 -9378 24187 -9352
rect 24213 -9378 24347 -9352
rect 24373 -9378 24507 -9352
rect 24533 -9378 24667 -9352
rect 24693 -9378 25000 -9352
rect 21000 -9500 25000 -9378
rect 3000 -11624 7000 -11500
rect 3000 -11650 3307 -11624
rect 3333 -11650 3467 -11624
rect 3493 -11650 3627 -11624
rect 3653 -11650 3787 -11624
rect 3813 -11650 3947 -11624
rect 3973 -11650 4107 -11624
rect 4133 -11650 4267 -11624
rect 4293 -11650 4427 -11624
rect 4453 -11650 4587 -11624
rect 4613 -11650 4747 -11624
rect 4773 -11650 4907 -11624
rect 4933 -11650 5067 -11624
rect 5093 -11650 5227 -11624
rect 5253 -11650 5387 -11624
rect 5413 -11650 5547 -11624
rect 5573 -11650 5707 -11624
rect 5733 -11650 5867 -11624
rect 5893 -11650 6027 -11624
rect 6053 -11650 6187 -11624
rect 6213 -11650 6347 -11624
rect 6373 -11650 6507 -11624
rect 6533 -11650 6667 -11624
rect 6693 -11650 7000 -11624
rect 3000 -11727 7000 -11650
rect 3000 -11753 3122 -11727
rect 3148 -11753 6855 -11727
rect 6881 -11753 7000 -11727
rect 3000 -11770 7000 -11753
rect 3000 -11887 3270 -11770
rect 3000 -11913 3122 -11887
rect 3148 -11913 3270 -11887
rect 3000 -12047 3270 -11913
rect 3000 -12073 3122 -12047
rect 3148 -12073 3270 -12047
rect 3000 -12207 3270 -12073
rect 3000 -12233 3122 -12207
rect 3148 -12233 3270 -12207
rect 3000 -12367 3270 -12233
rect 3000 -12393 3122 -12367
rect 3148 -12393 3270 -12367
rect 3000 -12527 3270 -12393
rect 3000 -12553 3122 -12527
rect 3148 -12553 3270 -12527
rect 3000 -12687 3270 -12553
rect 3000 -12713 3122 -12687
rect 3148 -12713 3270 -12687
rect 3000 -12847 3270 -12713
rect 3000 -12873 3122 -12847
rect 3148 -12873 3270 -12847
rect 3000 -13007 3270 -12873
rect 3000 -13033 3122 -13007
rect 3148 -13033 3270 -13007
rect 3000 -13167 3270 -13033
rect 3000 -13193 3122 -13167
rect 3148 -13193 3270 -13167
rect 3000 -13327 3270 -13193
rect 3000 -13353 3122 -13327
rect 3148 -13353 3270 -13327
rect 3000 -13487 3270 -13353
rect 3000 -13513 3122 -13487
rect 3148 -13513 3270 -13487
rect 3000 -13647 3270 -13513
rect 3000 -13673 3122 -13647
rect 3148 -13673 3270 -13647
rect 3000 -13807 3270 -13673
rect 3000 -13833 3122 -13807
rect 3148 -13833 3270 -13807
rect 3000 -13967 3270 -13833
rect 3000 -13993 3122 -13967
rect 3148 -13993 3270 -13967
rect 3000 -14127 3270 -13993
rect 3000 -14153 3122 -14127
rect 3148 -14153 3270 -14127
rect 3000 -14287 3270 -14153
rect 3000 -14313 3122 -14287
rect 3148 -14313 3270 -14287
rect 3000 -14447 3270 -14313
rect 3000 -14473 3122 -14447
rect 3148 -14473 3270 -14447
rect 3000 -14607 3270 -14473
rect 3000 -14633 3122 -14607
rect 3148 -14633 3270 -14607
rect 3000 -14767 3270 -14633
rect 3000 -14793 3122 -14767
rect 3148 -14793 3270 -14767
rect 3000 -14927 3270 -14793
rect 3000 -14953 3122 -14927
rect 3148 -14953 3270 -14927
rect 3000 -15087 3270 -14953
rect 3000 -15113 3122 -15087
rect 3148 -15113 3270 -15087
rect 3000 -15230 3270 -15113
rect 6730 -11887 7000 -11770
rect 6730 -11913 6855 -11887
rect 6881 -11913 7000 -11887
rect 6730 -12047 7000 -11913
rect 6730 -12073 6855 -12047
rect 6881 -12073 7000 -12047
rect 6730 -12207 7000 -12073
rect 6730 -12233 6855 -12207
rect 6881 -12233 7000 -12207
rect 6730 -12367 7000 -12233
rect 6730 -12393 6855 -12367
rect 6881 -12393 7000 -12367
rect 6730 -12527 7000 -12393
rect 6730 -12553 6855 -12527
rect 6881 -12553 7000 -12527
rect 6730 -12687 7000 -12553
rect 6730 -12713 6855 -12687
rect 6881 -12713 7000 -12687
rect 6730 -12847 7000 -12713
rect 6730 -12873 6855 -12847
rect 6881 -12873 7000 -12847
rect 6730 -13007 7000 -12873
rect 6730 -13033 6855 -13007
rect 6881 -13033 7000 -13007
rect 6730 -13167 7000 -13033
rect 6730 -13193 6855 -13167
rect 6881 -13193 7000 -13167
rect 6730 -13327 7000 -13193
rect 6730 -13353 6855 -13327
rect 6881 -13353 7000 -13327
rect 6730 -13487 7000 -13353
rect 6730 -13513 6855 -13487
rect 6881 -13513 7000 -13487
rect 6730 -13647 7000 -13513
rect 6730 -13673 6855 -13647
rect 6881 -13673 7000 -13647
rect 6730 -13807 7000 -13673
rect 6730 -13833 6855 -13807
rect 6881 -13833 7000 -13807
rect 6730 -13967 7000 -13833
rect 6730 -13993 6855 -13967
rect 6881 -13993 7000 -13967
rect 6730 -14127 7000 -13993
rect 6730 -14153 6855 -14127
rect 6881 -14153 7000 -14127
rect 6730 -14287 7000 -14153
rect 6730 -14313 6855 -14287
rect 6881 -14313 7000 -14287
rect 6730 -14447 7000 -14313
rect 6730 -14473 6855 -14447
rect 6881 -14473 7000 -14447
rect 6730 -14607 7000 -14473
rect 6730 -14633 6855 -14607
rect 6881 -14633 7000 -14607
rect 6730 -14767 7000 -14633
rect 6730 -14793 6855 -14767
rect 6881 -14793 7000 -14767
rect 6730 -14927 7000 -14793
rect 6730 -14953 6855 -14927
rect 6881 -14953 7000 -14927
rect 6730 -15087 7000 -14953
rect 6730 -15113 6855 -15087
rect 6881 -15113 7000 -15087
rect 6730 -15230 7000 -15113
rect 3000 -15247 7000 -15230
rect 3000 -15273 3122 -15247
rect 3148 -15273 6855 -15247
rect 6881 -15273 7000 -15247
rect 3000 -15352 7000 -15273
rect 3000 -15378 3307 -15352
rect 3333 -15378 3467 -15352
rect 3493 -15378 3627 -15352
rect 3653 -15378 3787 -15352
rect 3813 -15378 3947 -15352
rect 3973 -15378 4107 -15352
rect 4133 -15378 4267 -15352
rect 4293 -15378 4427 -15352
rect 4453 -15378 4587 -15352
rect 4613 -15378 4747 -15352
rect 4773 -15378 4907 -15352
rect 4933 -15378 5067 -15352
rect 5093 -15378 5227 -15352
rect 5253 -15378 5387 -15352
rect 5413 -15378 5547 -15352
rect 5573 -15378 5707 -15352
rect 5733 -15378 5867 -15352
rect 5893 -15378 6027 -15352
rect 6053 -15378 6187 -15352
rect 6213 -15378 6347 -15352
rect 6373 -15378 6507 -15352
rect 6533 -15378 6667 -15352
rect 6693 -15378 7000 -15352
rect 3000 -15500 7000 -15378
rect 9000 -11624 13000 -11500
rect 9000 -11650 9307 -11624
rect 9333 -11650 9467 -11624
rect 9493 -11650 9627 -11624
rect 9653 -11650 9787 -11624
rect 9813 -11650 9947 -11624
rect 9973 -11650 10107 -11624
rect 10133 -11650 10267 -11624
rect 10293 -11650 10427 -11624
rect 10453 -11650 10587 -11624
rect 10613 -11650 10747 -11624
rect 10773 -11650 10907 -11624
rect 10933 -11650 11067 -11624
rect 11093 -11650 11227 -11624
rect 11253 -11650 11387 -11624
rect 11413 -11650 11547 -11624
rect 11573 -11650 11707 -11624
rect 11733 -11650 11867 -11624
rect 11893 -11650 12027 -11624
rect 12053 -11650 12187 -11624
rect 12213 -11650 12347 -11624
rect 12373 -11650 12507 -11624
rect 12533 -11650 12667 -11624
rect 12693 -11650 13000 -11624
rect 9000 -11727 13000 -11650
rect 9000 -11753 9122 -11727
rect 9148 -11753 12855 -11727
rect 12881 -11753 13000 -11727
rect 9000 -11770 13000 -11753
rect 9000 -11887 9270 -11770
rect 9000 -11913 9122 -11887
rect 9148 -11913 9270 -11887
rect 9000 -12047 9270 -11913
rect 9000 -12073 9122 -12047
rect 9148 -12073 9270 -12047
rect 9000 -12207 9270 -12073
rect 9000 -12233 9122 -12207
rect 9148 -12233 9270 -12207
rect 9000 -12367 9270 -12233
rect 9000 -12393 9122 -12367
rect 9148 -12393 9270 -12367
rect 9000 -12527 9270 -12393
rect 9000 -12553 9122 -12527
rect 9148 -12553 9270 -12527
rect 9000 -12687 9270 -12553
rect 9000 -12713 9122 -12687
rect 9148 -12713 9270 -12687
rect 9000 -12847 9270 -12713
rect 9000 -12873 9122 -12847
rect 9148 -12873 9270 -12847
rect 9000 -13007 9270 -12873
rect 9000 -13033 9122 -13007
rect 9148 -13033 9270 -13007
rect 9000 -13167 9270 -13033
rect 9000 -13193 9122 -13167
rect 9148 -13193 9270 -13167
rect 9000 -13327 9270 -13193
rect 9000 -13353 9122 -13327
rect 9148 -13353 9270 -13327
rect 9000 -13487 9270 -13353
rect 9000 -13513 9122 -13487
rect 9148 -13513 9270 -13487
rect 9000 -13647 9270 -13513
rect 9000 -13673 9122 -13647
rect 9148 -13673 9270 -13647
rect 9000 -13807 9270 -13673
rect 9000 -13833 9122 -13807
rect 9148 -13833 9270 -13807
rect 9000 -13967 9270 -13833
rect 9000 -13993 9122 -13967
rect 9148 -13993 9270 -13967
rect 9000 -14127 9270 -13993
rect 9000 -14153 9122 -14127
rect 9148 -14153 9270 -14127
rect 9000 -14287 9270 -14153
rect 9000 -14313 9122 -14287
rect 9148 -14313 9270 -14287
rect 9000 -14447 9270 -14313
rect 9000 -14473 9122 -14447
rect 9148 -14473 9270 -14447
rect 9000 -14607 9270 -14473
rect 9000 -14633 9122 -14607
rect 9148 -14633 9270 -14607
rect 9000 -14767 9270 -14633
rect 9000 -14793 9122 -14767
rect 9148 -14793 9270 -14767
rect 9000 -14927 9270 -14793
rect 9000 -14953 9122 -14927
rect 9148 -14953 9270 -14927
rect 9000 -15087 9270 -14953
rect 9000 -15113 9122 -15087
rect 9148 -15113 9270 -15087
rect 9000 -15230 9270 -15113
rect 12730 -11887 13000 -11770
rect 12730 -11913 12855 -11887
rect 12881 -11913 13000 -11887
rect 12730 -12047 13000 -11913
rect 12730 -12073 12855 -12047
rect 12881 -12073 13000 -12047
rect 12730 -12207 13000 -12073
rect 12730 -12233 12855 -12207
rect 12881 -12233 13000 -12207
rect 12730 -12367 13000 -12233
rect 12730 -12393 12855 -12367
rect 12881 -12393 13000 -12367
rect 12730 -12527 13000 -12393
rect 12730 -12553 12855 -12527
rect 12881 -12553 13000 -12527
rect 12730 -12687 13000 -12553
rect 12730 -12713 12855 -12687
rect 12881 -12713 13000 -12687
rect 12730 -12847 13000 -12713
rect 12730 -12873 12855 -12847
rect 12881 -12873 13000 -12847
rect 12730 -13007 13000 -12873
rect 12730 -13033 12855 -13007
rect 12881 -13033 13000 -13007
rect 12730 -13167 13000 -13033
rect 12730 -13193 12855 -13167
rect 12881 -13193 13000 -13167
rect 12730 -13327 13000 -13193
rect 12730 -13353 12855 -13327
rect 12881 -13353 13000 -13327
rect 12730 -13487 13000 -13353
rect 12730 -13513 12855 -13487
rect 12881 -13513 13000 -13487
rect 12730 -13647 13000 -13513
rect 12730 -13673 12855 -13647
rect 12881 -13673 13000 -13647
rect 12730 -13807 13000 -13673
rect 12730 -13833 12855 -13807
rect 12881 -13833 13000 -13807
rect 12730 -13967 13000 -13833
rect 12730 -13993 12855 -13967
rect 12881 -13993 13000 -13967
rect 12730 -14127 13000 -13993
rect 12730 -14153 12855 -14127
rect 12881 -14153 13000 -14127
rect 12730 -14287 13000 -14153
rect 12730 -14313 12855 -14287
rect 12881 -14313 13000 -14287
rect 12730 -14447 13000 -14313
rect 12730 -14473 12855 -14447
rect 12881 -14473 13000 -14447
rect 12730 -14607 13000 -14473
rect 12730 -14633 12855 -14607
rect 12881 -14633 13000 -14607
rect 12730 -14767 13000 -14633
rect 12730 -14793 12855 -14767
rect 12881 -14793 13000 -14767
rect 12730 -14927 13000 -14793
rect 12730 -14953 12855 -14927
rect 12881 -14953 13000 -14927
rect 12730 -15087 13000 -14953
rect 12730 -15113 12855 -15087
rect 12881 -15113 13000 -15087
rect 12730 -15230 13000 -15113
rect 9000 -15247 13000 -15230
rect 9000 -15273 9122 -15247
rect 9148 -15273 12855 -15247
rect 12881 -15273 13000 -15247
rect 9000 -15352 13000 -15273
rect 9000 -15378 9307 -15352
rect 9333 -15378 9467 -15352
rect 9493 -15378 9627 -15352
rect 9653 -15378 9787 -15352
rect 9813 -15378 9947 -15352
rect 9973 -15378 10107 -15352
rect 10133 -15378 10267 -15352
rect 10293 -15378 10427 -15352
rect 10453 -15378 10587 -15352
rect 10613 -15378 10747 -15352
rect 10773 -15378 10907 -15352
rect 10933 -15378 11067 -15352
rect 11093 -15378 11227 -15352
rect 11253 -15378 11387 -15352
rect 11413 -15378 11547 -15352
rect 11573 -15378 11707 -15352
rect 11733 -15378 11867 -15352
rect 11893 -15378 12027 -15352
rect 12053 -15378 12187 -15352
rect 12213 -15378 12347 -15352
rect 12373 -15378 12507 -15352
rect 12533 -15378 12667 -15352
rect 12693 -15378 13000 -15352
rect 9000 -15500 13000 -15378
rect 15000 -11624 19000 -11500
rect 15000 -11650 15307 -11624
rect 15333 -11650 15467 -11624
rect 15493 -11650 15627 -11624
rect 15653 -11650 15787 -11624
rect 15813 -11650 15947 -11624
rect 15973 -11650 16107 -11624
rect 16133 -11650 16267 -11624
rect 16293 -11650 16427 -11624
rect 16453 -11650 16587 -11624
rect 16613 -11650 16747 -11624
rect 16773 -11650 16907 -11624
rect 16933 -11650 17067 -11624
rect 17093 -11650 17227 -11624
rect 17253 -11650 17387 -11624
rect 17413 -11650 17547 -11624
rect 17573 -11650 17707 -11624
rect 17733 -11650 17867 -11624
rect 17893 -11650 18027 -11624
rect 18053 -11650 18187 -11624
rect 18213 -11650 18347 -11624
rect 18373 -11650 18507 -11624
rect 18533 -11650 18667 -11624
rect 18693 -11650 19000 -11624
rect 15000 -11727 19000 -11650
rect 15000 -11753 15122 -11727
rect 15148 -11753 18855 -11727
rect 18881 -11753 19000 -11727
rect 15000 -11770 19000 -11753
rect 15000 -11887 15270 -11770
rect 15000 -11913 15122 -11887
rect 15148 -11913 15270 -11887
rect 15000 -12047 15270 -11913
rect 15000 -12073 15122 -12047
rect 15148 -12073 15270 -12047
rect 15000 -12207 15270 -12073
rect 15000 -12233 15122 -12207
rect 15148 -12233 15270 -12207
rect 15000 -12367 15270 -12233
rect 15000 -12393 15122 -12367
rect 15148 -12393 15270 -12367
rect 15000 -12527 15270 -12393
rect 15000 -12553 15122 -12527
rect 15148 -12553 15270 -12527
rect 15000 -12687 15270 -12553
rect 15000 -12713 15122 -12687
rect 15148 -12713 15270 -12687
rect 15000 -12847 15270 -12713
rect 15000 -12873 15122 -12847
rect 15148 -12873 15270 -12847
rect 15000 -13007 15270 -12873
rect 15000 -13033 15122 -13007
rect 15148 -13033 15270 -13007
rect 15000 -13167 15270 -13033
rect 15000 -13193 15122 -13167
rect 15148 -13193 15270 -13167
rect 15000 -13327 15270 -13193
rect 15000 -13353 15122 -13327
rect 15148 -13353 15270 -13327
rect 15000 -13487 15270 -13353
rect 15000 -13513 15122 -13487
rect 15148 -13513 15270 -13487
rect 15000 -13647 15270 -13513
rect 15000 -13673 15122 -13647
rect 15148 -13673 15270 -13647
rect 15000 -13807 15270 -13673
rect 15000 -13833 15122 -13807
rect 15148 -13833 15270 -13807
rect 15000 -13967 15270 -13833
rect 15000 -13993 15122 -13967
rect 15148 -13993 15270 -13967
rect 15000 -14127 15270 -13993
rect 15000 -14153 15122 -14127
rect 15148 -14153 15270 -14127
rect 15000 -14287 15270 -14153
rect 15000 -14313 15122 -14287
rect 15148 -14313 15270 -14287
rect 15000 -14447 15270 -14313
rect 15000 -14473 15122 -14447
rect 15148 -14473 15270 -14447
rect 15000 -14607 15270 -14473
rect 15000 -14633 15122 -14607
rect 15148 -14633 15270 -14607
rect 15000 -14767 15270 -14633
rect 15000 -14793 15122 -14767
rect 15148 -14793 15270 -14767
rect 15000 -14927 15270 -14793
rect 15000 -14953 15122 -14927
rect 15148 -14953 15270 -14927
rect 15000 -15087 15270 -14953
rect 15000 -15113 15122 -15087
rect 15148 -15113 15270 -15087
rect 15000 -15230 15270 -15113
rect 18730 -11887 19000 -11770
rect 18730 -11913 18855 -11887
rect 18881 -11913 19000 -11887
rect 18730 -12047 19000 -11913
rect 18730 -12073 18855 -12047
rect 18881 -12073 19000 -12047
rect 18730 -12207 19000 -12073
rect 18730 -12233 18855 -12207
rect 18881 -12233 19000 -12207
rect 18730 -12367 19000 -12233
rect 18730 -12393 18855 -12367
rect 18881 -12393 19000 -12367
rect 18730 -12527 19000 -12393
rect 18730 -12553 18855 -12527
rect 18881 -12553 19000 -12527
rect 18730 -12687 19000 -12553
rect 18730 -12713 18855 -12687
rect 18881 -12713 19000 -12687
rect 18730 -12847 19000 -12713
rect 18730 -12873 18855 -12847
rect 18881 -12873 19000 -12847
rect 18730 -13007 19000 -12873
rect 18730 -13033 18855 -13007
rect 18881 -13033 19000 -13007
rect 18730 -13167 19000 -13033
rect 18730 -13193 18855 -13167
rect 18881 -13193 19000 -13167
rect 18730 -13327 19000 -13193
rect 18730 -13353 18855 -13327
rect 18881 -13353 19000 -13327
rect 18730 -13487 19000 -13353
rect 18730 -13513 18855 -13487
rect 18881 -13513 19000 -13487
rect 18730 -13647 19000 -13513
rect 18730 -13673 18855 -13647
rect 18881 -13673 19000 -13647
rect 18730 -13807 19000 -13673
rect 18730 -13833 18855 -13807
rect 18881 -13833 19000 -13807
rect 18730 -13967 19000 -13833
rect 18730 -13993 18855 -13967
rect 18881 -13993 19000 -13967
rect 18730 -14127 19000 -13993
rect 18730 -14153 18855 -14127
rect 18881 -14153 19000 -14127
rect 18730 -14287 19000 -14153
rect 18730 -14313 18855 -14287
rect 18881 -14313 19000 -14287
rect 18730 -14447 19000 -14313
rect 18730 -14473 18855 -14447
rect 18881 -14473 19000 -14447
rect 18730 -14607 19000 -14473
rect 18730 -14633 18855 -14607
rect 18881 -14633 19000 -14607
rect 18730 -14767 19000 -14633
rect 18730 -14793 18855 -14767
rect 18881 -14793 19000 -14767
rect 18730 -14927 19000 -14793
rect 18730 -14953 18855 -14927
rect 18881 -14953 19000 -14927
rect 18730 -15087 19000 -14953
rect 18730 -15113 18855 -15087
rect 18881 -15113 19000 -15087
rect 18730 -15230 19000 -15113
rect 15000 -15247 19000 -15230
rect 15000 -15273 15122 -15247
rect 15148 -15273 18855 -15247
rect 18881 -15273 19000 -15247
rect 15000 -15352 19000 -15273
rect 15000 -15378 15307 -15352
rect 15333 -15378 15467 -15352
rect 15493 -15378 15627 -15352
rect 15653 -15378 15787 -15352
rect 15813 -15378 15947 -15352
rect 15973 -15378 16107 -15352
rect 16133 -15378 16267 -15352
rect 16293 -15378 16427 -15352
rect 16453 -15378 16587 -15352
rect 16613 -15378 16747 -15352
rect 16773 -15378 16907 -15352
rect 16933 -15378 17067 -15352
rect 17093 -15378 17227 -15352
rect 17253 -15378 17387 -15352
rect 17413 -15378 17547 -15352
rect 17573 -15378 17707 -15352
rect 17733 -15378 17867 -15352
rect 17893 -15378 18027 -15352
rect 18053 -15378 18187 -15352
rect 18213 -15378 18347 -15352
rect 18373 -15378 18507 -15352
rect 18533 -15378 18667 -15352
rect 18693 -15378 19000 -15352
rect 15000 -15500 19000 -15378
rect 21000 -11624 25000 -11500
rect 21000 -11650 21307 -11624
rect 21333 -11650 21467 -11624
rect 21493 -11650 21627 -11624
rect 21653 -11650 21787 -11624
rect 21813 -11650 21947 -11624
rect 21973 -11650 22107 -11624
rect 22133 -11650 22267 -11624
rect 22293 -11650 22427 -11624
rect 22453 -11650 22587 -11624
rect 22613 -11650 22747 -11624
rect 22773 -11650 22907 -11624
rect 22933 -11650 23067 -11624
rect 23093 -11650 23227 -11624
rect 23253 -11650 23387 -11624
rect 23413 -11650 23547 -11624
rect 23573 -11650 23707 -11624
rect 23733 -11650 23867 -11624
rect 23893 -11650 24027 -11624
rect 24053 -11650 24187 -11624
rect 24213 -11650 24347 -11624
rect 24373 -11650 24507 -11624
rect 24533 -11650 24667 -11624
rect 24693 -11650 25000 -11624
rect 21000 -11727 25000 -11650
rect 21000 -11753 21122 -11727
rect 21148 -11753 24855 -11727
rect 24881 -11753 25000 -11727
rect 21000 -11770 25000 -11753
rect 21000 -11887 21270 -11770
rect 21000 -11913 21122 -11887
rect 21148 -11913 21270 -11887
rect 21000 -12047 21270 -11913
rect 21000 -12073 21122 -12047
rect 21148 -12073 21270 -12047
rect 21000 -12207 21270 -12073
rect 21000 -12233 21122 -12207
rect 21148 -12233 21270 -12207
rect 21000 -12367 21270 -12233
rect 21000 -12393 21122 -12367
rect 21148 -12393 21270 -12367
rect 21000 -12527 21270 -12393
rect 21000 -12553 21122 -12527
rect 21148 -12553 21270 -12527
rect 21000 -12687 21270 -12553
rect 21000 -12713 21122 -12687
rect 21148 -12713 21270 -12687
rect 21000 -12847 21270 -12713
rect 21000 -12873 21122 -12847
rect 21148 -12873 21270 -12847
rect 21000 -13007 21270 -12873
rect 21000 -13033 21122 -13007
rect 21148 -13033 21270 -13007
rect 21000 -13167 21270 -13033
rect 21000 -13193 21122 -13167
rect 21148 -13193 21270 -13167
rect 21000 -13327 21270 -13193
rect 21000 -13353 21122 -13327
rect 21148 -13353 21270 -13327
rect 21000 -13487 21270 -13353
rect 21000 -13513 21122 -13487
rect 21148 -13513 21270 -13487
rect 21000 -13647 21270 -13513
rect 21000 -13673 21122 -13647
rect 21148 -13673 21270 -13647
rect 21000 -13807 21270 -13673
rect 21000 -13833 21122 -13807
rect 21148 -13833 21270 -13807
rect 21000 -13967 21270 -13833
rect 21000 -13993 21122 -13967
rect 21148 -13993 21270 -13967
rect 21000 -14127 21270 -13993
rect 21000 -14153 21122 -14127
rect 21148 -14153 21270 -14127
rect 21000 -14287 21270 -14153
rect 21000 -14313 21122 -14287
rect 21148 -14313 21270 -14287
rect 21000 -14447 21270 -14313
rect 21000 -14473 21122 -14447
rect 21148 -14473 21270 -14447
rect 21000 -14607 21270 -14473
rect 21000 -14633 21122 -14607
rect 21148 -14633 21270 -14607
rect 21000 -14767 21270 -14633
rect 21000 -14793 21122 -14767
rect 21148 -14793 21270 -14767
rect 21000 -14927 21270 -14793
rect 21000 -14953 21122 -14927
rect 21148 -14953 21270 -14927
rect 21000 -15087 21270 -14953
rect 21000 -15113 21122 -15087
rect 21148 -15113 21270 -15087
rect 21000 -15230 21270 -15113
rect 24730 -11887 25000 -11770
rect 24730 -11913 24855 -11887
rect 24881 -11913 25000 -11887
rect 24730 -12047 25000 -11913
rect 24730 -12073 24855 -12047
rect 24881 -12073 25000 -12047
rect 24730 -12207 25000 -12073
rect 24730 -12233 24855 -12207
rect 24881 -12233 25000 -12207
rect 24730 -12367 25000 -12233
rect 24730 -12393 24855 -12367
rect 24881 -12393 25000 -12367
rect 24730 -12527 25000 -12393
rect 24730 -12553 24855 -12527
rect 24881 -12553 25000 -12527
rect 24730 -12687 25000 -12553
rect 24730 -12713 24855 -12687
rect 24881 -12713 25000 -12687
rect 24730 -12847 25000 -12713
rect 24730 -12873 24855 -12847
rect 24881 -12873 25000 -12847
rect 24730 -13007 25000 -12873
rect 24730 -13033 24855 -13007
rect 24881 -13033 25000 -13007
rect 24730 -13167 25000 -13033
rect 24730 -13193 24855 -13167
rect 24881 -13193 25000 -13167
rect 24730 -13327 25000 -13193
rect 24730 -13353 24855 -13327
rect 24881 -13353 25000 -13327
rect 24730 -13487 25000 -13353
rect 24730 -13513 24855 -13487
rect 24881 -13513 25000 -13487
rect 24730 -13647 25000 -13513
rect 24730 -13673 24855 -13647
rect 24881 -13673 25000 -13647
rect 24730 -13807 25000 -13673
rect 24730 -13833 24855 -13807
rect 24881 -13833 25000 -13807
rect 24730 -13967 25000 -13833
rect 24730 -13993 24855 -13967
rect 24881 -13993 25000 -13967
rect 24730 -14127 25000 -13993
rect 24730 -14153 24855 -14127
rect 24881 -14153 25000 -14127
rect 24730 -14287 25000 -14153
rect 24730 -14313 24855 -14287
rect 24881 -14313 25000 -14287
rect 24730 -14447 25000 -14313
rect 24730 -14473 24855 -14447
rect 24881 -14473 25000 -14447
rect 24730 -14607 25000 -14473
rect 24730 -14633 24855 -14607
rect 24881 -14633 25000 -14607
rect 24730 -14767 25000 -14633
rect 24730 -14793 24855 -14767
rect 24881 -14793 25000 -14767
rect 24730 -14927 25000 -14793
rect 24730 -14953 24855 -14927
rect 24881 -14953 25000 -14927
rect 24730 -15087 25000 -14953
rect 24730 -15113 24855 -15087
rect 24881 -15113 25000 -15087
rect 24730 -15230 25000 -15113
rect 21000 -15247 25000 -15230
rect 21000 -15273 21122 -15247
rect 21148 -15273 24855 -15247
rect 24881 -15273 25000 -15247
rect 21000 -15352 25000 -15273
rect 21000 -15378 21307 -15352
rect 21333 -15378 21467 -15352
rect 21493 -15378 21627 -15352
rect 21653 -15378 21787 -15352
rect 21813 -15378 21947 -15352
rect 21973 -15378 22107 -15352
rect 22133 -15378 22267 -15352
rect 22293 -15378 22427 -15352
rect 22453 -15378 22587 -15352
rect 22613 -15378 22747 -15352
rect 22773 -15378 22907 -15352
rect 22933 -15378 23067 -15352
rect 23093 -15378 23227 -15352
rect 23253 -15378 23387 -15352
rect 23413 -15378 23547 -15352
rect 23573 -15378 23707 -15352
rect 23733 -15378 23867 -15352
rect 23893 -15378 24027 -15352
rect 24053 -15378 24187 -15352
rect 24213 -15378 24347 -15352
rect 24373 -15378 24507 -15352
rect 24533 -15378 24667 -15352
rect 24693 -15378 25000 -15352
rect 21000 -15500 25000 -15378
<< via1 >>
rect 11650 -3700 11750 -3600
rect 11635 -3860 11705 -3820
rect 11775 -3860 11845 -3820
rect 11650 -4050 11750 -3950
rect 8200 -4790 8230 -4760
rect 8235 -4860 8265 -4830
rect 8355 -5425 8400 -5255
rect 8515 -5370 8565 -5310
rect 8710 -5425 8755 -5255
rect 3307 -5650 3333 -5624
rect 3467 -5650 3493 -5624
rect 3627 -5650 3653 -5624
rect 3787 -5650 3813 -5624
rect 3947 -5650 3973 -5624
rect 4107 -5650 4133 -5624
rect 4267 -5650 4293 -5624
rect 4427 -5650 4453 -5624
rect 4587 -5650 4613 -5624
rect 4747 -5650 4773 -5624
rect 4907 -5650 4933 -5624
rect 5067 -5650 5093 -5624
rect 5227 -5650 5253 -5624
rect 5387 -5650 5413 -5624
rect 5547 -5650 5573 -5624
rect 5707 -5650 5733 -5624
rect 5867 -5650 5893 -5624
rect 6027 -5650 6053 -5624
rect 6187 -5650 6213 -5624
rect 6347 -5650 6373 -5624
rect 6507 -5650 6533 -5624
rect 6667 -5650 6693 -5624
rect 3122 -5753 3148 -5727
rect 6855 -5753 6881 -5727
rect 3122 -5913 3148 -5887
rect 3122 -6073 3148 -6047
rect 3122 -6233 3148 -6207
rect 3122 -6393 3148 -6367
rect 3122 -6553 3148 -6527
rect 3122 -6713 3148 -6687
rect 3122 -6873 3148 -6847
rect 3122 -7033 3148 -7007
rect 3122 -7193 3148 -7167
rect 3122 -7353 3148 -7327
rect 3122 -7513 3148 -7487
rect 3122 -7673 3148 -7647
rect 3122 -7833 3148 -7807
rect 3122 -7993 3148 -7967
rect 3122 -8153 3148 -8127
rect 3122 -8313 3148 -8287
rect 3122 -8473 3148 -8447
rect 3122 -8633 3148 -8607
rect 3122 -8793 3148 -8767
rect 3122 -8953 3148 -8927
rect 3122 -9113 3148 -9087
rect 6855 -5913 6881 -5887
rect 6855 -6073 6881 -6047
rect 6855 -6233 6881 -6207
rect 6855 -6393 6881 -6367
rect 6855 -6553 6881 -6527
rect 6855 -6713 6881 -6687
rect 6855 -6873 6881 -6847
rect 6855 -7033 6881 -7007
rect 6855 -7193 6881 -7167
rect 6855 -7353 6881 -7327
rect 6855 -7513 6881 -7487
rect 6855 -7673 6881 -7647
rect 6855 -7833 6881 -7807
rect 6855 -7993 6881 -7967
rect 6855 -8153 6881 -8127
rect 6855 -8313 6881 -8287
rect 6855 -8473 6881 -8447
rect 6855 -8633 6881 -8607
rect 6855 -8793 6881 -8767
rect 6855 -8953 6881 -8927
rect 6855 -9113 6881 -9087
rect 3122 -9273 3148 -9247
rect 6855 -9273 6881 -9247
rect 3307 -9378 3333 -9352
rect 3467 -9378 3493 -9352
rect 3627 -9378 3653 -9352
rect 3787 -9378 3813 -9352
rect 3947 -9378 3973 -9352
rect 4107 -9378 4133 -9352
rect 4267 -9378 4293 -9352
rect 4427 -9378 4453 -9352
rect 4587 -9378 4613 -9352
rect 4747 -9378 4773 -9352
rect 4907 -9378 4933 -9352
rect 5067 -9378 5093 -9352
rect 5227 -9378 5253 -9352
rect 5387 -9378 5413 -9352
rect 5547 -9378 5573 -9352
rect 5707 -9378 5733 -9352
rect 5867 -9378 5893 -9352
rect 6027 -9378 6053 -9352
rect 6187 -9378 6213 -9352
rect 6347 -9378 6373 -9352
rect 6507 -9378 6533 -9352
rect 6667 -9378 6693 -9352
rect 9307 -5650 9333 -5624
rect 9467 -5650 9493 -5624
rect 9627 -5650 9653 -5624
rect 9787 -5650 9813 -5624
rect 9947 -5650 9973 -5624
rect 10107 -5650 10133 -5624
rect 10267 -5650 10293 -5624
rect 10427 -5650 10453 -5624
rect 10587 -5650 10613 -5624
rect 10747 -5650 10773 -5624
rect 10907 -5650 10933 -5624
rect 11067 -5650 11093 -5624
rect 11227 -5650 11253 -5624
rect 11387 -5650 11413 -5624
rect 11547 -5650 11573 -5624
rect 11707 -5650 11733 -5624
rect 11867 -5650 11893 -5624
rect 12027 -5650 12053 -5624
rect 12187 -5650 12213 -5624
rect 12347 -5650 12373 -5624
rect 12507 -5650 12533 -5624
rect 12667 -5650 12693 -5624
rect 9122 -5753 9148 -5727
rect 12855 -5753 12881 -5727
rect 9122 -5913 9148 -5887
rect 9122 -6073 9148 -6047
rect 9122 -6233 9148 -6207
rect 9122 -6393 9148 -6367
rect 9122 -6553 9148 -6527
rect 9122 -6713 9148 -6687
rect 9122 -6873 9148 -6847
rect 9122 -7033 9148 -7007
rect 9122 -7193 9148 -7167
rect 9122 -7353 9148 -7327
rect 9122 -7513 9148 -7487
rect 9122 -7673 9148 -7647
rect 9122 -7833 9148 -7807
rect 9122 -7993 9148 -7967
rect 9122 -8153 9148 -8127
rect 9122 -8313 9148 -8287
rect 9122 -8473 9148 -8447
rect 9122 -8633 9148 -8607
rect 9122 -8793 9148 -8767
rect 9122 -8953 9148 -8927
rect 9122 -9113 9148 -9087
rect 12855 -5913 12881 -5887
rect 12855 -6073 12881 -6047
rect 12855 -6233 12881 -6207
rect 12855 -6393 12881 -6367
rect 12855 -6553 12881 -6527
rect 12855 -6713 12881 -6687
rect 12855 -6873 12881 -6847
rect 12855 -7033 12881 -7007
rect 12855 -7193 12881 -7167
rect 12855 -7353 12881 -7327
rect 12855 -7513 12881 -7487
rect 12855 -7673 12881 -7647
rect 12855 -7833 12881 -7807
rect 12855 -7993 12881 -7967
rect 12855 -8153 12881 -8127
rect 12855 -8313 12881 -8287
rect 12855 -8473 12881 -8447
rect 12855 -8633 12881 -8607
rect 12855 -8793 12881 -8767
rect 12855 -8953 12881 -8927
rect 12855 -9113 12881 -9087
rect 9122 -9273 9148 -9247
rect 12855 -9273 12881 -9247
rect 9307 -9378 9333 -9352
rect 9467 -9378 9493 -9352
rect 9627 -9378 9653 -9352
rect 9787 -9378 9813 -9352
rect 9947 -9378 9973 -9352
rect 10107 -9378 10133 -9352
rect 10267 -9378 10293 -9352
rect 10427 -9378 10453 -9352
rect 10587 -9378 10613 -9352
rect 10747 -9378 10773 -9352
rect 10907 -9378 10933 -9352
rect 11067 -9378 11093 -9352
rect 11227 -9378 11253 -9352
rect 11387 -9378 11413 -9352
rect 11547 -9378 11573 -9352
rect 11707 -9378 11733 -9352
rect 11867 -9378 11893 -9352
rect 12027 -9378 12053 -9352
rect 12187 -9378 12213 -9352
rect 12347 -9378 12373 -9352
rect 12507 -9378 12533 -9352
rect 12667 -9378 12693 -9352
rect 15307 -5650 15333 -5624
rect 15467 -5650 15493 -5624
rect 15627 -5650 15653 -5624
rect 15787 -5650 15813 -5624
rect 15947 -5650 15973 -5624
rect 16107 -5650 16133 -5624
rect 16267 -5650 16293 -5624
rect 16427 -5650 16453 -5624
rect 16587 -5650 16613 -5624
rect 16747 -5650 16773 -5624
rect 16907 -5650 16933 -5624
rect 17067 -5650 17093 -5624
rect 17227 -5650 17253 -5624
rect 17387 -5650 17413 -5624
rect 17547 -5650 17573 -5624
rect 17707 -5650 17733 -5624
rect 17867 -5650 17893 -5624
rect 18027 -5650 18053 -5624
rect 18187 -5650 18213 -5624
rect 18347 -5650 18373 -5624
rect 18507 -5650 18533 -5624
rect 18667 -5650 18693 -5624
rect 15122 -5753 15148 -5727
rect 18855 -5753 18881 -5727
rect 15122 -5913 15148 -5887
rect 15122 -6073 15148 -6047
rect 15122 -6233 15148 -6207
rect 15122 -6393 15148 -6367
rect 15122 -6553 15148 -6527
rect 15122 -6713 15148 -6687
rect 15122 -6873 15148 -6847
rect 15122 -7033 15148 -7007
rect 15122 -7193 15148 -7167
rect 15122 -7353 15148 -7327
rect 15122 -7513 15148 -7487
rect 15122 -7673 15148 -7647
rect 15122 -7833 15148 -7807
rect 15122 -7993 15148 -7967
rect 15122 -8153 15148 -8127
rect 15122 -8313 15148 -8287
rect 15122 -8473 15148 -8447
rect 15122 -8633 15148 -8607
rect 15122 -8793 15148 -8767
rect 15122 -8953 15148 -8927
rect 15122 -9113 15148 -9087
rect 18855 -5913 18881 -5887
rect 18855 -6073 18881 -6047
rect 18855 -6233 18881 -6207
rect 18855 -6393 18881 -6367
rect 18855 -6553 18881 -6527
rect 18855 -6713 18881 -6687
rect 18855 -6873 18881 -6847
rect 18855 -7033 18881 -7007
rect 18855 -7193 18881 -7167
rect 18855 -7353 18881 -7327
rect 18855 -7513 18881 -7487
rect 18855 -7673 18881 -7647
rect 18855 -7833 18881 -7807
rect 18855 -7993 18881 -7967
rect 18855 -8153 18881 -8127
rect 18855 -8313 18881 -8287
rect 18855 -8473 18881 -8447
rect 18855 -8633 18881 -8607
rect 18855 -8793 18881 -8767
rect 18855 -8953 18881 -8927
rect 18855 -9113 18881 -9087
rect 15122 -9273 15148 -9247
rect 18855 -9273 18881 -9247
rect 15307 -9378 15333 -9352
rect 15467 -9378 15493 -9352
rect 15627 -9378 15653 -9352
rect 15787 -9378 15813 -9352
rect 15947 -9378 15973 -9352
rect 16107 -9378 16133 -9352
rect 16267 -9378 16293 -9352
rect 16427 -9378 16453 -9352
rect 16587 -9378 16613 -9352
rect 16747 -9378 16773 -9352
rect 16907 -9378 16933 -9352
rect 17067 -9378 17093 -9352
rect 17227 -9378 17253 -9352
rect 17387 -9378 17413 -9352
rect 17547 -9378 17573 -9352
rect 17707 -9378 17733 -9352
rect 17867 -9378 17893 -9352
rect 18027 -9378 18053 -9352
rect 18187 -9378 18213 -9352
rect 18347 -9378 18373 -9352
rect 18507 -9378 18533 -9352
rect 18667 -9378 18693 -9352
rect 21307 -5650 21333 -5624
rect 21467 -5650 21493 -5624
rect 21627 -5650 21653 -5624
rect 21787 -5650 21813 -5624
rect 21947 -5650 21973 -5624
rect 22107 -5650 22133 -5624
rect 22267 -5650 22293 -5624
rect 22427 -5650 22453 -5624
rect 22587 -5650 22613 -5624
rect 22747 -5650 22773 -5624
rect 22907 -5650 22933 -5624
rect 23067 -5650 23093 -5624
rect 23227 -5650 23253 -5624
rect 23387 -5650 23413 -5624
rect 23547 -5650 23573 -5624
rect 23707 -5650 23733 -5624
rect 23867 -5650 23893 -5624
rect 24027 -5650 24053 -5624
rect 24187 -5650 24213 -5624
rect 24347 -5650 24373 -5624
rect 24507 -5650 24533 -5624
rect 24667 -5650 24693 -5624
rect 21122 -5753 21148 -5727
rect 24855 -5753 24881 -5727
rect 21122 -5913 21148 -5887
rect 21122 -6073 21148 -6047
rect 21122 -6233 21148 -6207
rect 21122 -6393 21148 -6367
rect 21122 -6553 21148 -6527
rect 21122 -6713 21148 -6687
rect 21122 -6873 21148 -6847
rect 21122 -7033 21148 -7007
rect 21122 -7193 21148 -7167
rect 21122 -7353 21148 -7327
rect 21122 -7513 21148 -7487
rect 21122 -7673 21148 -7647
rect 21122 -7833 21148 -7807
rect 21122 -7993 21148 -7967
rect 21122 -8153 21148 -8127
rect 21122 -8313 21148 -8287
rect 21122 -8473 21148 -8447
rect 21122 -8633 21148 -8607
rect 21122 -8793 21148 -8767
rect 21122 -8953 21148 -8927
rect 21122 -9113 21148 -9087
rect 24855 -5913 24881 -5887
rect 24855 -6073 24881 -6047
rect 24855 -6233 24881 -6207
rect 24855 -6393 24881 -6367
rect 24855 -6553 24881 -6527
rect 24855 -6713 24881 -6687
rect 24855 -6873 24881 -6847
rect 24855 -7033 24881 -7007
rect 24855 -7193 24881 -7167
rect 24855 -7353 24881 -7327
rect 24855 -7513 24881 -7487
rect 24855 -7673 24881 -7647
rect 24855 -7833 24881 -7807
rect 24855 -7993 24881 -7967
rect 24855 -8153 24881 -8127
rect 24855 -8313 24881 -8287
rect 24855 -8473 24881 -8447
rect 24855 -8633 24881 -8607
rect 24855 -8793 24881 -8767
rect 24855 -8953 24881 -8927
rect 24855 -9113 24881 -9087
rect 21122 -9273 21148 -9247
rect 24855 -9273 24881 -9247
rect 21307 -9378 21333 -9352
rect 21467 -9378 21493 -9352
rect 21627 -9378 21653 -9352
rect 21787 -9378 21813 -9352
rect 21947 -9378 21973 -9352
rect 22107 -9378 22133 -9352
rect 22267 -9378 22293 -9352
rect 22427 -9378 22453 -9352
rect 22587 -9378 22613 -9352
rect 22747 -9378 22773 -9352
rect 22907 -9378 22933 -9352
rect 23067 -9378 23093 -9352
rect 23227 -9378 23253 -9352
rect 23387 -9378 23413 -9352
rect 23547 -9378 23573 -9352
rect 23707 -9378 23733 -9352
rect 23867 -9378 23893 -9352
rect 24027 -9378 24053 -9352
rect 24187 -9378 24213 -9352
rect 24347 -9378 24373 -9352
rect 24507 -9378 24533 -9352
rect 24667 -9378 24693 -9352
rect 3307 -11650 3333 -11624
rect 3467 -11650 3493 -11624
rect 3627 -11650 3653 -11624
rect 3787 -11650 3813 -11624
rect 3947 -11650 3973 -11624
rect 4107 -11650 4133 -11624
rect 4267 -11650 4293 -11624
rect 4427 -11650 4453 -11624
rect 4587 -11650 4613 -11624
rect 4747 -11650 4773 -11624
rect 4907 -11650 4933 -11624
rect 5067 -11650 5093 -11624
rect 5227 -11650 5253 -11624
rect 5387 -11650 5413 -11624
rect 5547 -11650 5573 -11624
rect 5707 -11650 5733 -11624
rect 5867 -11650 5893 -11624
rect 6027 -11650 6053 -11624
rect 6187 -11650 6213 -11624
rect 6347 -11650 6373 -11624
rect 6507 -11650 6533 -11624
rect 6667 -11650 6693 -11624
rect 3122 -11753 3148 -11727
rect 6855 -11753 6881 -11727
rect 3122 -11913 3148 -11887
rect 3122 -12073 3148 -12047
rect 3122 -12233 3148 -12207
rect 3122 -12393 3148 -12367
rect 3122 -12553 3148 -12527
rect 3122 -12713 3148 -12687
rect 3122 -12873 3148 -12847
rect 3122 -13033 3148 -13007
rect 3122 -13193 3148 -13167
rect 3122 -13353 3148 -13327
rect 3122 -13513 3148 -13487
rect 3122 -13673 3148 -13647
rect 3122 -13833 3148 -13807
rect 3122 -13993 3148 -13967
rect 3122 -14153 3148 -14127
rect 3122 -14313 3148 -14287
rect 3122 -14473 3148 -14447
rect 3122 -14633 3148 -14607
rect 3122 -14793 3148 -14767
rect 3122 -14953 3148 -14927
rect 3122 -15113 3148 -15087
rect 6855 -11913 6881 -11887
rect 6855 -12073 6881 -12047
rect 6855 -12233 6881 -12207
rect 6855 -12393 6881 -12367
rect 6855 -12553 6881 -12527
rect 6855 -12713 6881 -12687
rect 6855 -12873 6881 -12847
rect 6855 -13033 6881 -13007
rect 6855 -13193 6881 -13167
rect 6855 -13353 6881 -13327
rect 6855 -13513 6881 -13487
rect 6855 -13673 6881 -13647
rect 6855 -13833 6881 -13807
rect 6855 -13993 6881 -13967
rect 6855 -14153 6881 -14127
rect 6855 -14313 6881 -14287
rect 6855 -14473 6881 -14447
rect 6855 -14633 6881 -14607
rect 6855 -14793 6881 -14767
rect 6855 -14953 6881 -14927
rect 6855 -15113 6881 -15087
rect 3122 -15273 3148 -15247
rect 6855 -15273 6881 -15247
rect 3307 -15378 3333 -15352
rect 3467 -15378 3493 -15352
rect 3627 -15378 3653 -15352
rect 3787 -15378 3813 -15352
rect 3947 -15378 3973 -15352
rect 4107 -15378 4133 -15352
rect 4267 -15378 4293 -15352
rect 4427 -15378 4453 -15352
rect 4587 -15378 4613 -15352
rect 4747 -15378 4773 -15352
rect 4907 -15378 4933 -15352
rect 5067 -15378 5093 -15352
rect 5227 -15378 5253 -15352
rect 5387 -15378 5413 -15352
rect 5547 -15378 5573 -15352
rect 5707 -15378 5733 -15352
rect 5867 -15378 5893 -15352
rect 6027 -15378 6053 -15352
rect 6187 -15378 6213 -15352
rect 6347 -15378 6373 -15352
rect 6507 -15378 6533 -15352
rect 6667 -15378 6693 -15352
rect 9307 -11650 9333 -11624
rect 9467 -11650 9493 -11624
rect 9627 -11650 9653 -11624
rect 9787 -11650 9813 -11624
rect 9947 -11650 9973 -11624
rect 10107 -11650 10133 -11624
rect 10267 -11650 10293 -11624
rect 10427 -11650 10453 -11624
rect 10587 -11650 10613 -11624
rect 10747 -11650 10773 -11624
rect 10907 -11650 10933 -11624
rect 11067 -11650 11093 -11624
rect 11227 -11650 11253 -11624
rect 11387 -11650 11413 -11624
rect 11547 -11650 11573 -11624
rect 11707 -11650 11733 -11624
rect 11867 -11650 11893 -11624
rect 12027 -11650 12053 -11624
rect 12187 -11650 12213 -11624
rect 12347 -11650 12373 -11624
rect 12507 -11650 12533 -11624
rect 12667 -11650 12693 -11624
rect 9122 -11753 9148 -11727
rect 12855 -11753 12881 -11727
rect 9122 -11913 9148 -11887
rect 9122 -12073 9148 -12047
rect 9122 -12233 9148 -12207
rect 9122 -12393 9148 -12367
rect 9122 -12553 9148 -12527
rect 9122 -12713 9148 -12687
rect 9122 -12873 9148 -12847
rect 9122 -13033 9148 -13007
rect 9122 -13193 9148 -13167
rect 9122 -13353 9148 -13327
rect 9122 -13513 9148 -13487
rect 9122 -13673 9148 -13647
rect 9122 -13833 9148 -13807
rect 9122 -13993 9148 -13967
rect 9122 -14153 9148 -14127
rect 9122 -14313 9148 -14287
rect 9122 -14473 9148 -14447
rect 9122 -14633 9148 -14607
rect 9122 -14793 9148 -14767
rect 9122 -14953 9148 -14927
rect 9122 -15113 9148 -15087
rect 12855 -11913 12881 -11887
rect 12855 -12073 12881 -12047
rect 12855 -12233 12881 -12207
rect 12855 -12393 12881 -12367
rect 12855 -12553 12881 -12527
rect 12855 -12713 12881 -12687
rect 12855 -12873 12881 -12847
rect 12855 -13033 12881 -13007
rect 12855 -13193 12881 -13167
rect 12855 -13353 12881 -13327
rect 12855 -13513 12881 -13487
rect 12855 -13673 12881 -13647
rect 12855 -13833 12881 -13807
rect 12855 -13993 12881 -13967
rect 12855 -14153 12881 -14127
rect 12855 -14313 12881 -14287
rect 12855 -14473 12881 -14447
rect 12855 -14633 12881 -14607
rect 12855 -14793 12881 -14767
rect 12855 -14953 12881 -14927
rect 12855 -15113 12881 -15087
rect 9122 -15273 9148 -15247
rect 12855 -15273 12881 -15247
rect 9307 -15378 9333 -15352
rect 9467 -15378 9493 -15352
rect 9627 -15378 9653 -15352
rect 9787 -15378 9813 -15352
rect 9947 -15378 9973 -15352
rect 10107 -15378 10133 -15352
rect 10267 -15378 10293 -15352
rect 10427 -15378 10453 -15352
rect 10587 -15378 10613 -15352
rect 10747 -15378 10773 -15352
rect 10907 -15378 10933 -15352
rect 11067 -15378 11093 -15352
rect 11227 -15378 11253 -15352
rect 11387 -15378 11413 -15352
rect 11547 -15378 11573 -15352
rect 11707 -15378 11733 -15352
rect 11867 -15378 11893 -15352
rect 12027 -15378 12053 -15352
rect 12187 -15378 12213 -15352
rect 12347 -15378 12373 -15352
rect 12507 -15378 12533 -15352
rect 12667 -15378 12693 -15352
rect 15307 -11650 15333 -11624
rect 15467 -11650 15493 -11624
rect 15627 -11650 15653 -11624
rect 15787 -11650 15813 -11624
rect 15947 -11650 15973 -11624
rect 16107 -11650 16133 -11624
rect 16267 -11650 16293 -11624
rect 16427 -11650 16453 -11624
rect 16587 -11650 16613 -11624
rect 16747 -11650 16773 -11624
rect 16907 -11650 16933 -11624
rect 17067 -11650 17093 -11624
rect 17227 -11650 17253 -11624
rect 17387 -11650 17413 -11624
rect 17547 -11650 17573 -11624
rect 17707 -11650 17733 -11624
rect 17867 -11650 17893 -11624
rect 18027 -11650 18053 -11624
rect 18187 -11650 18213 -11624
rect 18347 -11650 18373 -11624
rect 18507 -11650 18533 -11624
rect 18667 -11650 18693 -11624
rect 15122 -11753 15148 -11727
rect 18855 -11753 18881 -11727
rect 15122 -11913 15148 -11887
rect 15122 -12073 15148 -12047
rect 15122 -12233 15148 -12207
rect 15122 -12393 15148 -12367
rect 15122 -12553 15148 -12527
rect 15122 -12713 15148 -12687
rect 15122 -12873 15148 -12847
rect 15122 -13033 15148 -13007
rect 15122 -13193 15148 -13167
rect 15122 -13353 15148 -13327
rect 15122 -13513 15148 -13487
rect 15122 -13673 15148 -13647
rect 15122 -13833 15148 -13807
rect 15122 -13993 15148 -13967
rect 15122 -14153 15148 -14127
rect 15122 -14313 15148 -14287
rect 15122 -14473 15148 -14447
rect 15122 -14633 15148 -14607
rect 15122 -14793 15148 -14767
rect 15122 -14953 15148 -14927
rect 15122 -15113 15148 -15087
rect 18855 -11913 18881 -11887
rect 18855 -12073 18881 -12047
rect 18855 -12233 18881 -12207
rect 18855 -12393 18881 -12367
rect 18855 -12553 18881 -12527
rect 18855 -12713 18881 -12687
rect 18855 -12873 18881 -12847
rect 18855 -13033 18881 -13007
rect 18855 -13193 18881 -13167
rect 18855 -13353 18881 -13327
rect 18855 -13513 18881 -13487
rect 18855 -13673 18881 -13647
rect 18855 -13833 18881 -13807
rect 18855 -13993 18881 -13967
rect 18855 -14153 18881 -14127
rect 18855 -14313 18881 -14287
rect 18855 -14473 18881 -14447
rect 18855 -14633 18881 -14607
rect 18855 -14793 18881 -14767
rect 18855 -14953 18881 -14927
rect 18855 -15113 18881 -15087
rect 15122 -15273 15148 -15247
rect 18855 -15273 18881 -15247
rect 15307 -15378 15333 -15352
rect 15467 -15378 15493 -15352
rect 15627 -15378 15653 -15352
rect 15787 -15378 15813 -15352
rect 15947 -15378 15973 -15352
rect 16107 -15378 16133 -15352
rect 16267 -15378 16293 -15352
rect 16427 -15378 16453 -15352
rect 16587 -15378 16613 -15352
rect 16747 -15378 16773 -15352
rect 16907 -15378 16933 -15352
rect 17067 -15378 17093 -15352
rect 17227 -15378 17253 -15352
rect 17387 -15378 17413 -15352
rect 17547 -15378 17573 -15352
rect 17707 -15378 17733 -15352
rect 17867 -15378 17893 -15352
rect 18027 -15378 18053 -15352
rect 18187 -15378 18213 -15352
rect 18347 -15378 18373 -15352
rect 18507 -15378 18533 -15352
rect 18667 -15378 18693 -15352
rect 21307 -11650 21333 -11624
rect 21467 -11650 21493 -11624
rect 21627 -11650 21653 -11624
rect 21787 -11650 21813 -11624
rect 21947 -11650 21973 -11624
rect 22107 -11650 22133 -11624
rect 22267 -11650 22293 -11624
rect 22427 -11650 22453 -11624
rect 22587 -11650 22613 -11624
rect 22747 -11650 22773 -11624
rect 22907 -11650 22933 -11624
rect 23067 -11650 23093 -11624
rect 23227 -11650 23253 -11624
rect 23387 -11650 23413 -11624
rect 23547 -11650 23573 -11624
rect 23707 -11650 23733 -11624
rect 23867 -11650 23893 -11624
rect 24027 -11650 24053 -11624
rect 24187 -11650 24213 -11624
rect 24347 -11650 24373 -11624
rect 24507 -11650 24533 -11624
rect 24667 -11650 24693 -11624
rect 21122 -11753 21148 -11727
rect 24855 -11753 24881 -11727
rect 21122 -11913 21148 -11887
rect 21122 -12073 21148 -12047
rect 21122 -12233 21148 -12207
rect 21122 -12393 21148 -12367
rect 21122 -12553 21148 -12527
rect 21122 -12713 21148 -12687
rect 21122 -12873 21148 -12847
rect 21122 -13033 21148 -13007
rect 21122 -13193 21148 -13167
rect 21122 -13353 21148 -13327
rect 21122 -13513 21148 -13487
rect 21122 -13673 21148 -13647
rect 21122 -13833 21148 -13807
rect 21122 -13993 21148 -13967
rect 21122 -14153 21148 -14127
rect 21122 -14313 21148 -14287
rect 21122 -14473 21148 -14447
rect 21122 -14633 21148 -14607
rect 21122 -14793 21148 -14767
rect 21122 -14953 21148 -14927
rect 21122 -15113 21148 -15087
rect 24855 -11913 24881 -11887
rect 24855 -12073 24881 -12047
rect 24855 -12233 24881 -12207
rect 24855 -12393 24881 -12367
rect 24855 -12553 24881 -12527
rect 24855 -12713 24881 -12687
rect 24855 -12873 24881 -12847
rect 24855 -13033 24881 -13007
rect 24855 -13193 24881 -13167
rect 24855 -13353 24881 -13327
rect 24855 -13513 24881 -13487
rect 24855 -13673 24881 -13647
rect 24855 -13833 24881 -13807
rect 24855 -13993 24881 -13967
rect 24855 -14153 24881 -14127
rect 24855 -14313 24881 -14287
rect 24855 -14473 24881 -14447
rect 24855 -14633 24881 -14607
rect 24855 -14793 24881 -14767
rect 24855 -14953 24881 -14927
rect 24855 -15113 24881 -15087
rect 21122 -15273 21148 -15247
rect 24855 -15273 24881 -15247
rect 21307 -15378 21333 -15352
rect 21467 -15378 21493 -15352
rect 21627 -15378 21653 -15352
rect 21787 -15378 21813 -15352
rect 21947 -15378 21973 -15352
rect 22107 -15378 22133 -15352
rect 22267 -15378 22293 -15352
rect 22427 -15378 22453 -15352
rect 22587 -15378 22613 -15352
rect 22747 -15378 22773 -15352
rect 22907 -15378 22933 -15352
rect 23067 -15378 23093 -15352
rect 23227 -15378 23253 -15352
rect 23387 -15378 23413 -15352
rect 23547 -15378 23573 -15352
rect 23707 -15378 23733 -15352
rect 23867 -15378 23893 -15352
rect 24027 -15378 24053 -15352
rect 24187 -15378 24213 -15352
rect 24347 -15378 24373 -15352
rect 24507 -15378 24533 -15352
rect 24667 -15378 24693 -15352
<< metal2 >>
rect 10900 -1500 11700 -1400
rect 11600 -3600 11700 -1500
rect 11600 -3700 11650 -3600
rect 11750 -3700 11800 -3600
rect 11630 -3740 11710 -3735
rect 11630 -3770 11635 -3740
rect 11705 -3770 11710 -3740
rect 11630 -3820 11710 -3770
rect 11630 -3860 11635 -3820
rect 11705 -3860 11710 -3820
rect 11770 -3860 11775 -3820
rect 11845 -3860 11850 -3820
rect 11770 -3900 11850 -3860
rect 11770 -3930 11775 -3900
rect 11845 -3930 11850 -3900
rect 11770 -3935 11850 -3930
rect 11600 -4050 11650 -3950
rect 11750 -4050 11800 -3950
rect 11600 -4150 11700 -4050
rect 11050 -4250 11700 -4150
rect 8195 -4760 8235 -4755
rect 8195 -4790 8200 -4760
rect 8230 -4790 8235 -4760
rect 8195 -4795 8235 -4790
rect 8230 -4830 8270 -4825
rect 8230 -4860 8235 -4830
rect 8265 -4860 8270 -4830
rect 8230 -4865 8270 -4860
rect 7975 -5255 8405 -5250
rect 7975 -5425 8355 -5255
rect 8400 -5425 8405 -5255
rect 8705 -5255 8760 -4750
rect 8510 -5310 8570 -5305
rect 8510 -5370 8515 -5310
rect 8565 -5370 8570 -5310
rect 8510 -5375 8570 -5370
rect 7975 -5430 8405 -5425
rect 8705 -5425 8710 -5255
rect 8755 -5425 8760 -5255
rect 8705 -5430 8760 -5425
rect 3000 -5555 7000 -5500
rect 7975 -5555 8085 -5430
rect 3000 -5623 8085 -5555
rect 3000 -5651 3306 -5623
rect 3334 -5651 3466 -5623
rect 3494 -5651 3626 -5623
rect 3654 -5651 3786 -5623
rect 3814 -5651 3946 -5623
rect 3974 -5651 4106 -5623
rect 4134 -5651 4266 -5623
rect 4294 -5651 4426 -5623
rect 4454 -5651 4586 -5623
rect 4614 -5651 4746 -5623
rect 4774 -5651 4906 -5623
rect 4934 -5651 5066 -5623
rect 5094 -5651 5226 -5623
rect 5254 -5651 5386 -5623
rect 5414 -5651 5546 -5623
rect 5574 -5651 5706 -5623
rect 5734 -5651 5866 -5623
rect 5894 -5651 6026 -5623
rect 6054 -5651 6186 -5623
rect 6214 -5651 6346 -5623
rect 6374 -5651 6506 -5623
rect 6534 -5651 6666 -5623
rect 6694 -5651 8085 -5623
rect 3000 -5655 8085 -5651
rect 9000 -5623 13000 -5500
rect 9000 -5651 9306 -5623
rect 9334 -5651 9466 -5623
rect 9494 -5651 9626 -5623
rect 9654 -5651 9786 -5623
rect 9814 -5651 9946 -5623
rect 9974 -5651 10106 -5623
rect 10134 -5651 10266 -5623
rect 10294 -5651 10426 -5623
rect 10454 -5651 10586 -5623
rect 10614 -5651 10746 -5623
rect 10774 -5651 10906 -5623
rect 10934 -5651 11066 -5623
rect 11094 -5651 11226 -5623
rect 11254 -5651 11386 -5623
rect 11414 -5651 11546 -5623
rect 11574 -5651 11706 -5623
rect 11734 -5651 11866 -5623
rect 11894 -5651 12026 -5623
rect 12054 -5651 12186 -5623
rect 12214 -5651 12346 -5623
rect 12374 -5651 12506 -5623
rect 12534 -5651 12666 -5623
rect 12694 -5651 13000 -5623
rect 3000 -5726 7000 -5655
rect 3000 -5754 3121 -5726
rect 3149 -5754 6854 -5726
rect 6882 -5754 7000 -5726
rect 3000 -5770 7000 -5754
rect 3000 -5886 3270 -5770
rect 3000 -5914 3121 -5886
rect 3149 -5914 3270 -5886
rect 3000 -6046 3270 -5914
rect 3000 -6074 3121 -6046
rect 3149 -6074 3270 -6046
rect 3000 -6206 3270 -6074
rect 3000 -6234 3121 -6206
rect 3149 -6234 3270 -6206
rect 3000 -6366 3270 -6234
rect 3000 -6394 3121 -6366
rect 3149 -6394 3270 -6366
rect 3000 -6526 3270 -6394
rect 3000 -6554 3121 -6526
rect 3149 -6554 3270 -6526
rect 3000 -6686 3270 -6554
rect 3000 -6714 3121 -6686
rect 3149 -6714 3270 -6686
rect 3000 -6846 3270 -6714
rect 3000 -6874 3121 -6846
rect 3149 -6874 3270 -6846
rect 3000 -7006 3270 -6874
rect 3000 -7034 3121 -7006
rect 3149 -7034 3270 -7006
rect 3000 -7166 3270 -7034
rect 3000 -7194 3121 -7166
rect 3149 -7194 3270 -7166
rect 3000 -7326 3270 -7194
rect 3000 -7354 3121 -7326
rect 3149 -7354 3270 -7326
rect 3000 -7486 3270 -7354
rect 3000 -7514 3121 -7486
rect 3149 -7514 3270 -7486
rect 3000 -7646 3270 -7514
rect 3000 -7674 3121 -7646
rect 3149 -7674 3270 -7646
rect 3000 -7806 3270 -7674
rect 3000 -7834 3121 -7806
rect 3149 -7834 3270 -7806
rect 3000 -7966 3270 -7834
rect 3000 -7994 3121 -7966
rect 3149 -7994 3270 -7966
rect 3000 -8126 3270 -7994
rect 3000 -8154 3121 -8126
rect 3149 -8154 3270 -8126
rect 3000 -8286 3270 -8154
rect 3000 -8314 3121 -8286
rect 3149 -8314 3270 -8286
rect 3000 -8446 3270 -8314
rect 3000 -8474 3121 -8446
rect 3149 -8474 3270 -8446
rect 3000 -8606 3270 -8474
rect 3000 -8634 3121 -8606
rect 3149 -8634 3270 -8606
rect 3000 -8766 3270 -8634
rect 3000 -8794 3121 -8766
rect 3149 -8794 3270 -8766
rect 3000 -8926 3270 -8794
rect 3000 -8954 3121 -8926
rect 3149 -8954 3270 -8926
rect 3000 -9086 3270 -8954
rect 3000 -9114 3121 -9086
rect 3149 -9114 3270 -9086
rect 3000 -9230 3270 -9114
rect 6730 -5886 7000 -5770
rect 6730 -5914 6854 -5886
rect 6882 -5914 7000 -5886
rect 6730 -6046 7000 -5914
rect 6730 -6074 6854 -6046
rect 6882 -6074 7000 -6046
rect 6730 -6206 7000 -6074
rect 6730 -6234 6854 -6206
rect 6882 -6234 7000 -6206
rect 6730 -6366 7000 -6234
rect 6730 -6394 6854 -6366
rect 6882 -6394 7000 -6366
rect 6730 -6526 7000 -6394
rect 6730 -6554 6854 -6526
rect 6882 -6554 7000 -6526
rect 6730 -6686 7000 -6554
rect 6730 -6714 6854 -6686
rect 6882 -6714 7000 -6686
rect 6730 -6846 7000 -6714
rect 6730 -6874 6854 -6846
rect 6882 -6874 7000 -6846
rect 6730 -7006 7000 -6874
rect 6730 -7034 6854 -7006
rect 6882 -7034 7000 -7006
rect 6730 -7166 7000 -7034
rect 6730 -7194 6854 -7166
rect 6882 -7194 7000 -7166
rect 6730 -7326 7000 -7194
rect 6730 -7354 6854 -7326
rect 6882 -7354 7000 -7326
rect 6730 -7486 7000 -7354
rect 6730 -7514 6854 -7486
rect 6882 -7514 7000 -7486
rect 6730 -7646 7000 -7514
rect 6730 -7674 6854 -7646
rect 6882 -7674 7000 -7646
rect 6730 -7806 7000 -7674
rect 6730 -7834 6854 -7806
rect 6882 -7834 7000 -7806
rect 6730 -7966 7000 -7834
rect 6730 -7994 6854 -7966
rect 6882 -7994 7000 -7966
rect 6730 -8126 7000 -7994
rect 6730 -8154 6854 -8126
rect 6882 -8154 7000 -8126
rect 6730 -8286 7000 -8154
rect 6730 -8314 6854 -8286
rect 6882 -8314 7000 -8286
rect 6730 -8446 7000 -8314
rect 6730 -8474 6854 -8446
rect 6882 -8474 7000 -8446
rect 6730 -8606 7000 -8474
rect 6730 -8634 6854 -8606
rect 6882 -8634 7000 -8606
rect 6730 -8766 7000 -8634
rect 6730 -8794 6854 -8766
rect 6882 -8794 7000 -8766
rect 6730 -8926 7000 -8794
rect 6730 -8954 6854 -8926
rect 6882 -8954 7000 -8926
rect 6730 -9086 7000 -8954
rect 6730 -9114 6854 -9086
rect 6882 -9114 7000 -9086
rect 6730 -9230 7000 -9114
rect 3000 -9246 7000 -9230
rect 3000 -9274 3121 -9246
rect 3149 -9274 6854 -9246
rect 6882 -9274 7000 -9246
rect 3000 -9351 7000 -9274
rect 3000 -9379 3306 -9351
rect 3334 -9379 3466 -9351
rect 3494 -9379 3626 -9351
rect 3654 -9379 3786 -9351
rect 3814 -9379 3946 -9351
rect 3974 -9379 4106 -9351
rect 4134 -9379 4266 -9351
rect 4294 -9379 4426 -9351
rect 4454 -9379 4586 -9351
rect 4614 -9379 4746 -9351
rect 4774 -9379 4906 -9351
rect 4934 -9379 5066 -9351
rect 5094 -9379 5226 -9351
rect 5254 -9379 5386 -9351
rect 5414 -9379 5546 -9351
rect 5574 -9379 5706 -9351
rect 5734 -9379 5866 -9351
rect 5894 -9379 6026 -9351
rect 6054 -9379 6186 -9351
rect 6214 -9379 6346 -9351
rect 6374 -9379 6506 -9351
rect 6534 -9379 6666 -9351
rect 6694 -9379 7000 -9351
rect 3000 -9500 7000 -9379
rect 9000 -5726 13000 -5651
rect 9000 -5754 9121 -5726
rect 9149 -5754 12854 -5726
rect 12882 -5754 13000 -5726
rect 9000 -5770 13000 -5754
rect 9000 -5886 9270 -5770
rect 9000 -5914 9121 -5886
rect 9149 -5914 9270 -5886
rect 9000 -6046 9270 -5914
rect 9000 -6074 9121 -6046
rect 9149 -6074 9270 -6046
rect 9000 -6206 9270 -6074
rect 9000 -6234 9121 -6206
rect 9149 -6234 9270 -6206
rect 9000 -6366 9270 -6234
rect 9000 -6394 9121 -6366
rect 9149 -6394 9270 -6366
rect 9000 -6526 9270 -6394
rect 9000 -6554 9121 -6526
rect 9149 -6554 9270 -6526
rect 9000 -6686 9270 -6554
rect 9000 -6714 9121 -6686
rect 9149 -6714 9270 -6686
rect 9000 -6846 9270 -6714
rect 9000 -6874 9121 -6846
rect 9149 -6874 9270 -6846
rect 9000 -7006 9270 -6874
rect 9000 -7034 9121 -7006
rect 9149 -7034 9270 -7006
rect 9000 -7166 9270 -7034
rect 9000 -7194 9121 -7166
rect 9149 -7194 9270 -7166
rect 9000 -7326 9270 -7194
rect 9000 -7354 9121 -7326
rect 9149 -7354 9270 -7326
rect 9000 -7486 9270 -7354
rect 9000 -7514 9121 -7486
rect 9149 -7514 9270 -7486
rect 9000 -7646 9270 -7514
rect 9000 -7674 9121 -7646
rect 9149 -7674 9270 -7646
rect 9000 -7806 9270 -7674
rect 9000 -7834 9121 -7806
rect 9149 -7834 9270 -7806
rect 9000 -7966 9270 -7834
rect 9000 -7994 9121 -7966
rect 9149 -7994 9270 -7966
rect 9000 -8126 9270 -7994
rect 9000 -8154 9121 -8126
rect 9149 -8154 9270 -8126
rect 9000 -8286 9270 -8154
rect 9000 -8314 9121 -8286
rect 9149 -8314 9270 -8286
rect 9000 -8446 9270 -8314
rect 9000 -8474 9121 -8446
rect 9149 -8474 9270 -8446
rect 9000 -8606 9270 -8474
rect 9000 -8634 9121 -8606
rect 9149 -8634 9270 -8606
rect 9000 -8766 9270 -8634
rect 9000 -8794 9121 -8766
rect 9149 -8794 9270 -8766
rect 9000 -8926 9270 -8794
rect 9000 -8954 9121 -8926
rect 9149 -8954 9270 -8926
rect 9000 -9086 9270 -8954
rect 9000 -9114 9121 -9086
rect 9149 -9114 9270 -9086
rect 9000 -9230 9270 -9114
rect 12730 -5886 13000 -5770
rect 12730 -5914 12854 -5886
rect 12882 -5914 13000 -5886
rect 12730 -6046 13000 -5914
rect 12730 -6074 12854 -6046
rect 12882 -6074 13000 -6046
rect 12730 -6206 13000 -6074
rect 12730 -6234 12854 -6206
rect 12882 -6234 13000 -6206
rect 12730 -6366 13000 -6234
rect 12730 -6394 12854 -6366
rect 12882 -6394 13000 -6366
rect 12730 -6526 13000 -6394
rect 12730 -6554 12854 -6526
rect 12882 -6554 13000 -6526
rect 12730 -6686 13000 -6554
rect 12730 -6714 12854 -6686
rect 12882 -6714 13000 -6686
rect 12730 -6846 13000 -6714
rect 12730 -6874 12854 -6846
rect 12882 -6874 13000 -6846
rect 12730 -7006 13000 -6874
rect 12730 -7034 12854 -7006
rect 12882 -7034 13000 -7006
rect 12730 -7166 13000 -7034
rect 12730 -7194 12854 -7166
rect 12882 -7194 13000 -7166
rect 12730 -7326 13000 -7194
rect 12730 -7354 12854 -7326
rect 12882 -7354 13000 -7326
rect 12730 -7486 13000 -7354
rect 12730 -7514 12854 -7486
rect 12882 -7514 13000 -7486
rect 12730 -7646 13000 -7514
rect 12730 -7674 12854 -7646
rect 12882 -7674 13000 -7646
rect 12730 -7806 13000 -7674
rect 12730 -7834 12854 -7806
rect 12882 -7834 13000 -7806
rect 12730 -7966 13000 -7834
rect 12730 -7994 12854 -7966
rect 12882 -7994 13000 -7966
rect 12730 -8126 13000 -7994
rect 12730 -8154 12854 -8126
rect 12882 -8154 13000 -8126
rect 12730 -8286 13000 -8154
rect 12730 -8314 12854 -8286
rect 12882 -8314 13000 -8286
rect 12730 -8446 13000 -8314
rect 12730 -8474 12854 -8446
rect 12882 -8474 13000 -8446
rect 12730 -8606 13000 -8474
rect 12730 -8634 12854 -8606
rect 12882 -8634 13000 -8606
rect 12730 -8766 13000 -8634
rect 12730 -8794 12854 -8766
rect 12882 -8794 13000 -8766
rect 12730 -8926 13000 -8794
rect 12730 -8954 12854 -8926
rect 12882 -8954 13000 -8926
rect 12730 -9086 13000 -8954
rect 12730 -9114 12854 -9086
rect 12882 -9114 13000 -9086
rect 12730 -9230 13000 -9114
rect 9000 -9246 13000 -9230
rect 9000 -9274 9121 -9246
rect 9149 -9274 12854 -9246
rect 12882 -9274 13000 -9246
rect 9000 -9351 13000 -9274
rect 9000 -9379 9306 -9351
rect 9334 -9379 9466 -9351
rect 9494 -9379 9626 -9351
rect 9654 -9379 9786 -9351
rect 9814 -9379 9946 -9351
rect 9974 -9379 10106 -9351
rect 10134 -9379 10266 -9351
rect 10294 -9379 10426 -9351
rect 10454 -9379 10586 -9351
rect 10614 -9379 10746 -9351
rect 10774 -9379 10906 -9351
rect 10934 -9379 11066 -9351
rect 11094 -9379 11226 -9351
rect 11254 -9379 11386 -9351
rect 11414 -9379 11546 -9351
rect 11574 -9379 11706 -9351
rect 11734 -9379 11866 -9351
rect 11894 -9379 12026 -9351
rect 12054 -9379 12186 -9351
rect 12214 -9379 12346 -9351
rect 12374 -9379 12506 -9351
rect 12534 -9379 12666 -9351
rect 12694 -9379 13000 -9351
rect 9000 -9500 13000 -9379
rect 15000 -5623 19000 -5500
rect 15000 -5651 15306 -5623
rect 15334 -5651 15466 -5623
rect 15494 -5651 15626 -5623
rect 15654 -5651 15786 -5623
rect 15814 -5651 15946 -5623
rect 15974 -5651 16106 -5623
rect 16134 -5651 16266 -5623
rect 16294 -5651 16426 -5623
rect 16454 -5651 16586 -5623
rect 16614 -5651 16746 -5623
rect 16774 -5651 16906 -5623
rect 16934 -5651 17066 -5623
rect 17094 -5651 17226 -5623
rect 17254 -5651 17386 -5623
rect 17414 -5651 17546 -5623
rect 17574 -5651 17706 -5623
rect 17734 -5651 17866 -5623
rect 17894 -5651 18026 -5623
rect 18054 -5651 18186 -5623
rect 18214 -5651 18346 -5623
rect 18374 -5651 18506 -5623
rect 18534 -5651 18666 -5623
rect 18694 -5651 19000 -5623
rect 15000 -5726 19000 -5651
rect 15000 -5754 15121 -5726
rect 15149 -5754 18854 -5726
rect 18882 -5754 19000 -5726
rect 15000 -5770 19000 -5754
rect 15000 -5886 15270 -5770
rect 15000 -5914 15121 -5886
rect 15149 -5914 15270 -5886
rect 15000 -6046 15270 -5914
rect 15000 -6074 15121 -6046
rect 15149 -6074 15270 -6046
rect 15000 -6206 15270 -6074
rect 15000 -6234 15121 -6206
rect 15149 -6234 15270 -6206
rect 15000 -6366 15270 -6234
rect 15000 -6394 15121 -6366
rect 15149 -6394 15270 -6366
rect 15000 -6526 15270 -6394
rect 15000 -6554 15121 -6526
rect 15149 -6554 15270 -6526
rect 15000 -6686 15270 -6554
rect 15000 -6714 15121 -6686
rect 15149 -6714 15270 -6686
rect 15000 -6846 15270 -6714
rect 15000 -6874 15121 -6846
rect 15149 -6874 15270 -6846
rect 15000 -7006 15270 -6874
rect 15000 -7034 15121 -7006
rect 15149 -7034 15270 -7006
rect 15000 -7166 15270 -7034
rect 15000 -7194 15121 -7166
rect 15149 -7194 15270 -7166
rect 15000 -7326 15270 -7194
rect 15000 -7354 15121 -7326
rect 15149 -7354 15270 -7326
rect 15000 -7486 15270 -7354
rect 15000 -7514 15121 -7486
rect 15149 -7514 15270 -7486
rect 15000 -7646 15270 -7514
rect 15000 -7674 15121 -7646
rect 15149 -7674 15270 -7646
rect 15000 -7806 15270 -7674
rect 15000 -7834 15121 -7806
rect 15149 -7834 15270 -7806
rect 15000 -7966 15270 -7834
rect 15000 -7994 15121 -7966
rect 15149 -7994 15270 -7966
rect 15000 -8126 15270 -7994
rect 15000 -8154 15121 -8126
rect 15149 -8154 15270 -8126
rect 15000 -8286 15270 -8154
rect 15000 -8314 15121 -8286
rect 15149 -8314 15270 -8286
rect 15000 -8446 15270 -8314
rect 15000 -8474 15121 -8446
rect 15149 -8474 15270 -8446
rect 15000 -8606 15270 -8474
rect 15000 -8634 15121 -8606
rect 15149 -8634 15270 -8606
rect 15000 -8766 15270 -8634
rect 15000 -8794 15121 -8766
rect 15149 -8794 15270 -8766
rect 15000 -8926 15270 -8794
rect 15000 -8954 15121 -8926
rect 15149 -8954 15270 -8926
rect 15000 -9086 15270 -8954
rect 15000 -9114 15121 -9086
rect 15149 -9114 15270 -9086
rect 15000 -9230 15270 -9114
rect 18730 -5886 19000 -5770
rect 18730 -5914 18854 -5886
rect 18882 -5914 19000 -5886
rect 18730 -6046 19000 -5914
rect 18730 -6074 18854 -6046
rect 18882 -6074 19000 -6046
rect 18730 -6206 19000 -6074
rect 18730 -6234 18854 -6206
rect 18882 -6234 19000 -6206
rect 18730 -6366 19000 -6234
rect 18730 -6394 18854 -6366
rect 18882 -6394 19000 -6366
rect 18730 -6526 19000 -6394
rect 18730 -6554 18854 -6526
rect 18882 -6554 19000 -6526
rect 18730 -6686 19000 -6554
rect 18730 -6714 18854 -6686
rect 18882 -6714 19000 -6686
rect 18730 -6846 19000 -6714
rect 18730 -6874 18854 -6846
rect 18882 -6874 19000 -6846
rect 18730 -7006 19000 -6874
rect 18730 -7034 18854 -7006
rect 18882 -7034 19000 -7006
rect 18730 -7166 19000 -7034
rect 18730 -7194 18854 -7166
rect 18882 -7194 19000 -7166
rect 18730 -7326 19000 -7194
rect 18730 -7354 18854 -7326
rect 18882 -7354 19000 -7326
rect 18730 -7486 19000 -7354
rect 18730 -7514 18854 -7486
rect 18882 -7514 19000 -7486
rect 18730 -7646 19000 -7514
rect 18730 -7674 18854 -7646
rect 18882 -7674 19000 -7646
rect 18730 -7806 19000 -7674
rect 18730 -7834 18854 -7806
rect 18882 -7834 19000 -7806
rect 18730 -7966 19000 -7834
rect 18730 -7994 18854 -7966
rect 18882 -7994 19000 -7966
rect 18730 -8126 19000 -7994
rect 18730 -8154 18854 -8126
rect 18882 -8154 19000 -8126
rect 18730 -8286 19000 -8154
rect 18730 -8314 18854 -8286
rect 18882 -8314 19000 -8286
rect 18730 -8446 19000 -8314
rect 18730 -8474 18854 -8446
rect 18882 -8474 19000 -8446
rect 18730 -8606 19000 -8474
rect 18730 -8634 18854 -8606
rect 18882 -8634 19000 -8606
rect 18730 -8766 19000 -8634
rect 18730 -8794 18854 -8766
rect 18882 -8794 19000 -8766
rect 18730 -8926 19000 -8794
rect 18730 -8954 18854 -8926
rect 18882 -8954 19000 -8926
rect 18730 -9086 19000 -8954
rect 18730 -9114 18854 -9086
rect 18882 -9114 19000 -9086
rect 18730 -9230 19000 -9114
rect 15000 -9246 19000 -9230
rect 15000 -9274 15121 -9246
rect 15149 -9274 18854 -9246
rect 18882 -9274 19000 -9246
rect 15000 -9351 19000 -9274
rect 15000 -9379 15306 -9351
rect 15334 -9379 15466 -9351
rect 15494 -9379 15626 -9351
rect 15654 -9379 15786 -9351
rect 15814 -9379 15946 -9351
rect 15974 -9379 16106 -9351
rect 16134 -9379 16266 -9351
rect 16294 -9379 16426 -9351
rect 16454 -9379 16586 -9351
rect 16614 -9379 16746 -9351
rect 16774 -9379 16906 -9351
rect 16934 -9379 17066 -9351
rect 17094 -9379 17226 -9351
rect 17254 -9379 17386 -9351
rect 17414 -9379 17546 -9351
rect 17574 -9379 17706 -9351
rect 17734 -9379 17866 -9351
rect 17894 -9379 18026 -9351
rect 18054 -9379 18186 -9351
rect 18214 -9379 18346 -9351
rect 18374 -9379 18506 -9351
rect 18534 -9379 18666 -9351
rect 18694 -9379 19000 -9351
rect 15000 -9500 19000 -9379
rect 21000 -5623 25000 -5500
rect 21000 -5651 21306 -5623
rect 21334 -5651 21466 -5623
rect 21494 -5651 21626 -5623
rect 21654 -5651 21786 -5623
rect 21814 -5651 21946 -5623
rect 21974 -5651 22106 -5623
rect 22134 -5651 22266 -5623
rect 22294 -5651 22426 -5623
rect 22454 -5651 22586 -5623
rect 22614 -5651 22746 -5623
rect 22774 -5651 22906 -5623
rect 22934 -5651 23066 -5623
rect 23094 -5651 23226 -5623
rect 23254 -5651 23386 -5623
rect 23414 -5651 23546 -5623
rect 23574 -5651 23706 -5623
rect 23734 -5651 23866 -5623
rect 23894 -5651 24026 -5623
rect 24054 -5651 24186 -5623
rect 24214 -5651 24346 -5623
rect 24374 -5651 24506 -5623
rect 24534 -5651 24666 -5623
rect 24694 -5651 25000 -5623
rect 21000 -5726 25000 -5651
rect 21000 -5754 21121 -5726
rect 21149 -5754 24854 -5726
rect 24882 -5754 25000 -5726
rect 21000 -5770 25000 -5754
rect 21000 -5886 21270 -5770
rect 21000 -5914 21121 -5886
rect 21149 -5914 21270 -5886
rect 21000 -6046 21270 -5914
rect 21000 -6074 21121 -6046
rect 21149 -6074 21270 -6046
rect 21000 -6206 21270 -6074
rect 21000 -6234 21121 -6206
rect 21149 -6234 21270 -6206
rect 21000 -6366 21270 -6234
rect 21000 -6394 21121 -6366
rect 21149 -6394 21270 -6366
rect 21000 -6526 21270 -6394
rect 21000 -6554 21121 -6526
rect 21149 -6554 21270 -6526
rect 21000 -6686 21270 -6554
rect 21000 -6714 21121 -6686
rect 21149 -6714 21270 -6686
rect 21000 -6846 21270 -6714
rect 21000 -6874 21121 -6846
rect 21149 -6874 21270 -6846
rect 21000 -7006 21270 -6874
rect 21000 -7034 21121 -7006
rect 21149 -7034 21270 -7006
rect 21000 -7166 21270 -7034
rect 21000 -7194 21121 -7166
rect 21149 -7194 21270 -7166
rect 21000 -7326 21270 -7194
rect 21000 -7354 21121 -7326
rect 21149 -7354 21270 -7326
rect 21000 -7486 21270 -7354
rect 21000 -7514 21121 -7486
rect 21149 -7514 21270 -7486
rect 21000 -7646 21270 -7514
rect 21000 -7674 21121 -7646
rect 21149 -7674 21270 -7646
rect 21000 -7806 21270 -7674
rect 21000 -7834 21121 -7806
rect 21149 -7834 21270 -7806
rect 21000 -7966 21270 -7834
rect 21000 -7994 21121 -7966
rect 21149 -7994 21270 -7966
rect 21000 -8126 21270 -7994
rect 21000 -8154 21121 -8126
rect 21149 -8154 21270 -8126
rect 21000 -8286 21270 -8154
rect 21000 -8314 21121 -8286
rect 21149 -8314 21270 -8286
rect 21000 -8446 21270 -8314
rect 21000 -8474 21121 -8446
rect 21149 -8474 21270 -8446
rect 21000 -8606 21270 -8474
rect 21000 -8634 21121 -8606
rect 21149 -8634 21270 -8606
rect 21000 -8766 21270 -8634
rect 21000 -8794 21121 -8766
rect 21149 -8794 21270 -8766
rect 21000 -8926 21270 -8794
rect 21000 -8954 21121 -8926
rect 21149 -8954 21270 -8926
rect 21000 -9086 21270 -8954
rect 21000 -9114 21121 -9086
rect 21149 -9114 21270 -9086
rect 21000 -9230 21270 -9114
rect 24730 -5886 25000 -5770
rect 24730 -5914 24854 -5886
rect 24882 -5914 25000 -5886
rect 24730 -6046 25000 -5914
rect 24730 -6074 24854 -6046
rect 24882 -6074 25000 -6046
rect 24730 -6206 25000 -6074
rect 24730 -6234 24854 -6206
rect 24882 -6234 25000 -6206
rect 24730 -6366 25000 -6234
rect 24730 -6394 24854 -6366
rect 24882 -6394 25000 -6366
rect 24730 -6526 25000 -6394
rect 24730 -6554 24854 -6526
rect 24882 -6554 25000 -6526
rect 24730 -6686 25000 -6554
rect 24730 -6714 24854 -6686
rect 24882 -6714 25000 -6686
rect 24730 -6846 25000 -6714
rect 24730 -6874 24854 -6846
rect 24882 -6874 25000 -6846
rect 24730 -7006 25000 -6874
rect 24730 -7034 24854 -7006
rect 24882 -7034 25000 -7006
rect 24730 -7166 25000 -7034
rect 24730 -7194 24854 -7166
rect 24882 -7194 25000 -7166
rect 24730 -7326 25000 -7194
rect 24730 -7354 24854 -7326
rect 24882 -7354 25000 -7326
rect 24730 -7486 25000 -7354
rect 24730 -7514 24854 -7486
rect 24882 -7514 25000 -7486
rect 24730 -7646 25000 -7514
rect 24730 -7674 24854 -7646
rect 24882 -7674 25000 -7646
rect 24730 -7806 25000 -7674
rect 24730 -7834 24854 -7806
rect 24882 -7834 25000 -7806
rect 24730 -7966 25000 -7834
rect 24730 -7994 24854 -7966
rect 24882 -7994 25000 -7966
rect 24730 -8126 25000 -7994
rect 24730 -8154 24854 -8126
rect 24882 -8154 25000 -8126
rect 24730 -8286 25000 -8154
rect 24730 -8314 24854 -8286
rect 24882 -8314 25000 -8286
rect 24730 -8446 25000 -8314
rect 24730 -8474 24854 -8446
rect 24882 -8474 25000 -8446
rect 24730 -8606 25000 -8474
rect 24730 -8634 24854 -8606
rect 24882 -8634 25000 -8606
rect 24730 -8766 25000 -8634
rect 24730 -8794 24854 -8766
rect 24882 -8794 25000 -8766
rect 24730 -8926 25000 -8794
rect 24730 -8954 24854 -8926
rect 24882 -8954 25000 -8926
rect 24730 -9086 25000 -8954
rect 24730 -9114 24854 -9086
rect 24882 -9114 25000 -9086
rect 24730 -9230 25000 -9114
rect 21000 -9246 25000 -9230
rect 21000 -9274 21121 -9246
rect 21149 -9274 24854 -9246
rect 24882 -9274 25000 -9246
rect 21000 -9351 25000 -9274
rect 21000 -9379 21306 -9351
rect 21334 -9379 21466 -9351
rect 21494 -9379 21626 -9351
rect 21654 -9379 21786 -9351
rect 21814 -9379 21946 -9351
rect 21974 -9379 22106 -9351
rect 22134 -9379 22266 -9351
rect 22294 -9379 22426 -9351
rect 22454 -9379 22586 -9351
rect 22614 -9379 22746 -9351
rect 22774 -9379 22906 -9351
rect 22934 -9379 23066 -9351
rect 23094 -9379 23226 -9351
rect 23254 -9379 23386 -9351
rect 23414 -9379 23546 -9351
rect 23574 -9379 23706 -9351
rect 23734 -9379 23866 -9351
rect 23894 -9379 24026 -9351
rect 24054 -9379 24186 -9351
rect 24214 -9379 24346 -9351
rect 24374 -9379 24506 -9351
rect 24534 -9379 24666 -9351
rect 24694 -9379 25000 -9351
rect 21000 -9500 25000 -9379
rect 3000 -11623 7000 -11500
rect 3000 -11651 3306 -11623
rect 3334 -11651 3466 -11623
rect 3494 -11651 3626 -11623
rect 3654 -11651 3786 -11623
rect 3814 -11651 3946 -11623
rect 3974 -11651 4106 -11623
rect 4134 -11651 4266 -11623
rect 4294 -11651 4426 -11623
rect 4454 -11651 4586 -11623
rect 4614 -11651 4746 -11623
rect 4774 -11651 4906 -11623
rect 4934 -11651 5066 -11623
rect 5094 -11651 5226 -11623
rect 5254 -11651 5386 -11623
rect 5414 -11651 5546 -11623
rect 5574 -11651 5706 -11623
rect 5734 -11651 5866 -11623
rect 5894 -11651 6026 -11623
rect 6054 -11651 6186 -11623
rect 6214 -11651 6346 -11623
rect 6374 -11651 6506 -11623
rect 6534 -11651 6666 -11623
rect 6694 -11651 7000 -11623
rect 3000 -11726 7000 -11651
rect 3000 -11754 3121 -11726
rect 3149 -11754 6854 -11726
rect 6882 -11754 7000 -11726
rect 3000 -11770 7000 -11754
rect 3000 -11886 3270 -11770
rect 3000 -11914 3121 -11886
rect 3149 -11914 3270 -11886
rect 3000 -12046 3270 -11914
rect 3000 -12074 3121 -12046
rect 3149 -12074 3270 -12046
rect 3000 -12206 3270 -12074
rect 3000 -12234 3121 -12206
rect 3149 -12234 3270 -12206
rect 3000 -12366 3270 -12234
rect 3000 -12394 3121 -12366
rect 3149 -12394 3270 -12366
rect 3000 -12526 3270 -12394
rect 3000 -12554 3121 -12526
rect 3149 -12554 3270 -12526
rect 3000 -12686 3270 -12554
rect 3000 -12714 3121 -12686
rect 3149 -12714 3270 -12686
rect 3000 -12846 3270 -12714
rect 3000 -12874 3121 -12846
rect 3149 -12874 3270 -12846
rect 3000 -13006 3270 -12874
rect 3000 -13034 3121 -13006
rect 3149 -13034 3270 -13006
rect 3000 -13166 3270 -13034
rect 3000 -13194 3121 -13166
rect 3149 -13194 3270 -13166
rect 3000 -13326 3270 -13194
rect 3000 -13354 3121 -13326
rect 3149 -13354 3270 -13326
rect 3000 -13486 3270 -13354
rect 3000 -13514 3121 -13486
rect 3149 -13514 3270 -13486
rect 3000 -13646 3270 -13514
rect 3000 -13674 3121 -13646
rect 3149 -13674 3270 -13646
rect 3000 -13806 3270 -13674
rect 3000 -13834 3121 -13806
rect 3149 -13834 3270 -13806
rect 3000 -13966 3270 -13834
rect 3000 -13994 3121 -13966
rect 3149 -13994 3270 -13966
rect 3000 -14126 3270 -13994
rect 3000 -14154 3121 -14126
rect 3149 -14154 3270 -14126
rect 3000 -14286 3270 -14154
rect 3000 -14314 3121 -14286
rect 3149 -14314 3270 -14286
rect 3000 -14446 3270 -14314
rect 3000 -14474 3121 -14446
rect 3149 -14474 3270 -14446
rect 3000 -14606 3270 -14474
rect 3000 -14634 3121 -14606
rect 3149 -14634 3270 -14606
rect 3000 -14766 3270 -14634
rect 3000 -14794 3121 -14766
rect 3149 -14794 3270 -14766
rect 3000 -14926 3270 -14794
rect 3000 -14954 3121 -14926
rect 3149 -14954 3270 -14926
rect 3000 -15086 3270 -14954
rect 3000 -15114 3121 -15086
rect 3149 -15114 3270 -15086
rect 3000 -15230 3270 -15114
rect 6730 -11886 7000 -11770
rect 6730 -11914 6854 -11886
rect 6882 -11914 7000 -11886
rect 6730 -12046 7000 -11914
rect 6730 -12074 6854 -12046
rect 6882 -12074 7000 -12046
rect 6730 -12206 7000 -12074
rect 6730 -12234 6854 -12206
rect 6882 -12234 7000 -12206
rect 6730 -12366 7000 -12234
rect 6730 -12394 6854 -12366
rect 6882 -12394 7000 -12366
rect 6730 -12526 7000 -12394
rect 6730 -12554 6854 -12526
rect 6882 -12554 7000 -12526
rect 6730 -12686 7000 -12554
rect 6730 -12714 6854 -12686
rect 6882 -12714 7000 -12686
rect 6730 -12846 7000 -12714
rect 6730 -12874 6854 -12846
rect 6882 -12874 7000 -12846
rect 6730 -13006 7000 -12874
rect 6730 -13034 6854 -13006
rect 6882 -13034 7000 -13006
rect 6730 -13166 7000 -13034
rect 6730 -13194 6854 -13166
rect 6882 -13194 7000 -13166
rect 6730 -13326 7000 -13194
rect 6730 -13354 6854 -13326
rect 6882 -13354 7000 -13326
rect 6730 -13486 7000 -13354
rect 6730 -13514 6854 -13486
rect 6882 -13514 7000 -13486
rect 6730 -13646 7000 -13514
rect 6730 -13674 6854 -13646
rect 6882 -13674 7000 -13646
rect 6730 -13806 7000 -13674
rect 6730 -13834 6854 -13806
rect 6882 -13834 7000 -13806
rect 6730 -13966 7000 -13834
rect 6730 -13994 6854 -13966
rect 6882 -13994 7000 -13966
rect 6730 -14126 7000 -13994
rect 6730 -14154 6854 -14126
rect 6882 -14154 7000 -14126
rect 6730 -14286 7000 -14154
rect 6730 -14314 6854 -14286
rect 6882 -14314 7000 -14286
rect 6730 -14446 7000 -14314
rect 6730 -14474 6854 -14446
rect 6882 -14474 7000 -14446
rect 6730 -14606 7000 -14474
rect 6730 -14634 6854 -14606
rect 6882 -14634 7000 -14606
rect 6730 -14766 7000 -14634
rect 6730 -14794 6854 -14766
rect 6882 -14794 7000 -14766
rect 6730 -14926 7000 -14794
rect 6730 -14954 6854 -14926
rect 6882 -14954 7000 -14926
rect 6730 -15086 7000 -14954
rect 6730 -15114 6854 -15086
rect 6882 -15114 7000 -15086
rect 6730 -15230 7000 -15114
rect 3000 -15246 7000 -15230
rect 3000 -15274 3121 -15246
rect 3149 -15274 6854 -15246
rect 6882 -15274 7000 -15246
rect 3000 -15351 7000 -15274
rect 3000 -15379 3306 -15351
rect 3334 -15379 3466 -15351
rect 3494 -15379 3626 -15351
rect 3654 -15379 3786 -15351
rect 3814 -15379 3946 -15351
rect 3974 -15379 4106 -15351
rect 4134 -15379 4266 -15351
rect 4294 -15379 4426 -15351
rect 4454 -15379 4586 -15351
rect 4614 -15379 4746 -15351
rect 4774 -15379 4906 -15351
rect 4934 -15379 5066 -15351
rect 5094 -15379 5226 -15351
rect 5254 -15379 5386 -15351
rect 5414 -15379 5546 -15351
rect 5574 -15379 5706 -15351
rect 5734 -15379 5866 -15351
rect 5894 -15379 6026 -15351
rect 6054 -15379 6186 -15351
rect 6214 -15379 6346 -15351
rect 6374 -15379 6506 -15351
rect 6534 -15379 6666 -15351
rect 6694 -15379 7000 -15351
rect 3000 -15500 7000 -15379
rect 9000 -11623 13000 -11500
rect 9000 -11651 9306 -11623
rect 9334 -11651 9466 -11623
rect 9494 -11651 9626 -11623
rect 9654 -11651 9786 -11623
rect 9814 -11651 9946 -11623
rect 9974 -11651 10106 -11623
rect 10134 -11651 10266 -11623
rect 10294 -11651 10426 -11623
rect 10454 -11651 10586 -11623
rect 10614 -11651 10746 -11623
rect 10774 -11651 10906 -11623
rect 10934 -11651 11066 -11623
rect 11094 -11651 11226 -11623
rect 11254 -11651 11386 -11623
rect 11414 -11651 11546 -11623
rect 11574 -11651 11706 -11623
rect 11734 -11651 11866 -11623
rect 11894 -11651 12026 -11623
rect 12054 -11651 12186 -11623
rect 12214 -11651 12346 -11623
rect 12374 -11651 12506 -11623
rect 12534 -11651 12666 -11623
rect 12694 -11651 13000 -11623
rect 9000 -11726 13000 -11651
rect 9000 -11754 9121 -11726
rect 9149 -11754 12854 -11726
rect 12882 -11754 13000 -11726
rect 9000 -11770 13000 -11754
rect 9000 -11886 9270 -11770
rect 9000 -11914 9121 -11886
rect 9149 -11914 9270 -11886
rect 9000 -12046 9270 -11914
rect 9000 -12074 9121 -12046
rect 9149 -12074 9270 -12046
rect 9000 -12206 9270 -12074
rect 9000 -12234 9121 -12206
rect 9149 -12234 9270 -12206
rect 9000 -12366 9270 -12234
rect 9000 -12394 9121 -12366
rect 9149 -12394 9270 -12366
rect 9000 -12526 9270 -12394
rect 9000 -12554 9121 -12526
rect 9149 -12554 9270 -12526
rect 9000 -12686 9270 -12554
rect 9000 -12714 9121 -12686
rect 9149 -12714 9270 -12686
rect 9000 -12846 9270 -12714
rect 9000 -12874 9121 -12846
rect 9149 -12874 9270 -12846
rect 9000 -13006 9270 -12874
rect 9000 -13034 9121 -13006
rect 9149 -13034 9270 -13006
rect 9000 -13166 9270 -13034
rect 9000 -13194 9121 -13166
rect 9149 -13194 9270 -13166
rect 9000 -13326 9270 -13194
rect 9000 -13354 9121 -13326
rect 9149 -13354 9270 -13326
rect 9000 -13486 9270 -13354
rect 9000 -13514 9121 -13486
rect 9149 -13514 9270 -13486
rect 9000 -13646 9270 -13514
rect 9000 -13674 9121 -13646
rect 9149 -13674 9270 -13646
rect 9000 -13806 9270 -13674
rect 9000 -13834 9121 -13806
rect 9149 -13834 9270 -13806
rect 9000 -13966 9270 -13834
rect 9000 -13994 9121 -13966
rect 9149 -13994 9270 -13966
rect 9000 -14126 9270 -13994
rect 9000 -14154 9121 -14126
rect 9149 -14154 9270 -14126
rect 9000 -14286 9270 -14154
rect 9000 -14314 9121 -14286
rect 9149 -14314 9270 -14286
rect 9000 -14446 9270 -14314
rect 9000 -14474 9121 -14446
rect 9149 -14474 9270 -14446
rect 9000 -14606 9270 -14474
rect 9000 -14634 9121 -14606
rect 9149 -14634 9270 -14606
rect 9000 -14766 9270 -14634
rect 9000 -14794 9121 -14766
rect 9149 -14794 9270 -14766
rect 9000 -14926 9270 -14794
rect 9000 -14954 9121 -14926
rect 9149 -14954 9270 -14926
rect 9000 -15086 9270 -14954
rect 9000 -15114 9121 -15086
rect 9149 -15114 9270 -15086
rect 9000 -15230 9270 -15114
rect 12730 -11886 13000 -11770
rect 12730 -11914 12854 -11886
rect 12882 -11914 13000 -11886
rect 12730 -12046 13000 -11914
rect 12730 -12074 12854 -12046
rect 12882 -12074 13000 -12046
rect 12730 -12206 13000 -12074
rect 12730 -12234 12854 -12206
rect 12882 -12234 13000 -12206
rect 12730 -12366 13000 -12234
rect 12730 -12394 12854 -12366
rect 12882 -12394 13000 -12366
rect 12730 -12526 13000 -12394
rect 12730 -12554 12854 -12526
rect 12882 -12554 13000 -12526
rect 12730 -12686 13000 -12554
rect 12730 -12714 12854 -12686
rect 12882 -12714 13000 -12686
rect 12730 -12846 13000 -12714
rect 12730 -12874 12854 -12846
rect 12882 -12874 13000 -12846
rect 12730 -13006 13000 -12874
rect 12730 -13034 12854 -13006
rect 12882 -13034 13000 -13006
rect 12730 -13166 13000 -13034
rect 12730 -13194 12854 -13166
rect 12882 -13194 13000 -13166
rect 12730 -13326 13000 -13194
rect 12730 -13354 12854 -13326
rect 12882 -13354 13000 -13326
rect 12730 -13486 13000 -13354
rect 12730 -13514 12854 -13486
rect 12882 -13514 13000 -13486
rect 12730 -13646 13000 -13514
rect 12730 -13674 12854 -13646
rect 12882 -13674 13000 -13646
rect 12730 -13806 13000 -13674
rect 12730 -13834 12854 -13806
rect 12882 -13834 13000 -13806
rect 12730 -13966 13000 -13834
rect 12730 -13994 12854 -13966
rect 12882 -13994 13000 -13966
rect 12730 -14126 13000 -13994
rect 12730 -14154 12854 -14126
rect 12882 -14154 13000 -14126
rect 12730 -14286 13000 -14154
rect 12730 -14314 12854 -14286
rect 12882 -14314 13000 -14286
rect 12730 -14446 13000 -14314
rect 12730 -14474 12854 -14446
rect 12882 -14474 13000 -14446
rect 12730 -14606 13000 -14474
rect 12730 -14634 12854 -14606
rect 12882 -14634 13000 -14606
rect 12730 -14766 13000 -14634
rect 12730 -14794 12854 -14766
rect 12882 -14794 13000 -14766
rect 12730 -14926 13000 -14794
rect 12730 -14954 12854 -14926
rect 12882 -14954 13000 -14926
rect 12730 -15086 13000 -14954
rect 12730 -15114 12854 -15086
rect 12882 -15114 13000 -15086
rect 12730 -15230 13000 -15114
rect 9000 -15246 13000 -15230
rect 9000 -15274 9121 -15246
rect 9149 -15274 12854 -15246
rect 12882 -15274 13000 -15246
rect 9000 -15351 13000 -15274
rect 9000 -15379 9306 -15351
rect 9334 -15379 9466 -15351
rect 9494 -15379 9626 -15351
rect 9654 -15379 9786 -15351
rect 9814 -15379 9946 -15351
rect 9974 -15379 10106 -15351
rect 10134 -15379 10266 -15351
rect 10294 -15379 10426 -15351
rect 10454 -15379 10586 -15351
rect 10614 -15379 10746 -15351
rect 10774 -15379 10906 -15351
rect 10934 -15379 11066 -15351
rect 11094 -15379 11226 -15351
rect 11254 -15379 11386 -15351
rect 11414 -15379 11546 -15351
rect 11574 -15379 11706 -15351
rect 11734 -15379 11866 -15351
rect 11894 -15379 12026 -15351
rect 12054 -15379 12186 -15351
rect 12214 -15379 12346 -15351
rect 12374 -15379 12506 -15351
rect 12534 -15379 12666 -15351
rect 12694 -15379 13000 -15351
rect 9000 -15500 13000 -15379
rect 15000 -11623 19000 -11500
rect 15000 -11651 15306 -11623
rect 15334 -11651 15466 -11623
rect 15494 -11651 15626 -11623
rect 15654 -11651 15786 -11623
rect 15814 -11651 15946 -11623
rect 15974 -11651 16106 -11623
rect 16134 -11651 16266 -11623
rect 16294 -11651 16426 -11623
rect 16454 -11651 16586 -11623
rect 16614 -11651 16746 -11623
rect 16774 -11651 16906 -11623
rect 16934 -11651 17066 -11623
rect 17094 -11651 17226 -11623
rect 17254 -11651 17386 -11623
rect 17414 -11651 17546 -11623
rect 17574 -11651 17706 -11623
rect 17734 -11651 17866 -11623
rect 17894 -11651 18026 -11623
rect 18054 -11651 18186 -11623
rect 18214 -11651 18346 -11623
rect 18374 -11651 18506 -11623
rect 18534 -11651 18666 -11623
rect 18694 -11651 19000 -11623
rect 15000 -11726 19000 -11651
rect 15000 -11754 15121 -11726
rect 15149 -11754 18854 -11726
rect 18882 -11754 19000 -11726
rect 15000 -11770 19000 -11754
rect 15000 -11886 15270 -11770
rect 15000 -11914 15121 -11886
rect 15149 -11914 15270 -11886
rect 15000 -12046 15270 -11914
rect 15000 -12074 15121 -12046
rect 15149 -12074 15270 -12046
rect 15000 -12206 15270 -12074
rect 15000 -12234 15121 -12206
rect 15149 -12234 15270 -12206
rect 15000 -12366 15270 -12234
rect 15000 -12394 15121 -12366
rect 15149 -12394 15270 -12366
rect 15000 -12526 15270 -12394
rect 15000 -12554 15121 -12526
rect 15149 -12554 15270 -12526
rect 15000 -12686 15270 -12554
rect 15000 -12714 15121 -12686
rect 15149 -12714 15270 -12686
rect 15000 -12846 15270 -12714
rect 15000 -12874 15121 -12846
rect 15149 -12874 15270 -12846
rect 15000 -13006 15270 -12874
rect 15000 -13034 15121 -13006
rect 15149 -13034 15270 -13006
rect 15000 -13166 15270 -13034
rect 15000 -13194 15121 -13166
rect 15149 -13194 15270 -13166
rect 15000 -13326 15270 -13194
rect 15000 -13354 15121 -13326
rect 15149 -13354 15270 -13326
rect 15000 -13486 15270 -13354
rect 15000 -13514 15121 -13486
rect 15149 -13514 15270 -13486
rect 15000 -13646 15270 -13514
rect 15000 -13674 15121 -13646
rect 15149 -13674 15270 -13646
rect 15000 -13806 15270 -13674
rect 15000 -13834 15121 -13806
rect 15149 -13834 15270 -13806
rect 15000 -13966 15270 -13834
rect 15000 -13994 15121 -13966
rect 15149 -13994 15270 -13966
rect 15000 -14126 15270 -13994
rect 15000 -14154 15121 -14126
rect 15149 -14154 15270 -14126
rect 15000 -14286 15270 -14154
rect 15000 -14314 15121 -14286
rect 15149 -14314 15270 -14286
rect 15000 -14446 15270 -14314
rect 15000 -14474 15121 -14446
rect 15149 -14474 15270 -14446
rect 15000 -14606 15270 -14474
rect 15000 -14634 15121 -14606
rect 15149 -14634 15270 -14606
rect 15000 -14766 15270 -14634
rect 15000 -14794 15121 -14766
rect 15149 -14794 15270 -14766
rect 15000 -14926 15270 -14794
rect 15000 -14954 15121 -14926
rect 15149 -14954 15270 -14926
rect 15000 -15086 15270 -14954
rect 15000 -15114 15121 -15086
rect 15149 -15114 15270 -15086
rect 15000 -15230 15270 -15114
rect 18730 -11886 19000 -11770
rect 18730 -11914 18854 -11886
rect 18882 -11914 19000 -11886
rect 18730 -12046 19000 -11914
rect 18730 -12074 18854 -12046
rect 18882 -12074 19000 -12046
rect 18730 -12206 19000 -12074
rect 18730 -12234 18854 -12206
rect 18882 -12234 19000 -12206
rect 18730 -12366 19000 -12234
rect 18730 -12394 18854 -12366
rect 18882 -12394 19000 -12366
rect 18730 -12526 19000 -12394
rect 18730 -12554 18854 -12526
rect 18882 -12554 19000 -12526
rect 18730 -12686 19000 -12554
rect 18730 -12714 18854 -12686
rect 18882 -12714 19000 -12686
rect 18730 -12846 19000 -12714
rect 18730 -12874 18854 -12846
rect 18882 -12874 19000 -12846
rect 18730 -13006 19000 -12874
rect 18730 -13034 18854 -13006
rect 18882 -13034 19000 -13006
rect 18730 -13166 19000 -13034
rect 18730 -13194 18854 -13166
rect 18882 -13194 19000 -13166
rect 18730 -13326 19000 -13194
rect 18730 -13354 18854 -13326
rect 18882 -13354 19000 -13326
rect 18730 -13486 19000 -13354
rect 18730 -13514 18854 -13486
rect 18882 -13514 19000 -13486
rect 18730 -13646 19000 -13514
rect 18730 -13674 18854 -13646
rect 18882 -13674 19000 -13646
rect 18730 -13806 19000 -13674
rect 18730 -13834 18854 -13806
rect 18882 -13834 19000 -13806
rect 18730 -13966 19000 -13834
rect 18730 -13994 18854 -13966
rect 18882 -13994 19000 -13966
rect 18730 -14126 19000 -13994
rect 18730 -14154 18854 -14126
rect 18882 -14154 19000 -14126
rect 18730 -14286 19000 -14154
rect 18730 -14314 18854 -14286
rect 18882 -14314 19000 -14286
rect 18730 -14446 19000 -14314
rect 18730 -14474 18854 -14446
rect 18882 -14474 19000 -14446
rect 18730 -14606 19000 -14474
rect 18730 -14634 18854 -14606
rect 18882 -14634 19000 -14606
rect 18730 -14766 19000 -14634
rect 18730 -14794 18854 -14766
rect 18882 -14794 19000 -14766
rect 18730 -14926 19000 -14794
rect 18730 -14954 18854 -14926
rect 18882 -14954 19000 -14926
rect 18730 -15086 19000 -14954
rect 18730 -15114 18854 -15086
rect 18882 -15114 19000 -15086
rect 18730 -15230 19000 -15114
rect 15000 -15246 19000 -15230
rect 15000 -15274 15121 -15246
rect 15149 -15274 18854 -15246
rect 18882 -15274 19000 -15246
rect 15000 -15351 19000 -15274
rect 15000 -15379 15306 -15351
rect 15334 -15379 15466 -15351
rect 15494 -15379 15626 -15351
rect 15654 -15379 15786 -15351
rect 15814 -15379 15946 -15351
rect 15974 -15379 16106 -15351
rect 16134 -15379 16266 -15351
rect 16294 -15379 16426 -15351
rect 16454 -15379 16586 -15351
rect 16614 -15379 16746 -15351
rect 16774 -15379 16906 -15351
rect 16934 -15379 17066 -15351
rect 17094 -15379 17226 -15351
rect 17254 -15379 17386 -15351
rect 17414 -15379 17546 -15351
rect 17574 -15379 17706 -15351
rect 17734 -15379 17866 -15351
rect 17894 -15379 18026 -15351
rect 18054 -15379 18186 -15351
rect 18214 -15379 18346 -15351
rect 18374 -15379 18506 -15351
rect 18534 -15379 18666 -15351
rect 18694 -15379 19000 -15351
rect 15000 -15500 19000 -15379
rect 21000 -11623 25000 -11500
rect 21000 -11651 21306 -11623
rect 21334 -11651 21466 -11623
rect 21494 -11651 21626 -11623
rect 21654 -11651 21786 -11623
rect 21814 -11651 21946 -11623
rect 21974 -11651 22106 -11623
rect 22134 -11651 22266 -11623
rect 22294 -11651 22426 -11623
rect 22454 -11651 22586 -11623
rect 22614 -11651 22746 -11623
rect 22774 -11651 22906 -11623
rect 22934 -11651 23066 -11623
rect 23094 -11651 23226 -11623
rect 23254 -11651 23386 -11623
rect 23414 -11651 23546 -11623
rect 23574 -11651 23706 -11623
rect 23734 -11651 23866 -11623
rect 23894 -11651 24026 -11623
rect 24054 -11651 24186 -11623
rect 24214 -11651 24346 -11623
rect 24374 -11651 24506 -11623
rect 24534 -11651 24666 -11623
rect 24694 -11651 25000 -11623
rect 21000 -11726 25000 -11651
rect 21000 -11754 21121 -11726
rect 21149 -11754 24854 -11726
rect 24882 -11754 25000 -11726
rect 21000 -11770 25000 -11754
rect 21000 -11886 21270 -11770
rect 21000 -11914 21121 -11886
rect 21149 -11914 21270 -11886
rect 21000 -12046 21270 -11914
rect 21000 -12074 21121 -12046
rect 21149 -12074 21270 -12046
rect 21000 -12206 21270 -12074
rect 21000 -12234 21121 -12206
rect 21149 -12234 21270 -12206
rect 21000 -12366 21270 -12234
rect 21000 -12394 21121 -12366
rect 21149 -12394 21270 -12366
rect 21000 -12526 21270 -12394
rect 21000 -12554 21121 -12526
rect 21149 -12554 21270 -12526
rect 21000 -12686 21270 -12554
rect 21000 -12714 21121 -12686
rect 21149 -12714 21270 -12686
rect 21000 -12846 21270 -12714
rect 21000 -12874 21121 -12846
rect 21149 -12874 21270 -12846
rect 21000 -13006 21270 -12874
rect 21000 -13034 21121 -13006
rect 21149 -13034 21270 -13006
rect 21000 -13166 21270 -13034
rect 21000 -13194 21121 -13166
rect 21149 -13194 21270 -13166
rect 21000 -13326 21270 -13194
rect 21000 -13354 21121 -13326
rect 21149 -13354 21270 -13326
rect 21000 -13486 21270 -13354
rect 21000 -13514 21121 -13486
rect 21149 -13514 21270 -13486
rect 21000 -13646 21270 -13514
rect 21000 -13674 21121 -13646
rect 21149 -13674 21270 -13646
rect 21000 -13806 21270 -13674
rect 21000 -13834 21121 -13806
rect 21149 -13834 21270 -13806
rect 21000 -13966 21270 -13834
rect 21000 -13994 21121 -13966
rect 21149 -13994 21270 -13966
rect 21000 -14126 21270 -13994
rect 21000 -14154 21121 -14126
rect 21149 -14154 21270 -14126
rect 21000 -14286 21270 -14154
rect 21000 -14314 21121 -14286
rect 21149 -14314 21270 -14286
rect 21000 -14446 21270 -14314
rect 21000 -14474 21121 -14446
rect 21149 -14474 21270 -14446
rect 21000 -14606 21270 -14474
rect 21000 -14634 21121 -14606
rect 21149 -14634 21270 -14606
rect 21000 -14766 21270 -14634
rect 21000 -14794 21121 -14766
rect 21149 -14794 21270 -14766
rect 21000 -14926 21270 -14794
rect 21000 -14954 21121 -14926
rect 21149 -14954 21270 -14926
rect 21000 -15086 21270 -14954
rect 21000 -15114 21121 -15086
rect 21149 -15114 21270 -15086
rect 21000 -15230 21270 -15114
rect 24730 -11886 25000 -11770
rect 24730 -11914 24854 -11886
rect 24882 -11914 25000 -11886
rect 24730 -12046 25000 -11914
rect 24730 -12074 24854 -12046
rect 24882 -12074 25000 -12046
rect 24730 -12206 25000 -12074
rect 24730 -12234 24854 -12206
rect 24882 -12234 25000 -12206
rect 24730 -12366 25000 -12234
rect 24730 -12394 24854 -12366
rect 24882 -12394 25000 -12366
rect 24730 -12526 25000 -12394
rect 24730 -12554 24854 -12526
rect 24882 -12554 25000 -12526
rect 24730 -12686 25000 -12554
rect 24730 -12714 24854 -12686
rect 24882 -12714 25000 -12686
rect 24730 -12846 25000 -12714
rect 24730 -12874 24854 -12846
rect 24882 -12874 25000 -12846
rect 24730 -13006 25000 -12874
rect 24730 -13034 24854 -13006
rect 24882 -13034 25000 -13006
rect 24730 -13166 25000 -13034
rect 24730 -13194 24854 -13166
rect 24882 -13194 25000 -13166
rect 24730 -13326 25000 -13194
rect 24730 -13354 24854 -13326
rect 24882 -13354 25000 -13326
rect 24730 -13486 25000 -13354
rect 24730 -13514 24854 -13486
rect 24882 -13514 25000 -13486
rect 24730 -13646 25000 -13514
rect 24730 -13674 24854 -13646
rect 24882 -13674 25000 -13646
rect 24730 -13806 25000 -13674
rect 24730 -13834 24854 -13806
rect 24882 -13834 25000 -13806
rect 24730 -13966 25000 -13834
rect 24730 -13994 24854 -13966
rect 24882 -13994 25000 -13966
rect 24730 -14126 25000 -13994
rect 24730 -14154 24854 -14126
rect 24882 -14154 25000 -14126
rect 24730 -14286 25000 -14154
rect 24730 -14314 24854 -14286
rect 24882 -14314 25000 -14286
rect 24730 -14446 25000 -14314
rect 24730 -14474 24854 -14446
rect 24882 -14474 25000 -14446
rect 24730 -14606 25000 -14474
rect 24730 -14634 24854 -14606
rect 24882 -14634 25000 -14606
rect 24730 -14766 25000 -14634
rect 24730 -14794 24854 -14766
rect 24882 -14794 25000 -14766
rect 24730 -14926 25000 -14794
rect 24730 -14954 24854 -14926
rect 24882 -14954 25000 -14926
rect 24730 -15086 25000 -14954
rect 24730 -15114 24854 -15086
rect 24882 -15114 25000 -15086
rect 24730 -15230 25000 -15114
rect 21000 -15246 25000 -15230
rect 21000 -15274 21121 -15246
rect 21149 -15274 24854 -15246
rect 24882 -15274 25000 -15246
rect 21000 -15351 25000 -15274
rect 21000 -15379 21306 -15351
rect 21334 -15379 21466 -15351
rect 21494 -15379 21626 -15351
rect 21654 -15379 21786 -15351
rect 21814 -15379 21946 -15351
rect 21974 -15379 22106 -15351
rect 22134 -15379 22266 -15351
rect 22294 -15379 22426 -15351
rect 22454 -15379 22586 -15351
rect 22614 -15379 22746 -15351
rect 22774 -15379 22906 -15351
rect 22934 -15379 23066 -15351
rect 23094 -15379 23226 -15351
rect 23254 -15379 23386 -15351
rect 23414 -15379 23546 -15351
rect 23574 -15379 23706 -15351
rect 23734 -15379 23866 -15351
rect 23894 -15379 24026 -15351
rect 24054 -15379 24186 -15351
rect 24214 -15379 24346 -15351
rect 24374 -15379 24506 -15351
rect 24534 -15379 24666 -15351
rect 24694 -15379 25000 -15351
rect 21000 -15500 25000 -15379
<< via2 >>
rect 11635 -3770 11705 -3740
rect 11775 -3930 11845 -3900
rect 8200 -4790 8230 -4760
rect 8305 -4785 8335 -4755
rect 8235 -4860 8265 -4830
rect 8520 -5370 8560 -5310
rect 3306 -5624 3334 -5623
rect 3306 -5650 3307 -5624
rect 3307 -5650 3333 -5624
rect 3333 -5650 3334 -5624
rect 3306 -5651 3334 -5650
rect 3466 -5624 3494 -5623
rect 3466 -5650 3467 -5624
rect 3467 -5650 3493 -5624
rect 3493 -5650 3494 -5624
rect 3466 -5651 3494 -5650
rect 3626 -5624 3654 -5623
rect 3626 -5650 3627 -5624
rect 3627 -5650 3653 -5624
rect 3653 -5650 3654 -5624
rect 3626 -5651 3654 -5650
rect 3786 -5624 3814 -5623
rect 3786 -5650 3787 -5624
rect 3787 -5650 3813 -5624
rect 3813 -5650 3814 -5624
rect 3786 -5651 3814 -5650
rect 3946 -5624 3974 -5623
rect 3946 -5650 3947 -5624
rect 3947 -5650 3973 -5624
rect 3973 -5650 3974 -5624
rect 3946 -5651 3974 -5650
rect 4106 -5624 4134 -5623
rect 4106 -5650 4107 -5624
rect 4107 -5650 4133 -5624
rect 4133 -5650 4134 -5624
rect 4106 -5651 4134 -5650
rect 4266 -5624 4294 -5623
rect 4266 -5650 4267 -5624
rect 4267 -5650 4293 -5624
rect 4293 -5650 4294 -5624
rect 4266 -5651 4294 -5650
rect 4426 -5624 4454 -5623
rect 4426 -5650 4427 -5624
rect 4427 -5650 4453 -5624
rect 4453 -5650 4454 -5624
rect 4426 -5651 4454 -5650
rect 4586 -5624 4614 -5623
rect 4586 -5650 4587 -5624
rect 4587 -5650 4613 -5624
rect 4613 -5650 4614 -5624
rect 4586 -5651 4614 -5650
rect 4746 -5624 4774 -5623
rect 4746 -5650 4747 -5624
rect 4747 -5650 4773 -5624
rect 4773 -5650 4774 -5624
rect 4746 -5651 4774 -5650
rect 4906 -5624 4934 -5623
rect 4906 -5650 4907 -5624
rect 4907 -5650 4933 -5624
rect 4933 -5650 4934 -5624
rect 4906 -5651 4934 -5650
rect 5066 -5624 5094 -5623
rect 5066 -5650 5067 -5624
rect 5067 -5650 5093 -5624
rect 5093 -5650 5094 -5624
rect 5066 -5651 5094 -5650
rect 5226 -5624 5254 -5623
rect 5226 -5650 5227 -5624
rect 5227 -5650 5253 -5624
rect 5253 -5650 5254 -5624
rect 5226 -5651 5254 -5650
rect 5386 -5624 5414 -5623
rect 5386 -5650 5387 -5624
rect 5387 -5650 5413 -5624
rect 5413 -5650 5414 -5624
rect 5386 -5651 5414 -5650
rect 5546 -5624 5574 -5623
rect 5546 -5650 5547 -5624
rect 5547 -5650 5573 -5624
rect 5573 -5650 5574 -5624
rect 5546 -5651 5574 -5650
rect 5706 -5624 5734 -5623
rect 5706 -5650 5707 -5624
rect 5707 -5650 5733 -5624
rect 5733 -5650 5734 -5624
rect 5706 -5651 5734 -5650
rect 5866 -5624 5894 -5623
rect 5866 -5650 5867 -5624
rect 5867 -5650 5893 -5624
rect 5893 -5650 5894 -5624
rect 5866 -5651 5894 -5650
rect 6026 -5624 6054 -5623
rect 6026 -5650 6027 -5624
rect 6027 -5650 6053 -5624
rect 6053 -5650 6054 -5624
rect 6026 -5651 6054 -5650
rect 6186 -5624 6214 -5623
rect 6186 -5650 6187 -5624
rect 6187 -5650 6213 -5624
rect 6213 -5650 6214 -5624
rect 6186 -5651 6214 -5650
rect 6346 -5624 6374 -5623
rect 6346 -5650 6347 -5624
rect 6347 -5650 6373 -5624
rect 6373 -5650 6374 -5624
rect 6346 -5651 6374 -5650
rect 6506 -5624 6534 -5623
rect 6506 -5650 6507 -5624
rect 6507 -5650 6533 -5624
rect 6533 -5650 6534 -5624
rect 6506 -5651 6534 -5650
rect 6666 -5624 6694 -5623
rect 6666 -5650 6667 -5624
rect 6667 -5650 6693 -5624
rect 6693 -5650 6694 -5624
rect 6666 -5651 6694 -5650
rect 9306 -5624 9334 -5623
rect 9306 -5650 9307 -5624
rect 9307 -5650 9333 -5624
rect 9333 -5650 9334 -5624
rect 9306 -5651 9334 -5650
rect 9466 -5624 9494 -5623
rect 9466 -5650 9467 -5624
rect 9467 -5650 9493 -5624
rect 9493 -5650 9494 -5624
rect 9466 -5651 9494 -5650
rect 9626 -5624 9654 -5623
rect 9626 -5650 9627 -5624
rect 9627 -5650 9653 -5624
rect 9653 -5650 9654 -5624
rect 9626 -5651 9654 -5650
rect 9786 -5624 9814 -5623
rect 9786 -5650 9787 -5624
rect 9787 -5650 9813 -5624
rect 9813 -5650 9814 -5624
rect 9786 -5651 9814 -5650
rect 9946 -5624 9974 -5623
rect 9946 -5650 9947 -5624
rect 9947 -5650 9973 -5624
rect 9973 -5650 9974 -5624
rect 9946 -5651 9974 -5650
rect 10106 -5624 10134 -5623
rect 10106 -5650 10107 -5624
rect 10107 -5650 10133 -5624
rect 10133 -5650 10134 -5624
rect 10106 -5651 10134 -5650
rect 10266 -5624 10294 -5623
rect 10266 -5650 10267 -5624
rect 10267 -5650 10293 -5624
rect 10293 -5650 10294 -5624
rect 10266 -5651 10294 -5650
rect 10426 -5624 10454 -5623
rect 10426 -5650 10427 -5624
rect 10427 -5650 10453 -5624
rect 10453 -5650 10454 -5624
rect 10426 -5651 10454 -5650
rect 10586 -5624 10614 -5623
rect 10586 -5650 10587 -5624
rect 10587 -5650 10613 -5624
rect 10613 -5650 10614 -5624
rect 10586 -5651 10614 -5650
rect 10746 -5624 10774 -5623
rect 10746 -5650 10747 -5624
rect 10747 -5650 10773 -5624
rect 10773 -5650 10774 -5624
rect 10746 -5651 10774 -5650
rect 10906 -5624 10934 -5623
rect 10906 -5650 10907 -5624
rect 10907 -5650 10933 -5624
rect 10933 -5650 10934 -5624
rect 10906 -5651 10934 -5650
rect 11066 -5624 11094 -5623
rect 11066 -5650 11067 -5624
rect 11067 -5650 11093 -5624
rect 11093 -5650 11094 -5624
rect 11066 -5651 11094 -5650
rect 11226 -5624 11254 -5623
rect 11226 -5650 11227 -5624
rect 11227 -5650 11253 -5624
rect 11253 -5650 11254 -5624
rect 11226 -5651 11254 -5650
rect 11386 -5624 11414 -5623
rect 11386 -5650 11387 -5624
rect 11387 -5650 11413 -5624
rect 11413 -5650 11414 -5624
rect 11386 -5651 11414 -5650
rect 11546 -5624 11574 -5623
rect 11546 -5650 11547 -5624
rect 11547 -5650 11573 -5624
rect 11573 -5650 11574 -5624
rect 11546 -5651 11574 -5650
rect 11706 -5624 11734 -5623
rect 11706 -5650 11707 -5624
rect 11707 -5650 11733 -5624
rect 11733 -5650 11734 -5624
rect 11706 -5651 11734 -5650
rect 11866 -5624 11894 -5623
rect 11866 -5650 11867 -5624
rect 11867 -5650 11893 -5624
rect 11893 -5650 11894 -5624
rect 11866 -5651 11894 -5650
rect 12026 -5624 12054 -5623
rect 12026 -5650 12027 -5624
rect 12027 -5650 12053 -5624
rect 12053 -5650 12054 -5624
rect 12026 -5651 12054 -5650
rect 12186 -5624 12214 -5623
rect 12186 -5650 12187 -5624
rect 12187 -5650 12213 -5624
rect 12213 -5650 12214 -5624
rect 12186 -5651 12214 -5650
rect 12346 -5624 12374 -5623
rect 12346 -5650 12347 -5624
rect 12347 -5650 12373 -5624
rect 12373 -5650 12374 -5624
rect 12346 -5651 12374 -5650
rect 12506 -5624 12534 -5623
rect 12506 -5650 12507 -5624
rect 12507 -5650 12533 -5624
rect 12533 -5650 12534 -5624
rect 12506 -5651 12534 -5650
rect 12666 -5624 12694 -5623
rect 12666 -5650 12667 -5624
rect 12667 -5650 12693 -5624
rect 12693 -5650 12694 -5624
rect 12666 -5651 12694 -5650
rect 3121 -5727 3149 -5726
rect 3121 -5753 3122 -5727
rect 3122 -5753 3148 -5727
rect 3148 -5753 3149 -5727
rect 3121 -5754 3149 -5753
rect 6854 -5727 6882 -5726
rect 6854 -5753 6855 -5727
rect 6855 -5753 6881 -5727
rect 6881 -5753 6882 -5727
rect 6854 -5754 6882 -5753
rect 3121 -5887 3149 -5886
rect 3121 -5913 3122 -5887
rect 3122 -5913 3148 -5887
rect 3148 -5913 3149 -5887
rect 3121 -5914 3149 -5913
rect 3121 -6047 3149 -6046
rect 3121 -6073 3122 -6047
rect 3122 -6073 3148 -6047
rect 3148 -6073 3149 -6047
rect 3121 -6074 3149 -6073
rect 3121 -6207 3149 -6206
rect 3121 -6233 3122 -6207
rect 3122 -6233 3148 -6207
rect 3148 -6233 3149 -6207
rect 3121 -6234 3149 -6233
rect 3121 -6367 3149 -6366
rect 3121 -6393 3122 -6367
rect 3122 -6393 3148 -6367
rect 3148 -6393 3149 -6367
rect 3121 -6394 3149 -6393
rect 3121 -6527 3149 -6526
rect 3121 -6553 3122 -6527
rect 3122 -6553 3148 -6527
rect 3148 -6553 3149 -6527
rect 3121 -6554 3149 -6553
rect 3121 -6687 3149 -6686
rect 3121 -6713 3122 -6687
rect 3122 -6713 3148 -6687
rect 3148 -6713 3149 -6687
rect 3121 -6714 3149 -6713
rect 3121 -6847 3149 -6846
rect 3121 -6873 3122 -6847
rect 3122 -6873 3148 -6847
rect 3148 -6873 3149 -6847
rect 3121 -6874 3149 -6873
rect 3121 -7007 3149 -7006
rect 3121 -7033 3122 -7007
rect 3122 -7033 3148 -7007
rect 3148 -7033 3149 -7007
rect 3121 -7034 3149 -7033
rect 3121 -7167 3149 -7166
rect 3121 -7193 3122 -7167
rect 3122 -7193 3148 -7167
rect 3148 -7193 3149 -7167
rect 3121 -7194 3149 -7193
rect 3121 -7327 3149 -7326
rect 3121 -7353 3122 -7327
rect 3122 -7353 3148 -7327
rect 3148 -7353 3149 -7327
rect 3121 -7354 3149 -7353
rect 3121 -7487 3149 -7486
rect 3121 -7513 3122 -7487
rect 3122 -7513 3148 -7487
rect 3148 -7513 3149 -7487
rect 3121 -7514 3149 -7513
rect 3121 -7647 3149 -7646
rect 3121 -7673 3122 -7647
rect 3122 -7673 3148 -7647
rect 3148 -7673 3149 -7647
rect 3121 -7674 3149 -7673
rect 3121 -7807 3149 -7806
rect 3121 -7833 3122 -7807
rect 3122 -7833 3148 -7807
rect 3148 -7833 3149 -7807
rect 3121 -7834 3149 -7833
rect 3121 -7967 3149 -7966
rect 3121 -7993 3122 -7967
rect 3122 -7993 3148 -7967
rect 3148 -7993 3149 -7967
rect 3121 -7994 3149 -7993
rect 3121 -8127 3149 -8126
rect 3121 -8153 3122 -8127
rect 3122 -8153 3148 -8127
rect 3148 -8153 3149 -8127
rect 3121 -8154 3149 -8153
rect 3121 -8287 3149 -8286
rect 3121 -8313 3122 -8287
rect 3122 -8313 3148 -8287
rect 3148 -8313 3149 -8287
rect 3121 -8314 3149 -8313
rect 3121 -8447 3149 -8446
rect 3121 -8473 3122 -8447
rect 3122 -8473 3148 -8447
rect 3148 -8473 3149 -8447
rect 3121 -8474 3149 -8473
rect 3121 -8607 3149 -8606
rect 3121 -8633 3122 -8607
rect 3122 -8633 3148 -8607
rect 3148 -8633 3149 -8607
rect 3121 -8634 3149 -8633
rect 3121 -8767 3149 -8766
rect 3121 -8793 3122 -8767
rect 3122 -8793 3148 -8767
rect 3148 -8793 3149 -8767
rect 3121 -8794 3149 -8793
rect 3121 -8927 3149 -8926
rect 3121 -8953 3122 -8927
rect 3122 -8953 3148 -8927
rect 3148 -8953 3149 -8927
rect 3121 -8954 3149 -8953
rect 3121 -9087 3149 -9086
rect 3121 -9113 3122 -9087
rect 3122 -9113 3148 -9087
rect 3148 -9113 3149 -9087
rect 3121 -9114 3149 -9113
rect 6854 -5887 6882 -5886
rect 6854 -5913 6855 -5887
rect 6855 -5913 6881 -5887
rect 6881 -5913 6882 -5887
rect 6854 -5914 6882 -5913
rect 6854 -6047 6882 -6046
rect 6854 -6073 6855 -6047
rect 6855 -6073 6881 -6047
rect 6881 -6073 6882 -6047
rect 6854 -6074 6882 -6073
rect 6854 -6207 6882 -6206
rect 6854 -6233 6855 -6207
rect 6855 -6233 6881 -6207
rect 6881 -6233 6882 -6207
rect 6854 -6234 6882 -6233
rect 6854 -6367 6882 -6366
rect 6854 -6393 6855 -6367
rect 6855 -6393 6881 -6367
rect 6881 -6393 6882 -6367
rect 6854 -6394 6882 -6393
rect 6854 -6527 6882 -6526
rect 6854 -6553 6855 -6527
rect 6855 -6553 6881 -6527
rect 6881 -6553 6882 -6527
rect 6854 -6554 6882 -6553
rect 6854 -6687 6882 -6686
rect 6854 -6713 6855 -6687
rect 6855 -6713 6881 -6687
rect 6881 -6713 6882 -6687
rect 6854 -6714 6882 -6713
rect 6854 -6847 6882 -6846
rect 6854 -6873 6855 -6847
rect 6855 -6873 6881 -6847
rect 6881 -6873 6882 -6847
rect 6854 -6874 6882 -6873
rect 6854 -7007 6882 -7006
rect 6854 -7033 6855 -7007
rect 6855 -7033 6881 -7007
rect 6881 -7033 6882 -7007
rect 6854 -7034 6882 -7033
rect 6854 -7167 6882 -7166
rect 6854 -7193 6855 -7167
rect 6855 -7193 6881 -7167
rect 6881 -7193 6882 -7167
rect 6854 -7194 6882 -7193
rect 6854 -7327 6882 -7326
rect 6854 -7353 6855 -7327
rect 6855 -7353 6881 -7327
rect 6881 -7353 6882 -7327
rect 6854 -7354 6882 -7353
rect 6854 -7487 6882 -7486
rect 6854 -7513 6855 -7487
rect 6855 -7513 6881 -7487
rect 6881 -7513 6882 -7487
rect 6854 -7514 6882 -7513
rect 6854 -7647 6882 -7646
rect 6854 -7673 6855 -7647
rect 6855 -7673 6881 -7647
rect 6881 -7673 6882 -7647
rect 6854 -7674 6882 -7673
rect 6854 -7807 6882 -7806
rect 6854 -7833 6855 -7807
rect 6855 -7833 6881 -7807
rect 6881 -7833 6882 -7807
rect 6854 -7834 6882 -7833
rect 6854 -7967 6882 -7966
rect 6854 -7993 6855 -7967
rect 6855 -7993 6881 -7967
rect 6881 -7993 6882 -7967
rect 6854 -7994 6882 -7993
rect 6854 -8127 6882 -8126
rect 6854 -8153 6855 -8127
rect 6855 -8153 6881 -8127
rect 6881 -8153 6882 -8127
rect 6854 -8154 6882 -8153
rect 6854 -8287 6882 -8286
rect 6854 -8313 6855 -8287
rect 6855 -8313 6881 -8287
rect 6881 -8313 6882 -8287
rect 6854 -8314 6882 -8313
rect 6854 -8447 6882 -8446
rect 6854 -8473 6855 -8447
rect 6855 -8473 6881 -8447
rect 6881 -8473 6882 -8447
rect 6854 -8474 6882 -8473
rect 6854 -8607 6882 -8606
rect 6854 -8633 6855 -8607
rect 6855 -8633 6881 -8607
rect 6881 -8633 6882 -8607
rect 6854 -8634 6882 -8633
rect 6854 -8767 6882 -8766
rect 6854 -8793 6855 -8767
rect 6855 -8793 6881 -8767
rect 6881 -8793 6882 -8767
rect 6854 -8794 6882 -8793
rect 6854 -8927 6882 -8926
rect 6854 -8953 6855 -8927
rect 6855 -8953 6881 -8927
rect 6881 -8953 6882 -8927
rect 6854 -8954 6882 -8953
rect 6854 -9087 6882 -9086
rect 6854 -9113 6855 -9087
rect 6855 -9113 6881 -9087
rect 6881 -9113 6882 -9087
rect 6854 -9114 6882 -9113
rect 3121 -9247 3149 -9246
rect 3121 -9273 3122 -9247
rect 3122 -9273 3148 -9247
rect 3148 -9273 3149 -9247
rect 3121 -9274 3149 -9273
rect 6854 -9247 6882 -9246
rect 6854 -9273 6855 -9247
rect 6855 -9273 6881 -9247
rect 6881 -9273 6882 -9247
rect 6854 -9274 6882 -9273
rect 3306 -9352 3334 -9351
rect 3306 -9378 3307 -9352
rect 3307 -9378 3333 -9352
rect 3333 -9378 3334 -9352
rect 3306 -9379 3334 -9378
rect 3466 -9352 3494 -9351
rect 3466 -9378 3467 -9352
rect 3467 -9378 3493 -9352
rect 3493 -9378 3494 -9352
rect 3466 -9379 3494 -9378
rect 3626 -9352 3654 -9351
rect 3626 -9378 3627 -9352
rect 3627 -9378 3653 -9352
rect 3653 -9378 3654 -9352
rect 3626 -9379 3654 -9378
rect 3786 -9352 3814 -9351
rect 3786 -9378 3787 -9352
rect 3787 -9378 3813 -9352
rect 3813 -9378 3814 -9352
rect 3786 -9379 3814 -9378
rect 3946 -9352 3974 -9351
rect 3946 -9378 3947 -9352
rect 3947 -9378 3973 -9352
rect 3973 -9378 3974 -9352
rect 3946 -9379 3974 -9378
rect 4106 -9352 4134 -9351
rect 4106 -9378 4107 -9352
rect 4107 -9378 4133 -9352
rect 4133 -9378 4134 -9352
rect 4106 -9379 4134 -9378
rect 4266 -9352 4294 -9351
rect 4266 -9378 4267 -9352
rect 4267 -9378 4293 -9352
rect 4293 -9378 4294 -9352
rect 4266 -9379 4294 -9378
rect 4426 -9352 4454 -9351
rect 4426 -9378 4427 -9352
rect 4427 -9378 4453 -9352
rect 4453 -9378 4454 -9352
rect 4426 -9379 4454 -9378
rect 4586 -9352 4614 -9351
rect 4586 -9378 4587 -9352
rect 4587 -9378 4613 -9352
rect 4613 -9378 4614 -9352
rect 4586 -9379 4614 -9378
rect 4746 -9352 4774 -9351
rect 4746 -9378 4747 -9352
rect 4747 -9378 4773 -9352
rect 4773 -9378 4774 -9352
rect 4746 -9379 4774 -9378
rect 4906 -9352 4934 -9351
rect 4906 -9378 4907 -9352
rect 4907 -9378 4933 -9352
rect 4933 -9378 4934 -9352
rect 4906 -9379 4934 -9378
rect 5066 -9352 5094 -9351
rect 5066 -9378 5067 -9352
rect 5067 -9378 5093 -9352
rect 5093 -9378 5094 -9352
rect 5066 -9379 5094 -9378
rect 5226 -9352 5254 -9351
rect 5226 -9378 5227 -9352
rect 5227 -9378 5253 -9352
rect 5253 -9378 5254 -9352
rect 5226 -9379 5254 -9378
rect 5386 -9352 5414 -9351
rect 5386 -9378 5387 -9352
rect 5387 -9378 5413 -9352
rect 5413 -9378 5414 -9352
rect 5386 -9379 5414 -9378
rect 5546 -9352 5574 -9351
rect 5546 -9378 5547 -9352
rect 5547 -9378 5573 -9352
rect 5573 -9378 5574 -9352
rect 5546 -9379 5574 -9378
rect 5706 -9352 5734 -9351
rect 5706 -9378 5707 -9352
rect 5707 -9378 5733 -9352
rect 5733 -9378 5734 -9352
rect 5706 -9379 5734 -9378
rect 5866 -9352 5894 -9351
rect 5866 -9378 5867 -9352
rect 5867 -9378 5893 -9352
rect 5893 -9378 5894 -9352
rect 5866 -9379 5894 -9378
rect 6026 -9352 6054 -9351
rect 6026 -9378 6027 -9352
rect 6027 -9378 6053 -9352
rect 6053 -9378 6054 -9352
rect 6026 -9379 6054 -9378
rect 6186 -9352 6214 -9351
rect 6186 -9378 6187 -9352
rect 6187 -9378 6213 -9352
rect 6213 -9378 6214 -9352
rect 6186 -9379 6214 -9378
rect 6346 -9352 6374 -9351
rect 6346 -9378 6347 -9352
rect 6347 -9378 6373 -9352
rect 6373 -9378 6374 -9352
rect 6346 -9379 6374 -9378
rect 6506 -9352 6534 -9351
rect 6506 -9378 6507 -9352
rect 6507 -9378 6533 -9352
rect 6533 -9378 6534 -9352
rect 6506 -9379 6534 -9378
rect 6666 -9352 6694 -9351
rect 6666 -9378 6667 -9352
rect 6667 -9378 6693 -9352
rect 6693 -9378 6694 -9352
rect 6666 -9379 6694 -9378
rect 9121 -5727 9149 -5726
rect 9121 -5753 9122 -5727
rect 9122 -5753 9148 -5727
rect 9148 -5753 9149 -5727
rect 9121 -5754 9149 -5753
rect 12854 -5727 12882 -5726
rect 12854 -5753 12855 -5727
rect 12855 -5753 12881 -5727
rect 12881 -5753 12882 -5727
rect 12854 -5754 12882 -5753
rect 9121 -5887 9149 -5886
rect 9121 -5913 9122 -5887
rect 9122 -5913 9148 -5887
rect 9148 -5913 9149 -5887
rect 9121 -5914 9149 -5913
rect 9121 -6047 9149 -6046
rect 9121 -6073 9122 -6047
rect 9122 -6073 9148 -6047
rect 9148 -6073 9149 -6047
rect 9121 -6074 9149 -6073
rect 9121 -6207 9149 -6206
rect 9121 -6233 9122 -6207
rect 9122 -6233 9148 -6207
rect 9148 -6233 9149 -6207
rect 9121 -6234 9149 -6233
rect 9121 -6367 9149 -6366
rect 9121 -6393 9122 -6367
rect 9122 -6393 9148 -6367
rect 9148 -6393 9149 -6367
rect 9121 -6394 9149 -6393
rect 9121 -6527 9149 -6526
rect 9121 -6553 9122 -6527
rect 9122 -6553 9148 -6527
rect 9148 -6553 9149 -6527
rect 9121 -6554 9149 -6553
rect 9121 -6687 9149 -6686
rect 9121 -6713 9122 -6687
rect 9122 -6713 9148 -6687
rect 9148 -6713 9149 -6687
rect 9121 -6714 9149 -6713
rect 9121 -6847 9149 -6846
rect 9121 -6873 9122 -6847
rect 9122 -6873 9148 -6847
rect 9148 -6873 9149 -6847
rect 9121 -6874 9149 -6873
rect 9121 -7007 9149 -7006
rect 9121 -7033 9122 -7007
rect 9122 -7033 9148 -7007
rect 9148 -7033 9149 -7007
rect 9121 -7034 9149 -7033
rect 9121 -7167 9149 -7166
rect 9121 -7193 9122 -7167
rect 9122 -7193 9148 -7167
rect 9148 -7193 9149 -7167
rect 9121 -7194 9149 -7193
rect 9121 -7327 9149 -7326
rect 9121 -7353 9122 -7327
rect 9122 -7353 9148 -7327
rect 9148 -7353 9149 -7327
rect 9121 -7354 9149 -7353
rect 9121 -7487 9149 -7486
rect 9121 -7513 9122 -7487
rect 9122 -7513 9148 -7487
rect 9148 -7513 9149 -7487
rect 9121 -7514 9149 -7513
rect 9121 -7647 9149 -7646
rect 9121 -7673 9122 -7647
rect 9122 -7673 9148 -7647
rect 9148 -7673 9149 -7647
rect 9121 -7674 9149 -7673
rect 9121 -7807 9149 -7806
rect 9121 -7833 9122 -7807
rect 9122 -7833 9148 -7807
rect 9148 -7833 9149 -7807
rect 9121 -7834 9149 -7833
rect 9121 -7967 9149 -7966
rect 9121 -7993 9122 -7967
rect 9122 -7993 9148 -7967
rect 9148 -7993 9149 -7967
rect 9121 -7994 9149 -7993
rect 9121 -8127 9149 -8126
rect 9121 -8153 9122 -8127
rect 9122 -8153 9148 -8127
rect 9148 -8153 9149 -8127
rect 9121 -8154 9149 -8153
rect 9121 -8287 9149 -8286
rect 9121 -8313 9122 -8287
rect 9122 -8313 9148 -8287
rect 9148 -8313 9149 -8287
rect 9121 -8314 9149 -8313
rect 9121 -8447 9149 -8446
rect 9121 -8473 9122 -8447
rect 9122 -8473 9148 -8447
rect 9148 -8473 9149 -8447
rect 9121 -8474 9149 -8473
rect 9121 -8607 9149 -8606
rect 9121 -8633 9122 -8607
rect 9122 -8633 9148 -8607
rect 9148 -8633 9149 -8607
rect 9121 -8634 9149 -8633
rect 9121 -8767 9149 -8766
rect 9121 -8793 9122 -8767
rect 9122 -8793 9148 -8767
rect 9148 -8793 9149 -8767
rect 9121 -8794 9149 -8793
rect 9121 -8927 9149 -8926
rect 9121 -8953 9122 -8927
rect 9122 -8953 9148 -8927
rect 9148 -8953 9149 -8927
rect 9121 -8954 9149 -8953
rect 9121 -9087 9149 -9086
rect 9121 -9113 9122 -9087
rect 9122 -9113 9148 -9087
rect 9148 -9113 9149 -9087
rect 9121 -9114 9149 -9113
rect 12854 -5887 12882 -5886
rect 12854 -5913 12855 -5887
rect 12855 -5913 12881 -5887
rect 12881 -5913 12882 -5887
rect 12854 -5914 12882 -5913
rect 12854 -6047 12882 -6046
rect 12854 -6073 12855 -6047
rect 12855 -6073 12881 -6047
rect 12881 -6073 12882 -6047
rect 12854 -6074 12882 -6073
rect 12854 -6207 12882 -6206
rect 12854 -6233 12855 -6207
rect 12855 -6233 12881 -6207
rect 12881 -6233 12882 -6207
rect 12854 -6234 12882 -6233
rect 12854 -6367 12882 -6366
rect 12854 -6393 12855 -6367
rect 12855 -6393 12881 -6367
rect 12881 -6393 12882 -6367
rect 12854 -6394 12882 -6393
rect 12854 -6527 12882 -6526
rect 12854 -6553 12855 -6527
rect 12855 -6553 12881 -6527
rect 12881 -6553 12882 -6527
rect 12854 -6554 12882 -6553
rect 12854 -6687 12882 -6686
rect 12854 -6713 12855 -6687
rect 12855 -6713 12881 -6687
rect 12881 -6713 12882 -6687
rect 12854 -6714 12882 -6713
rect 12854 -6847 12882 -6846
rect 12854 -6873 12855 -6847
rect 12855 -6873 12881 -6847
rect 12881 -6873 12882 -6847
rect 12854 -6874 12882 -6873
rect 12854 -7007 12882 -7006
rect 12854 -7033 12855 -7007
rect 12855 -7033 12881 -7007
rect 12881 -7033 12882 -7007
rect 12854 -7034 12882 -7033
rect 12854 -7167 12882 -7166
rect 12854 -7193 12855 -7167
rect 12855 -7193 12881 -7167
rect 12881 -7193 12882 -7167
rect 12854 -7194 12882 -7193
rect 12854 -7327 12882 -7326
rect 12854 -7353 12855 -7327
rect 12855 -7353 12881 -7327
rect 12881 -7353 12882 -7327
rect 12854 -7354 12882 -7353
rect 12854 -7487 12882 -7486
rect 12854 -7513 12855 -7487
rect 12855 -7513 12881 -7487
rect 12881 -7513 12882 -7487
rect 12854 -7514 12882 -7513
rect 12854 -7647 12882 -7646
rect 12854 -7673 12855 -7647
rect 12855 -7673 12881 -7647
rect 12881 -7673 12882 -7647
rect 12854 -7674 12882 -7673
rect 12854 -7807 12882 -7806
rect 12854 -7833 12855 -7807
rect 12855 -7833 12881 -7807
rect 12881 -7833 12882 -7807
rect 12854 -7834 12882 -7833
rect 12854 -7967 12882 -7966
rect 12854 -7993 12855 -7967
rect 12855 -7993 12881 -7967
rect 12881 -7993 12882 -7967
rect 12854 -7994 12882 -7993
rect 12854 -8127 12882 -8126
rect 12854 -8153 12855 -8127
rect 12855 -8153 12881 -8127
rect 12881 -8153 12882 -8127
rect 12854 -8154 12882 -8153
rect 12854 -8287 12882 -8286
rect 12854 -8313 12855 -8287
rect 12855 -8313 12881 -8287
rect 12881 -8313 12882 -8287
rect 12854 -8314 12882 -8313
rect 12854 -8447 12882 -8446
rect 12854 -8473 12855 -8447
rect 12855 -8473 12881 -8447
rect 12881 -8473 12882 -8447
rect 12854 -8474 12882 -8473
rect 12854 -8607 12882 -8606
rect 12854 -8633 12855 -8607
rect 12855 -8633 12881 -8607
rect 12881 -8633 12882 -8607
rect 12854 -8634 12882 -8633
rect 12854 -8767 12882 -8766
rect 12854 -8793 12855 -8767
rect 12855 -8793 12881 -8767
rect 12881 -8793 12882 -8767
rect 12854 -8794 12882 -8793
rect 12854 -8927 12882 -8926
rect 12854 -8953 12855 -8927
rect 12855 -8953 12881 -8927
rect 12881 -8953 12882 -8927
rect 12854 -8954 12882 -8953
rect 12854 -9087 12882 -9086
rect 12854 -9113 12855 -9087
rect 12855 -9113 12881 -9087
rect 12881 -9113 12882 -9087
rect 12854 -9114 12882 -9113
rect 9121 -9247 9149 -9246
rect 9121 -9273 9122 -9247
rect 9122 -9273 9148 -9247
rect 9148 -9273 9149 -9247
rect 9121 -9274 9149 -9273
rect 12854 -9247 12882 -9246
rect 12854 -9273 12855 -9247
rect 12855 -9273 12881 -9247
rect 12881 -9273 12882 -9247
rect 12854 -9274 12882 -9273
rect 9306 -9352 9334 -9351
rect 9306 -9378 9307 -9352
rect 9307 -9378 9333 -9352
rect 9333 -9378 9334 -9352
rect 9306 -9379 9334 -9378
rect 9466 -9352 9494 -9351
rect 9466 -9378 9467 -9352
rect 9467 -9378 9493 -9352
rect 9493 -9378 9494 -9352
rect 9466 -9379 9494 -9378
rect 9626 -9352 9654 -9351
rect 9626 -9378 9627 -9352
rect 9627 -9378 9653 -9352
rect 9653 -9378 9654 -9352
rect 9626 -9379 9654 -9378
rect 9786 -9352 9814 -9351
rect 9786 -9378 9787 -9352
rect 9787 -9378 9813 -9352
rect 9813 -9378 9814 -9352
rect 9786 -9379 9814 -9378
rect 9946 -9352 9974 -9351
rect 9946 -9378 9947 -9352
rect 9947 -9378 9973 -9352
rect 9973 -9378 9974 -9352
rect 9946 -9379 9974 -9378
rect 10106 -9352 10134 -9351
rect 10106 -9378 10107 -9352
rect 10107 -9378 10133 -9352
rect 10133 -9378 10134 -9352
rect 10106 -9379 10134 -9378
rect 10266 -9352 10294 -9351
rect 10266 -9378 10267 -9352
rect 10267 -9378 10293 -9352
rect 10293 -9378 10294 -9352
rect 10266 -9379 10294 -9378
rect 10426 -9352 10454 -9351
rect 10426 -9378 10427 -9352
rect 10427 -9378 10453 -9352
rect 10453 -9378 10454 -9352
rect 10426 -9379 10454 -9378
rect 10586 -9352 10614 -9351
rect 10586 -9378 10587 -9352
rect 10587 -9378 10613 -9352
rect 10613 -9378 10614 -9352
rect 10586 -9379 10614 -9378
rect 10746 -9352 10774 -9351
rect 10746 -9378 10747 -9352
rect 10747 -9378 10773 -9352
rect 10773 -9378 10774 -9352
rect 10746 -9379 10774 -9378
rect 10906 -9352 10934 -9351
rect 10906 -9378 10907 -9352
rect 10907 -9378 10933 -9352
rect 10933 -9378 10934 -9352
rect 10906 -9379 10934 -9378
rect 11066 -9352 11094 -9351
rect 11066 -9378 11067 -9352
rect 11067 -9378 11093 -9352
rect 11093 -9378 11094 -9352
rect 11066 -9379 11094 -9378
rect 11226 -9352 11254 -9351
rect 11226 -9378 11227 -9352
rect 11227 -9378 11253 -9352
rect 11253 -9378 11254 -9352
rect 11226 -9379 11254 -9378
rect 11386 -9352 11414 -9351
rect 11386 -9378 11387 -9352
rect 11387 -9378 11413 -9352
rect 11413 -9378 11414 -9352
rect 11386 -9379 11414 -9378
rect 11546 -9352 11574 -9351
rect 11546 -9378 11547 -9352
rect 11547 -9378 11573 -9352
rect 11573 -9378 11574 -9352
rect 11546 -9379 11574 -9378
rect 11706 -9352 11734 -9351
rect 11706 -9378 11707 -9352
rect 11707 -9378 11733 -9352
rect 11733 -9378 11734 -9352
rect 11706 -9379 11734 -9378
rect 11866 -9352 11894 -9351
rect 11866 -9378 11867 -9352
rect 11867 -9378 11893 -9352
rect 11893 -9378 11894 -9352
rect 11866 -9379 11894 -9378
rect 12026 -9352 12054 -9351
rect 12026 -9378 12027 -9352
rect 12027 -9378 12053 -9352
rect 12053 -9378 12054 -9352
rect 12026 -9379 12054 -9378
rect 12186 -9352 12214 -9351
rect 12186 -9378 12187 -9352
rect 12187 -9378 12213 -9352
rect 12213 -9378 12214 -9352
rect 12186 -9379 12214 -9378
rect 12346 -9352 12374 -9351
rect 12346 -9378 12347 -9352
rect 12347 -9378 12373 -9352
rect 12373 -9378 12374 -9352
rect 12346 -9379 12374 -9378
rect 12506 -9352 12534 -9351
rect 12506 -9378 12507 -9352
rect 12507 -9378 12533 -9352
rect 12533 -9378 12534 -9352
rect 12506 -9379 12534 -9378
rect 12666 -9352 12694 -9351
rect 12666 -9378 12667 -9352
rect 12667 -9378 12693 -9352
rect 12693 -9378 12694 -9352
rect 12666 -9379 12694 -9378
rect 15306 -5624 15334 -5623
rect 15306 -5650 15307 -5624
rect 15307 -5650 15333 -5624
rect 15333 -5650 15334 -5624
rect 15306 -5651 15334 -5650
rect 15466 -5624 15494 -5623
rect 15466 -5650 15467 -5624
rect 15467 -5650 15493 -5624
rect 15493 -5650 15494 -5624
rect 15466 -5651 15494 -5650
rect 15626 -5624 15654 -5623
rect 15626 -5650 15627 -5624
rect 15627 -5650 15653 -5624
rect 15653 -5650 15654 -5624
rect 15626 -5651 15654 -5650
rect 15786 -5624 15814 -5623
rect 15786 -5650 15787 -5624
rect 15787 -5650 15813 -5624
rect 15813 -5650 15814 -5624
rect 15786 -5651 15814 -5650
rect 15946 -5624 15974 -5623
rect 15946 -5650 15947 -5624
rect 15947 -5650 15973 -5624
rect 15973 -5650 15974 -5624
rect 15946 -5651 15974 -5650
rect 16106 -5624 16134 -5623
rect 16106 -5650 16107 -5624
rect 16107 -5650 16133 -5624
rect 16133 -5650 16134 -5624
rect 16106 -5651 16134 -5650
rect 16266 -5624 16294 -5623
rect 16266 -5650 16267 -5624
rect 16267 -5650 16293 -5624
rect 16293 -5650 16294 -5624
rect 16266 -5651 16294 -5650
rect 16426 -5624 16454 -5623
rect 16426 -5650 16427 -5624
rect 16427 -5650 16453 -5624
rect 16453 -5650 16454 -5624
rect 16426 -5651 16454 -5650
rect 16586 -5624 16614 -5623
rect 16586 -5650 16587 -5624
rect 16587 -5650 16613 -5624
rect 16613 -5650 16614 -5624
rect 16586 -5651 16614 -5650
rect 16746 -5624 16774 -5623
rect 16746 -5650 16747 -5624
rect 16747 -5650 16773 -5624
rect 16773 -5650 16774 -5624
rect 16746 -5651 16774 -5650
rect 16906 -5624 16934 -5623
rect 16906 -5650 16907 -5624
rect 16907 -5650 16933 -5624
rect 16933 -5650 16934 -5624
rect 16906 -5651 16934 -5650
rect 17066 -5624 17094 -5623
rect 17066 -5650 17067 -5624
rect 17067 -5650 17093 -5624
rect 17093 -5650 17094 -5624
rect 17066 -5651 17094 -5650
rect 17226 -5624 17254 -5623
rect 17226 -5650 17227 -5624
rect 17227 -5650 17253 -5624
rect 17253 -5650 17254 -5624
rect 17226 -5651 17254 -5650
rect 17386 -5624 17414 -5623
rect 17386 -5650 17387 -5624
rect 17387 -5650 17413 -5624
rect 17413 -5650 17414 -5624
rect 17386 -5651 17414 -5650
rect 17546 -5624 17574 -5623
rect 17546 -5650 17547 -5624
rect 17547 -5650 17573 -5624
rect 17573 -5650 17574 -5624
rect 17546 -5651 17574 -5650
rect 17706 -5624 17734 -5623
rect 17706 -5650 17707 -5624
rect 17707 -5650 17733 -5624
rect 17733 -5650 17734 -5624
rect 17706 -5651 17734 -5650
rect 17866 -5624 17894 -5623
rect 17866 -5650 17867 -5624
rect 17867 -5650 17893 -5624
rect 17893 -5650 17894 -5624
rect 17866 -5651 17894 -5650
rect 18026 -5624 18054 -5623
rect 18026 -5650 18027 -5624
rect 18027 -5650 18053 -5624
rect 18053 -5650 18054 -5624
rect 18026 -5651 18054 -5650
rect 18186 -5624 18214 -5623
rect 18186 -5650 18187 -5624
rect 18187 -5650 18213 -5624
rect 18213 -5650 18214 -5624
rect 18186 -5651 18214 -5650
rect 18346 -5624 18374 -5623
rect 18346 -5650 18347 -5624
rect 18347 -5650 18373 -5624
rect 18373 -5650 18374 -5624
rect 18346 -5651 18374 -5650
rect 18506 -5624 18534 -5623
rect 18506 -5650 18507 -5624
rect 18507 -5650 18533 -5624
rect 18533 -5650 18534 -5624
rect 18506 -5651 18534 -5650
rect 18666 -5624 18694 -5623
rect 18666 -5650 18667 -5624
rect 18667 -5650 18693 -5624
rect 18693 -5650 18694 -5624
rect 18666 -5651 18694 -5650
rect 15121 -5727 15149 -5726
rect 15121 -5753 15122 -5727
rect 15122 -5753 15148 -5727
rect 15148 -5753 15149 -5727
rect 15121 -5754 15149 -5753
rect 18854 -5727 18882 -5726
rect 18854 -5753 18855 -5727
rect 18855 -5753 18881 -5727
rect 18881 -5753 18882 -5727
rect 18854 -5754 18882 -5753
rect 15121 -5887 15149 -5886
rect 15121 -5913 15122 -5887
rect 15122 -5913 15148 -5887
rect 15148 -5913 15149 -5887
rect 15121 -5914 15149 -5913
rect 15121 -6047 15149 -6046
rect 15121 -6073 15122 -6047
rect 15122 -6073 15148 -6047
rect 15148 -6073 15149 -6047
rect 15121 -6074 15149 -6073
rect 15121 -6207 15149 -6206
rect 15121 -6233 15122 -6207
rect 15122 -6233 15148 -6207
rect 15148 -6233 15149 -6207
rect 15121 -6234 15149 -6233
rect 15121 -6367 15149 -6366
rect 15121 -6393 15122 -6367
rect 15122 -6393 15148 -6367
rect 15148 -6393 15149 -6367
rect 15121 -6394 15149 -6393
rect 15121 -6527 15149 -6526
rect 15121 -6553 15122 -6527
rect 15122 -6553 15148 -6527
rect 15148 -6553 15149 -6527
rect 15121 -6554 15149 -6553
rect 15121 -6687 15149 -6686
rect 15121 -6713 15122 -6687
rect 15122 -6713 15148 -6687
rect 15148 -6713 15149 -6687
rect 15121 -6714 15149 -6713
rect 15121 -6847 15149 -6846
rect 15121 -6873 15122 -6847
rect 15122 -6873 15148 -6847
rect 15148 -6873 15149 -6847
rect 15121 -6874 15149 -6873
rect 15121 -7007 15149 -7006
rect 15121 -7033 15122 -7007
rect 15122 -7033 15148 -7007
rect 15148 -7033 15149 -7007
rect 15121 -7034 15149 -7033
rect 15121 -7167 15149 -7166
rect 15121 -7193 15122 -7167
rect 15122 -7193 15148 -7167
rect 15148 -7193 15149 -7167
rect 15121 -7194 15149 -7193
rect 15121 -7327 15149 -7326
rect 15121 -7353 15122 -7327
rect 15122 -7353 15148 -7327
rect 15148 -7353 15149 -7327
rect 15121 -7354 15149 -7353
rect 15121 -7487 15149 -7486
rect 15121 -7513 15122 -7487
rect 15122 -7513 15148 -7487
rect 15148 -7513 15149 -7487
rect 15121 -7514 15149 -7513
rect 15121 -7647 15149 -7646
rect 15121 -7673 15122 -7647
rect 15122 -7673 15148 -7647
rect 15148 -7673 15149 -7647
rect 15121 -7674 15149 -7673
rect 15121 -7807 15149 -7806
rect 15121 -7833 15122 -7807
rect 15122 -7833 15148 -7807
rect 15148 -7833 15149 -7807
rect 15121 -7834 15149 -7833
rect 15121 -7967 15149 -7966
rect 15121 -7993 15122 -7967
rect 15122 -7993 15148 -7967
rect 15148 -7993 15149 -7967
rect 15121 -7994 15149 -7993
rect 15121 -8127 15149 -8126
rect 15121 -8153 15122 -8127
rect 15122 -8153 15148 -8127
rect 15148 -8153 15149 -8127
rect 15121 -8154 15149 -8153
rect 15121 -8287 15149 -8286
rect 15121 -8313 15122 -8287
rect 15122 -8313 15148 -8287
rect 15148 -8313 15149 -8287
rect 15121 -8314 15149 -8313
rect 15121 -8447 15149 -8446
rect 15121 -8473 15122 -8447
rect 15122 -8473 15148 -8447
rect 15148 -8473 15149 -8447
rect 15121 -8474 15149 -8473
rect 15121 -8607 15149 -8606
rect 15121 -8633 15122 -8607
rect 15122 -8633 15148 -8607
rect 15148 -8633 15149 -8607
rect 15121 -8634 15149 -8633
rect 15121 -8767 15149 -8766
rect 15121 -8793 15122 -8767
rect 15122 -8793 15148 -8767
rect 15148 -8793 15149 -8767
rect 15121 -8794 15149 -8793
rect 15121 -8927 15149 -8926
rect 15121 -8953 15122 -8927
rect 15122 -8953 15148 -8927
rect 15148 -8953 15149 -8927
rect 15121 -8954 15149 -8953
rect 15121 -9087 15149 -9086
rect 15121 -9113 15122 -9087
rect 15122 -9113 15148 -9087
rect 15148 -9113 15149 -9087
rect 15121 -9114 15149 -9113
rect 18854 -5887 18882 -5886
rect 18854 -5913 18855 -5887
rect 18855 -5913 18881 -5887
rect 18881 -5913 18882 -5887
rect 18854 -5914 18882 -5913
rect 18854 -6047 18882 -6046
rect 18854 -6073 18855 -6047
rect 18855 -6073 18881 -6047
rect 18881 -6073 18882 -6047
rect 18854 -6074 18882 -6073
rect 18854 -6207 18882 -6206
rect 18854 -6233 18855 -6207
rect 18855 -6233 18881 -6207
rect 18881 -6233 18882 -6207
rect 18854 -6234 18882 -6233
rect 18854 -6367 18882 -6366
rect 18854 -6393 18855 -6367
rect 18855 -6393 18881 -6367
rect 18881 -6393 18882 -6367
rect 18854 -6394 18882 -6393
rect 18854 -6527 18882 -6526
rect 18854 -6553 18855 -6527
rect 18855 -6553 18881 -6527
rect 18881 -6553 18882 -6527
rect 18854 -6554 18882 -6553
rect 18854 -6687 18882 -6686
rect 18854 -6713 18855 -6687
rect 18855 -6713 18881 -6687
rect 18881 -6713 18882 -6687
rect 18854 -6714 18882 -6713
rect 18854 -6847 18882 -6846
rect 18854 -6873 18855 -6847
rect 18855 -6873 18881 -6847
rect 18881 -6873 18882 -6847
rect 18854 -6874 18882 -6873
rect 18854 -7007 18882 -7006
rect 18854 -7033 18855 -7007
rect 18855 -7033 18881 -7007
rect 18881 -7033 18882 -7007
rect 18854 -7034 18882 -7033
rect 18854 -7167 18882 -7166
rect 18854 -7193 18855 -7167
rect 18855 -7193 18881 -7167
rect 18881 -7193 18882 -7167
rect 18854 -7194 18882 -7193
rect 18854 -7327 18882 -7326
rect 18854 -7353 18855 -7327
rect 18855 -7353 18881 -7327
rect 18881 -7353 18882 -7327
rect 18854 -7354 18882 -7353
rect 18854 -7487 18882 -7486
rect 18854 -7513 18855 -7487
rect 18855 -7513 18881 -7487
rect 18881 -7513 18882 -7487
rect 18854 -7514 18882 -7513
rect 18854 -7647 18882 -7646
rect 18854 -7673 18855 -7647
rect 18855 -7673 18881 -7647
rect 18881 -7673 18882 -7647
rect 18854 -7674 18882 -7673
rect 18854 -7807 18882 -7806
rect 18854 -7833 18855 -7807
rect 18855 -7833 18881 -7807
rect 18881 -7833 18882 -7807
rect 18854 -7834 18882 -7833
rect 18854 -7967 18882 -7966
rect 18854 -7993 18855 -7967
rect 18855 -7993 18881 -7967
rect 18881 -7993 18882 -7967
rect 18854 -7994 18882 -7993
rect 18854 -8127 18882 -8126
rect 18854 -8153 18855 -8127
rect 18855 -8153 18881 -8127
rect 18881 -8153 18882 -8127
rect 18854 -8154 18882 -8153
rect 18854 -8287 18882 -8286
rect 18854 -8313 18855 -8287
rect 18855 -8313 18881 -8287
rect 18881 -8313 18882 -8287
rect 18854 -8314 18882 -8313
rect 18854 -8447 18882 -8446
rect 18854 -8473 18855 -8447
rect 18855 -8473 18881 -8447
rect 18881 -8473 18882 -8447
rect 18854 -8474 18882 -8473
rect 18854 -8607 18882 -8606
rect 18854 -8633 18855 -8607
rect 18855 -8633 18881 -8607
rect 18881 -8633 18882 -8607
rect 18854 -8634 18882 -8633
rect 18854 -8767 18882 -8766
rect 18854 -8793 18855 -8767
rect 18855 -8793 18881 -8767
rect 18881 -8793 18882 -8767
rect 18854 -8794 18882 -8793
rect 18854 -8927 18882 -8926
rect 18854 -8953 18855 -8927
rect 18855 -8953 18881 -8927
rect 18881 -8953 18882 -8927
rect 18854 -8954 18882 -8953
rect 18854 -9087 18882 -9086
rect 18854 -9113 18855 -9087
rect 18855 -9113 18881 -9087
rect 18881 -9113 18882 -9087
rect 18854 -9114 18882 -9113
rect 15121 -9247 15149 -9246
rect 15121 -9273 15122 -9247
rect 15122 -9273 15148 -9247
rect 15148 -9273 15149 -9247
rect 15121 -9274 15149 -9273
rect 18854 -9247 18882 -9246
rect 18854 -9273 18855 -9247
rect 18855 -9273 18881 -9247
rect 18881 -9273 18882 -9247
rect 18854 -9274 18882 -9273
rect 15306 -9352 15334 -9351
rect 15306 -9378 15307 -9352
rect 15307 -9378 15333 -9352
rect 15333 -9378 15334 -9352
rect 15306 -9379 15334 -9378
rect 15466 -9352 15494 -9351
rect 15466 -9378 15467 -9352
rect 15467 -9378 15493 -9352
rect 15493 -9378 15494 -9352
rect 15466 -9379 15494 -9378
rect 15626 -9352 15654 -9351
rect 15626 -9378 15627 -9352
rect 15627 -9378 15653 -9352
rect 15653 -9378 15654 -9352
rect 15626 -9379 15654 -9378
rect 15786 -9352 15814 -9351
rect 15786 -9378 15787 -9352
rect 15787 -9378 15813 -9352
rect 15813 -9378 15814 -9352
rect 15786 -9379 15814 -9378
rect 15946 -9352 15974 -9351
rect 15946 -9378 15947 -9352
rect 15947 -9378 15973 -9352
rect 15973 -9378 15974 -9352
rect 15946 -9379 15974 -9378
rect 16106 -9352 16134 -9351
rect 16106 -9378 16107 -9352
rect 16107 -9378 16133 -9352
rect 16133 -9378 16134 -9352
rect 16106 -9379 16134 -9378
rect 16266 -9352 16294 -9351
rect 16266 -9378 16267 -9352
rect 16267 -9378 16293 -9352
rect 16293 -9378 16294 -9352
rect 16266 -9379 16294 -9378
rect 16426 -9352 16454 -9351
rect 16426 -9378 16427 -9352
rect 16427 -9378 16453 -9352
rect 16453 -9378 16454 -9352
rect 16426 -9379 16454 -9378
rect 16586 -9352 16614 -9351
rect 16586 -9378 16587 -9352
rect 16587 -9378 16613 -9352
rect 16613 -9378 16614 -9352
rect 16586 -9379 16614 -9378
rect 16746 -9352 16774 -9351
rect 16746 -9378 16747 -9352
rect 16747 -9378 16773 -9352
rect 16773 -9378 16774 -9352
rect 16746 -9379 16774 -9378
rect 16906 -9352 16934 -9351
rect 16906 -9378 16907 -9352
rect 16907 -9378 16933 -9352
rect 16933 -9378 16934 -9352
rect 16906 -9379 16934 -9378
rect 17066 -9352 17094 -9351
rect 17066 -9378 17067 -9352
rect 17067 -9378 17093 -9352
rect 17093 -9378 17094 -9352
rect 17066 -9379 17094 -9378
rect 17226 -9352 17254 -9351
rect 17226 -9378 17227 -9352
rect 17227 -9378 17253 -9352
rect 17253 -9378 17254 -9352
rect 17226 -9379 17254 -9378
rect 17386 -9352 17414 -9351
rect 17386 -9378 17387 -9352
rect 17387 -9378 17413 -9352
rect 17413 -9378 17414 -9352
rect 17386 -9379 17414 -9378
rect 17546 -9352 17574 -9351
rect 17546 -9378 17547 -9352
rect 17547 -9378 17573 -9352
rect 17573 -9378 17574 -9352
rect 17546 -9379 17574 -9378
rect 17706 -9352 17734 -9351
rect 17706 -9378 17707 -9352
rect 17707 -9378 17733 -9352
rect 17733 -9378 17734 -9352
rect 17706 -9379 17734 -9378
rect 17866 -9352 17894 -9351
rect 17866 -9378 17867 -9352
rect 17867 -9378 17893 -9352
rect 17893 -9378 17894 -9352
rect 17866 -9379 17894 -9378
rect 18026 -9352 18054 -9351
rect 18026 -9378 18027 -9352
rect 18027 -9378 18053 -9352
rect 18053 -9378 18054 -9352
rect 18026 -9379 18054 -9378
rect 18186 -9352 18214 -9351
rect 18186 -9378 18187 -9352
rect 18187 -9378 18213 -9352
rect 18213 -9378 18214 -9352
rect 18186 -9379 18214 -9378
rect 18346 -9352 18374 -9351
rect 18346 -9378 18347 -9352
rect 18347 -9378 18373 -9352
rect 18373 -9378 18374 -9352
rect 18346 -9379 18374 -9378
rect 18506 -9352 18534 -9351
rect 18506 -9378 18507 -9352
rect 18507 -9378 18533 -9352
rect 18533 -9378 18534 -9352
rect 18506 -9379 18534 -9378
rect 18666 -9352 18694 -9351
rect 18666 -9378 18667 -9352
rect 18667 -9378 18693 -9352
rect 18693 -9378 18694 -9352
rect 18666 -9379 18694 -9378
rect 21306 -5624 21334 -5623
rect 21306 -5650 21307 -5624
rect 21307 -5650 21333 -5624
rect 21333 -5650 21334 -5624
rect 21306 -5651 21334 -5650
rect 21466 -5624 21494 -5623
rect 21466 -5650 21467 -5624
rect 21467 -5650 21493 -5624
rect 21493 -5650 21494 -5624
rect 21466 -5651 21494 -5650
rect 21626 -5624 21654 -5623
rect 21626 -5650 21627 -5624
rect 21627 -5650 21653 -5624
rect 21653 -5650 21654 -5624
rect 21626 -5651 21654 -5650
rect 21786 -5624 21814 -5623
rect 21786 -5650 21787 -5624
rect 21787 -5650 21813 -5624
rect 21813 -5650 21814 -5624
rect 21786 -5651 21814 -5650
rect 21946 -5624 21974 -5623
rect 21946 -5650 21947 -5624
rect 21947 -5650 21973 -5624
rect 21973 -5650 21974 -5624
rect 21946 -5651 21974 -5650
rect 22106 -5624 22134 -5623
rect 22106 -5650 22107 -5624
rect 22107 -5650 22133 -5624
rect 22133 -5650 22134 -5624
rect 22106 -5651 22134 -5650
rect 22266 -5624 22294 -5623
rect 22266 -5650 22267 -5624
rect 22267 -5650 22293 -5624
rect 22293 -5650 22294 -5624
rect 22266 -5651 22294 -5650
rect 22426 -5624 22454 -5623
rect 22426 -5650 22427 -5624
rect 22427 -5650 22453 -5624
rect 22453 -5650 22454 -5624
rect 22426 -5651 22454 -5650
rect 22586 -5624 22614 -5623
rect 22586 -5650 22587 -5624
rect 22587 -5650 22613 -5624
rect 22613 -5650 22614 -5624
rect 22586 -5651 22614 -5650
rect 22746 -5624 22774 -5623
rect 22746 -5650 22747 -5624
rect 22747 -5650 22773 -5624
rect 22773 -5650 22774 -5624
rect 22746 -5651 22774 -5650
rect 22906 -5624 22934 -5623
rect 22906 -5650 22907 -5624
rect 22907 -5650 22933 -5624
rect 22933 -5650 22934 -5624
rect 22906 -5651 22934 -5650
rect 23066 -5624 23094 -5623
rect 23066 -5650 23067 -5624
rect 23067 -5650 23093 -5624
rect 23093 -5650 23094 -5624
rect 23066 -5651 23094 -5650
rect 23226 -5624 23254 -5623
rect 23226 -5650 23227 -5624
rect 23227 -5650 23253 -5624
rect 23253 -5650 23254 -5624
rect 23226 -5651 23254 -5650
rect 23386 -5624 23414 -5623
rect 23386 -5650 23387 -5624
rect 23387 -5650 23413 -5624
rect 23413 -5650 23414 -5624
rect 23386 -5651 23414 -5650
rect 23546 -5624 23574 -5623
rect 23546 -5650 23547 -5624
rect 23547 -5650 23573 -5624
rect 23573 -5650 23574 -5624
rect 23546 -5651 23574 -5650
rect 23706 -5624 23734 -5623
rect 23706 -5650 23707 -5624
rect 23707 -5650 23733 -5624
rect 23733 -5650 23734 -5624
rect 23706 -5651 23734 -5650
rect 23866 -5624 23894 -5623
rect 23866 -5650 23867 -5624
rect 23867 -5650 23893 -5624
rect 23893 -5650 23894 -5624
rect 23866 -5651 23894 -5650
rect 24026 -5624 24054 -5623
rect 24026 -5650 24027 -5624
rect 24027 -5650 24053 -5624
rect 24053 -5650 24054 -5624
rect 24026 -5651 24054 -5650
rect 24186 -5624 24214 -5623
rect 24186 -5650 24187 -5624
rect 24187 -5650 24213 -5624
rect 24213 -5650 24214 -5624
rect 24186 -5651 24214 -5650
rect 24346 -5624 24374 -5623
rect 24346 -5650 24347 -5624
rect 24347 -5650 24373 -5624
rect 24373 -5650 24374 -5624
rect 24346 -5651 24374 -5650
rect 24506 -5624 24534 -5623
rect 24506 -5650 24507 -5624
rect 24507 -5650 24533 -5624
rect 24533 -5650 24534 -5624
rect 24506 -5651 24534 -5650
rect 24666 -5624 24694 -5623
rect 24666 -5650 24667 -5624
rect 24667 -5650 24693 -5624
rect 24693 -5650 24694 -5624
rect 24666 -5651 24694 -5650
rect 21121 -5727 21149 -5726
rect 21121 -5753 21122 -5727
rect 21122 -5753 21148 -5727
rect 21148 -5753 21149 -5727
rect 21121 -5754 21149 -5753
rect 24854 -5727 24882 -5726
rect 24854 -5753 24855 -5727
rect 24855 -5753 24881 -5727
rect 24881 -5753 24882 -5727
rect 24854 -5754 24882 -5753
rect 21121 -5887 21149 -5886
rect 21121 -5913 21122 -5887
rect 21122 -5913 21148 -5887
rect 21148 -5913 21149 -5887
rect 21121 -5914 21149 -5913
rect 21121 -6047 21149 -6046
rect 21121 -6073 21122 -6047
rect 21122 -6073 21148 -6047
rect 21148 -6073 21149 -6047
rect 21121 -6074 21149 -6073
rect 21121 -6207 21149 -6206
rect 21121 -6233 21122 -6207
rect 21122 -6233 21148 -6207
rect 21148 -6233 21149 -6207
rect 21121 -6234 21149 -6233
rect 21121 -6367 21149 -6366
rect 21121 -6393 21122 -6367
rect 21122 -6393 21148 -6367
rect 21148 -6393 21149 -6367
rect 21121 -6394 21149 -6393
rect 21121 -6527 21149 -6526
rect 21121 -6553 21122 -6527
rect 21122 -6553 21148 -6527
rect 21148 -6553 21149 -6527
rect 21121 -6554 21149 -6553
rect 21121 -6687 21149 -6686
rect 21121 -6713 21122 -6687
rect 21122 -6713 21148 -6687
rect 21148 -6713 21149 -6687
rect 21121 -6714 21149 -6713
rect 21121 -6847 21149 -6846
rect 21121 -6873 21122 -6847
rect 21122 -6873 21148 -6847
rect 21148 -6873 21149 -6847
rect 21121 -6874 21149 -6873
rect 21121 -7007 21149 -7006
rect 21121 -7033 21122 -7007
rect 21122 -7033 21148 -7007
rect 21148 -7033 21149 -7007
rect 21121 -7034 21149 -7033
rect 21121 -7167 21149 -7166
rect 21121 -7193 21122 -7167
rect 21122 -7193 21148 -7167
rect 21148 -7193 21149 -7167
rect 21121 -7194 21149 -7193
rect 21121 -7327 21149 -7326
rect 21121 -7353 21122 -7327
rect 21122 -7353 21148 -7327
rect 21148 -7353 21149 -7327
rect 21121 -7354 21149 -7353
rect 21121 -7487 21149 -7486
rect 21121 -7513 21122 -7487
rect 21122 -7513 21148 -7487
rect 21148 -7513 21149 -7487
rect 21121 -7514 21149 -7513
rect 21121 -7647 21149 -7646
rect 21121 -7673 21122 -7647
rect 21122 -7673 21148 -7647
rect 21148 -7673 21149 -7647
rect 21121 -7674 21149 -7673
rect 21121 -7807 21149 -7806
rect 21121 -7833 21122 -7807
rect 21122 -7833 21148 -7807
rect 21148 -7833 21149 -7807
rect 21121 -7834 21149 -7833
rect 21121 -7967 21149 -7966
rect 21121 -7993 21122 -7967
rect 21122 -7993 21148 -7967
rect 21148 -7993 21149 -7967
rect 21121 -7994 21149 -7993
rect 21121 -8127 21149 -8126
rect 21121 -8153 21122 -8127
rect 21122 -8153 21148 -8127
rect 21148 -8153 21149 -8127
rect 21121 -8154 21149 -8153
rect 21121 -8287 21149 -8286
rect 21121 -8313 21122 -8287
rect 21122 -8313 21148 -8287
rect 21148 -8313 21149 -8287
rect 21121 -8314 21149 -8313
rect 21121 -8447 21149 -8446
rect 21121 -8473 21122 -8447
rect 21122 -8473 21148 -8447
rect 21148 -8473 21149 -8447
rect 21121 -8474 21149 -8473
rect 21121 -8607 21149 -8606
rect 21121 -8633 21122 -8607
rect 21122 -8633 21148 -8607
rect 21148 -8633 21149 -8607
rect 21121 -8634 21149 -8633
rect 21121 -8767 21149 -8766
rect 21121 -8793 21122 -8767
rect 21122 -8793 21148 -8767
rect 21148 -8793 21149 -8767
rect 21121 -8794 21149 -8793
rect 21121 -8927 21149 -8926
rect 21121 -8953 21122 -8927
rect 21122 -8953 21148 -8927
rect 21148 -8953 21149 -8927
rect 21121 -8954 21149 -8953
rect 21121 -9087 21149 -9086
rect 21121 -9113 21122 -9087
rect 21122 -9113 21148 -9087
rect 21148 -9113 21149 -9087
rect 21121 -9114 21149 -9113
rect 24854 -5887 24882 -5886
rect 24854 -5913 24855 -5887
rect 24855 -5913 24881 -5887
rect 24881 -5913 24882 -5887
rect 24854 -5914 24882 -5913
rect 24854 -6047 24882 -6046
rect 24854 -6073 24855 -6047
rect 24855 -6073 24881 -6047
rect 24881 -6073 24882 -6047
rect 24854 -6074 24882 -6073
rect 24854 -6207 24882 -6206
rect 24854 -6233 24855 -6207
rect 24855 -6233 24881 -6207
rect 24881 -6233 24882 -6207
rect 24854 -6234 24882 -6233
rect 24854 -6367 24882 -6366
rect 24854 -6393 24855 -6367
rect 24855 -6393 24881 -6367
rect 24881 -6393 24882 -6367
rect 24854 -6394 24882 -6393
rect 24854 -6527 24882 -6526
rect 24854 -6553 24855 -6527
rect 24855 -6553 24881 -6527
rect 24881 -6553 24882 -6527
rect 24854 -6554 24882 -6553
rect 24854 -6687 24882 -6686
rect 24854 -6713 24855 -6687
rect 24855 -6713 24881 -6687
rect 24881 -6713 24882 -6687
rect 24854 -6714 24882 -6713
rect 24854 -6847 24882 -6846
rect 24854 -6873 24855 -6847
rect 24855 -6873 24881 -6847
rect 24881 -6873 24882 -6847
rect 24854 -6874 24882 -6873
rect 24854 -7007 24882 -7006
rect 24854 -7033 24855 -7007
rect 24855 -7033 24881 -7007
rect 24881 -7033 24882 -7007
rect 24854 -7034 24882 -7033
rect 24854 -7167 24882 -7166
rect 24854 -7193 24855 -7167
rect 24855 -7193 24881 -7167
rect 24881 -7193 24882 -7167
rect 24854 -7194 24882 -7193
rect 24854 -7327 24882 -7326
rect 24854 -7353 24855 -7327
rect 24855 -7353 24881 -7327
rect 24881 -7353 24882 -7327
rect 24854 -7354 24882 -7353
rect 24854 -7487 24882 -7486
rect 24854 -7513 24855 -7487
rect 24855 -7513 24881 -7487
rect 24881 -7513 24882 -7487
rect 24854 -7514 24882 -7513
rect 24854 -7647 24882 -7646
rect 24854 -7673 24855 -7647
rect 24855 -7673 24881 -7647
rect 24881 -7673 24882 -7647
rect 24854 -7674 24882 -7673
rect 24854 -7807 24882 -7806
rect 24854 -7833 24855 -7807
rect 24855 -7833 24881 -7807
rect 24881 -7833 24882 -7807
rect 24854 -7834 24882 -7833
rect 24854 -7967 24882 -7966
rect 24854 -7993 24855 -7967
rect 24855 -7993 24881 -7967
rect 24881 -7993 24882 -7967
rect 24854 -7994 24882 -7993
rect 24854 -8127 24882 -8126
rect 24854 -8153 24855 -8127
rect 24855 -8153 24881 -8127
rect 24881 -8153 24882 -8127
rect 24854 -8154 24882 -8153
rect 24854 -8287 24882 -8286
rect 24854 -8313 24855 -8287
rect 24855 -8313 24881 -8287
rect 24881 -8313 24882 -8287
rect 24854 -8314 24882 -8313
rect 24854 -8447 24882 -8446
rect 24854 -8473 24855 -8447
rect 24855 -8473 24881 -8447
rect 24881 -8473 24882 -8447
rect 24854 -8474 24882 -8473
rect 24854 -8607 24882 -8606
rect 24854 -8633 24855 -8607
rect 24855 -8633 24881 -8607
rect 24881 -8633 24882 -8607
rect 24854 -8634 24882 -8633
rect 24854 -8767 24882 -8766
rect 24854 -8793 24855 -8767
rect 24855 -8793 24881 -8767
rect 24881 -8793 24882 -8767
rect 24854 -8794 24882 -8793
rect 24854 -8927 24882 -8926
rect 24854 -8953 24855 -8927
rect 24855 -8953 24881 -8927
rect 24881 -8953 24882 -8927
rect 24854 -8954 24882 -8953
rect 24854 -9087 24882 -9086
rect 24854 -9113 24855 -9087
rect 24855 -9113 24881 -9087
rect 24881 -9113 24882 -9087
rect 24854 -9114 24882 -9113
rect 21121 -9247 21149 -9246
rect 21121 -9273 21122 -9247
rect 21122 -9273 21148 -9247
rect 21148 -9273 21149 -9247
rect 21121 -9274 21149 -9273
rect 24854 -9247 24882 -9246
rect 24854 -9273 24855 -9247
rect 24855 -9273 24881 -9247
rect 24881 -9273 24882 -9247
rect 24854 -9274 24882 -9273
rect 21306 -9352 21334 -9351
rect 21306 -9378 21307 -9352
rect 21307 -9378 21333 -9352
rect 21333 -9378 21334 -9352
rect 21306 -9379 21334 -9378
rect 21466 -9352 21494 -9351
rect 21466 -9378 21467 -9352
rect 21467 -9378 21493 -9352
rect 21493 -9378 21494 -9352
rect 21466 -9379 21494 -9378
rect 21626 -9352 21654 -9351
rect 21626 -9378 21627 -9352
rect 21627 -9378 21653 -9352
rect 21653 -9378 21654 -9352
rect 21626 -9379 21654 -9378
rect 21786 -9352 21814 -9351
rect 21786 -9378 21787 -9352
rect 21787 -9378 21813 -9352
rect 21813 -9378 21814 -9352
rect 21786 -9379 21814 -9378
rect 21946 -9352 21974 -9351
rect 21946 -9378 21947 -9352
rect 21947 -9378 21973 -9352
rect 21973 -9378 21974 -9352
rect 21946 -9379 21974 -9378
rect 22106 -9352 22134 -9351
rect 22106 -9378 22107 -9352
rect 22107 -9378 22133 -9352
rect 22133 -9378 22134 -9352
rect 22106 -9379 22134 -9378
rect 22266 -9352 22294 -9351
rect 22266 -9378 22267 -9352
rect 22267 -9378 22293 -9352
rect 22293 -9378 22294 -9352
rect 22266 -9379 22294 -9378
rect 22426 -9352 22454 -9351
rect 22426 -9378 22427 -9352
rect 22427 -9378 22453 -9352
rect 22453 -9378 22454 -9352
rect 22426 -9379 22454 -9378
rect 22586 -9352 22614 -9351
rect 22586 -9378 22587 -9352
rect 22587 -9378 22613 -9352
rect 22613 -9378 22614 -9352
rect 22586 -9379 22614 -9378
rect 22746 -9352 22774 -9351
rect 22746 -9378 22747 -9352
rect 22747 -9378 22773 -9352
rect 22773 -9378 22774 -9352
rect 22746 -9379 22774 -9378
rect 22906 -9352 22934 -9351
rect 22906 -9378 22907 -9352
rect 22907 -9378 22933 -9352
rect 22933 -9378 22934 -9352
rect 22906 -9379 22934 -9378
rect 23066 -9352 23094 -9351
rect 23066 -9378 23067 -9352
rect 23067 -9378 23093 -9352
rect 23093 -9378 23094 -9352
rect 23066 -9379 23094 -9378
rect 23226 -9352 23254 -9351
rect 23226 -9378 23227 -9352
rect 23227 -9378 23253 -9352
rect 23253 -9378 23254 -9352
rect 23226 -9379 23254 -9378
rect 23386 -9352 23414 -9351
rect 23386 -9378 23387 -9352
rect 23387 -9378 23413 -9352
rect 23413 -9378 23414 -9352
rect 23386 -9379 23414 -9378
rect 23546 -9352 23574 -9351
rect 23546 -9378 23547 -9352
rect 23547 -9378 23573 -9352
rect 23573 -9378 23574 -9352
rect 23546 -9379 23574 -9378
rect 23706 -9352 23734 -9351
rect 23706 -9378 23707 -9352
rect 23707 -9378 23733 -9352
rect 23733 -9378 23734 -9352
rect 23706 -9379 23734 -9378
rect 23866 -9352 23894 -9351
rect 23866 -9378 23867 -9352
rect 23867 -9378 23893 -9352
rect 23893 -9378 23894 -9352
rect 23866 -9379 23894 -9378
rect 24026 -9352 24054 -9351
rect 24026 -9378 24027 -9352
rect 24027 -9378 24053 -9352
rect 24053 -9378 24054 -9352
rect 24026 -9379 24054 -9378
rect 24186 -9352 24214 -9351
rect 24186 -9378 24187 -9352
rect 24187 -9378 24213 -9352
rect 24213 -9378 24214 -9352
rect 24186 -9379 24214 -9378
rect 24346 -9352 24374 -9351
rect 24346 -9378 24347 -9352
rect 24347 -9378 24373 -9352
rect 24373 -9378 24374 -9352
rect 24346 -9379 24374 -9378
rect 24506 -9352 24534 -9351
rect 24506 -9378 24507 -9352
rect 24507 -9378 24533 -9352
rect 24533 -9378 24534 -9352
rect 24506 -9379 24534 -9378
rect 24666 -9352 24694 -9351
rect 24666 -9378 24667 -9352
rect 24667 -9378 24693 -9352
rect 24693 -9378 24694 -9352
rect 24666 -9379 24694 -9378
rect 3306 -11624 3334 -11623
rect 3306 -11650 3307 -11624
rect 3307 -11650 3333 -11624
rect 3333 -11650 3334 -11624
rect 3306 -11651 3334 -11650
rect 3466 -11624 3494 -11623
rect 3466 -11650 3467 -11624
rect 3467 -11650 3493 -11624
rect 3493 -11650 3494 -11624
rect 3466 -11651 3494 -11650
rect 3626 -11624 3654 -11623
rect 3626 -11650 3627 -11624
rect 3627 -11650 3653 -11624
rect 3653 -11650 3654 -11624
rect 3626 -11651 3654 -11650
rect 3786 -11624 3814 -11623
rect 3786 -11650 3787 -11624
rect 3787 -11650 3813 -11624
rect 3813 -11650 3814 -11624
rect 3786 -11651 3814 -11650
rect 3946 -11624 3974 -11623
rect 3946 -11650 3947 -11624
rect 3947 -11650 3973 -11624
rect 3973 -11650 3974 -11624
rect 3946 -11651 3974 -11650
rect 4106 -11624 4134 -11623
rect 4106 -11650 4107 -11624
rect 4107 -11650 4133 -11624
rect 4133 -11650 4134 -11624
rect 4106 -11651 4134 -11650
rect 4266 -11624 4294 -11623
rect 4266 -11650 4267 -11624
rect 4267 -11650 4293 -11624
rect 4293 -11650 4294 -11624
rect 4266 -11651 4294 -11650
rect 4426 -11624 4454 -11623
rect 4426 -11650 4427 -11624
rect 4427 -11650 4453 -11624
rect 4453 -11650 4454 -11624
rect 4426 -11651 4454 -11650
rect 4586 -11624 4614 -11623
rect 4586 -11650 4587 -11624
rect 4587 -11650 4613 -11624
rect 4613 -11650 4614 -11624
rect 4586 -11651 4614 -11650
rect 4746 -11624 4774 -11623
rect 4746 -11650 4747 -11624
rect 4747 -11650 4773 -11624
rect 4773 -11650 4774 -11624
rect 4746 -11651 4774 -11650
rect 4906 -11624 4934 -11623
rect 4906 -11650 4907 -11624
rect 4907 -11650 4933 -11624
rect 4933 -11650 4934 -11624
rect 4906 -11651 4934 -11650
rect 5066 -11624 5094 -11623
rect 5066 -11650 5067 -11624
rect 5067 -11650 5093 -11624
rect 5093 -11650 5094 -11624
rect 5066 -11651 5094 -11650
rect 5226 -11624 5254 -11623
rect 5226 -11650 5227 -11624
rect 5227 -11650 5253 -11624
rect 5253 -11650 5254 -11624
rect 5226 -11651 5254 -11650
rect 5386 -11624 5414 -11623
rect 5386 -11650 5387 -11624
rect 5387 -11650 5413 -11624
rect 5413 -11650 5414 -11624
rect 5386 -11651 5414 -11650
rect 5546 -11624 5574 -11623
rect 5546 -11650 5547 -11624
rect 5547 -11650 5573 -11624
rect 5573 -11650 5574 -11624
rect 5546 -11651 5574 -11650
rect 5706 -11624 5734 -11623
rect 5706 -11650 5707 -11624
rect 5707 -11650 5733 -11624
rect 5733 -11650 5734 -11624
rect 5706 -11651 5734 -11650
rect 5866 -11624 5894 -11623
rect 5866 -11650 5867 -11624
rect 5867 -11650 5893 -11624
rect 5893 -11650 5894 -11624
rect 5866 -11651 5894 -11650
rect 6026 -11624 6054 -11623
rect 6026 -11650 6027 -11624
rect 6027 -11650 6053 -11624
rect 6053 -11650 6054 -11624
rect 6026 -11651 6054 -11650
rect 6186 -11624 6214 -11623
rect 6186 -11650 6187 -11624
rect 6187 -11650 6213 -11624
rect 6213 -11650 6214 -11624
rect 6186 -11651 6214 -11650
rect 6346 -11624 6374 -11623
rect 6346 -11650 6347 -11624
rect 6347 -11650 6373 -11624
rect 6373 -11650 6374 -11624
rect 6346 -11651 6374 -11650
rect 6506 -11624 6534 -11623
rect 6506 -11650 6507 -11624
rect 6507 -11650 6533 -11624
rect 6533 -11650 6534 -11624
rect 6506 -11651 6534 -11650
rect 6666 -11624 6694 -11623
rect 6666 -11650 6667 -11624
rect 6667 -11650 6693 -11624
rect 6693 -11650 6694 -11624
rect 6666 -11651 6694 -11650
rect 3121 -11727 3149 -11726
rect 3121 -11753 3122 -11727
rect 3122 -11753 3148 -11727
rect 3148 -11753 3149 -11727
rect 3121 -11754 3149 -11753
rect 6854 -11727 6882 -11726
rect 6854 -11753 6855 -11727
rect 6855 -11753 6881 -11727
rect 6881 -11753 6882 -11727
rect 6854 -11754 6882 -11753
rect 3121 -11887 3149 -11886
rect 3121 -11913 3122 -11887
rect 3122 -11913 3148 -11887
rect 3148 -11913 3149 -11887
rect 3121 -11914 3149 -11913
rect 3121 -12047 3149 -12046
rect 3121 -12073 3122 -12047
rect 3122 -12073 3148 -12047
rect 3148 -12073 3149 -12047
rect 3121 -12074 3149 -12073
rect 3121 -12207 3149 -12206
rect 3121 -12233 3122 -12207
rect 3122 -12233 3148 -12207
rect 3148 -12233 3149 -12207
rect 3121 -12234 3149 -12233
rect 3121 -12367 3149 -12366
rect 3121 -12393 3122 -12367
rect 3122 -12393 3148 -12367
rect 3148 -12393 3149 -12367
rect 3121 -12394 3149 -12393
rect 3121 -12527 3149 -12526
rect 3121 -12553 3122 -12527
rect 3122 -12553 3148 -12527
rect 3148 -12553 3149 -12527
rect 3121 -12554 3149 -12553
rect 3121 -12687 3149 -12686
rect 3121 -12713 3122 -12687
rect 3122 -12713 3148 -12687
rect 3148 -12713 3149 -12687
rect 3121 -12714 3149 -12713
rect 3121 -12847 3149 -12846
rect 3121 -12873 3122 -12847
rect 3122 -12873 3148 -12847
rect 3148 -12873 3149 -12847
rect 3121 -12874 3149 -12873
rect 3121 -13007 3149 -13006
rect 3121 -13033 3122 -13007
rect 3122 -13033 3148 -13007
rect 3148 -13033 3149 -13007
rect 3121 -13034 3149 -13033
rect 3121 -13167 3149 -13166
rect 3121 -13193 3122 -13167
rect 3122 -13193 3148 -13167
rect 3148 -13193 3149 -13167
rect 3121 -13194 3149 -13193
rect 3121 -13327 3149 -13326
rect 3121 -13353 3122 -13327
rect 3122 -13353 3148 -13327
rect 3148 -13353 3149 -13327
rect 3121 -13354 3149 -13353
rect 3121 -13487 3149 -13486
rect 3121 -13513 3122 -13487
rect 3122 -13513 3148 -13487
rect 3148 -13513 3149 -13487
rect 3121 -13514 3149 -13513
rect 3121 -13647 3149 -13646
rect 3121 -13673 3122 -13647
rect 3122 -13673 3148 -13647
rect 3148 -13673 3149 -13647
rect 3121 -13674 3149 -13673
rect 3121 -13807 3149 -13806
rect 3121 -13833 3122 -13807
rect 3122 -13833 3148 -13807
rect 3148 -13833 3149 -13807
rect 3121 -13834 3149 -13833
rect 3121 -13967 3149 -13966
rect 3121 -13993 3122 -13967
rect 3122 -13993 3148 -13967
rect 3148 -13993 3149 -13967
rect 3121 -13994 3149 -13993
rect 3121 -14127 3149 -14126
rect 3121 -14153 3122 -14127
rect 3122 -14153 3148 -14127
rect 3148 -14153 3149 -14127
rect 3121 -14154 3149 -14153
rect 3121 -14287 3149 -14286
rect 3121 -14313 3122 -14287
rect 3122 -14313 3148 -14287
rect 3148 -14313 3149 -14287
rect 3121 -14314 3149 -14313
rect 3121 -14447 3149 -14446
rect 3121 -14473 3122 -14447
rect 3122 -14473 3148 -14447
rect 3148 -14473 3149 -14447
rect 3121 -14474 3149 -14473
rect 3121 -14607 3149 -14606
rect 3121 -14633 3122 -14607
rect 3122 -14633 3148 -14607
rect 3148 -14633 3149 -14607
rect 3121 -14634 3149 -14633
rect 3121 -14767 3149 -14766
rect 3121 -14793 3122 -14767
rect 3122 -14793 3148 -14767
rect 3148 -14793 3149 -14767
rect 3121 -14794 3149 -14793
rect 3121 -14927 3149 -14926
rect 3121 -14953 3122 -14927
rect 3122 -14953 3148 -14927
rect 3148 -14953 3149 -14927
rect 3121 -14954 3149 -14953
rect 3121 -15087 3149 -15086
rect 3121 -15113 3122 -15087
rect 3122 -15113 3148 -15087
rect 3148 -15113 3149 -15087
rect 3121 -15114 3149 -15113
rect 6854 -11887 6882 -11886
rect 6854 -11913 6855 -11887
rect 6855 -11913 6881 -11887
rect 6881 -11913 6882 -11887
rect 6854 -11914 6882 -11913
rect 6854 -12047 6882 -12046
rect 6854 -12073 6855 -12047
rect 6855 -12073 6881 -12047
rect 6881 -12073 6882 -12047
rect 6854 -12074 6882 -12073
rect 6854 -12207 6882 -12206
rect 6854 -12233 6855 -12207
rect 6855 -12233 6881 -12207
rect 6881 -12233 6882 -12207
rect 6854 -12234 6882 -12233
rect 6854 -12367 6882 -12366
rect 6854 -12393 6855 -12367
rect 6855 -12393 6881 -12367
rect 6881 -12393 6882 -12367
rect 6854 -12394 6882 -12393
rect 6854 -12527 6882 -12526
rect 6854 -12553 6855 -12527
rect 6855 -12553 6881 -12527
rect 6881 -12553 6882 -12527
rect 6854 -12554 6882 -12553
rect 6854 -12687 6882 -12686
rect 6854 -12713 6855 -12687
rect 6855 -12713 6881 -12687
rect 6881 -12713 6882 -12687
rect 6854 -12714 6882 -12713
rect 6854 -12847 6882 -12846
rect 6854 -12873 6855 -12847
rect 6855 -12873 6881 -12847
rect 6881 -12873 6882 -12847
rect 6854 -12874 6882 -12873
rect 6854 -13007 6882 -13006
rect 6854 -13033 6855 -13007
rect 6855 -13033 6881 -13007
rect 6881 -13033 6882 -13007
rect 6854 -13034 6882 -13033
rect 6854 -13167 6882 -13166
rect 6854 -13193 6855 -13167
rect 6855 -13193 6881 -13167
rect 6881 -13193 6882 -13167
rect 6854 -13194 6882 -13193
rect 6854 -13327 6882 -13326
rect 6854 -13353 6855 -13327
rect 6855 -13353 6881 -13327
rect 6881 -13353 6882 -13327
rect 6854 -13354 6882 -13353
rect 6854 -13487 6882 -13486
rect 6854 -13513 6855 -13487
rect 6855 -13513 6881 -13487
rect 6881 -13513 6882 -13487
rect 6854 -13514 6882 -13513
rect 6854 -13647 6882 -13646
rect 6854 -13673 6855 -13647
rect 6855 -13673 6881 -13647
rect 6881 -13673 6882 -13647
rect 6854 -13674 6882 -13673
rect 6854 -13807 6882 -13806
rect 6854 -13833 6855 -13807
rect 6855 -13833 6881 -13807
rect 6881 -13833 6882 -13807
rect 6854 -13834 6882 -13833
rect 6854 -13967 6882 -13966
rect 6854 -13993 6855 -13967
rect 6855 -13993 6881 -13967
rect 6881 -13993 6882 -13967
rect 6854 -13994 6882 -13993
rect 6854 -14127 6882 -14126
rect 6854 -14153 6855 -14127
rect 6855 -14153 6881 -14127
rect 6881 -14153 6882 -14127
rect 6854 -14154 6882 -14153
rect 6854 -14287 6882 -14286
rect 6854 -14313 6855 -14287
rect 6855 -14313 6881 -14287
rect 6881 -14313 6882 -14287
rect 6854 -14314 6882 -14313
rect 6854 -14447 6882 -14446
rect 6854 -14473 6855 -14447
rect 6855 -14473 6881 -14447
rect 6881 -14473 6882 -14447
rect 6854 -14474 6882 -14473
rect 6854 -14607 6882 -14606
rect 6854 -14633 6855 -14607
rect 6855 -14633 6881 -14607
rect 6881 -14633 6882 -14607
rect 6854 -14634 6882 -14633
rect 6854 -14767 6882 -14766
rect 6854 -14793 6855 -14767
rect 6855 -14793 6881 -14767
rect 6881 -14793 6882 -14767
rect 6854 -14794 6882 -14793
rect 6854 -14927 6882 -14926
rect 6854 -14953 6855 -14927
rect 6855 -14953 6881 -14927
rect 6881 -14953 6882 -14927
rect 6854 -14954 6882 -14953
rect 6854 -15087 6882 -15086
rect 6854 -15113 6855 -15087
rect 6855 -15113 6881 -15087
rect 6881 -15113 6882 -15087
rect 6854 -15114 6882 -15113
rect 3121 -15247 3149 -15246
rect 3121 -15273 3122 -15247
rect 3122 -15273 3148 -15247
rect 3148 -15273 3149 -15247
rect 3121 -15274 3149 -15273
rect 6854 -15247 6882 -15246
rect 6854 -15273 6855 -15247
rect 6855 -15273 6881 -15247
rect 6881 -15273 6882 -15247
rect 6854 -15274 6882 -15273
rect 3306 -15352 3334 -15351
rect 3306 -15378 3307 -15352
rect 3307 -15378 3333 -15352
rect 3333 -15378 3334 -15352
rect 3306 -15379 3334 -15378
rect 3466 -15352 3494 -15351
rect 3466 -15378 3467 -15352
rect 3467 -15378 3493 -15352
rect 3493 -15378 3494 -15352
rect 3466 -15379 3494 -15378
rect 3626 -15352 3654 -15351
rect 3626 -15378 3627 -15352
rect 3627 -15378 3653 -15352
rect 3653 -15378 3654 -15352
rect 3626 -15379 3654 -15378
rect 3786 -15352 3814 -15351
rect 3786 -15378 3787 -15352
rect 3787 -15378 3813 -15352
rect 3813 -15378 3814 -15352
rect 3786 -15379 3814 -15378
rect 3946 -15352 3974 -15351
rect 3946 -15378 3947 -15352
rect 3947 -15378 3973 -15352
rect 3973 -15378 3974 -15352
rect 3946 -15379 3974 -15378
rect 4106 -15352 4134 -15351
rect 4106 -15378 4107 -15352
rect 4107 -15378 4133 -15352
rect 4133 -15378 4134 -15352
rect 4106 -15379 4134 -15378
rect 4266 -15352 4294 -15351
rect 4266 -15378 4267 -15352
rect 4267 -15378 4293 -15352
rect 4293 -15378 4294 -15352
rect 4266 -15379 4294 -15378
rect 4426 -15352 4454 -15351
rect 4426 -15378 4427 -15352
rect 4427 -15378 4453 -15352
rect 4453 -15378 4454 -15352
rect 4426 -15379 4454 -15378
rect 4586 -15352 4614 -15351
rect 4586 -15378 4587 -15352
rect 4587 -15378 4613 -15352
rect 4613 -15378 4614 -15352
rect 4586 -15379 4614 -15378
rect 4746 -15352 4774 -15351
rect 4746 -15378 4747 -15352
rect 4747 -15378 4773 -15352
rect 4773 -15378 4774 -15352
rect 4746 -15379 4774 -15378
rect 4906 -15352 4934 -15351
rect 4906 -15378 4907 -15352
rect 4907 -15378 4933 -15352
rect 4933 -15378 4934 -15352
rect 4906 -15379 4934 -15378
rect 5066 -15352 5094 -15351
rect 5066 -15378 5067 -15352
rect 5067 -15378 5093 -15352
rect 5093 -15378 5094 -15352
rect 5066 -15379 5094 -15378
rect 5226 -15352 5254 -15351
rect 5226 -15378 5227 -15352
rect 5227 -15378 5253 -15352
rect 5253 -15378 5254 -15352
rect 5226 -15379 5254 -15378
rect 5386 -15352 5414 -15351
rect 5386 -15378 5387 -15352
rect 5387 -15378 5413 -15352
rect 5413 -15378 5414 -15352
rect 5386 -15379 5414 -15378
rect 5546 -15352 5574 -15351
rect 5546 -15378 5547 -15352
rect 5547 -15378 5573 -15352
rect 5573 -15378 5574 -15352
rect 5546 -15379 5574 -15378
rect 5706 -15352 5734 -15351
rect 5706 -15378 5707 -15352
rect 5707 -15378 5733 -15352
rect 5733 -15378 5734 -15352
rect 5706 -15379 5734 -15378
rect 5866 -15352 5894 -15351
rect 5866 -15378 5867 -15352
rect 5867 -15378 5893 -15352
rect 5893 -15378 5894 -15352
rect 5866 -15379 5894 -15378
rect 6026 -15352 6054 -15351
rect 6026 -15378 6027 -15352
rect 6027 -15378 6053 -15352
rect 6053 -15378 6054 -15352
rect 6026 -15379 6054 -15378
rect 6186 -15352 6214 -15351
rect 6186 -15378 6187 -15352
rect 6187 -15378 6213 -15352
rect 6213 -15378 6214 -15352
rect 6186 -15379 6214 -15378
rect 6346 -15352 6374 -15351
rect 6346 -15378 6347 -15352
rect 6347 -15378 6373 -15352
rect 6373 -15378 6374 -15352
rect 6346 -15379 6374 -15378
rect 6506 -15352 6534 -15351
rect 6506 -15378 6507 -15352
rect 6507 -15378 6533 -15352
rect 6533 -15378 6534 -15352
rect 6506 -15379 6534 -15378
rect 6666 -15352 6694 -15351
rect 6666 -15378 6667 -15352
rect 6667 -15378 6693 -15352
rect 6693 -15378 6694 -15352
rect 6666 -15379 6694 -15378
rect 9306 -11624 9334 -11623
rect 9306 -11650 9307 -11624
rect 9307 -11650 9333 -11624
rect 9333 -11650 9334 -11624
rect 9306 -11651 9334 -11650
rect 9466 -11624 9494 -11623
rect 9466 -11650 9467 -11624
rect 9467 -11650 9493 -11624
rect 9493 -11650 9494 -11624
rect 9466 -11651 9494 -11650
rect 9626 -11624 9654 -11623
rect 9626 -11650 9627 -11624
rect 9627 -11650 9653 -11624
rect 9653 -11650 9654 -11624
rect 9626 -11651 9654 -11650
rect 9786 -11624 9814 -11623
rect 9786 -11650 9787 -11624
rect 9787 -11650 9813 -11624
rect 9813 -11650 9814 -11624
rect 9786 -11651 9814 -11650
rect 9946 -11624 9974 -11623
rect 9946 -11650 9947 -11624
rect 9947 -11650 9973 -11624
rect 9973 -11650 9974 -11624
rect 9946 -11651 9974 -11650
rect 10106 -11624 10134 -11623
rect 10106 -11650 10107 -11624
rect 10107 -11650 10133 -11624
rect 10133 -11650 10134 -11624
rect 10106 -11651 10134 -11650
rect 10266 -11624 10294 -11623
rect 10266 -11650 10267 -11624
rect 10267 -11650 10293 -11624
rect 10293 -11650 10294 -11624
rect 10266 -11651 10294 -11650
rect 10426 -11624 10454 -11623
rect 10426 -11650 10427 -11624
rect 10427 -11650 10453 -11624
rect 10453 -11650 10454 -11624
rect 10426 -11651 10454 -11650
rect 10586 -11624 10614 -11623
rect 10586 -11650 10587 -11624
rect 10587 -11650 10613 -11624
rect 10613 -11650 10614 -11624
rect 10586 -11651 10614 -11650
rect 10746 -11624 10774 -11623
rect 10746 -11650 10747 -11624
rect 10747 -11650 10773 -11624
rect 10773 -11650 10774 -11624
rect 10746 -11651 10774 -11650
rect 10906 -11624 10934 -11623
rect 10906 -11650 10907 -11624
rect 10907 -11650 10933 -11624
rect 10933 -11650 10934 -11624
rect 10906 -11651 10934 -11650
rect 11066 -11624 11094 -11623
rect 11066 -11650 11067 -11624
rect 11067 -11650 11093 -11624
rect 11093 -11650 11094 -11624
rect 11066 -11651 11094 -11650
rect 11226 -11624 11254 -11623
rect 11226 -11650 11227 -11624
rect 11227 -11650 11253 -11624
rect 11253 -11650 11254 -11624
rect 11226 -11651 11254 -11650
rect 11386 -11624 11414 -11623
rect 11386 -11650 11387 -11624
rect 11387 -11650 11413 -11624
rect 11413 -11650 11414 -11624
rect 11386 -11651 11414 -11650
rect 11546 -11624 11574 -11623
rect 11546 -11650 11547 -11624
rect 11547 -11650 11573 -11624
rect 11573 -11650 11574 -11624
rect 11546 -11651 11574 -11650
rect 11706 -11624 11734 -11623
rect 11706 -11650 11707 -11624
rect 11707 -11650 11733 -11624
rect 11733 -11650 11734 -11624
rect 11706 -11651 11734 -11650
rect 11866 -11624 11894 -11623
rect 11866 -11650 11867 -11624
rect 11867 -11650 11893 -11624
rect 11893 -11650 11894 -11624
rect 11866 -11651 11894 -11650
rect 12026 -11624 12054 -11623
rect 12026 -11650 12027 -11624
rect 12027 -11650 12053 -11624
rect 12053 -11650 12054 -11624
rect 12026 -11651 12054 -11650
rect 12186 -11624 12214 -11623
rect 12186 -11650 12187 -11624
rect 12187 -11650 12213 -11624
rect 12213 -11650 12214 -11624
rect 12186 -11651 12214 -11650
rect 12346 -11624 12374 -11623
rect 12346 -11650 12347 -11624
rect 12347 -11650 12373 -11624
rect 12373 -11650 12374 -11624
rect 12346 -11651 12374 -11650
rect 12506 -11624 12534 -11623
rect 12506 -11650 12507 -11624
rect 12507 -11650 12533 -11624
rect 12533 -11650 12534 -11624
rect 12506 -11651 12534 -11650
rect 12666 -11624 12694 -11623
rect 12666 -11650 12667 -11624
rect 12667 -11650 12693 -11624
rect 12693 -11650 12694 -11624
rect 12666 -11651 12694 -11650
rect 9121 -11727 9149 -11726
rect 9121 -11753 9122 -11727
rect 9122 -11753 9148 -11727
rect 9148 -11753 9149 -11727
rect 9121 -11754 9149 -11753
rect 12854 -11727 12882 -11726
rect 12854 -11753 12855 -11727
rect 12855 -11753 12881 -11727
rect 12881 -11753 12882 -11727
rect 12854 -11754 12882 -11753
rect 9121 -11887 9149 -11886
rect 9121 -11913 9122 -11887
rect 9122 -11913 9148 -11887
rect 9148 -11913 9149 -11887
rect 9121 -11914 9149 -11913
rect 9121 -12047 9149 -12046
rect 9121 -12073 9122 -12047
rect 9122 -12073 9148 -12047
rect 9148 -12073 9149 -12047
rect 9121 -12074 9149 -12073
rect 9121 -12207 9149 -12206
rect 9121 -12233 9122 -12207
rect 9122 -12233 9148 -12207
rect 9148 -12233 9149 -12207
rect 9121 -12234 9149 -12233
rect 9121 -12367 9149 -12366
rect 9121 -12393 9122 -12367
rect 9122 -12393 9148 -12367
rect 9148 -12393 9149 -12367
rect 9121 -12394 9149 -12393
rect 9121 -12527 9149 -12526
rect 9121 -12553 9122 -12527
rect 9122 -12553 9148 -12527
rect 9148 -12553 9149 -12527
rect 9121 -12554 9149 -12553
rect 9121 -12687 9149 -12686
rect 9121 -12713 9122 -12687
rect 9122 -12713 9148 -12687
rect 9148 -12713 9149 -12687
rect 9121 -12714 9149 -12713
rect 9121 -12847 9149 -12846
rect 9121 -12873 9122 -12847
rect 9122 -12873 9148 -12847
rect 9148 -12873 9149 -12847
rect 9121 -12874 9149 -12873
rect 9121 -13007 9149 -13006
rect 9121 -13033 9122 -13007
rect 9122 -13033 9148 -13007
rect 9148 -13033 9149 -13007
rect 9121 -13034 9149 -13033
rect 9121 -13167 9149 -13166
rect 9121 -13193 9122 -13167
rect 9122 -13193 9148 -13167
rect 9148 -13193 9149 -13167
rect 9121 -13194 9149 -13193
rect 9121 -13327 9149 -13326
rect 9121 -13353 9122 -13327
rect 9122 -13353 9148 -13327
rect 9148 -13353 9149 -13327
rect 9121 -13354 9149 -13353
rect 9121 -13487 9149 -13486
rect 9121 -13513 9122 -13487
rect 9122 -13513 9148 -13487
rect 9148 -13513 9149 -13487
rect 9121 -13514 9149 -13513
rect 9121 -13647 9149 -13646
rect 9121 -13673 9122 -13647
rect 9122 -13673 9148 -13647
rect 9148 -13673 9149 -13647
rect 9121 -13674 9149 -13673
rect 9121 -13807 9149 -13806
rect 9121 -13833 9122 -13807
rect 9122 -13833 9148 -13807
rect 9148 -13833 9149 -13807
rect 9121 -13834 9149 -13833
rect 9121 -13967 9149 -13966
rect 9121 -13993 9122 -13967
rect 9122 -13993 9148 -13967
rect 9148 -13993 9149 -13967
rect 9121 -13994 9149 -13993
rect 9121 -14127 9149 -14126
rect 9121 -14153 9122 -14127
rect 9122 -14153 9148 -14127
rect 9148 -14153 9149 -14127
rect 9121 -14154 9149 -14153
rect 9121 -14287 9149 -14286
rect 9121 -14313 9122 -14287
rect 9122 -14313 9148 -14287
rect 9148 -14313 9149 -14287
rect 9121 -14314 9149 -14313
rect 9121 -14447 9149 -14446
rect 9121 -14473 9122 -14447
rect 9122 -14473 9148 -14447
rect 9148 -14473 9149 -14447
rect 9121 -14474 9149 -14473
rect 9121 -14607 9149 -14606
rect 9121 -14633 9122 -14607
rect 9122 -14633 9148 -14607
rect 9148 -14633 9149 -14607
rect 9121 -14634 9149 -14633
rect 9121 -14767 9149 -14766
rect 9121 -14793 9122 -14767
rect 9122 -14793 9148 -14767
rect 9148 -14793 9149 -14767
rect 9121 -14794 9149 -14793
rect 9121 -14927 9149 -14926
rect 9121 -14953 9122 -14927
rect 9122 -14953 9148 -14927
rect 9148 -14953 9149 -14927
rect 9121 -14954 9149 -14953
rect 9121 -15087 9149 -15086
rect 9121 -15113 9122 -15087
rect 9122 -15113 9148 -15087
rect 9148 -15113 9149 -15087
rect 9121 -15114 9149 -15113
rect 12854 -11887 12882 -11886
rect 12854 -11913 12855 -11887
rect 12855 -11913 12881 -11887
rect 12881 -11913 12882 -11887
rect 12854 -11914 12882 -11913
rect 12854 -12047 12882 -12046
rect 12854 -12073 12855 -12047
rect 12855 -12073 12881 -12047
rect 12881 -12073 12882 -12047
rect 12854 -12074 12882 -12073
rect 12854 -12207 12882 -12206
rect 12854 -12233 12855 -12207
rect 12855 -12233 12881 -12207
rect 12881 -12233 12882 -12207
rect 12854 -12234 12882 -12233
rect 12854 -12367 12882 -12366
rect 12854 -12393 12855 -12367
rect 12855 -12393 12881 -12367
rect 12881 -12393 12882 -12367
rect 12854 -12394 12882 -12393
rect 12854 -12527 12882 -12526
rect 12854 -12553 12855 -12527
rect 12855 -12553 12881 -12527
rect 12881 -12553 12882 -12527
rect 12854 -12554 12882 -12553
rect 12854 -12687 12882 -12686
rect 12854 -12713 12855 -12687
rect 12855 -12713 12881 -12687
rect 12881 -12713 12882 -12687
rect 12854 -12714 12882 -12713
rect 12854 -12847 12882 -12846
rect 12854 -12873 12855 -12847
rect 12855 -12873 12881 -12847
rect 12881 -12873 12882 -12847
rect 12854 -12874 12882 -12873
rect 12854 -13007 12882 -13006
rect 12854 -13033 12855 -13007
rect 12855 -13033 12881 -13007
rect 12881 -13033 12882 -13007
rect 12854 -13034 12882 -13033
rect 12854 -13167 12882 -13166
rect 12854 -13193 12855 -13167
rect 12855 -13193 12881 -13167
rect 12881 -13193 12882 -13167
rect 12854 -13194 12882 -13193
rect 12854 -13327 12882 -13326
rect 12854 -13353 12855 -13327
rect 12855 -13353 12881 -13327
rect 12881 -13353 12882 -13327
rect 12854 -13354 12882 -13353
rect 12854 -13487 12882 -13486
rect 12854 -13513 12855 -13487
rect 12855 -13513 12881 -13487
rect 12881 -13513 12882 -13487
rect 12854 -13514 12882 -13513
rect 12854 -13647 12882 -13646
rect 12854 -13673 12855 -13647
rect 12855 -13673 12881 -13647
rect 12881 -13673 12882 -13647
rect 12854 -13674 12882 -13673
rect 12854 -13807 12882 -13806
rect 12854 -13833 12855 -13807
rect 12855 -13833 12881 -13807
rect 12881 -13833 12882 -13807
rect 12854 -13834 12882 -13833
rect 12854 -13967 12882 -13966
rect 12854 -13993 12855 -13967
rect 12855 -13993 12881 -13967
rect 12881 -13993 12882 -13967
rect 12854 -13994 12882 -13993
rect 12854 -14127 12882 -14126
rect 12854 -14153 12855 -14127
rect 12855 -14153 12881 -14127
rect 12881 -14153 12882 -14127
rect 12854 -14154 12882 -14153
rect 12854 -14287 12882 -14286
rect 12854 -14313 12855 -14287
rect 12855 -14313 12881 -14287
rect 12881 -14313 12882 -14287
rect 12854 -14314 12882 -14313
rect 12854 -14447 12882 -14446
rect 12854 -14473 12855 -14447
rect 12855 -14473 12881 -14447
rect 12881 -14473 12882 -14447
rect 12854 -14474 12882 -14473
rect 12854 -14607 12882 -14606
rect 12854 -14633 12855 -14607
rect 12855 -14633 12881 -14607
rect 12881 -14633 12882 -14607
rect 12854 -14634 12882 -14633
rect 12854 -14767 12882 -14766
rect 12854 -14793 12855 -14767
rect 12855 -14793 12881 -14767
rect 12881 -14793 12882 -14767
rect 12854 -14794 12882 -14793
rect 12854 -14927 12882 -14926
rect 12854 -14953 12855 -14927
rect 12855 -14953 12881 -14927
rect 12881 -14953 12882 -14927
rect 12854 -14954 12882 -14953
rect 12854 -15087 12882 -15086
rect 12854 -15113 12855 -15087
rect 12855 -15113 12881 -15087
rect 12881 -15113 12882 -15087
rect 12854 -15114 12882 -15113
rect 9121 -15247 9149 -15246
rect 9121 -15273 9122 -15247
rect 9122 -15273 9148 -15247
rect 9148 -15273 9149 -15247
rect 9121 -15274 9149 -15273
rect 12854 -15247 12882 -15246
rect 12854 -15273 12855 -15247
rect 12855 -15273 12881 -15247
rect 12881 -15273 12882 -15247
rect 12854 -15274 12882 -15273
rect 9306 -15352 9334 -15351
rect 9306 -15378 9307 -15352
rect 9307 -15378 9333 -15352
rect 9333 -15378 9334 -15352
rect 9306 -15379 9334 -15378
rect 9466 -15352 9494 -15351
rect 9466 -15378 9467 -15352
rect 9467 -15378 9493 -15352
rect 9493 -15378 9494 -15352
rect 9466 -15379 9494 -15378
rect 9626 -15352 9654 -15351
rect 9626 -15378 9627 -15352
rect 9627 -15378 9653 -15352
rect 9653 -15378 9654 -15352
rect 9626 -15379 9654 -15378
rect 9786 -15352 9814 -15351
rect 9786 -15378 9787 -15352
rect 9787 -15378 9813 -15352
rect 9813 -15378 9814 -15352
rect 9786 -15379 9814 -15378
rect 9946 -15352 9974 -15351
rect 9946 -15378 9947 -15352
rect 9947 -15378 9973 -15352
rect 9973 -15378 9974 -15352
rect 9946 -15379 9974 -15378
rect 10106 -15352 10134 -15351
rect 10106 -15378 10107 -15352
rect 10107 -15378 10133 -15352
rect 10133 -15378 10134 -15352
rect 10106 -15379 10134 -15378
rect 10266 -15352 10294 -15351
rect 10266 -15378 10267 -15352
rect 10267 -15378 10293 -15352
rect 10293 -15378 10294 -15352
rect 10266 -15379 10294 -15378
rect 10426 -15352 10454 -15351
rect 10426 -15378 10427 -15352
rect 10427 -15378 10453 -15352
rect 10453 -15378 10454 -15352
rect 10426 -15379 10454 -15378
rect 10586 -15352 10614 -15351
rect 10586 -15378 10587 -15352
rect 10587 -15378 10613 -15352
rect 10613 -15378 10614 -15352
rect 10586 -15379 10614 -15378
rect 10746 -15352 10774 -15351
rect 10746 -15378 10747 -15352
rect 10747 -15378 10773 -15352
rect 10773 -15378 10774 -15352
rect 10746 -15379 10774 -15378
rect 10906 -15352 10934 -15351
rect 10906 -15378 10907 -15352
rect 10907 -15378 10933 -15352
rect 10933 -15378 10934 -15352
rect 10906 -15379 10934 -15378
rect 11066 -15352 11094 -15351
rect 11066 -15378 11067 -15352
rect 11067 -15378 11093 -15352
rect 11093 -15378 11094 -15352
rect 11066 -15379 11094 -15378
rect 11226 -15352 11254 -15351
rect 11226 -15378 11227 -15352
rect 11227 -15378 11253 -15352
rect 11253 -15378 11254 -15352
rect 11226 -15379 11254 -15378
rect 11386 -15352 11414 -15351
rect 11386 -15378 11387 -15352
rect 11387 -15378 11413 -15352
rect 11413 -15378 11414 -15352
rect 11386 -15379 11414 -15378
rect 11546 -15352 11574 -15351
rect 11546 -15378 11547 -15352
rect 11547 -15378 11573 -15352
rect 11573 -15378 11574 -15352
rect 11546 -15379 11574 -15378
rect 11706 -15352 11734 -15351
rect 11706 -15378 11707 -15352
rect 11707 -15378 11733 -15352
rect 11733 -15378 11734 -15352
rect 11706 -15379 11734 -15378
rect 11866 -15352 11894 -15351
rect 11866 -15378 11867 -15352
rect 11867 -15378 11893 -15352
rect 11893 -15378 11894 -15352
rect 11866 -15379 11894 -15378
rect 12026 -15352 12054 -15351
rect 12026 -15378 12027 -15352
rect 12027 -15378 12053 -15352
rect 12053 -15378 12054 -15352
rect 12026 -15379 12054 -15378
rect 12186 -15352 12214 -15351
rect 12186 -15378 12187 -15352
rect 12187 -15378 12213 -15352
rect 12213 -15378 12214 -15352
rect 12186 -15379 12214 -15378
rect 12346 -15352 12374 -15351
rect 12346 -15378 12347 -15352
rect 12347 -15378 12373 -15352
rect 12373 -15378 12374 -15352
rect 12346 -15379 12374 -15378
rect 12506 -15352 12534 -15351
rect 12506 -15378 12507 -15352
rect 12507 -15378 12533 -15352
rect 12533 -15378 12534 -15352
rect 12506 -15379 12534 -15378
rect 12666 -15352 12694 -15351
rect 12666 -15378 12667 -15352
rect 12667 -15378 12693 -15352
rect 12693 -15378 12694 -15352
rect 12666 -15379 12694 -15378
rect 15306 -11624 15334 -11623
rect 15306 -11650 15307 -11624
rect 15307 -11650 15333 -11624
rect 15333 -11650 15334 -11624
rect 15306 -11651 15334 -11650
rect 15466 -11624 15494 -11623
rect 15466 -11650 15467 -11624
rect 15467 -11650 15493 -11624
rect 15493 -11650 15494 -11624
rect 15466 -11651 15494 -11650
rect 15626 -11624 15654 -11623
rect 15626 -11650 15627 -11624
rect 15627 -11650 15653 -11624
rect 15653 -11650 15654 -11624
rect 15626 -11651 15654 -11650
rect 15786 -11624 15814 -11623
rect 15786 -11650 15787 -11624
rect 15787 -11650 15813 -11624
rect 15813 -11650 15814 -11624
rect 15786 -11651 15814 -11650
rect 15946 -11624 15974 -11623
rect 15946 -11650 15947 -11624
rect 15947 -11650 15973 -11624
rect 15973 -11650 15974 -11624
rect 15946 -11651 15974 -11650
rect 16106 -11624 16134 -11623
rect 16106 -11650 16107 -11624
rect 16107 -11650 16133 -11624
rect 16133 -11650 16134 -11624
rect 16106 -11651 16134 -11650
rect 16266 -11624 16294 -11623
rect 16266 -11650 16267 -11624
rect 16267 -11650 16293 -11624
rect 16293 -11650 16294 -11624
rect 16266 -11651 16294 -11650
rect 16426 -11624 16454 -11623
rect 16426 -11650 16427 -11624
rect 16427 -11650 16453 -11624
rect 16453 -11650 16454 -11624
rect 16426 -11651 16454 -11650
rect 16586 -11624 16614 -11623
rect 16586 -11650 16587 -11624
rect 16587 -11650 16613 -11624
rect 16613 -11650 16614 -11624
rect 16586 -11651 16614 -11650
rect 16746 -11624 16774 -11623
rect 16746 -11650 16747 -11624
rect 16747 -11650 16773 -11624
rect 16773 -11650 16774 -11624
rect 16746 -11651 16774 -11650
rect 16906 -11624 16934 -11623
rect 16906 -11650 16907 -11624
rect 16907 -11650 16933 -11624
rect 16933 -11650 16934 -11624
rect 16906 -11651 16934 -11650
rect 17066 -11624 17094 -11623
rect 17066 -11650 17067 -11624
rect 17067 -11650 17093 -11624
rect 17093 -11650 17094 -11624
rect 17066 -11651 17094 -11650
rect 17226 -11624 17254 -11623
rect 17226 -11650 17227 -11624
rect 17227 -11650 17253 -11624
rect 17253 -11650 17254 -11624
rect 17226 -11651 17254 -11650
rect 17386 -11624 17414 -11623
rect 17386 -11650 17387 -11624
rect 17387 -11650 17413 -11624
rect 17413 -11650 17414 -11624
rect 17386 -11651 17414 -11650
rect 17546 -11624 17574 -11623
rect 17546 -11650 17547 -11624
rect 17547 -11650 17573 -11624
rect 17573 -11650 17574 -11624
rect 17546 -11651 17574 -11650
rect 17706 -11624 17734 -11623
rect 17706 -11650 17707 -11624
rect 17707 -11650 17733 -11624
rect 17733 -11650 17734 -11624
rect 17706 -11651 17734 -11650
rect 17866 -11624 17894 -11623
rect 17866 -11650 17867 -11624
rect 17867 -11650 17893 -11624
rect 17893 -11650 17894 -11624
rect 17866 -11651 17894 -11650
rect 18026 -11624 18054 -11623
rect 18026 -11650 18027 -11624
rect 18027 -11650 18053 -11624
rect 18053 -11650 18054 -11624
rect 18026 -11651 18054 -11650
rect 18186 -11624 18214 -11623
rect 18186 -11650 18187 -11624
rect 18187 -11650 18213 -11624
rect 18213 -11650 18214 -11624
rect 18186 -11651 18214 -11650
rect 18346 -11624 18374 -11623
rect 18346 -11650 18347 -11624
rect 18347 -11650 18373 -11624
rect 18373 -11650 18374 -11624
rect 18346 -11651 18374 -11650
rect 18506 -11624 18534 -11623
rect 18506 -11650 18507 -11624
rect 18507 -11650 18533 -11624
rect 18533 -11650 18534 -11624
rect 18506 -11651 18534 -11650
rect 18666 -11624 18694 -11623
rect 18666 -11650 18667 -11624
rect 18667 -11650 18693 -11624
rect 18693 -11650 18694 -11624
rect 18666 -11651 18694 -11650
rect 15121 -11727 15149 -11726
rect 15121 -11753 15122 -11727
rect 15122 -11753 15148 -11727
rect 15148 -11753 15149 -11727
rect 15121 -11754 15149 -11753
rect 18854 -11727 18882 -11726
rect 18854 -11753 18855 -11727
rect 18855 -11753 18881 -11727
rect 18881 -11753 18882 -11727
rect 18854 -11754 18882 -11753
rect 15121 -11887 15149 -11886
rect 15121 -11913 15122 -11887
rect 15122 -11913 15148 -11887
rect 15148 -11913 15149 -11887
rect 15121 -11914 15149 -11913
rect 15121 -12047 15149 -12046
rect 15121 -12073 15122 -12047
rect 15122 -12073 15148 -12047
rect 15148 -12073 15149 -12047
rect 15121 -12074 15149 -12073
rect 15121 -12207 15149 -12206
rect 15121 -12233 15122 -12207
rect 15122 -12233 15148 -12207
rect 15148 -12233 15149 -12207
rect 15121 -12234 15149 -12233
rect 15121 -12367 15149 -12366
rect 15121 -12393 15122 -12367
rect 15122 -12393 15148 -12367
rect 15148 -12393 15149 -12367
rect 15121 -12394 15149 -12393
rect 15121 -12527 15149 -12526
rect 15121 -12553 15122 -12527
rect 15122 -12553 15148 -12527
rect 15148 -12553 15149 -12527
rect 15121 -12554 15149 -12553
rect 15121 -12687 15149 -12686
rect 15121 -12713 15122 -12687
rect 15122 -12713 15148 -12687
rect 15148 -12713 15149 -12687
rect 15121 -12714 15149 -12713
rect 15121 -12847 15149 -12846
rect 15121 -12873 15122 -12847
rect 15122 -12873 15148 -12847
rect 15148 -12873 15149 -12847
rect 15121 -12874 15149 -12873
rect 15121 -13007 15149 -13006
rect 15121 -13033 15122 -13007
rect 15122 -13033 15148 -13007
rect 15148 -13033 15149 -13007
rect 15121 -13034 15149 -13033
rect 15121 -13167 15149 -13166
rect 15121 -13193 15122 -13167
rect 15122 -13193 15148 -13167
rect 15148 -13193 15149 -13167
rect 15121 -13194 15149 -13193
rect 15121 -13327 15149 -13326
rect 15121 -13353 15122 -13327
rect 15122 -13353 15148 -13327
rect 15148 -13353 15149 -13327
rect 15121 -13354 15149 -13353
rect 15121 -13487 15149 -13486
rect 15121 -13513 15122 -13487
rect 15122 -13513 15148 -13487
rect 15148 -13513 15149 -13487
rect 15121 -13514 15149 -13513
rect 15121 -13647 15149 -13646
rect 15121 -13673 15122 -13647
rect 15122 -13673 15148 -13647
rect 15148 -13673 15149 -13647
rect 15121 -13674 15149 -13673
rect 15121 -13807 15149 -13806
rect 15121 -13833 15122 -13807
rect 15122 -13833 15148 -13807
rect 15148 -13833 15149 -13807
rect 15121 -13834 15149 -13833
rect 15121 -13967 15149 -13966
rect 15121 -13993 15122 -13967
rect 15122 -13993 15148 -13967
rect 15148 -13993 15149 -13967
rect 15121 -13994 15149 -13993
rect 15121 -14127 15149 -14126
rect 15121 -14153 15122 -14127
rect 15122 -14153 15148 -14127
rect 15148 -14153 15149 -14127
rect 15121 -14154 15149 -14153
rect 15121 -14287 15149 -14286
rect 15121 -14313 15122 -14287
rect 15122 -14313 15148 -14287
rect 15148 -14313 15149 -14287
rect 15121 -14314 15149 -14313
rect 15121 -14447 15149 -14446
rect 15121 -14473 15122 -14447
rect 15122 -14473 15148 -14447
rect 15148 -14473 15149 -14447
rect 15121 -14474 15149 -14473
rect 15121 -14607 15149 -14606
rect 15121 -14633 15122 -14607
rect 15122 -14633 15148 -14607
rect 15148 -14633 15149 -14607
rect 15121 -14634 15149 -14633
rect 15121 -14767 15149 -14766
rect 15121 -14793 15122 -14767
rect 15122 -14793 15148 -14767
rect 15148 -14793 15149 -14767
rect 15121 -14794 15149 -14793
rect 15121 -14927 15149 -14926
rect 15121 -14953 15122 -14927
rect 15122 -14953 15148 -14927
rect 15148 -14953 15149 -14927
rect 15121 -14954 15149 -14953
rect 15121 -15087 15149 -15086
rect 15121 -15113 15122 -15087
rect 15122 -15113 15148 -15087
rect 15148 -15113 15149 -15087
rect 15121 -15114 15149 -15113
rect 18854 -11887 18882 -11886
rect 18854 -11913 18855 -11887
rect 18855 -11913 18881 -11887
rect 18881 -11913 18882 -11887
rect 18854 -11914 18882 -11913
rect 18854 -12047 18882 -12046
rect 18854 -12073 18855 -12047
rect 18855 -12073 18881 -12047
rect 18881 -12073 18882 -12047
rect 18854 -12074 18882 -12073
rect 18854 -12207 18882 -12206
rect 18854 -12233 18855 -12207
rect 18855 -12233 18881 -12207
rect 18881 -12233 18882 -12207
rect 18854 -12234 18882 -12233
rect 18854 -12367 18882 -12366
rect 18854 -12393 18855 -12367
rect 18855 -12393 18881 -12367
rect 18881 -12393 18882 -12367
rect 18854 -12394 18882 -12393
rect 18854 -12527 18882 -12526
rect 18854 -12553 18855 -12527
rect 18855 -12553 18881 -12527
rect 18881 -12553 18882 -12527
rect 18854 -12554 18882 -12553
rect 18854 -12687 18882 -12686
rect 18854 -12713 18855 -12687
rect 18855 -12713 18881 -12687
rect 18881 -12713 18882 -12687
rect 18854 -12714 18882 -12713
rect 18854 -12847 18882 -12846
rect 18854 -12873 18855 -12847
rect 18855 -12873 18881 -12847
rect 18881 -12873 18882 -12847
rect 18854 -12874 18882 -12873
rect 18854 -13007 18882 -13006
rect 18854 -13033 18855 -13007
rect 18855 -13033 18881 -13007
rect 18881 -13033 18882 -13007
rect 18854 -13034 18882 -13033
rect 18854 -13167 18882 -13166
rect 18854 -13193 18855 -13167
rect 18855 -13193 18881 -13167
rect 18881 -13193 18882 -13167
rect 18854 -13194 18882 -13193
rect 18854 -13327 18882 -13326
rect 18854 -13353 18855 -13327
rect 18855 -13353 18881 -13327
rect 18881 -13353 18882 -13327
rect 18854 -13354 18882 -13353
rect 18854 -13487 18882 -13486
rect 18854 -13513 18855 -13487
rect 18855 -13513 18881 -13487
rect 18881 -13513 18882 -13487
rect 18854 -13514 18882 -13513
rect 18854 -13647 18882 -13646
rect 18854 -13673 18855 -13647
rect 18855 -13673 18881 -13647
rect 18881 -13673 18882 -13647
rect 18854 -13674 18882 -13673
rect 18854 -13807 18882 -13806
rect 18854 -13833 18855 -13807
rect 18855 -13833 18881 -13807
rect 18881 -13833 18882 -13807
rect 18854 -13834 18882 -13833
rect 18854 -13967 18882 -13966
rect 18854 -13993 18855 -13967
rect 18855 -13993 18881 -13967
rect 18881 -13993 18882 -13967
rect 18854 -13994 18882 -13993
rect 18854 -14127 18882 -14126
rect 18854 -14153 18855 -14127
rect 18855 -14153 18881 -14127
rect 18881 -14153 18882 -14127
rect 18854 -14154 18882 -14153
rect 18854 -14287 18882 -14286
rect 18854 -14313 18855 -14287
rect 18855 -14313 18881 -14287
rect 18881 -14313 18882 -14287
rect 18854 -14314 18882 -14313
rect 18854 -14447 18882 -14446
rect 18854 -14473 18855 -14447
rect 18855 -14473 18881 -14447
rect 18881 -14473 18882 -14447
rect 18854 -14474 18882 -14473
rect 18854 -14607 18882 -14606
rect 18854 -14633 18855 -14607
rect 18855 -14633 18881 -14607
rect 18881 -14633 18882 -14607
rect 18854 -14634 18882 -14633
rect 18854 -14767 18882 -14766
rect 18854 -14793 18855 -14767
rect 18855 -14793 18881 -14767
rect 18881 -14793 18882 -14767
rect 18854 -14794 18882 -14793
rect 18854 -14927 18882 -14926
rect 18854 -14953 18855 -14927
rect 18855 -14953 18881 -14927
rect 18881 -14953 18882 -14927
rect 18854 -14954 18882 -14953
rect 18854 -15087 18882 -15086
rect 18854 -15113 18855 -15087
rect 18855 -15113 18881 -15087
rect 18881 -15113 18882 -15087
rect 18854 -15114 18882 -15113
rect 15121 -15247 15149 -15246
rect 15121 -15273 15122 -15247
rect 15122 -15273 15148 -15247
rect 15148 -15273 15149 -15247
rect 15121 -15274 15149 -15273
rect 18854 -15247 18882 -15246
rect 18854 -15273 18855 -15247
rect 18855 -15273 18881 -15247
rect 18881 -15273 18882 -15247
rect 18854 -15274 18882 -15273
rect 15306 -15352 15334 -15351
rect 15306 -15378 15307 -15352
rect 15307 -15378 15333 -15352
rect 15333 -15378 15334 -15352
rect 15306 -15379 15334 -15378
rect 15466 -15352 15494 -15351
rect 15466 -15378 15467 -15352
rect 15467 -15378 15493 -15352
rect 15493 -15378 15494 -15352
rect 15466 -15379 15494 -15378
rect 15626 -15352 15654 -15351
rect 15626 -15378 15627 -15352
rect 15627 -15378 15653 -15352
rect 15653 -15378 15654 -15352
rect 15626 -15379 15654 -15378
rect 15786 -15352 15814 -15351
rect 15786 -15378 15787 -15352
rect 15787 -15378 15813 -15352
rect 15813 -15378 15814 -15352
rect 15786 -15379 15814 -15378
rect 15946 -15352 15974 -15351
rect 15946 -15378 15947 -15352
rect 15947 -15378 15973 -15352
rect 15973 -15378 15974 -15352
rect 15946 -15379 15974 -15378
rect 16106 -15352 16134 -15351
rect 16106 -15378 16107 -15352
rect 16107 -15378 16133 -15352
rect 16133 -15378 16134 -15352
rect 16106 -15379 16134 -15378
rect 16266 -15352 16294 -15351
rect 16266 -15378 16267 -15352
rect 16267 -15378 16293 -15352
rect 16293 -15378 16294 -15352
rect 16266 -15379 16294 -15378
rect 16426 -15352 16454 -15351
rect 16426 -15378 16427 -15352
rect 16427 -15378 16453 -15352
rect 16453 -15378 16454 -15352
rect 16426 -15379 16454 -15378
rect 16586 -15352 16614 -15351
rect 16586 -15378 16587 -15352
rect 16587 -15378 16613 -15352
rect 16613 -15378 16614 -15352
rect 16586 -15379 16614 -15378
rect 16746 -15352 16774 -15351
rect 16746 -15378 16747 -15352
rect 16747 -15378 16773 -15352
rect 16773 -15378 16774 -15352
rect 16746 -15379 16774 -15378
rect 16906 -15352 16934 -15351
rect 16906 -15378 16907 -15352
rect 16907 -15378 16933 -15352
rect 16933 -15378 16934 -15352
rect 16906 -15379 16934 -15378
rect 17066 -15352 17094 -15351
rect 17066 -15378 17067 -15352
rect 17067 -15378 17093 -15352
rect 17093 -15378 17094 -15352
rect 17066 -15379 17094 -15378
rect 17226 -15352 17254 -15351
rect 17226 -15378 17227 -15352
rect 17227 -15378 17253 -15352
rect 17253 -15378 17254 -15352
rect 17226 -15379 17254 -15378
rect 17386 -15352 17414 -15351
rect 17386 -15378 17387 -15352
rect 17387 -15378 17413 -15352
rect 17413 -15378 17414 -15352
rect 17386 -15379 17414 -15378
rect 17546 -15352 17574 -15351
rect 17546 -15378 17547 -15352
rect 17547 -15378 17573 -15352
rect 17573 -15378 17574 -15352
rect 17546 -15379 17574 -15378
rect 17706 -15352 17734 -15351
rect 17706 -15378 17707 -15352
rect 17707 -15378 17733 -15352
rect 17733 -15378 17734 -15352
rect 17706 -15379 17734 -15378
rect 17866 -15352 17894 -15351
rect 17866 -15378 17867 -15352
rect 17867 -15378 17893 -15352
rect 17893 -15378 17894 -15352
rect 17866 -15379 17894 -15378
rect 18026 -15352 18054 -15351
rect 18026 -15378 18027 -15352
rect 18027 -15378 18053 -15352
rect 18053 -15378 18054 -15352
rect 18026 -15379 18054 -15378
rect 18186 -15352 18214 -15351
rect 18186 -15378 18187 -15352
rect 18187 -15378 18213 -15352
rect 18213 -15378 18214 -15352
rect 18186 -15379 18214 -15378
rect 18346 -15352 18374 -15351
rect 18346 -15378 18347 -15352
rect 18347 -15378 18373 -15352
rect 18373 -15378 18374 -15352
rect 18346 -15379 18374 -15378
rect 18506 -15352 18534 -15351
rect 18506 -15378 18507 -15352
rect 18507 -15378 18533 -15352
rect 18533 -15378 18534 -15352
rect 18506 -15379 18534 -15378
rect 18666 -15352 18694 -15351
rect 18666 -15378 18667 -15352
rect 18667 -15378 18693 -15352
rect 18693 -15378 18694 -15352
rect 18666 -15379 18694 -15378
rect 21306 -11624 21334 -11623
rect 21306 -11650 21307 -11624
rect 21307 -11650 21333 -11624
rect 21333 -11650 21334 -11624
rect 21306 -11651 21334 -11650
rect 21466 -11624 21494 -11623
rect 21466 -11650 21467 -11624
rect 21467 -11650 21493 -11624
rect 21493 -11650 21494 -11624
rect 21466 -11651 21494 -11650
rect 21626 -11624 21654 -11623
rect 21626 -11650 21627 -11624
rect 21627 -11650 21653 -11624
rect 21653 -11650 21654 -11624
rect 21626 -11651 21654 -11650
rect 21786 -11624 21814 -11623
rect 21786 -11650 21787 -11624
rect 21787 -11650 21813 -11624
rect 21813 -11650 21814 -11624
rect 21786 -11651 21814 -11650
rect 21946 -11624 21974 -11623
rect 21946 -11650 21947 -11624
rect 21947 -11650 21973 -11624
rect 21973 -11650 21974 -11624
rect 21946 -11651 21974 -11650
rect 22106 -11624 22134 -11623
rect 22106 -11650 22107 -11624
rect 22107 -11650 22133 -11624
rect 22133 -11650 22134 -11624
rect 22106 -11651 22134 -11650
rect 22266 -11624 22294 -11623
rect 22266 -11650 22267 -11624
rect 22267 -11650 22293 -11624
rect 22293 -11650 22294 -11624
rect 22266 -11651 22294 -11650
rect 22426 -11624 22454 -11623
rect 22426 -11650 22427 -11624
rect 22427 -11650 22453 -11624
rect 22453 -11650 22454 -11624
rect 22426 -11651 22454 -11650
rect 22586 -11624 22614 -11623
rect 22586 -11650 22587 -11624
rect 22587 -11650 22613 -11624
rect 22613 -11650 22614 -11624
rect 22586 -11651 22614 -11650
rect 22746 -11624 22774 -11623
rect 22746 -11650 22747 -11624
rect 22747 -11650 22773 -11624
rect 22773 -11650 22774 -11624
rect 22746 -11651 22774 -11650
rect 22906 -11624 22934 -11623
rect 22906 -11650 22907 -11624
rect 22907 -11650 22933 -11624
rect 22933 -11650 22934 -11624
rect 22906 -11651 22934 -11650
rect 23066 -11624 23094 -11623
rect 23066 -11650 23067 -11624
rect 23067 -11650 23093 -11624
rect 23093 -11650 23094 -11624
rect 23066 -11651 23094 -11650
rect 23226 -11624 23254 -11623
rect 23226 -11650 23227 -11624
rect 23227 -11650 23253 -11624
rect 23253 -11650 23254 -11624
rect 23226 -11651 23254 -11650
rect 23386 -11624 23414 -11623
rect 23386 -11650 23387 -11624
rect 23387 -11650 23413 -11624
rect 23413 -11650 23414 -11624
rect 23386 -11651 23414 -11650
rect 23546 -11624 23574 -11623
rect 23546 -11650 23547 -11624
rect 23547 -11650 23573 -11624
rect 23573 -11650 23574 -11624
rect 23546 -11651 23574 -11650
rect 23706 -11624 23734 -11623
rect 23706 -11650 23707 -11624
rect 23707 -11650 23733 -11624
rect 23733 -11650 23734 -11624
rect 23706 -11651 23734 -11650
rect 23866 -11624 23894 -11623
rect 23866 -11650 23867 -11624
rect 23867 -11650 23893 -11624
rect 23893 -11650 23894 -11624
rect 23866 -11651 23894 -11650
rect 24026 -11624 24054 -11623
rect 24026 -11650 24027 -11624
rect 24027 -11650 24053 -11624
rect 24053 -11650 24054 -11624
rect 24026 -11651 24054 -11650
rect 24186 -11624 24214 -11623
rect 24186 -11650 24187 -11624
rect 24187 -11650 24213 -11624
rect 24213 -11650 24214 -11624
rect 24186 -11651 24214 -11650
rect 24346 -11624 24374 -11623
rect 24346 -11650 24347 -11624
rect 24347 -11650 24373 -11624
rect 24373 -11650 24374 -11624
rect 24346 -11651 24374 -11650
rect 24506 -11624 24534 -11623
rect 24506 -11650 24507 -11624
rect 24507 -11650 24533 -11624
rect 24533 -11650 24534 -11624
rect 24506 -11651 24534 -11650
rect 24666 -11624 24694 -11623
rect 24666 -11650 24667 -11624
rect 24667 -11650 24693 -11624
rect 24693 -11650 24694 -11624
rect 24666 -11651 24694 -11650
rect 21121 -11727 21149 -11726
rect 21121 -11753 21122 -11727
rect 21122 -11753 21148 -11727
rect 21148 -11753 21149 -11727
rect 21121 -11754 21149 -11753
rect 24854 -11727 24882 -11726
rect 24854 -11753 24855 -11727
rect 24855 -11753 24881 -11727
rect 24881 -11753 24882 -11727
rect 24854 -11754 24882 -11753
rect 21121 -11887 21149 -11886
rect 21121 -11913 21122 -11887
rect 21122 -11913 21148 -11887
rect 21148 -11913 21149 -11887
rect 21121 -11914 21149 -11913
rect 21121 -12047 21149 -12046
rect 21121 -12073 21122 -12047
rect 21122 -12073 21148 -12047
rect 21148 -12073 21149 -12047
rect 21121 -12074 21149 -12073
rect 21121 -12207 21149 -12206
rect 21121 -12233 21122 -12207
rect 21122 -12233 21148 -12207
rect 21148 -12233 21149 -12207
rect 21121 -12234 21149 -12233
rect 21121 -12367 21149 -12366
rect 21121 -12393 21122 -12367
rect 21122 -12393 21148 -12367
rect 21148 -12393 21149 -12367
rect 21121 -12394 21149 -12393
rect 21121 -12527 21149 -12526
rect 21121 -12553 21122 -12527
rect 21122 -12553 21148 -12527
rect 21148 -12553 21149 -12527
rect 21121 -12554 21149 -12553
rect 21121 -12687 21149 -12686
rect 21121 -12713 21122 -12687
rect 21122 -12713 21148 -12687
rect 21148 -12713 21149 -12687
rect 21121 -12714 21149 -12713
rect 21121 -12847 21149 -12846
rect 21121 -12873 21122 -12847
rect 21122 -12873 21148 -12847
rect 21148 -12873 21149 -12847
rect 21121 -12874 21149 -12873
rect 21121 -13007 21149 -13006
rect 21121 -13033 21122 -13007
rect 21122 -13033 21148 -13007
rect 21148 -13033 21149 -13007
rect 21121 -13034 21149 -13033
rect 21121 -13167 21149 -13166
rect 21121 -13193 21122 -13167
rect 21122 -13193 21148 -13167
rect 21148 -13193 21149 -13167
rect 21121 -13194 21149 -13193
rect 21121 -13327 21149 -13326
rect 21121 -13353 21122 -13327
rect 21122 -13353 21148 -13327
rect 21148 -13353 21149 -13327
rect 21121 -13354 21149 -13353
rect 21121 -13487 21149 -13486
rect 21121 -13513 21122 -13487
rect 21122 -13513 21148 -13487
rect 21148 -13513 21149 -13487
rect 21121 -13514 21149 -13513
rect 21121 -13647 21149 -13646
rect 21121 -13673 21122 -13647
rect 21122 -13673 21148 -13647
rect 21148 -13673 21149 -13647
rect 21121 -13674 21149 -13673
rect 21121 -13807 21149 -13806
rect 21121 -13833 21122 -13807
rect 21122 -13833 21148 -13807
rect 21148 -13833 21149 -13807
rect 21121 -13834 21149 -13833
rect 21121 -13967 21149 -13966
rect 21121 -13993 21122 -13967
rect 21122 -13993 21148 -13967
rect 21148 -13993 21149 -13967
rect 21121 -13994 21149 -13993
rect 21121 -14127 21149 -14126
rect 21121 -14153 21122 -14127
rect 21122 -14153 21148 -14127
rect 21148 -14153 21149 -14127
rect 21121 -14154 21149 -14153
rect 21121 -14287 21149 -14286
rect 21121 -14313 21122 -14287
rect 21122 -14313 21148 -14287
rect 21148 -14313 21149 -14287
rect 21121 -14314 21149 -14313
rect 21121 -14447 21149 -14446
rect 21121 -14473 21122 -14447
rect 21122 -14473 21148 -14447
rect 21148 -14473 21149 -14447
rect 21121 -14474 21149 -14473
rect 21121 -14607 21149 -14606
rect 21121 -14633 21122 -14607
rect 21122 -14633 21148 -14607
rect 21148 -14633 21149 -14607
rect 21121 -14634 21149 -14633
rect 21121 -14767 21149 -14766
rect 21121 -14793 21122 -14767
rect 21122 -14793 21148 -14767
rect 21148 -14793 21149 -14767
rect 21121 -14794 21149 -14793
rect 21121 -14927 21149 -14926
rect 21121 -14953 21122 -14927
rect 21122 -14953 21148 -14927
rect 21148 -14953 21149 -14927
rect 21121 -14954 21149 -14953
rect 21121 -15087 21149 -15086
rect 21121 -15113 21122 -15087
rect 21122 -15113 21148 -15087
rect 21148 -15113 21149 -15087
rect 21121 -15114 21149 -15113
rect 24854 -11887 24882 -11886
rect 24854 -11913 24855 -11887
rect 24855 -11913 24881 -11887
rect 24881 -11913 24882 -11887
rect 24854 -11914 24882 -11913
rect 24854 -12047 24882 -12046
rect 24854 -12073 24855 -12047
rect 24855 -12073 24881 -12047
rect 24881 -12073 24882 -12047
rect 24854 -12074 24882 -12073
rect 24854 -12207 24882 -12206
rect 24854 -12233 24855 -12207
rect 24855 -12233 24881 -12207
rect 24881 -12233 24882 -12207
rect 24854 -12234 24882 -12233
rect 24854 -12367 24882 -12366
rect 24854 -12393 24855 -12367
rect 24855 -12393 24881 -12367
rect 24881 -12393 24882 -12367
rect 24854 -12394 24882 -12393
rect 24854 -12527 24882 -12526
rect 24854 -12553 24855 -12527
rect 24855 -12553 24881 -12527
rect 24881 -12553 24882 -12527
rect 24854 -12554 24882 -12553
rect 24854 -12687 24882 -12686
rect 24854 -12713 24855 -12687
rect 24855 -12713 24881 -12687
rect 24881 -12713 24882 -12687
rect 24854 -12714 24882 -12713
rect 24854 -12847 24882 -12846
rect 24854 -12873 24855 -12847
rect 24855 -12873 24881 -12847
rect 24881 -12873 24882 -12847
rect 24854 -12874 24882 -12873
rect 24854 -13007 24882 -13006
rect 24854 -13033 24855 -13007
rect 24855 -13033 24881 -13007
rect 24881 -13033 24882 -13007
rect 24854 -13034 24882 -13033
rect 24854 -13167 24882 -13166
rect 24854 -13193 24855 -13167
rect 24855 -13193 24881 -13167
rect 24881 -13193 24882 -13167
rect 24854 -13194 24882 -13193
rect 24854 -13327 24882 -13326
rect 24854 -13353 24855 -13327
rect 24855 -13353 24881 -13327
rect 24881 -13353 24882 -13327
rect 24854 -13354 24882 -13353
rect 24854 -13487 24882 -13486
rect 24854 -13513 24855 -13487
rect 24855 -13513 24881 -13487
rect 24881 -13513 24882 -13487
rect 24854 -13514 24882 -13513
rect 24854 -13647 24882 -13646
rect 24854 -13673 24855 -13647
rect 24855 -13673 24881 -13647
rect 24881 -13673 24882 -13647
rect 24854 -13674 24882 -13673
rect 24854 -13807 24882 -13806
rect 24854 -13833 24855 -13807
rect 24855 -13833 24881 -13807
rect 24881 -13833 24882 -13807
rect 24854 -13834 24882 -13833
rect 24854 -13967 24882 -13966
rect 24854 -13993 24855 -13967
rect 24855 -13993 24881 -13967
rect 24881 -13993 24882 -13967
rect 24854 -13994 24882 -13993
rect 24854 -14127 24882 -14126
rect 24854 -14153 24855 -14127
rect 24855 -14153 24881 -14127
rect 24881 -14153 24882 -14127
rect 24854 -14154 24882 -14153
rect 24854 -14287 24882 -14286
rect 24854 -14313 24855 -14287
rect 24855 -14313 24881 -14287
rect 24881 -14313 24882 -14287
rect 24854 -14314 24882 -14313
rect 24854 -14447 24882 -14446
rect 24854 -14473 24855 -14447
rect 24855 -14473 24881 -14447
rect 24881 -14473 24882 -14447
rect 24854 -14474 24882 -14473
rect 24854 -14607 24882 -14606
rect 24854 -14633 24855 -14607
rect 24855 -14633 24881 -14607
rect 24881 -14633 24882 -14607
rect 24854 -14634 24882 -14633
rect 24854 -14767 24882 -14766
rect 24854 -14793 24855 -14767
rect 24855 -14793 24881 -14767
rect 24881 -14793 24882 -14767
rect 24854 -14794 24882 -14793
rect 24854 -14927 24882 -14926
rect 24854 -14953 24855 -14927
rect 24855 -14953 24881 -14927
rect 24881 -14953 24882 -14927
rect 24854 -14954 24882 -14953
rect 24854 -15087 24882 -15086
rect 24854 -15113 24855 -15087
rect 24855 -15113 24881 -15087
rect 24881 -15113 24882 -15087
rect 24854 -15114 24882 -15113
rect 21121 -15247 21149 -15246
rect 21121 -15273 21122 -15247
rect 21122 -15273 21148 -15247
rect 21148 -15273 21149 -15247
rect 21121 -15274 21149 -15273
rect 24854 -15247 24882 -15246
rect 24854 -15273 24855 -15247
rect 24855 -15273 24881 -15247
rect 24881 -15273 24882 -15247
rect 24854 -15274 24882 -15273
rect 21306 -15352 21334 -15351
rect 21306 -15378 21307 -15352
rect 21307 -15378 21333 -15352
rect 21333 -15378 21334 -15352
rect 21306 -15379 21334 -15378
rect 21466 -15352 21494 -15351
rect 21466 -15378 21467 -15352
rect 21467 -15378 21493 -15352
rect 21493 -15378 21494 -15352
rect 21466 -15379 21494 -15378
rect 21626 -15352 21654 -15351
rect 21626 -15378 21627 -15352
rect 21627 -15378 21653 -15352
rect 21653 -15378 21654 -15352
rect 21626 -15379 21654 -15378
rect 21786 -15352 21814 -15351
rect 21786 -15378 21787 -15352
rect 21787 -15378 21813 -15352
rect 21813 -15378 21814 -15352
rect 21786 -15379 21814 -15378
rect 21946 -15352 21974 -15351
rect 21946 -15378 21947 -15352
rect 21947 -15378 21973 -15352
rect 21973 -15378 21974 -15352
rect 21946 -15379 21974 -15378
rect 22106 -15352 22134 -15351
rect 22106 -15378 22107 -15352
rect 22107 -15378 22133 -15352
rect 22133 -15378 22134 -15352
rect 22106 -15379 22134 -15378
rect 22266 -15352 22294 -15351
rect 22266 -15378 22267 -15352
rect 22267 -15378 22293 -15352
rect 22293 -15378 22294 -15352
rect 22266 -15379 22294 -15378
rect 22426 -15352 22454 -15351
rect 22426 -15378 22427 -15352
rect 22427 -15378 22453 -15352
rect 22453 -15378 22454 -15352
rect 22426 -15379 22454 -15378
rect 22586 -15352 22614 -15351
rect 22586 -15378 22587 -15352
rect 22587 -15378 22613 -15352
rect 22613 -15378 22614 -15352
rect 22586 -15379 22614 -15378
rect 22746 -15352 22774 -15351
rect 22746 -15378 22747 -15352
rect 22747 -15378 22773 -15352
rect 22773 -15378 22774 -15352
rect 22746 -15379 22774 -15378
rect 22906 -15352 22934 -15351
rect 22906 -15378 22907 -15352
rect 22907 -15378 22933 -15352
rect 22933 -15378 22934 -15352
rect 22906 -15379 22934 -15378
rect 23066 -15352 23094 -15351
rect 23066 -15378 23067 -15352
rect 23067 -15378 23093 -15352
rect 23093 -15378 23094 -15352
rect 23066 -15379 23094 -15378
rect 23226 -15352 23254 -15351
rect 23226 -15378 23227 -15352
rect 23227 -15378 23253 -15352
rect 23253 -15378 23254 -15352
rect 23226 -15379 23254 -15378
rect 23386 -15352 23414 -15351
rect 23386 -15378 23387 -15352
rect 23387 -15378 23413 -15352
rect 23413 -15378 23414 -15352
rect 23386 -15379 23414 -15378
rect 23546 -15352 23574 -15351
rect 23546 -15378 23547 -15352
rect 23547 -15378 23573 -15352
rect 23573 -15378 23574 -15352
rect 23546 -15379 23574 -15378
rect 23706 -15352 23734 -15351
rect 23706 -15378 23707 -15352
rect 23707 -15378 23733 -15352
rect 23733 -15378 23734 -15352
rect 23706 -15379 23734 -15378
rect 23866 -15352 23894 -15351
rect 23866 -15378 23867 -15352
rect 23867 -15378 23893 -15352
rect 23893 -15378 23894 -15352
rect 23866 -15379 23894 -15378
rect 24026 -15352 24054 -15351
rect 24026 -15378 24027 -15352
rect 24027 -15378 24053 -15352
rect 24053 -15378 24054 -15352
rect 24026 -15379 24054 -15378
rect 24186 -15352 24214 -15351
rect 24186 -15378 24187 -15352
rect 24187 -15378 24213 -15352
rect 24213 -15378 24214 -15352
rect 24186 -15379 24214 -15378
rect 24346 -15352 24374 -15351
rect 24346 -15378 24347 -15352
rect 24347 -15378 24373 -15352
rect 24373 -15378 24374 -15352
rect 24346 -15379 24374 -15378
rect 24506 -15352 24534 -15351
rect 24506 -15378 24507 -15352
rect 24507 -15378 24533 -15352
rect 24533 -15378 24534 -15352
rect 24506 -15379 24534 -15378
rect 24666 -15352 24694 -15351
rect 24666 -15378 24667 -15352
rect 24667 -15378 24693 -15352
rect 24693 -15378 24694 -15352
rect 24666 -15379 24694 -15378
<< metal3 >>
rect 9930 -3465 9970 -3325
rect 10030 -3390 10070 -3325
rect 10030 -3430 10600 -3390
rect 9930 -3505 10520 -3465
rect 10480 -4130 10520 -3505
rect 10560 -4050 10600 -3430
rect 11540 -3740 12205 -3735
rect 11540 -3770 11635 -3740
rect 11705 -3770 12205 -3740
rect 11540 -3775 12205 -3770
rect 11540 -4050 11580 -3775
rect 10560 -4090 11580 -4050
rect 11645 -3900 12100 -3895
rect 11645 -3930 11775 -3900
rect 11845 -3930 12100 -3900
rect 11645 -3935 12100 -3930
rect 11645 -4130 11685 -3935
rect 10480 -4170 11685 -4130
rect 8300 -4755 8340 -4750
rect 8165 -4760 8235 -4755
rect 8165 -4790 8200 -4760
rect 8230 -4790 8235 -4760
rect 8165 -4795 8235 -4790
rect 8300 -4785 8305 -4755
rect 8335 -4785 8340 -4755
rect 8300 -4790 8340 -4785
rect 3000 -5621 7000 -5500
rect 3000 -5653 3304 -5621
rect 3336 -5653 3464 -5621
rect 3496 -5653 3624 -5621
rect 3656 -5653 3784 -5621
rect 3816 -5653 3944 -5621
rect 3976 -5653 4104 -5621
rect 4136 -5653 4264 -5621
rect 4296 -5653 4424 -5621
rect 4456 -5653 4584 -5621
rect 4616 -5653 4744 -5621
rect 4776 -5653 4904 -5621
rect 4936 -5653 5064 -5621
rect 5096 -5653 5224 -5621
rect 5256 -5653 5384 -5621
rect 5416 -5653 5544 -5621
rect 5576 -5653 5704 -5621
rect 5736 -5653 5864 -5621
rect 5896 -5653 6024 -5621
rect 6056 -5653 6184 -5621
rect 6216 -5653 6344 -5621
rect 6376 -5653 6504 -5621
rect 6536 -5653 6664 -5621
rect 6696 -5653 7000 -5621
rect 3000 -5724 7000 -5653
rect 3000 -5756 3119 -5724
rect 3151 -5756 6852 -5724
rect 6884 -5756 7000 -5724
rect 3000 -5770 7000 -5756
rect 3000 -5884 3270 -5770
rect 3000 -5916 3119 -5884
rect 3151 -5916 3270 -5884
rect 3000 -6044 3270 -5916
rect 3000 -6076 3119 -6044
rect 3151 -6076 3270 -6044
rect 3000 -6204 3270 -6076
rect 3000 -6236 3119 -6204
rect 3151 -6236 3270 -6204
rect 3000 -6364 3270 -6236
rect 3000 -6396 3119 -6364
rect 3151 -6396 3270 -6364
rect 3000 -6524 3270 -6396
rect 3000 -6556 3119 -6524
rect 3151 -6556 3270 -6524
rect 3000 -6684 3270 -6556
rect 3000 -6716 3119 -6684
rect 3151 -6716 3270 -6684
rect 3000 -6844 3270 -6716
rect 3000 -6876 3119 -6844
rect 3151 -6876 3270 -6844
rect 3000 -7004 3270 -6876
rect 3000 -7036 3119 -7004
rect 3151 -7036 3270 -7004
rect 3000 -7164 3270 -7036
rect 3000 -7196 3119 -7164
rect 3151 -7196 3270 -7164
rect 3000 -7324 3270 -7196
rect 3000 -7356 3119 -7324
rect 3151 -7356 3270 -7324
rect 3000 -7484 3270 -7356
rect 3000 -7516 3119 -7484
rect 3151 -7516 3270 -7484
rect 3000 -7644 3270 -7516
rect 3000 -7676 3119 -7644
rect 3151 -7676 3270 -7644
rect 3000 -7804 3270 -7676
rect 3000 -7836 3119 -7804
rect 3151 -7836 3270 -7804
rect 3000 -7964 3270 -7836
rect 3000 -7996 3119 -7964
rect 3151 -7996 3270 -7964
rect 3000 -8124 3270 -7996
rect 3000 -8156 3119 -8124
rect 3151 -8156 3270 -8124
rect 3000 -8284 3270 -8156
rect 3000 -8316 3119 -8284
rect 3151 -8316 3270 -8284
rect 3000 -8444 3270 -8316
rect 3000 -8476 3119 -8444
rect 3151 -8476 3270 -8444
rect 3000 -8604 3270 -8476
rect 3000 -8636 3119 -8604
rect 3151 -8636 3270 -8604
rect 3000 -8764 3270 -8636
rect 3000 -8796 3119 -8764
rect 3151 -8796 3270 -8764
rect 3000 -8924 3270 -8796
rect 3000 -8956 3119 -8924
rect 3151 -8956 3270 -8924
rect 3000 -9084 3270 -8956
rect 3000 -9116 3119 -9084
rect 3151 -9116 3270 -9084
rect 3000 -9230 3270 -9116
rect 6730 -5884 7000 -5770
rect 6730 -5916 6852 -5884
rect 6884 -5916 7000 -5884
rect 6730 -6044 7000 -5916
rect 6730 -6076 6852 -6044
rect 6884 -6076 7000 -6044
rect 6730 -6204 7000 -6076
rect 6730 -6236 6852 -6204
rect 6884 -6236 7000 -6204
rect 6730 -6364 7000 -6236
rect 6730 -6396 6852 -6364
rect 6884 -6396 7000 -6364
rect 6730 -6524 7000 -6396
rect 6730 -6556 6852 -6524
rect 6884 -6556 7000 -6524
rect 6730 -6684 7000 -6556
rect 6730 -6716 6852 -6684
rect 6884 -6716 7000 -6684
rect 6730 -6844 7000 -6716
rect 6730 -6876 6852 -6844
rect 6884 -6876 7000 -6844
rect 6730 -7004 7000 -6876
rect 6730 -7036 6852 -7004
rect 6884 -7036 7000 -7004
rect 6730 -7164 7000 -7036
rect 6730 -7196 6852 -7164
rect 6884 -7196 7000 -7164
rect 6730 -7324 7000 -7196
rect 6730 -7356 6852 -7324
rect 6884 -7356 7000 -7324
rect 6730 -7484 7000 -7356
rect 6730 -7516 6852 -7484
rect 6884 -7516 7000 -7484
rect 6730 -7644 7000 -7516
rect 6730 -7676 6852 -7644
rect 6884 -7676 7000 -7644
rect 6730 -7804 7000 -7676
rect 6730 -7836 6852 -7804
rect 6884 -7836 7000 -7804
rect 6730 -7964 7000 -7836
rect 6730 -7996 6852 -7964
rect 6884 -7996 7000 -7964
rect 6730 -8124 7000 -7996
rect 6730 -8156 6852 -8124
rect 6884 -8156 7000 -8124
rect 6730 -8284 7000 -8156
rect 6730 -8316 6852 -8284
rect 6884 -8316 7000 -8284
rect 6730 -8444 7000 -8316
rect 6730 -8476 6852 -8444
rect 6884 -8476 7000 -8444
rect 6730 -8604 7000 -8476
rect 6730 -8636 6852 -8604
rect 6884 -8636 7000 -8604
rect 6730 -8764 7000 -8636
rect 6730 -8796 6852 -8764
rect 6884 -8796 7000 -8764
rect 6730 -8924 7000 -8796
rect 6730 -8956 6852 -8924
rect 6884 -8956 7000 -8924
rect 6730 -9084 7000 -8956
rect 6730 -9116 6852 -9084
rect 6884 -9116 7000 -9084
rect 6730 -9230 7000 -9116
rect 3000 -9244 7000 -9230
rect 3000 -9276 3119 -9244
rect 3151 -9276 6852 -9244
rect 6884 -9276 7000 -9244
rect 3000 -9349 7000 -9276
rect 3000 -9381 3304 -9349
rect 3336 -9381 3464 -9349
rect 3496 -9381 3624 -9349
rect 3656 -9381 3784 -9349
rect 3816 -9381 3944 -9349
rect 3976 -9381 4104 -9349
rect 4136 -9381 4264 -9349
rect 4296 -9381 4424 -9349
rect 4456 -9381 4584 -9349
rect 4616 -9381 4744 -9349
rect 4776 -9381 4904 -9349
rect 4936 -9381 5064 -9349
rect 5096 -9381 5224 -9349
rect 5256 -9381 5384 -9349
rect 5416 -9381 5544 -9349
rect 5576 -9381 5704 -9349
rect 5736 -9381 5864 -9349
rect 5896 -9381 6024 -9349
rect 6056 -9381 6184 -9349
rect 6216 -9381 6344 -9349
rect 6376 -9381 6504 -9349
rect 6536 -9381 6664 -9349
rect 6696 -9381 7000 -9349
rect 3000 -9500 7000 -9381
rect 3000 -11621 7000 -11500
rect 3000 -11653 3304 -11621
rect 3336 -11653 3464 -11621
rect 3496 -11653 3624 -11621
rect 3656 -11653 3784 -11621
rect 3816 -11653 3944 -11621
rect 3976 -11653 4104 -11621
rect 4136 -11653 4264 -11621
rect 4296 -11653 4424 -11621
rect 4456 -11653 4584 -11621
rect 4616 -11653 4744 -11621
rect 4776 -11653 4904 -11621
rect 4936 -11653 5064 -11621
rect 5096 -11653 5224 -11621
rect 5256 -11653 5384 -11621
rect 5416 -11653 5544 -11621
rect 5576 -11653 5704 -11621
rect 5736 -11653 5864 -11621
rect 5896 -11653 6024 -11621
rect 6056 -11653 6184 -11621
rect 6216 -11653 6344 -11621
rect 6376 -11653 6504 -11621
rect 6536 -11653 6664 -11621
rect 6696 -11653 7000 -11621
rect 3000 -11724 7000 -11653
rect 3000 -11756 3119 -11724
rect 3151 -11756 6852 -11724
rect 6884 -11756 7000 -11724
rect 3000 -11770 7000 -11756
rect 3000 -11884 3270 -11770
rect 3000 -11916 3119 -11884
rect 3151 -11916 3270 -11884
rect 3000 -12044 3270 -11916
rect 3000 -12076 3119 -12044
rect 3151 -12076 3270 -12044
rect 3000 -12204 3270 -12076
rect 3000 -12236 3119 -12204
rect 3151 -12236 3270 -12204
rect 3000 -12364 3270 -12236
rect 3000 -12396 3119 -12364
rect 3151 -12396 3270 -12364
rect 3000 -12524 3270 -12396
rect 3000 -12556 3119 -12524
rect 3151 -12556 3270 -12524
rect 3000 -12684 3270 -12556
rect 3000 -12716 3119 -12684
rect 3151 -12716 3270 -12684
rect 3000 -12844 3270 -12716
rect 3000 -12876 3119 -12844
rect 3151 -12876 3270 -12844
rect 3000 -13004 3270 -12876
rect 3000 -13036 3119 -13004
rect 3151 -13036 3270 -13004
rect 3000 -13164 3270 -13036
rect 3000 -13196 3119 -13164
rect 3151 -13196 3270 -13164
rect 3000 -13324 3270 -13196
rect 3000 -13356 3119 -13324
rect 3151 -13356 3270 -13324
rect 3000 -13484 3270 -13356
rect 3000 -13516 3119 -13484
rect 3151 -13516 3270 -13484
rect 3000 -13644 3270 -13516
rect 3000 -13676 3119 -13644
rect 3151 -13676 3270 -13644
rect 3000 -13804 3270 -13676
rect 3000 -13836 3119 -13804
rect 3151 -13836 3270 -13804
rect 3000 -13964 3270 -13836
rect 3000 -13996 3119 -13964
rect 3151 -13996 3270 -13964
rect 3000 -14124 3270 -13996
rect 3000 -14156 3119 -14124
rect 3151 -14156 3270 -14124
rect 3000 -14284 3270 -14156
rect 3000 -14316 3119 -14284
rect 3151 -14316 3270 -14284
rect 3000 -14444 3270 -14316
rect 3000 -14476 3119 -14444
rect 3151 -14476 3270 -14444
rect 3000 -14604 3270 -14476
rect 3000 -14636 3119 -14604
rect 3151 -14636 3270 -14604
rect 3000 -14764 3270 -14636
rect 3000 -14796 3119 -14764
rect 3151 -14796 3270 -14764
rect 3000 -14924 3270 -14796
rect 3000 -14956 3119 -14924
rect 3151 -14956 3270 -14924
rect 3000 -15084 3270 -14956
rect 3000 -15116 3119 -15084
rect 3151 -15116 3270 -15084
rect 3000 -15230 3270 -15116
rect 6730 -11884 7000 -11770
rect 6730 -11916 6852 -11884
rect 6884 -11916 7000 -11884
rect 6730 -12044 7000 -11916
rect 6730 -12076 6852 -12044
rect 6884 -12076 7000 -12044
rect 6730 -12204 7000 -12076
rect 6730 -12236 6852 -12204
rect 6884 -12236 7000 -12204
rect 6730 -12364 7000 -12236
rect 6730 -12396 6852 -12364
rect 6884 -12396 7000 -12364
rect 6730 -12524 7000 -12396
rect 6730 -12556 6852 -12524
rect 6884 -12556 7000 -12524
rect 6730 -12684 7000 -12556
rect 6730 -12716 6852 -12684
rect 6884 -12716 7000 -12684
rect 6730 -12844 7000 -12716
rect 6730 -12876 6852 -12844
rect 6884 -12870 7000 -12844
rect 8165 -12870 8195 -4795
rect 6884 -12876 8195 -12870
rect 6730 -12900 8195 -12876
rect 8230 -4830 8270 -4825
rect 8230 -4860 8235 -4830
rect 8265 -4860 8270 -4830
rect 8230 -4865 8270 -4860
rect 8230 -12875 8260 -4865
rect 8300 -5305 8330 -4790
rect 8300 -5310 8570 -5305
rect 8300 -5370 8520 -5310
rect 8560 -5370 8570 -5310
rect 8300 -5375 8570 -5370
rect 8300 -11330 8330 -5375
rect 12060 -5400 12100 -3935
rect 12165 -5300 12205 -3775
rect 12165 -5340 13340 -5300
rect 12060 -5440 13240 -5400
rect 9000 -5621 13000 -5500
rect 9000 -5653 9304 -5621
rect 9336 -5653 9464 -5621
rect 9496 -5653 9624 -5621
rect 9656 -5653 9784 -5621
rect 9816 -5653 9944 -5621
rect 9976 -5653 10104 -5621
rect 10136 -5653 10264 -5621
rect 10296 -5653 10424 -5621
rect 10456 -5653 10584 -5621
rect 10616 -5653 10744 -5621
rect 10776 -5653 10904 -5621
rect 10936 -5653 11064 -5621
rect 11096 -5653 11224 -5621
rect 11256 -5653 11384 -5621
rect 11416 -5653 11544 -5621
rect 11576 -5653 11704 -5621
rect 11736 -5653 11864 -5621
rect 11896 -5653 12024 -5621
rect 12056 -5653 12184 -5621
rect 12216 -5653 12344 -5621
rect 12376 -5653 12504 -5621
rect 12536 -5653 12664 -5621
rect 12696 -5653 13000 -5621
rect 9000 -5724 13000 -5653
rect 9000 -5756 9119 -5724
rect 9151 -5756 12852 -5724
rect 12884 -5756 13000 -5724
rect 9000 -5770 13000 -5756
rect 9000 -5884 9270 -5770
rect 9000 -5916 9119 -5884
rect 9151 -5916 9270 -5884
rect 9000 -6044 9270 -5916
rect 9000 -6076 9119 -6044
rect 9151 -6076 9270 -6044
rect 9000 -6204 9270 -6076
rect 9000 -6236 9119 -6204
rect 9151 -6236 9270 -6204
rect 9000 -6364 9270 -6236
rect 9000 -6396 9119 -6364
rect 9151 -6396 9270 -6364
rect 9000 -6524 9270 -6396
rect 9000 -6556 9119 -6524
rect 9151 -6556 9270 -6524
rect 9000 -6684 9270 -6556
rect 9000 -6716 9119 -6684
rect 9151 -6716 9270 -6684
rect 9000 -6844 9270 -6716
rect 9000 -6876 9119 -6844
rect 9151 -6876 9270 -6844
rect 9000 -7004 9270 -6876
rect 9000 -7036 9119 -7004
rect 9151 -7036 9270 -7004
rect 9000 -7164 9270 -7036
rect 9000 -7196 9119 -7164
rect 9151 -7196 9270 -7164
rect 9000 -7324 9270 -7196
rect 9000 -7356 9119 -7324
rect 9151 -7356 9270 -7324
rect 9000 -7484 9270 -7356
rect 9000 -7516 9119 -7484
rect 9151 -7516 9270 -7484
rect 9000 -7644 9270 -7516
rect 9000 -7676 9119 -7644
rect 9151 -7676 9270 -7644
rect 9000 -7804 9270 -7676
rect 9000 -7836 9119 -7804
rect 9151 -7836 9270 -7804
rect 9000 -7964 9270 -7836
rect 9000 -7996 9119 -7964
rect 9151 -7996 9270 -7964
rect 9000 -8124 9270 -7996
rect 9000 -8156 9119 -8124
rect 9151 -8156 9270 -8124
rect 9000 -8284 9270 -8156
rect 9000 -8316 9119 -8284
rect 9151 -8316 9270 -8284
rect 9000 -8444 9270 -8316
rect 9000 -8476 9119 -8444
rect 9151 -8476 9270 -8444
rect 9000 -8604 9270 -8476
rect 9000 -8636 9119 -8604
rect 9151 -8636 9270 -8604
rect 9000 -8764 9270 -8636
rect 9000 -8796 9119 -8764
rect 9151 -8796 9270 -8764
rect 9000 -8924 9270 -8796
rect 9000 -8956 9119 -8924
rect 9151 -8956 9270 -8924
rect 9000 -9084 9270 -8956
rect 9000 -9116 9119 -9084
rect 9151 -9116 9270 -9084
rect 9000 -9230 9270 -9116
rect 12730 -5884 13000 -5770
rect 12730 -5916 12852 -5884
rect 12884 -5916 13000 -5884
rect 12730 -6044 13000 -5916
rect 12730 -6076 12852 -6044
rect 12884 -6076 13000 -6044
rect 12730 -6204 13000 -6076
rect 12730 -6236 12852 -6204
rect 12884 -6236 13000 -6204
rect 12730 -6364 13000 -6236
rect 12730 -6396 12852 -6364
rect 12884 -6396 13000 -6364
rect 12730 -6524 13000 -6396
rect 12730 -6556 12852 -6524
rect 12884 -6556 13000 -6524
rect 12730 -6684 13000 -6556
rect 12730 -6716 12852 -6684
rect 12884 -6716 13000 -6684
rect 12730 -6844 13000 -6716
rect 12730 -6876 12852 -6844
rect 12884 -6876 13000 -6844
rect 12730 -7004 13000 -6876
rect 12730 -7036 12852 -7004
rect 12884 -7036 13000 -7004
rect 12730 -7164 13000 -7036
rect 12730 -7196 12852 -7164
rect 12884 -7196 13000 -7164
rect 12730 -7324 13000 -7196
rect 12730 -7356 12852 -7324
rect 12884 -7356 13000 -7324
rect 12730 -7484 13000 -7356
rect 12730 -7516 12852 -7484
rect 12884 -7516 13000 -7484
rect 12730 -7644 13000 -7516
rect 12730 -7676 12852 -7644
rect 12884 -7676 13000 -7644
rect 12730 -7804 13000 -7676
rect 12730 -7836 12852 -7804
rect 12884 -7836 13000 -7804
rect 13200 -7795 13240 -5440
rect 13300 -7675 13340 -5340
rect 15000 -5621 19000 -5500
rect 15000 -5653 15304 -5621
rect 15336 -5653 15464 -5621
rect 15496 -5653 15624 -5621
rect 15656 -5653 15784 -5621
rect 15816 -5653 15944 -5621
rect 15976 -5653 16104 -5621
rect 16136 -5653 16264 -5621
rect 16296 -5653 16424 -5621
rect 16456 -5653 16584 -5621
rect 16616 -5653 16744 -5621
rect 16776 -5653 16904 -5621
rect 16936 -5653 17064 -5621
rect 17096 -5653 17224 -5621
rect 17256 -5653 17384 -5621
rect 17416 -5653 17544 -5621
rect 17576 -5653 17704 -5621
rect 17736 -5653 17864 -5621
rect 17896 -5653 18024 -5621
rect 18056 -5653 18184 -5621
rect 18216 -5653 18344 -5621
rect 18376 -5653 18504 -5621
rect 18536 -5653 18664 -5621
rect 18696 -5653 19000 -5621
rect 15000 -5724 19000 -5653
rect 15000 -5756 15119 -5724
rect 15151 -5756 18852 -5724
rect 18884 -5756 19000 -5724
rect 15000 -5770 19000 -5756
rect 15000 -5884 15270 -5770
rect 15000 -5916 15119 -5884
rect 15151 -5916 15270 -5884
rect 15000 -6044 15270 -5916
rect 15000 -6076 15119 -6044
rect 15151 -6076 15270 -6044
rect 15000 -6204 15270 -6076
rect 15000 -6236 15119 -6204
rect 15151 -6236 15270 -6204
rect 15000 -6364 15270 -6236
rect 15000 -6396 15119 -6364
rect 15151 -6396 15270 -6364
rect 15000 -6524 15270 -6396
rect 15000 -6556 15119 -6524
rect 15151 -6556 15270 -6524
rect 15000 -6684 15270 -6556
rect 15000 -6716 15119 -6684
rect 15151 -6716 15270 -6684
rect 15000 -6844 15270 -6716
rect 15000 -6876 15119 -6844
rect 15151 -6876 15270 -6844
rect 15000 -7004 15270 -6876
rect 15000 -7036 15119 -7004
rect 15151 -7036 15270 -7004
rect 15000 -7164 15270 -7036
rect 15000 -7196 15119 -7164
rect 15151 -7196 15270 -7164
rect 15000 -7324 15270 -7196
rect 15000 -7356 15119 -7324
rect 15151 -7356 15270 -7324
rect 15000 -7484 15270 -7356
rect 15000 -7516 15119 -7484
rect 15151 -7516 15270 -7484
rect 15000 -7644 15270 -7516
rect 15000 -7675 15119 -7644
rect 13300 -7676 15119 -7675
rect 15151 -7676 15270 -7644
rect 13300 -7715 15270 -7676
rect 13200 -7835 14585 -7795
rect 12730 -7964 13000 -7836
rect 12730 -7996 12852 -7964
rect 12884 -7996 13000 -7964
rect 12730 -8124 13000 -7996
rect 12730 -8156 12852 -8124
rect 12884 -8156 13000 -8124
rect 12730 -8284 13000 -8156
rect 12730 -8316 12852 -8284
rect 12884 -8316 13000 -8284
rect 12730 -8444 13000 -8316
rect 12730 -8476 12852 -8444
rect 12884 -8476 13000 -8444
rect 12730 -8604 13000 -8476
rect 12730 -8636 12852 -8604
rect 12884 -8636 13000 -8604
rect 12730 -8764 13000 -8636
rect 12730 -8796 12852 -8764
rect 12884 -8796 13000 -8764
rect 12730 -8924 13000 -8796
rect 12730 -8956 12852 -8924
rect 12884 -8956 13000 -8924
rect 12730 -9084 13000 -8956
rect 12730 -9116 12852 -9084
rect 12884 -9116 13000 -9084
rect 12730 -9230 13000 -9116
rect 9000 -9244 13000 -9230
rect 9000 -9276 9119 -9244
rect 9151 -9276 12852 -9244
rect 12884 -9276 13000 -9244
rect 9000 -9349 13000 -9276
rect 9000 -9381 9304 -9349
rect 9336 -9381 9464 -9349
rect 9496 -9381 9624 -9349
rect 9656 -9381 9784 -9349
rect 9816 -9381 9944 -9349
rect 9976 -9381 10104 -9349
rect 10136 -9381 10264 -9349
rect 10296 -9381 10424 -9349
rect 10456 -9381 10584 -9349
rect 10616 -9381 10744 -9349
rect 10776 -9381 10904 -9349
rect 10936 -9381 11064 -9349
rect 11096 -9381 11224 -9349
rect 11256 -9381 11384 -9349
rect 11416 -9381 11544 -9349
rect 11576 -9381 11704 -9349
rect 11736 -9381 11864 -9349
rect 11896 -9381 12024 -9349
rect 12056 -9381 12184 -9349
rect 12216 -9381 12344 -9349
rect 12376 -9381 12504 -9349
rect 12536 -9381 12664 -9349
rect 12696 -9381 13000 -9349
rect 9000 -9500 13000 -9381
rect 14545 -11120 14585 -7835
rect 15000 -7804 15270 -7715
rect 15000 -7836 15119 -7804
rect 15151 -7836 15270 -7804
rect 15000 -7964 15270 -7836
rect 15000 -7996 15119 -7964
rect 15151 -7996 15270 -7964
rect 15000 -8124 15270 -7996
rect 15000 -8156 15119 -8124
rect 15151 -8156 15270 -8124
rect 15000 -8284 15270 -8156
rect 15000 -8316 15119 -8284
rect 15151 -8316 15270 -8284
rect 15000 -8444 15270 -8316
rect 15000 -8476 15119 -8444
rect 15151 -8476 15270 -8444
rect 15000 -8604 15270 -8476
rect 15000 -8636 15119 -8604
rect 15151 -8636 15270 -8604
rect 15000 -8764 15270 -8636
rect 15000 -8796 15119 -8764
rect 15151 -8796 15270 -8764
rect 15000 -8924 15270 -8796
rect 15000 -8956 15119 -8924
rect 15151 -8956 15270 -8924
rect 15000 -9084 15270 -8956
rect 15000 -9116 15119 -9084
rect 15151 -9116 15270 -9084
rect 15000 -9230 15270 -9116
rect 18730 -5884 19000 -5770
rect 18730 -5916 18852 -5884
rect 18884 -5916 19000 -5884
rect 18730 -6044 19000 -5916
rect 18730 -6076 18852 -6044
rect 18884 -6076 19000 -6044
rect 18730 -6204 19000 -6076
rect 18730 -6236 18852 -6204
rect 18884 -6236 19000 -6204
rect 18730 -6364 19000 -6236
rect 18730 -6396 18852 -6364
rect 18884 -6396 19000 -6364
rect 18730 -6524 19000 -6396
rect 18730 -6556 18852 -6524
rect 18884 -6556 19000 -6524
rect 18730 -6684 19000 -6556
rect 18730 -6716 18852 -6684
rect 18884 -6716 19000 -6684
rect 18730 -6844 19000 -6716
rect 18730 -6876 18852 -6844
rect 18884 -6876 19000 -6844
rect 18730 -7004 19000 -6876
rect 18730 -7036 18852 -7004
rect 18884 -7036 19000 -7004
rect 18730 -7164 19000 -7036
rect 18730 -7196 18852 -7164
rect 18884 -7196 19000 -7164
rect 18730 -7324 19000 -7196
rect 18730 -7356 18852 -7324
rect 18884 -7356 19000 -7324
rect 18730 -7484 19000 -7356
rect 18730 -7516 18852 -7484
rect 18884 -7516 19000 -7484
rect 18730 -7644 19000 -7516
rect 18730 -7676 18852 -7644
rect 18884 -7676 19000 -7644
rect 18730 -7804 19000 -7676
rect 18730 -7836 18852 -7804
rect 18884 -7836 19000 -7804
rect 18730 -7964 19000 -7836
rect 18730 -7996 18852 -7964
rect 18884 -7996 19000 -7964
rect 18730 -8124 19000 -7996
rect 18730 -8156 18852 -8124
rect 18884 -8156 19000 -8124
rect 18730 -8284 19000 -8156
rect 18730 -8316 18852 -8284
rect 18884 -8316 19000 -8284
rect 18730 -8444 19000 -8316
rect 18730 -8476 18852 -8444
rect 18884 -8476 19000 -8444
rect 18730 -8604 19000 -8476
rect 18730 -8636 18852 -8604
rect 18884 -8636 19000 -8604
rect 18730 -8764 19000 -8636
rect 18730 -8796 18852 -8764
rect 18884 -8796 19000 -8764
rect 18730 -8924 19000 -8796
rect 18730 -8956 18852 -8924
rect 18884 -8956 19000 -8924
rect 18730 -9084 19000 -8956
rect 18730 -9116 18852 -9084
rect 18884 -9116 19000 -9084
rect 18730 -9230 19000 -9116
rect 15000 -9244 19000 -9230
rect 15000 -9276 15119 -9244
rect 15151 -9276 18852 -9244
rect 18884 -9276 19000 -9244
rect 15000 -9349 19000 -9276
rect 15000 -9381 15304 -9349
rect 15336 -9381 15464 -9349
rect 15496 -9381 15624 -9349
rect 15656 -9381 15784 -9349
rect 15816 -9381 15944 -9349
rect 15976 -9381 16104 -9349
rect 16136 -9381 16264 -9349
rect 16296 -9381 16424 -9349
rect 16456 -9381 16584 -9349
rect 16616 -9381 16744 -9349
rect 16776 -9381 16904 -9349
rect 16936 -9381 17064 -9349
rect 17096 -9381 17224 -9349
rect 17256 -9381 17384 -9349
rect 17416 -9381 17544 -9349
rect 17576 -9381 17704 -9349
rect 17736 -9381 17864 -9349
rect 17896 -9381 18024 -9349
rect 18056 -9381 18184 -9349
rect 18216 -9381 18344 -9349
rect 18376 -9381 18504 -9349
rect 18536 -9381 18664 -9349
rect 18696 -9381 19000 -9349
rect 15000 -9500 19000 -9381
rect 21000 -5621 25000 -5500
rect 21000 -5653 21304 -5621
rect 21336 -5653 21464 -5621
rect 21496 -5653 21624 -5621
rect 21656 -5653 21784 -5621
rect 21816 -5653 21944 -5621
rect 21976 -5653 22104 -5621
rect 22136 -5653 22264 -5621
rect 22296 -5653 22424 -5621
rect 22456 -5653 22584 -5621
rect 22616 -5653 22744 -5621
rect 22776 -5653 22904 -5621
rect 22936 -5653 23064 -5621
rect 23096 -5653 23224 -5621
rect 23256 -5653 23384 -5621
rect 23416 -5653 23544 -5621
rect 23576 -5653 23704 -5621
rect 23736 -5653 23864 -5621
rect 23896 -5653 24024 -5621
rect 24056 -5653 24184 -5621
rect 24216 -5653 24344 -5621
rect 24376 -5653 24504 -5621
rect 24536 -5653 24664 -5621
rect 24696 -5653 25000 -5621
rect 21000 -5724 25000 -5653
rect 21000 -5756 21119 -5724
rect 21151 -5756 24852 -5724
rect 24884 -5756 25000 -5724
rect 21000 -5770 25000 -5756
rect 21000 -5884 21270 -5770
rect 21000 -5916 21119 -5884
rect 21151 -5916 21270 -5884
rect 21000 -6044 21270 -5916
rect 21000 -6076 21119 -6044
rect 21151 -6076 21270 -6044
rect 21000 -6204 21270 -6076
rect 21000 -6236 21119 -6204
rect 21151 -6236 21270 -6204
rect 21000 -6364 21270 -6236
rect 21000 -6396 21119 -6364
rect 21151 -6396 21270 -6364
rect 21000 -6524 21270 -6396
rect 21000 -6556 21119 -6524
rect 21151 -6556 21270 -6524
rect 21000 -6684 21270 -6556
rect 21000 -6716 21119 -6684
rect 21151 -6716 21270 -6684
rect 21000 -6844 21270 -6716
rect 21000 -6876 21119 -6844
rect 21151 -6876 21270 -6844
rect 21000 -7004 21270 -6876
rect 21000 -7036 21119 -7004
rect 21151 -7036 21270 -7004
rect 21000 -7164 21270 -7036
rect 21000 -7196 21119 -7164
rect 21151 -7196 21270 -7164
rect 21000 -7324 21270 -7196
rect 21000 -7356 21119 -7324
rect 21151 -7356 21270 -7324
rect 21000 -7484 21270 -7356
rect 21000 -7516 21119 -7484
rect 21151 -7516 21270 -7484
rect 21000 -7644 21270 -7516
rect 21000 -7676 21119 -7644
rect 21151 -7676 21270 -7644
rect 21000 -7804 21270 -7676
rect 21000 -7836 21119 -7804
rect 21151 -7836 21270 -7804
rect 21000 -7964 21270 -7836
rect 21000 -7996 21119 -7964
rect 21151 -7996 21270 -7964
rect 21000 -8124 21270 -7996
rect 21000 -8156 21119 -8124
rect 21151 -8156 21270 -8124
rect 21000 -8284 21270 -8156
rect 21000 -8316 21119 -8284
rect 21151 -8316 21270 -8284
rect 21000 -8444 21270 -8316
rect 21000 -8476 21119 -8444
rect 21151 -8476 21270 -8444
rect 21000 -8604 21270 -8476
rect 21000 -8636 21119 -8604
rect 21151 -8636 21270 -8604
rect 21000 -8764 21270 -8636
rect 21000 -8796 21119 -8764
rect 21151 -8796 21270 -8764
rect 21000 -8924 21270 -8796
rect 21000 -8956 21119 -8924
rect 21151 -8956 21270 -8924
rect 21000 -9084 21270 -8956
rect 21000 -9116 21119 -9084
rect 21151 -9116 21270 -9084
rect 21000 -9230 21270 -9116
rect 24730 -5884 25000 -5770
rect 24730 -5916 24852 -5884
rect 24884 -5916 25000 -5884
rect 24730 -6044 25000 -5916
rect 24730 -6076 24852 -6044
rect 24884 -6076 25000 -6044
rect 24730 -6204 25000 -6076
rect 24730 -6236 24852 -6204
rect 24884 -6236 25000 -6204
rect 24730 -6364 25000 -6236
rect 24730 -6396 24852 -6364
rect 24884 -6396 25000 -6364
rect 24730 -6524 25000 -6396
rect 24730 -6556 24852 -6524
rect 24884 -6556 25000 -6524
rect 24730 -6684 25000 -6556
rect 24730 -6716 24852 -6684
rect 24884 -6716 25000 -6684
rect 24730 -6844 25000 -6716
rect 24730 -6876 24852 -6844
rect 24884 -6876 25000 -6844
rect 24730 -7004 25000 -6876
rect 24730 -7036 24852 -7004
rect 24884 -7036 25000 -7004
rect 24730 -7164 25000 -7036
rect 24730 -7196 24852 -7164
rect 24884 -7196 25000 -7164
rect 24730 -7324 25000 -7196
rect 24730 -7356 24852 -7324
rect 24884 -7356 25000 -7324
rect 24730 -7484 25000 -7356
rect 24730 -7516 24852 -7484
rect 24884 -7516 25000 -7484
rect 24730 -7644 25000 -7516
rect 24730 -7676 24852 -7644
rect 24884 -7676 25000 -7644
rect 24730 -7804 25000 -7676
rect 24730 -7836 24852 -7804
rect 24884 -7836 25000 -7804
rect 24730 -7964 25000 -7836
rect 24730 -7996 24852 -7964
rect 24884 -7996 25000 -7964
rect 24730 -8124 25000 -7996
rect 24730 -8156 24852 -8124
rect 24884 -8156 25000 -8124
rect 24730 -8284 25000 -8156
rect 24730 -8316 24852 -8284
rect 24884 -8316 25000 -8284
rect 24730 -8444 25000 -8316
rect 24730 -8476 24852 -8444
rect 24884 -8476 25000 -8444
rect 24730 -8604 25000 -8476
rect 24730 -8636 24852 -8604
rect 24884 -8636 25000 -8604
rect 24730 -8764 25000 -8636
rect 24730 -8796 24852 -8764
rect 24884 -8796 25000 -8764
rect 24730 -8924 25000 -8796
rect 24730 -8956 24852 -8924
rect 24884 -8956 25000 -8924
rect 24730 -9084 25000 -8956
rect 24730 -9116 24852 -9084
rect 24884 -9116 25000 -9084
rect 24730 -9230 25000 -9116
rect 21000 -9244 25000 -9230
rect 21000 -9276 21119 -9244
rect 21151 -9276 24852 -9244
rect 24884 -9276 25000 -9244
rect 21000 -9349 25000 -9276
rect 21000 -9381 21304 -9349
rect 21336 -9381 21464 -9349
rect 21496 -9381 21624 -9349
rect 21656 -9381 21784 -9349
rect 21816 -9381 21944 -9349
rect 21976 -9381 22104 -9349
rect 22136 -9381 22264 -9349
rect 22296 -9381 22424 -9349
rect 22456 -9381 22584 -9349
rect 22616 -9381 22744 -9349
rect 22776 -9381 22904 -9349
rect 22936 -9381 23064 -9349
rect 23096 -9381 23224 -9349
rect 23256 -9381 23384 -9349
rect 23416 -9381 23544 -9349
rect 23576 -9381 23704 -9349
rect 23736 -9381 23864 -9349
rect 23896 -9381 24024 -9349
rect 24056 -9381 24184 -9349
rect 24216 -9381 24344 -9349
rect 24376 -9381 24504 -9349
rect 24536 -9381 24664 -9349
rect 24696 -9381 25000 -9349
rect 21000 -9500 25000 -9381
rect 14545 -11160 21375 -11120
rect 8300 -11360 14150 -11330
rect 9000 -11621 13000 -11500
rect 9000 -11653 9304 -11621
rect 9336 -11653 9464 -11621
rect 9496 -11653 9624 -11621
rect 9656 -11653 9784 -11621
rect 9816 -11653 9944 -11621
rect 9976 -11653 10104 -11621
rect 10136 -11653 10264 -11621
rect 10296 -11653 10424 -11621
rect 10456 -11653 10584 -11621
rect 10616 -11653 10744 -11621
rect 10776 -11653 10904 -11621
rect 10936 -11653 11064 -11621
rect 11096 -11653 11224 -11621
rect 11256 -11653 11384 -11621
rect 11416 -11653 11544 -11621
rect 11576 -11653 11704 -11621
rect 11736 -11653 11864 -11621
rect 11896 -11653 12024 -11621
rect 12056 -11653 12184 -11621
rect 12216 -11653 12344 -11621
rect 12376 -11653 12504 -11621
rect 12536 -11653 12664 -11621
rect 12696 -11653 13000 -11621
rect 9000 -11724 13000 -11653
rect 9000 -11756 9119 -11724
rect 9151 -11756 12852 -11724
rect 12884 -11756 13000 -11724
rect 9000 -11770 13000 -11756
rect 9000 -11884 9270 -11770
rect 9000 -11916 9119 -11884
rect 9151 -11916 9270 -11884
rect 9000 -12044 9270 -11916
rect 9000 -12076 9119 -12044
rect 9151 -12076 9270 -12044
rect 9000 -12204 9270 -12076
rect 9000 -12236 9119 -12204
rect 9151 -12236 9270 -12204
rect 9000 -12364 9270 -12236
rect 9000 -12396 9119 -12364
rect 9151 -12396 9270 -12364
rect 9000 -12524 9270 -12396
rect 9000 -12556 9119 -12524
rect 9151 -12556 9270 -12524
rect 9000 -12684 9270 -12556
rect 9000 -12716 9119 -12684
rect 9151 -12716 9270 -12684
rect 9000 -12844 9270 -12716
rect 9000 -12875 9119 -12844
rect 8230 -12876 9119 -12875
rect 9151 -12876 9270 -12844
rect 6730 -13004 7000 -12900
rect 8230 -12905 9270 -12876
rect 6730 -13036 6852 -13004
rect 6884 -13036 7000 -13004
rect 6730 -13164 7000 -13036
rect 6730 -13196 6852 -13164
rect 6884 -13196 7000 -13164
rect 6730 -13324 7000 -13196
rect 6730 -13356 6852 -13324
rect 6884 -13356 7000 -13324
rect 6730 -13484 7000 -13356
rect 6730 -13516 6852 -13484
rect 6884 -13516 7000 -13484
rect 6730 -13644 7000 -13516
rect 6730 -13676 6852 -13644
rect 6884 -13676 7000 -13644
rect 6730 -13804 7000 -13676
rect 6730 -13836 6852 -13804
rect 6884 -13836 7000 -13804
rect 6730 -13964 7000 -13836
rect 6730 -13996 6852 -13964
rect 6884 -13996 7000 -13964
rect 6730 -14124 7000 -13996
rect 6730 -14156 6852 -14124
rect 6884 -14156 7000 -14124
rect 6730 -14284 7000 -14156
rect 6730 -14316 6852 -14284
rect 6884 -14316 7000 -14284
rect 6730 -14444 7000 -14316
rect 6730 -14476 6852 -14444
rect 6884 -14476 7000 -14444
rect 6730 -14604 7000 -14476
rect 6730 -14636 6852 -14604
rect 6884 -14636 7000 -14604
rect 6730 -14764 7000 -14636
rect 6730 -14796 6852 -14764
rect 6884 -14796 7000 -14764
rect 6730 -14924 7000 -14796
rect 6730 -14956 6852 -14924
rect 6884 -14956 7000 -14924
rect 6730 -15084 7000 -14956
rect 6730 -15116 6852 -15084
rect 6884 -15116 7000 -15084
rect 6730 -15230 7000 -15116
rect 3000 -15244 7000 -15230
rect 3000 -15276 3119 -15244
rect 3151 -15276 6852 -15244
rect 6884 -15276 7000 -15244
rect 3000 -15349 7000 -15276
rect 3000 -15381 3304 -15349
rect 3336 -15381 3464 -15349
rect 3496 -15381 3624 -15349
rect 3656 -15381 3784 -15349
rect 3816 -15381 3944 -15349
rect 3976 -15381 4104 -15349
rect 4136 -15381 4264 -15349
rect 4296 -15381 4424 -15349
rect 4456 -15381 4584 -15349
rect 4616 -15381 4744 -15349
rect 4776 -15381 4904 -15349
rect 4936 -15381 5064 -15349
rect 5096 -15381 5224 -15349
rect 5256 -15381 5384 -15349
rect 5416 -15381 5544 -15349
rect 5576 -15381 5704 -15349
rect 5736 -15381 5864 -15349
rect 5896 -15381 6024 -15349
rect 6056 -15381 6184 -15349
rect 6216 -15381 6344 -15349
rect 6376 -15381 6504 -15349
rect 6536 -15381 6664 -15349
rect 6696 -15381 7000 -15349
rect 3000 -15500 7000 -15381
rect 9000 -13004 9270 -12905
rect 9000 -13036 9119 -13004
rect 9151 -13036 9270 -13004
rect 9000 -13164 9270 -13036
rect 9000 -13196 9119 -13164
rect 9151 -13196 9270 -13164
rect 9000 -13324 9270 -13196
rect 9000 -13356 9119 -13324
rect 9151 -13356 9270 -13324
rect 9000 -13484 9270 -13356
rect 9000 -13516 9119 -13484
rect 9151 -13516 9270 -13484
rect 9000 -13644 9270 -13516
rect 9000 -13676 9119 -13644
rect 9151 -13676 9270 -13644
rect 9000 -13804 9270 -13676
rect 9000 -13836 9119 -13804
rect 9151 -13836 9270 -13804
rect 9000 -13964 9270 -13836
rect 9000 -13996 9119 -13964
rect 9151 -13996 9270 -13964
rect 9000 -14124 9270 -13996
rect 9000 -14156 9119 -14124
rect 9151 -14156 9270 -14124
rect 9000 -14284 9270 -14156
rect 9000 -14316 9119 -14284
rect 9151 -14316 9270 -14284
rect 9000 -14444 9270 -14316
rect 9000 -14476 9119 -14444
rect 9151 -14476 9270 -14444
rect 9000 -14604 9270 -14476
rect 9000 -14636 9119 -14604
rect 9151 -14636 9270 -14604
rect 9000 -14764 9270 -14636
rect 9000 -14796 9119 -14764
rect 9151 -14796 9270 -14764
rect 9000 -14924 9270 -14796
rect 9000 -14956 9119 -14924
rect 9151 -14956 9270 -14924
rect 9000 -15084 9270 -14956
rect 9000 -15116 9119 -15084
rect 9151 -15116 9270 -15084
rect 9000 -15230 9270 -15116
rect 12730 -11884 13000 -11770
rect 12730 -11916 12852 -11884
rect 12884 -11916 13000 -11884
rect 12730 -12044 13000 -11916
rect 12730 -12076 12852 -12044
rect 12884 -12076 13000 -12044
rect 12730 -12204 13000 -12076
rect 12730 -12236 12852 -12204
rect 12884 -12236 13000 -12204
rect 12730 -12364 13000 -12236
rect 12730 -12396 12852 -12364
rect 12884 -12396 13000 -12364
rect 12730 -12524 13000 -12396
rect 12730 -12556 12852 -12524
rect 12884 -12556 13000 -12524
rect 12730 -12684 13000 -12556
rect 12730 -12716 12852 -12684
rect 12884 -12716 13000 -12684
rect 12730 -12844 13000 -12716
rect 12730 -12876 12852 -12844
rect 12884 -12876 13000 -12844
rect 12730 -13004 13000 -12876
rect 14120 -12870 14150 -11360
rect 21335 -11500 21375 -11160
rect 15000 -11621 19000 -11500
rect 15000 -11653 15304 -11621
rect 15336 -11653 15464 -11621
rect 15496 -11653 15624 -11621
rect 15656 -11653 15784 -11621
rect 15816 -11653 15944 -11621
rect 15976 -11653 16104 -11621
rect 16136 -11653 16264 -11621
rect 16296 -11653 16424 -11621
rect 16456 -11653 16584 -11621
rect 16616 -11653 16744 -11621
rect 16776 -11653 16904 -11621
rect 16936 -11653 17064 -11621
rect 17096 -11653 17224 -11621
rect 17256 -11653 17384 -11621
rect 17416 -11653 17544 -11621
rect 17576 -11653 17704 -11621
rect 17736 -11653 17864 -11621
rect 17896 -11653 18024 -11621
rect 18056 -11653 18184 -11621
rect 18216 -11653 18344 -11621
rect 18376 -11653 18504 -11621
rect 18536 -11653 18664 -11621
rect 18696 -11653 19000 -11621
rect 15000 -11724 19000 -11653
rect 15000 -11756 15119 -11724
rect 15151 -11756 18852 -11724
rect 18884 -11756 19000 -11724
rect 15000 -11770 19000 -11756
rect 15000 -11884 15270 -11770
rect 15000 -11916 15119 -11884
rect 15151 -11916 15270 -11884
rect 15000 -12044 15270 -11916
rect 15000 -12076 15119 -12044
rect 15151 -12076 15270 -12044
rect 15000 -12204 15270 -12076
rect 15000 -12236 15119 -12204
rect 15151 -12236 15270 -12204
rect 15000 -12364 15270 -12236
rect 15000 -12396 15119 -12364
rect 15151 -12396 15270 -12364
rect 15000 -12524 15270 -12396
rect 15000 -12556 15119 -12524
rect 15151 -12556 15270 -12524
rect 15000 -12684 15270 -12556
rect 15000 -12716 15119 -12684
rect 15151 -12716 15270 -12684
rect 15000 -12844 15270 -12716
rect 15000 -12870 15119 -12844
rect 14120 -12876 15119 -12870
rect 15151 -12876 15270 -12844
rect 14120 -12900 15270 -12876
rect 12730 -13036 12852 -13004
rect 12884 -13036 13000 -13004
rect 12730 -13164 13000 -13036
rect 12730 -13196 12852 -13164
rect 12884 -13196 13000 -13164
rect 12730 -13324 13000 -13196
rect 12730 -13356 12852 -13324
rect 12884 -13356 13000 -13324
rect 12730 -13484 13000 -13356
rect 12730 -13516 12852 -13484
rect 12884 -13516 13000 -13484
rect 12730 -13644 13000 -13516
rect 12730 -13676 12852 -13644
rect 12884 -13676 13000 -13644
rect 12730 -13804 13000 -13676
rect 12730 -13836 12852 -13804
rect 12884 -13836 13000 -13804
rect 12730 -13964 13000 -13836
rect 12730 -13996 12852 -13964
rect 12884 -13996 13000 -13964
rect 12730 -14124 13000 -13996
rect 12730 -14156 12852 -14124
rect 12884 -14156 13000 -14124
rect 12730 -14284 13000 -14156
rect 12730 -14316 12852 -14284
rect 12884 -14316 13000 -14284
rect 12730 -14444 13000 -14316
rect 12730 -14476 12852 -14444
rect 12884 -14476 13000 -14444
rect 12730 -14604 13000 -14476
rect 12730 -14636 12852 -14604
rect 12884 -14636 13000 -14604
rect 12730 -14764 13000 -14636
rect 12730 -14796 12852 -14764
rect 12884 -14796 13000 -14764
rect 12730 -14924 13000 -14796
rect 12730 -14956 12852 -14924
rect 12884 -14956 13000 -14924
rect 12730 -15084 13000 -14956
rect 12730 -15116 12852 -15084
rect 12884 -15116 13000 -15084
rect 12730 -15230 13000 -15116
rect 9000 -15244 13000 -15230
rect 9000 -15276 9119 -15244
rect 9151 -15276 12852 -15244
rect 12884 -15276 13000 -15244
rect 9000 -15349 13000 -15276
rect 9000 -15381 9304 -15349
rect 9336 -15381 9464 -15349
rect 9496 -15381 9624 -15349
rect 9656 -15381 9784 -15349
rect 9816 -15381 9944 -15349
rect 9976 -15381 10104 -15349
rect 10136 -15381 10264 -15349
rect 10296 -15381 10424 -15349
rect 10456 -15381 10584 -15349
rect 10616 -15381 10744 -15349
rect 10776 -15381 10904 -15349
rect 10936 -15381 11064 -15349
rect 11096 -15381 11224 -15349
rect 11256 -15381 11384 -15349
rect 11416 -15381 11544 -15349
rect 11576 -15381 11704 -15349
rect 11736 -15381 11864 -15349
rect 11896 -15381 12024 -15349
rect 12056 -15381 12184 -15349
rect 12216 -15381 12344 -15349
rect 12376 -15381 12504 -15349
rect 12536 -15381 12664 -15349
rect 12696 -15381 13000 -15349
rect 9000 -15500 13000 -15381
rect 15000 -13004 15270 -12900
rect 15000 -13036 15119 -13004
rect 15151 -13036 15270 -13004
rect 15000 -13164 15270 -13036
rect 15000 -13196 15119 -13164
rect 15151 -13196 15270 -13164
rect 15000 -13324 15270 -13196
rect 15000 -13356 15119 -13324
rect 15151 -13356 15270 -13324
rect 15000 -13484 15270 -13356
rect 15000 -13516 15119 -13484
rect 15151 -13516 15270 -13484
rect 15000 -13644 15270 -13516
rect 15000 -13676 15119 -13644
rect 15151 -13676 15270 -13644
rect 15000 -13804 15270 -13676
rect 15000 -13836 15119 -13804
rect 15151 -13836 15270 -13804
rect 15000 -13964 15270 -13836
rect 15000 -13996 15119 -13964
rect 15151 -13996 15270 -13964
rect 15000 -14124 15270 -13996
rect 15000 -14156 15119 -14124
rect 15151 -14156 15270 -14124
rect 15000 -14284 15270 -14156
rect 15000 -14316 15119 -14284
rect 15151 -14316 15270 -14284
rect 15000 -14444 15270 -14316
rect 15000 -14476 15119 -14444
rect 15151 -14476 15270 -14444
rect 15000 -14604 15270 -14476
rect 15000 -14636 15119 -14604
rect 15151 -14636 15270 -14604
rect 15000 -14764 15270 -14636
rect 15000 -14796 15119 -14764
rect 15151 -14796 15270 -14764
rect 15000 -14924 15270 -14796
rect 15000 -14956 15119 -14924
rect 15151 -14956 15270 -14924
rect 15000 -15084 15270 -14956
rect 15000 -15116 15119 -15084
rect 15151 -15116 15270 -15084
rect 15000 -15230 15270 -15116
rect 18730 -11884 19000 -11770
rect 18730 -11916 18852 -11884
rect 18884 -11916 19000 -11884
rect 18730 -12044 19000 -11916
rect 18730 -12076 18852 -12044
rect 18884 -12076 19000 -12044
rect 18730 -12204 19000 -12076
rect 18730 -12236 18852 -12204
rect 18884 -12236 19000 -12204
rect 18730 -12364 19000 -12236
rect 18730 -12396 18852 -12364
rect 18884 -12396 19000 -12364
rect 18730 -12524 19000 -12396
rect 18730 -12556 18852 -12524
rect 18884 -12556 19000 -12524
rect 18730 -12684 19000 -12556
rect 18730 -12716 18852 -12684
rect 18884 -12716 19000 -12684
rect 18730 -12844 19000 -12716
rect 18730 -12876 18852 -12844
rect 18884 -12876 19000 -12844
rect 18730 -13004 19000 -12876
rect 18730 -13036 18852 -13004
rect 18884 -13036 19000 -13004
rect 18730 -13164 19000 -13036
rect 18730 -13196 18852 -13164
rect 18884 -13196 19000 -13164
rect 18730 -13324 19000 -13196
rect 18730 -13356 18852 -13324
rect 18884 -13356 19000 -13324
rect 18730 -13484 19000 -13356
rect 18730 -13516 18852 -13484
rect 18884 -13516 19000 -13484
rect 18730 -13644 19000 -13516
rect 18730 -13676 18852 -13644
rect 18884 -13676 19000 -13644
rect 18730 -13804 19000 -13676
rect 18730 -13836 18852 -13804
rect 18884 -13836 19000 -13804
rect 18730 -13964 19000 -13836
rect 18730 -13996 18852 -13964
rect 18884 -13996 19000 -13964
rect 18730 -14124 19000 -13996
rect 18730 -14156 18852 -14124
rect 18884 -14156 19000 -14124
rect 18730 -14284 19000 -14156
rect 18730 -14316 18852 -14284
rect 18884 -14316 19000 -14284
rect 18730 -14444 19000 -14316
rect 18730 -14476 18852 -14444
rect 18884 -14476 19000 -14444
rect 18730 -14604 19000 -14476
rect 18730 -14636 18852 -14604
rect 18884 -14636 19000 -14604
rect 18730 -14764 19000 -14636
rect 18730 -14796 18852 -14764
rect 18884 -14796 19000 -14764
rect 18730 -14924 19000 -14796
rect 18730 -14956 18852 -14924
rect 18884 -14956 19000 -14924
rect 18730 -15084 19000 -14956
rect 18730 -15116 18852 -15084
rect 18884 -15116 19000 -15084
rect 18730 -15230 19000 -15116
rect 15000 -15244 19000 -15230
rect 15000 -15276 15119 -15244
rect 15151 -15276 18852 -15244
rect 18884 -15276 19000 -15244
rect 15000 -15349 19000 -15276
rect 15000 -15381 15304 -15349
rect 15336 -15381 15464 -15349
rect 15496 -15381 15624 -15349
rect 15656 -15381 15784 -15349
rect 15816 -15381 15944 -15349
rect 15976 -15381 16104 -15349
rect 16136 -15381 16264 -15349
rect 16296 -15381 16424 -15349
rect 16456 -15381 16584 -15349
rect 16616 -15381 16744 -15349
rect 16776 -15381 16904 -15349
rect 16936 -15381 17064 -15349
rect 17096 -15381 17224 -15349
rect 17256 -15381 17384 -15349
rect 17416 -15381 17544 -15349
rect 17576 -15381 17704 -15349
rect 17736 -15381 17864 -15349
rect 17896 -15381 18024 -15349
rect 18056 -15381 18184 -15349
rect 18216 -15381 18344 -15349
rect 18376 -15381 18504 -15349
rect 18536 -15381 18664 -15349
rect 18696 -15381 19000 -15349
rect 15000 -15500 19000 -15381
rect 21000 -11621 25000 -11500
rect 21000 -11653 21304 -11621
rect 21336 -11653 21464 -11621
rect 21496 -11653 21624 -11621
rect 21656 -11653 21784 -11621
rect 21816 -11653 21944 -11621
rect 21976 -11653 22104 -11621
rect 22136 -11653 22264 -11621
rect 22296 -11653 22424 -11621
rect 22456 -11653 22584 -11621
rect 22616 -11653 22744 -11621
rect 22776 -11653 22904 -11621
rect 22936 -11653 23064 -11621
rect 23096 -11653 23224 -11621
rect 23256 -11653 23384 -11621
rect 23416 -11653 23544 -11621
rect 23576 -11653 23704 -11621
rect 23736 -11653 23864 -11621
rect 23896 -11653 24024 -11621
rect 24056 -11653 24184 -11621
rect 24216 -11653 24344 -11621
rect 24376 -11653 24504 -11621
rect 24536 -11653 24664 -11621
rect 24696 -11653 25000 -11621
rect 21000 -11724 25000 -11653
rect 21000 -11756 21119 -11724
rect 21151 -11756 24852 -11724
rect 24884 -11756 25000 -11724
rect 21000 -11770 25000 -11756
rect 21000 -11884 21270 -11770
rect 21000 -11916 21119 -11884
rect 21151 -11916 21270 -11884
rect 21000 -12044 21270 -11916
rect 21000 -12076 21119 -12044
rect 21151 -12076 21270 -12044
rect 21000 -12204 21270 -12076
rect 21000 -12236 21119 -12204
rect 21151 -12236 21270 -12204
rect 21000 -12364 21270 -12236
rect 21000 -12396 21119 -12364
rect 21151 -12396 21270 -12364
rect 21000 -12524 21270 -12396
rect 21000 -12556 21119 -12524
rect 21151 -12556 21270 -12524
rect 21000 -12684 21270 -12556
rect 21000 -12716 21119 -12684
rect 21151 -12716 21270 -12684
rect 21000 -12844 21270 -12716
rect 21000 -12876 21119 -12844
rect 21151 -12876 21270 -12844
rect 21000 -13004 21270 -12876
rect 21000 -13036 21119 -13004
rect 21151 -13036 21270 -13004
rect 21000 -13164 21270 -13036
rect 21000 -13196 21119 -13164
rect 21151 -13196 21270 -13164
rect 21000 -13324 21270 -13196
rect 21000 -13356 21119 -13324
rect 21151 -13356 21270 -13324
rect 21000 -13484 21270 -13356
rect 21000 -13516 21119 -13484
rect 21151 -13516 21270 -13484
rect 21000 -13644 21270 -13516
rect 21000 -13676 21119 -13644
rect 21151 -13676 21270 -13644
rect 21000 -13804 21270 -13676
rect 21000 -13836 21119 -13804
rect 21151 -13836 21270 -13804
rect 21000 -13964 21270 -13836
rect 21000 -13996 21119 -13964
rect 21151 -13996 21270 -13964
rect 21000 -14124 21270 -13996
rect 21000 -14156 21119 -14124
rect 21151 -14156 21270 -14124
rect 21000 -14284 21270 -14156
rect 21000 -14316 21119 -14284
rect 21151 -14316 21270 -14284
rect 21000 -14444 21270 -14316
rect 21000 -14476 21119 -14444
rect 21151 -14476 21270 -14444
rect 21000 -14604 21270 -14476
rect 21000 -14636 21119 -14604
rect 21151 -14636 21270 -14604
rect 21000 -14764 21270 -14636
rect 21000 -14796 21119 -14764
rect 21151 -14796 21270 -14764
rect 21000 -14924 21270 -14796
rect 21000 -14956 21119 -14924
rect 21151 -14956 21270 -14924
rect 21000 -15084 21270 -14956
rect 21000 -15116 21119 -15084
rect 21151 -15116 21270 -15084
rect 21000 -15230 21270 -15116
rect 24730 -11884 25000 -11770
rect 24730 -11916 24852 -11884
rect 24884 -11916 25000 -11884
rect 24730 -12044 25000 -11916
rect 24730 -12076 24852 -12044
rect 24884 -12076 25000 -12044
rect 24730 -12204 25000 -12076
rect 24730 -12236 24852 -12204
rect 24884 -12236 25000 -12204
rect 24730 -12364 25000 -12236
rect 24730 -12396 24852 -12364
rect 24884 -12396 25000 -12364
rect 24730 -12524 25000 -12396
rect 24730 -12556 24852 -12524
rect 24884 -12556 25000 -12524
rect 24730 -12684 25000 -12556
rect 24730 -12716 24852 -12684
rect 24884 -12716 25000 -12684
rect 24730 -12844 25000 -12716
rect 24730 -12876 24852 -12844
rect 24884 -12876 25000 -12844
rect 24730 -13004 25000 -12876
rect 24730 -13036 24852 -13004
rect 24884 -13036 25000 -13004
rect 24730 -13164 25000 -13036
rect 24730 -13196 24852 -13164
rect 24884 -13196 25000 -13164
rect 24730 -13324 25000 -13196
rect 24730 -13356 24852 -13324
rect 24884 -13356 25000 -13324
rect 24730 -13484 25000 -13356
rect 24730 -13516 24852 -13484
rect 24884 -13516 25000 -13484
rect 24730 -13644 25000 -13516
rect 24730 -13676 24852 -13644
rect 24884 -13676 25000 -13644
rect 24730 -13804 25000 -13676
rect 24730 -13836 24852 -13804
rect 24884 -13836 25000 -13804
rect 24730 -13964 25000 -13836
rect 24730 -13996 24852 -13964
rect 24884 -13996 25000 -13964
rect 24730 -14124 25000 -13996
rect 24730 -14156 24852 -14124
rect 24884 -14156 25000 -14124
rect 24730 -14284 25000 -14156
rect 24730 -14316 24852 -14284
rect 24884 -14316 25000 -14284
rect 24730 -14444 25000 -14316
rect 24730 -14476 24852 -14444
rect 24884 -14476 25000 -14444
rect 24730 -14604 25000 -14476
rect 24730 -14636 24852 -14604
rect 24884 -14636 25000 -14604
rect 24730 -14764 25000 -14636
rect 24730 -14796 24852 -14764
rect 24884 -14796 25000 -14764
rect 24730 -14924 25000 -14796
rect 24730 -14956 24852 -14924
rect 24884 -14956 25000 -14924
rect 24730 -15084 25000 -14956
rect 24730 -15116 24852 -15084
rect 24884 -15116 25000 -15084
rect 24730 -15230 25000 -15116
rect 21000 -15244 25000 -15230
rect 21000 -15276 21119 -15244
rect 21151 -15276 24852 -15244
rect 24884 -15276 25000 -15244
rect 21000 -15349 25000 -15276
rect 21000 -15381 21304 -15349
rect 21336 -15381 21464 -15349
rect 21496 -15381 21624 -15349
rect 21656 -15381 21784 -15349
rect 21816 -15381 21944 -15349
rect 21976 -15381 22104 -15349
rect 22136 -15381 22264 -15349
rect 22296 -15381 22424 -15349
rect 22456 -15381 22584 -15349
rect 22616 -15381 22744 -15349
rect 22776 -15381 22904 -15349
rect 22936 -15381 23064 -15349
rect 23096 -15381 23224 -15349
rect 23256 -15381 23384 -15349
rect 23416 -15381 23544 -15349
rect 23576 -15381 23704 -15349
rect 23736 -15381 23864 -15349
rect 23896 -15381 24024 -15349
rect 24056 -15381 24184 -15349
rect 24216 -15381 24344 -15349
rect 24376 -15381 24504 -15349
rect 24536 -15381 24664 -15349
rect 24696 -15381 25000 -15349
rect 21000 -15500 25000 -15381
<< via3 >>
rect 3304 -5623 3336 -5621
rect 3304 -5651 3306 -5623
rect 3306 -5651 3334 -5623
rect 3334 -5651 3336 -5623
rect 3304 -5653 3336 -5651
rect 3464 -5623 3496 -5621
rect 3464 -5651 3466 -5623
rect 3466 -5651 3494 -5623
rect 3494 -5651 3496 -5623
rect 3464 -5653 3496 -5651
rect 3624 -5623 3656 -5621
rect 3624 -5651 3626 -5623
rect 3626 -5651 3654 -5623
rect 3654 -5651 3656 -5623
rect 3624 -5653 3656 -5651
rect 3784 -5623 3816 -5621
rect 3784 -5651 3786 -5623
rect 3786 -5651 3814 -5623
rect 3814 -5651 3816 -5623
rect 3784 -5653 3816 -5651
rect 3944 -5623 3976 -5621
rect 3944 -5651 3946 -5623
rect 3946 -5651 3974 -5623
rect 3974 -5651 3976 -5623
rect 3944 -5653 3976 -5651
rect 4104 -5623 4136 -5621
rect 4104 -5651 4106 -5623
rect 4106 -5651 4134 -5623
rect 4134 -5651 4136 -5623
rect 4104 -5653 4136 -5651
rect 4264 -5623 4296 -5621
rect 4264 -5651 4266 -5623
rect 4266 -5651 4294 -5623
rect 4294 -5651 4296 -5623
rect 4264 -5653 4296 -5651
rect 4424 -5623 4456 -5621
rect 4424 -5651 4426 -5623
rect 4426 -5651 4454 -5623
rect 4454 -5651 4456 -5623
rect 4424 -5653 4456 -5651
rect 4584 -5623 4616 -5621
rect 4584 -5651 4586 -5623
rect 4586 -5651 4614 -5623
rect 4614 -5651 4616 -5623
rect 4584 -5653 4616 -5651
rect 4744 -5623 4776 -5621
rect 4744 -5651 4746 -5623
rect 4746 -5651 4774 -5623
rect 4774 -5651 4776 -5623
rect 4744 -5653 4776 -5651
rect 4904 -5623 4936 -5621
rect 4904 -5651 4906 -5623
rect 4906 -5651 4934 -5623
rect 4934 -5651 4936 -5623
rect 4904 -5653 4936 -5651
rect 5064 -5623 5096 -5621
rect 5064 -5651 5066 -5623
rect 5066 -5651 5094 -5623
rect 5094 -5651 5096 -5623
rect 5064 -5653 5096 -5651
rect 5224 -5623 5256 -5621
rect 5224 -5651 5226 -5623
rect 5226 -5651 5254 -5623
rect 5254 -5651 5256 -5623
rect 5224 -5653 5256 -5651
rect 5384 -5623 5416 -5621
rect 5384 -5651 5386 -5623
rect 5386 -5651 5414 -5623
rect 5414 -5651 5416 -5623
rect 5384 -5653 5416 -5651
rect 5544 -5623 5576 -5621
rect 5544 -5651 5546 -5623
rect 5546 -5651 5574 -5623
rect 5574 -5651 5576 -5623
rect 5544 -5653 5576 -5651
rect 5704 -5623 5736 -5621
rect 5704 -5651 5706 -5623
rect 5706 -5651 5734 -5623
rect 5734 -5651 5736 -5623
rect 5704 -5653 5736 -5651
rect 5864 -5623 5896 -5621
rect 5864 -5651 5866 -5623
rect 5866 -5651 5894 -5623
rect 5894 -5651 5896 -5623
rect 5864 -5653 5896 -5651
rect 6024 -5623 6056 -5621
rect 6024 -5651 6026 -5623
rect 6026 -5651 6054 -5623
rect 6054 -5651 6056 -5623
rect 6024 -5653 6056 -5651
rect 6184 -5623 6216 -5621
rect 6184 -5651 6186 -5623
rect 6186 -5651 6214 -5623
rect 6214 -5651 6216 -5623
rect 6184 -5653 6216 -5651
rect 6344 -5623 6376 -5621
rect 6344 -5651 6346 -5623
rect 6346 -5651 6374 -5623
rect 6374 -5651 6376 -5623
rect 6344 -5653 6376 -5651
rect 6504 -5623 6536 -5621
rect 6504 -5651 6506 -5623
rect 6506 -5651 6534 -5623
rect 6534 -5651 6536 -5623
rect 6504 -5653 6536 -5651
rect 6664 -5623 6696 -5621
rect 6664 -5651 6666 -5623
rect 6666 -5651 6694 -5623
rect 6694 -5651 6696 -5623
rect 6664 -5653 6696 -5651
rect 3119 -5726 3151 -5724
rect 3119 -5754 3121 -5726
rect 3121 -5754 3149 -5726
rect 3149 -5754 3151 -5726
rect 3119 -5756 3151 -5754
rect 6852 -5726 6884 -5724
rect 6852 -5754 6854 -5726
rect 6854 -5754 6882 -5726
rect 6882 -5754 6884 -5726
rect 6852 -5756 6884 -5754
rect 3119 -5886 3151 -5884
rect 3119 -5914 3121 -5886
rect 3121 -5914 3149 -5886
rect 3149 -5914 3151 -5886
rect 3119 -5916 3151 -5914
rect 3119 -6046 3151 -6044
rect 3119 -6074 3121 -6046
rect 3121 -6074 3149 -6046
rect 3149 -6074 3151 -6046
rect 3119 -6076 3151 -6074
rect 3119 -6206 3151 -6204
rect 3119 -6234 3121 -6206
rect 3121 -6234 3149 -6206
rect 3149 -6234 3151 -6206
rect 3119 -6236 3151 -6234
rect 3119 -6366 3151 -6364
rect 3119 -6394 3121 -6366
rect 3121 -6394 3149 -6366
rect 3149 -6394 3151 -6366
rect 3119 -6396 3151 -6394
rect 3119 -6526 3151 -6524
rect 3119 -6554 3121 -6526
rect 3121 -6554 3149 -6526
rect 3149 -6554 3151 -6526
rect 3119 -6556 3151 -6554
rect 3119 -6686 3151 -6684
rect 3119 -6714 3121 -6686
rect 3121 -6714 3149 -6686
rect 3149 -6714 3151 -6686
rect 3119 -6716 3151 -6714
rect 3119 -6846 3151 -6844
rect 3119 -6874 3121 -6846
rect 3121 -6874 3149 -6846
rect 3149 -6874 3151 -6846
rect 3119 -6876 3151 -6874
rect 3119 -7006 3151 -7004
rect 3119 -7034 3121 -7006
rect 3121 -7034 3149 -7006
rect 3149 -7034 3151 -7006
rect 3119 -7036 3151 -7034
rect 3119 -7166 3151 -7164
rect 3119 -7194 3121 -7166
rect 3121 -7194 3149 -7166
rect 3149 -7194 3151 -7166
rect 3119 -7196 3151 -7194
rect 3119 -7326 3151 -7324
rect 3119 -7354 3121 -7326
rect 3121 -7354 3149 -7326
rect 3149 -7354 3151 -7326
rect 3119 -7356 3151 -7354
rect 3119 -7486 3151 -7484
rect 3119 -7514 3121 -7486
rect 3121 -7514 3149 -7486
rect 3149 -7514 3151 -7486
rect 3119 -7516 3151 -7514
rect 3119 -7646 3151 -7644
rect 3119 -7674 3121 -7646
rect 3121 -7674 3149 -7646
rect 3149 -7674 3151 -7646
rect 3119 -7676 3151 -7674
rect 3119 -7806 3151 -7804
rect 3119 -7834 3121 -7806
rect 3121 -7834 3149 -7806
rect 3149 -7834 3151 -7806
rect 3119 -7836 3151 -7834
rect 3119 -7966 3151 -7964
rect 3119 -7994 3121 -7966
rect 3121 -7994 3149 -7966
rect 3149 -7994 3151 -7966
rect 3119 -7996 3151 -7994
rect 3119 -8126 3151 -8124
rect 3119 -8154 3121 -8126
rect 3121 -8154 3149 -8126
rect 3149 -8154 3151 -8126
rect 3119 -8156 3151 -8154
rect 3119 -8286 3151 -8284
rect 3119 -8314 3121 -8286
rect 3121 -8314 3149 -8286
rect 3149 -8314 3151 -8286
rect 3119 -8316 3151 -8314
rect 3119 -8446 3151 -8444
rect 3119 -8474 3121 -8446
rect 3121 -8474 3149 -8446
rect 3149 -8474 3151 -8446
rect 3119 -8476 3151 -8474
rect 3119 -8606 3151 -8604
rect 3119 -8634 3121 -8606
rect 3121 -8634 3149 -8606
rect 3149 -8634 3151 -8606
rect 3119 -8636 3151 -8634
rect 3119 -8766 3151 -8764
rect 3119 -8794 3121 -8766
rect 3121 -8794 3149 -8766
rect 3149 -8794 3151 -8766
rect 3119 -8796 3151 -8794
rect 3119 -8926 3151 -8924
rect 3119 -8954 3121 -8926
rect 3121 -8954 3149 -8926
rect 3149 -8954 3151 -8926
rect 3119 -8956 3151 -8954
rect 3119 -9086 3151 -9084
rect 3119 -9114 3121 -9086
rect 3121 -9114 3149 -9086
rect 3149 -9114 3151 -9086
rect 3119 -9116 3151 -9114
rect 6852 -5886 6884 -5884
rect 6852 -5914 6854 -5886
rect 6854 -5914 6882 -5886
rect 6882 -5914 6884 -5886
rect 6852 -5916 6884 -5914
rect 6852 -6046 6884 -6044
rect 6852 -6074 6854 -6046
rect 6854 -6074 6882 -6046
rect 6882 -6074 6884 -6046
rect 6852 -6076 6884 -6074
rect 6852 -6206 6884 -6204
rect 6852 -6234 6854 -6206
rect 6854 -6234 6882 -6206
rect 6882 -6234 6884 -6206
rect 6852 -6236 6884 -6234
rect 6852 -6366 6884 -6364
rect 6852 -6394 6854 -6366
rect 6854 -6394 6882 -6366
rect 6882 -6394 6884 -6366
rect 6852 -6396 6884 -6394
rect 6852 -6526 6884 -6524
rect 6852 -6554 6854 -6526
rect 6854 -6554 6882 -6526
rect 6882 -6554 6884 -6526
rect 6852 -6556 6884 -6554
rect 6852 -6686 6884 -6684
rect 6852 -6714 6854 -6686
rect 6854 -6714 6882 -6686
rect 6882 -6714 6884 -6686
rect 6852 -6716 6884 -6714
rect 6852 -6846 6884 -6844
rect 6852 -6874 6854 -6846
rect 6854 -6874 6882 -6846
rect 6882 -6874 6884 -6846
rect 6852 -6876 6884 -6874
rect 6852 -7006 6884 -7004
rect 6852 -7034 6854 -7006
rect 6854 -7034 6882 -7006
rect 6882 -7034 6884 -7006
rect 6852 -7036 6884 -7034
rect 6852 -7166 6884 -7164
rect 6852 -7194 6854 -7166
rect 6854 -7194 6882 -7166
rect 6882 -7194 6884 -7166
rect 6852 -7196 6884 -7194
rect 6852 -7326 6884 -7324
rect 6852 -7354 6854 -7326
rect 6854 -7354 6882 -7326
rect 6882 -7354 6884 -7326
rect 6852 -7356 6884 -7354
rect 6852 -7486 6884 -7484
rect 6852 -7514 6854 -7486
rect 6854 -7514 6882 -7486
rect 6882 -7514 6884 -7486
rect 6852 -7516 6884 -7514
rect 6852 -7646 6884 -7644
rect 6852 -7674 6854 -7646
rect 6854 -7674 6882 -7646
rect 6882 -7674 6884 -7646
rect 6852 -7676 6884 -7674
rect 6852 -7806 6884 -7804
rect 6852 -7834 6854 -7806
rect 6854 -7834 6882 -7806
rect 6882 -7834 6884 -7806
rect 6852 -7836 6884 -7834
rect 6852 -7966 6884 -7964
rect 6852 -7994 6854 -7966
rect 6854 -7994 6882 -7966
rect 6882 -7994 6884 -7966
rect 6852 -7996 6884 -7994
rect 6852 -8126 6884 -8124
rect 6852 -8154 6854 -8126
rect 6854 -8154 6882 -8126
rect 6882 -8154 6884 -8126
rect 6852 -8156 6884 -8154
rect 6852 -8286 6884 -8284
rect 6852 -8314 6854 -8286
rect 6854 -8314 6882 -8286
rect 6882 -8314 6884 -8286
rect 6852 -8316 6884 -8314
rect 6852 -8446 6884 -8444
rect 6852 -8474 6854 -8446
rect 6854 -8474 6882 -8446
rect 6882 -8474 6884 -8446
rect 6852 -8476 6884 -8474
rect 6852 -8606 6884 -8604
rect 6852 -8634 6854 -8606
rect 6854 -8634 6882 -8606
rect 6882 -8634 6884 -8606
rect 6852 -8636 6884 -8634
rect 6852 -8766 6884 -8764
rect 6852 -8794 6854 -8766
rect 6854 -8794 6882 -8766
rect 6882 -8794 6884 -8766
rect 6852 -8796 6884 -8794
rect 6852 -8926 6884 -8924
rect 6852 -8954 6854 -8926
rect 6854 -8954 6882 -8926
rect 6882 -8954 6884 -8926
rect 6852 -8956 6884 -8954
rect 6852 -9086 6884 -9084
rect 6852 -9114 6854 -9086
rect 6854 -9114 6882 -9086
rect 6882 -9114 6884 -9086
rect 6852 -9116 6884 -9114
rect 3119 -9246 3151 -9244
rect 3119 -9274 3121 -9246
rect 3121 -9274 3149 -9246
rect 3149 -9274 3151 -9246
rect 3119 -9276 3151 -9274
rect 6852 -9246 6884 -9244
rect 6852 -9274 6854 -9246
rect 6854 -9274 6882 -9246
rect 6882 -9274 6884 -9246
rect 6852 -9276 6884 -9274
rect 3304 -9351 3336 -9349
rect 3304 -9379 3306 -9351
rect 3306 -9379 3334 -9351
rect 3334 -9379 3336 -9351
rect 3304 -9381 3336 -9379
rect 3464 -9351 3496 -9349
rect 3464 -9379 3466 -9351
rect 3466 -9379 3494 -9351
rect 3494 -9379 3496 -9351
rect 3464 -9381 3496 -9379
rect 3624 -9351 3656 -9349
rect 3624 -9379 3626 -9351
rect 3626 -9379 3654 -9351
rect 3654 -9379 3656 -9351
rect 3624 -9381 3656 -9379
rect 3784 -9351 3816 -9349
rect 3784 -9379 3786 -9351
rect 3786 -9379 3814 -9351
rect 3814 -9379 3816 -9351
rect 3784 -9381 3816 -9379
rect 3944 -9351 3976 -9349
rect 3944 -9379 3946 -9351
rect 3946 -9379 3974 -9351
rect 3974 -9379 3976 -9351
rect 3944 -9381 3976 -9379
rect 4104 -9351 4136 -9349
rect 4104 -9379 4106 -9351
rect 4106 -9379 4134 -9351
rect 4134 -9379 4136 -9351
rect 4104 -9381 4136 -9379
rect 4264 -9351 4296 -9349
rect 4264 -9379 4266 -9351
rect 4266 -9379 4294 -9351
rect 4294 -9379 4296 -9351
rect 4264 -9381 4296 -9379
rect 4424 -9351 4456 -9349
rect 4424 -9379 4426 -9351
rect 4426 -9379 4454 -9351
rect 4454 -9379 4456 -9351
rect 4424 -9381 4456 -9379
rect 4584 -9351 4616 -9349
rect 4584 -9379 4586 -9351
rect 4586 -9379 4614 -9351
rect 4614 -9379 4616 -9351
rect 4584 -9381 4616 -9379
rect 4744 -9351 4776 -9349
rect 4744 -9379 4746 -9351
rect 4746 -9379 4774 -9351
rect 4774 -9379 4776 -9351
rect 4744 -9381 4776 -9379
rect 4904 -9351 4936 -9349
rect 4904 -9379 4906 -9351
rect 4906 -9379 4934 -9351
rect 4934 -9379 4936 -9351
rect 4904 -9381 4936 -9379
rect 5064 -9351 5096 -9349
rect 5064 -9379 5066 -9351
rect 5066 -9379 5094 -9351
rect 5094 -9379 5096 -9351
rect 5064 -9381 5096 -9379
rect 5224 -9351 5256 -9349
rect 5224 -9379 5226 -9351
rect 5226 -9379 5254 -9351
rect 5254 -9379 5256 -9351
rect 5224 -9381 5256 -9379
rect 5384 -9351 5416 -9349
rect 5384 -9379 5386 -9351
rect 5386 -9379 5414 -9351
rect 5414 -9379 5416 -9351
rect 5384 -9381 5416 -9379
rect 5544 -9351 5576 -9349
rect 5544 -9379 5546 -9351
rect 5546 -9379 5574 -9351
rect 5574 -9379 5576 -9351
rect 5544 -9381 5576 -9379
rect 5704 -9351 5736 -9349
rect 5704 -9379 5706 -9351
rect 5706 -9379 5734 -9351
rect 5734 -9379 5736 -9351
rect 5704 -9381 5736 -9379
rect 5864 -9351 5896 -9349
rect 5864 -9379 5866 -9351
rect 5866 -9379 5894 -9351
rect 5894 -9379 5896 -9351
rect 5864 -9381 5896 -9379
rect 6024 -9351 6056 -9349
rect 6024 -9379 6026 -9351
rect 6026 -9379 6054 -9351
rect 6054 -9379 6056 -9351
rect 6024 -9381 6056 -9379
rect 6184 -9351 6216 -9349
rect 6184 -9379 6186 -9351
rect 6186 -9379 6214 -9351
rect 6214 -9379 6216 -9351
rect 6184 -9381 6216 -9379
rect 6344 -9351 6376 -9349
rect 6344 -9379 6346 -9351
rect 6346 -9379 6374 -9351
rect 6374 -9379 6376 -9351
rect 6344 -9381 6376 -9379
rect 6504 -9351 6536 -9349
rect 6504 -9379 6506 -9351
rect 6506 -9379 6534 -9351
rect 6534 -9379 6536 -9351
rect 6504 -9381 6536 -9379
rect 6664 -9351 6696 -9349
rect 6664 -9379 6666 -9351
rect 6666 -9379 6694 -9351
rect 6694 -9379 6696 -9351
rect 6664 -9381 6696 -9379
rect 3304 -11623 3336 -11621
rect 3304 -11651 3306 -11623
rect 3306 -11651 3334 -11623
rect 3334 -11651 3336 -11623
rect 3304 -11653 3336 -11651
rect 3464 -11623 3496 -11621
rect 3464 -11651 3466 -11623
rect 3466 -11651 3494 -11623
rect 3494 -11651 3496 -11623
rect 3464 -11653 3496 -11651
rect 3624 -11623 3656 -11621
rect 3624 -11651 3626 -11623
rect 3626 -11651 3654 -11623
rect 3654 -11651 3656 -11623
rect 3624 -11653 3656 -11651
rect 3784 -11623 3816 -11621
rect 3784 -11651 3786 -11623
rect 3786 -11651 3814 -11623
rect 3814 -11651 3816 -11623
rect 3784 -11653 3816 -11651
rect 3944 -11623 3976 -11621
rect 3944 -11651 3946 -11623
rect 3946 -11651 3974 -11623
rect 3974 -11651 3976 -11623
rect 3944 -11653 3976 -11651
rect 4104 -11623 4136 -11621
rect 4104 -11651 4106 -11623
rect 4106 -11651 4134 -11623
rect 4134 -11651 4136 -11623
rect 4104 -11653 4136 -11651
rect 4264 -11623 4296 -11621
rect 4264 -11651 4266 -11623
rect 4266 -11651 4294 -11623
rect 4294 -11651 4296 -11623
rect 4264 -11653 4296 -11651
rect 4424 -11623 4456 -11621
rect 4424 -11651 4426 -11623
rect 4426 -11651 4454 -11623
rect 4454 -11651 4456 -11623
rect 4424 -11653 4456 -11651
rect 4584 -11623 4616 -11621
rect 4584 -11651 4586 -11623
rect 4586 -11651 4614 -11623
rect 4614 -11651 4616 -11623
rect 4584 -11653 4616 -11651
rect 4744 -11623 4776 -11621
rect 4744 -11651 4746 -11623
rect 4746 -11651 4774 -11623
rect 4774 -11651 4776 -11623
rect 4744 -11653 4776 -11651
rect 4904 -11623 4936 -11621
rect 4904 -11651 4906 -11623
rect 4906 -11651 4934 -11623
rect 4934 -11651 4936 -11623
rect 4904 -11653 4936 -11651
rect 5064 -11623 5096 -11621
rect 5064 -11651 5066 -11623
rect 5066 -11651 5094 -11623
rect 5094 -11651 5096 -11623
rect 5064 -11653 5096 -11651
rect 5224 -11623 5256 -11621
rect 5224 -11651 5226 -11623
rect 5226 -11651 5254 -11623
rect 5254 -11651 5256 -11623
rect 5224 -11653 5256 -11651
rect 5384 -11623 5416 -11621
rect 5384 -11651 5386 -11623
rect 5386 -11651 5414 -11623
rect 5414 -11651 5416 -11623
rect 5384 -11653 5416 -11651
rect 5544 -11623 5576 -11621
rect 5544 -11651 5546 -11623
rect 5546 -11651 5574 -11623
rect 5574 -11651 5576 -11623
rect 5544 -11653 5576 -11651
rect 5704 -11623 5736 -11621
rect 5704 -11651 5706 -11623
rect 5706 -11651 5734 -11623
rect 5734 -11651 5736 -11623
rect 5704 -11653 5736 -11651
rect 5864 -11623 5896 -11621
rect 5864 -11651 5866 -11623
rect 5866 -11651 5894 -11623
rect 5894 -11651 5896 -11623
rect 5864 -11653 5896 -11651
rect 6024 -11623 6056 -11621
rect 6024 -11651 6026 -11623
rect 6026 -11651 6054 -11623
rect 6054 -11651 6056 -11623
rect 6024 -11653 6056 -11651
rect 6184 -11623 6216 -11621
rect 6184 -11651 6186 -11623
rect 6186 -11651 6214 -11623
rect 6214 -11651 6216 -11623
rect 6184 -11653 6216 -11651
rect 6344 -11623 6376 -11621
rect 6344 -11651 6346 -11623
rect 6346 -11651 6374 -11623
rect 6374 -11651 6376 -11623
rect 6344 -11653 6376 -11651
rect 6504 -11623 6536 -11621
rect 6504 -11651 6506 -11623
rect 6506 -11651 6534 -11623
rect 6534 -11651 6536 -11623
rect 6504 -11653 6536 -11651
rect 6664 -11623 6696 -11621
rect 6664 -11651 6666 -11623
rect 6666 -11651 6694 -11623
rect 6694 -11651 6696 -11623
rect 6664 -11653 6696 -11651
rect 3119 -11726 3151 -11724
rect 3119 -11754 3121 -11726
rect 3121 -11754 3149 -11726
rect 3149 -11754 3151 -11726
rect 3119 -11756 3151 -11754
rect 6852 -11726 6884 -11724
rect 6852 -11754 6854 -11726
rect 6854 -11754 6882 -11726
rect 6882 -11754 6884 -11726
rect 6852 -11756 6884 -11754
rect 3119 -11886 3151 -11884
rect 3119 -11914 3121 -11886
rect 3121 -11914 3149 -11886
rect 3149 -11914 3151 -11886
rect 3119 -11916 3151 -11914
rect 3119 -12046 3151 -12044
rect 3119 -12074 3121 -12046
rect 3121 -12074 3149 -12046
rect 3149 -12074 3151 -12046
rect 3119 -12076 3151 -12074
rect 3119 -12206 3151 -12204
rect 3119 -12234 3121 -12206
rect 3121 -12234 3149 -12206
rect 3149 -12234 3151 -12206
rect 3119 -12236 3151 -12234
rect 3119 -12366 3151 -12364
rect 3119 -12394 3121 -12366
rect 3121 -12394 3149 -12366
rect 3149 -12394 3151 -12366
rect 3119 -12396 3151 -12394
rect 3119 -12526 3151 -12524
rect 3119 -12554 3121 -12526
rect 3121 -12554 3149 -12526
rect 3149 -12554 3151 -12526
rect 3119 -12556 3151 -12554
rect 3119 -12686 3151 -12684
rect 3119 -12714 3121 -12686
rect 3121 -12714 3149 -12686
rect 3149 -12714 3151 -12686
rect 3119 -12716 3151 -12714
rect 3119 -12846 3151 -12844
rect 3119 -12874 3121 -12846
rect 3121 -12874 3149 -12846
rect 3149 -12874 3151 -12846
rect 3119 -12876 3151 -12874
rect 3119 -13006 3151 -13004
rect 3119 -13034 3121 -13006
rect 3121 -13034 3149 -13006
rect 3149 -13034 3151 -13006
rect 3119 -13036 3151 -13034
rect 3119 -13166 3151 -13164
rect 3119 -13194 3121 -13166
rect 3121 -13194 3149 -13166
rect 3149 -13194 3151 -13166
rect 3119 -13196 3151 -13194
rect 3119 -13326 3151 -13324
rect 3119 -13354 3121 -13326
rect 3121 -13354 3149 -13326
rect 3149 -13354 3151 -13326
rect 3119 -13356 3151 -13354
rect 3119 -13486 3151 -13484
rect 3119 -13514 3121 -13486
rect 3121 -13514 3149 -13486
rect 3149 -13514 3151 -13486
rect 3119 -13516 3151 -13514
rect 3119 -13646 3151 -13644
rect 3119 -13674 3121 -13646
rect 3121 -13674 3149 -13646
rect 3149 -13674 3151 -13646
rect 3119 -13676 3151 -13674
rect 3119 -13806 3151 -13804
rect 3119 -13834 3121 -13806
rect 3121 -13834 3149 -13806
rect 3149 -13834 3151 -13806
rect 3119 -13836 3151 -13834
rect 3119 -13966 3151 -13964
rect 3119 -13994 3121 -13966
rect 3121 -13994 3149 -13966
rect 3149 -13994 3151 -13966
rect 3119 -13996 3151 -13994
rect 3119 -14126 3151 -14124
rect 3119 -14154 3121 -14126
rect 3121 -14154 3149 -14126
rect 3149 -14154 3151 -14126
rect 3119 -14156 3151 -14154
rect 3119 -14286 3151 -14284
rect 3119 -14314 3121 -14286
rect 3121 -14314 3149 -14286
rect 3149 -14314 3151 -14286
rect 3119 -14316 3151 -14314
rect 3119 -14446 3151 -14444
rect 3119 -14474 3121 -14446
rect 3121 -14474 3149 -14446
rect 3149 -14474 3151 -14446
rect 3119 -14476 3151 -14474
rect 3119 -14606 3151 -14604
rect 3119 -14634 3121 -14606
rect 3121 -14634 3149 -14606
rect 3149 -14634 3151 -14606
rect 3119 -14636 3151 -14634
rect 3119 -14766 3151 -14764
rect 3119 -14794 3121 -14766
rect 3121 -14794 3149 -14766
rect 3149 -14794 3151 -14766
rect 3119 -14796 3151 -14794
rect 3119 -14926 3151 -14924
rect 3119 -14954 3121 -14926
rect 3121 -14954 3149 -14926
rect 3149 -14954 3151 -14926
rect 3119 -14956 3151 -14954
rect 3119 -15086 3151 -15084
rect 3119 -15114 3121 -15086
rect 3121 -15114 3149 -15086
rect 3149 -15114 3151 -15086
rect 3119 -15116 3151 -15114
rect 6852 -11886 6884 -11884
rect 6852 -11914 6854 -11886
rect 6854 -11914 6882 -11886
rect 6882 -11914 6884 -11886
rect 6852 -11916 6884 -11914
rect 6852 -12046 6884 -12044
rect 6852 -12074 6854 -12046
rect 6854 -12074 6882 -12046
rect 6882 -12074 6884 -12046
rect 6852 -12076 6884 -12074
rect 6852 -12206 6884 -12204
rect 6852 -12234 6854 -12206
rect 6854 -12234 6882 -12206
rect 6882 -12234 6884 -12206
rect 6852 -12236 6884 -12234
rect 6852 -12366 6884 -12364
rect 6852 -12394 6854 -12366
rect 6854 -12394 6882 -12366
rect 6882 -12394 6884 -12366
rect 6852 -12396 6884 -12394
rect 6852 -12526 6884 -12524
rect 6852 -12554 6854 -12526
rect 6854 -12554 6882 -12526
rect 6882 -12554 6884 -12526
rect 6852 -12556 6884 -12554
rect 6852 -12686 6884 -12684
rect 6852 -12714 6854 -12686
rect 6854 -12714 6882 -12686
rect 6882 -12714 6884 -12686
rect 6852 -12716 6884 -12714
rect 6852 -12846 6884 -12844
rect 6852 -12874 6854 -12846
rect 6854 -12874 6882 -12846
rect 6882 -12874 6884 -12846
rect 6852 -12876 6884 -12874
rect 9304 -5623 9336 -5621
rect 9304 -5651 9306 -5623
rect 9306 -5651 9334 -5623
rect 9334 -5651 9336 -5623
rect 9304 -5653 9336 -5651
rect 9464 -5623 9496 -5621
rect 9464 -5651 9466 -5623
rect 9466 -5651 9494 -5623
rect 9494 -5651 9496 -5623
rect 9464 -5653 9496 -5651
rect 9624 -5623 9656 -5621
rect 9624 -5651 9626 -5623
rect 9626 -5651 9654 -5623
rect 9654 -5651 9656 -5623
rect 9624 -5653 9656 -5651
rect 9784 -5623 9816 -5621
rect 9784 -5651 9786 -5623
rect 9786 -5651 9814 -5623
rect 9814 -5651 9816 -5623
rect 9784 -5653 9816 -5651
rect 9944 -5623 9976 -5621
rect 9944 -5651 9946 -5623
rect 9946 -5651 9974 -5623
rect 9974 -5651 9976 -5623
rect 9944 -5653 9976 -5651
rect 10104 -5623 10136 -5621
rect 10104 -5651 10106 -5623
rect 10106 -5651 10134 -5623
rect 10134 -5651 10136 -5623
rect 10104 -5653 10136 -5651
rect 10264 -5623 10296 -5621
rect 10264 -5651 10266 -5623
rect 10266 -5651 10294 -5623
rect 10294 -5651 10296 -5623
rect 10264 -5653 10296 -5651
rect 10424 -5623 10456 -5621
rect 10424 -5651 10426 -5623
rect 10426 -5651 10454 -5623
rect 10454 -5651 10456 -5623
rect 10424 -5653 10456 -5651
rect 10584 -5623 10616 -5621
rect 10584 -5651 10586 -5623
rect 10586 -5651 10614 -5623
rect 10614 -5651 10616 -5623
rect 10584 -5653 10616 -5651
rect 10744 -5623 10776 -5621
rect 10744 -5651 10746 -5623
rect 10746 -5651 10774 -5623
rect 10774 -5651 10776 -5623
rect 10744 -5653 10776 -5651
rect 10904 -5623 10936 -5621
rect 10904 -5651 10906 -5623
rect 10906 -5651 10934 -5623
rect 10934 -5651 10936 -5623
rect 10904 -5653 10936 -5651
rect 11064 -5623 11096 -5621
rect 11064 -5651 11066 -5623
rect 11066 -5651 11094 -5623
rect 11094 -5651 11096 -5623
rect 11064 -5653 11096 -5651
rect 11224 -5623 11256 -5621
rect 11224 -5651 11226 -5623
rect 11226 -5651 11254 -5623
rect 11254 -5651 11256 -5623
rect 11224 -5653 11256 -5651
rect 11384 -5623 11416 -5621
rect 11384 -5651 11386 -5623
rect 11386 -5651 11414 -5623
rect 11414 -5651 11416 -5623
rect 11384 -5653 11416 -5651
rect 11544 -5623 11576 -5621
rect 11544 -5651 11546 -5623
rect 11546 -5651 11574 -5623
rect 11574 -5651 11576 -5623
rect 11544 -5653 11576 -5651
rect 11704 -5623 11736 -5621
rect 11704 -5651 11706 -5623
rect 11706 -5651 11734 -5623
rect 11734 -5651 11736 -5623
rect 11704 -5653 11736 -5651
rect 11864 -5623 11896 -5621
rect 11864 -5651 11866 -5623
rect 11866 -5651 11894 -5623
rect 11894 -5651 11896 -5623
rect 11864 -5653 11896 -5651
rect 12024 -5623 12056 -5621
rect 12024 -5651 12026 -5623
rect 12026 -5651 12054 -5623
rect 12054 -5651 12056 -5623
rect 12024 -5653 12056 -5651
rect 12184 -5623 12216 -5621
rect 12184 -5651 12186 -5623
rect 12186 -5651 12214 -5623
rect 12214 -5651 12216 -5623
rect 12184 -5653 12216 -5651
rect 12344 -5623 12376 -5621
rect 12344 -5651 12346 -5623
rect 12346 -5651 12374 -5623
rect 12374 -5651 12376 -5623
rect 12344 -5653 12376 -5651
rect 12504 -5623 12536 -5621
rect 12504 -5651 12506 -5623
rect 12506 -5651 12534 -5623
rect 12534 -5651 12536 -5623
rect 12504 -5653 12536 -5651
rect 12664 -5623 12696 -5621
rect 12664 -5651 12666 -5623
rect 12666 -5651 12694 -5623
rect 12694 -5651 12696 -5623
rect 12664 -5653 12696 -5651
rect 9119 -5726 9151 -5724
rect 9119 -5754 9121 -5726
rect 9121 -5754 9149 -5726
rect 9149 -5754 9151 -5726
rect 9119 -5756 9151 -5754
rect 12852 -5726 12884 -5724
rect 12852 -5754 12854 -5726
rect 12854 -5754 12882 -5726
rect 12882 -5754 12884 -5726
rect 12852 -5756 12884 -5754
rect 9119 -5886 9151 -5884
rect 9119 -5914 9121 -5886
rect 9121 -5914 9149 -5886
rect 9149 -5914 9151 -5886
rect 9119 -5916 9151 -5914
rect 9119 -6046 9151 -6044
rect 9119 -6074 9121 -6046
rect 9121 -6074 9149 -6046
rect 9149 -6074 9151 -6046
rect 9119 -6076 9151 -6074
rect 9119 -6206 9151 -6204
rect 9119 -6234 9121 -6206
rect 9121 -6234 9149 -6206
rect 9149 -6234 9151 -6206
rect 9119 -6236 9151 -6234
rect 9119 -6366 9151 -6364
rect 9119 -6394 9121 -6366
rect 9121 -6394 9149 -6366
rect 9149 -6394 9151 -6366
rect 9119 -6396 9151 -6394
rect 9119 -6526 9151 -6524
rect 9119 -6554 9121 -6526
rect 9121 -6554 9149 -6526
rect 9149 -6554 9151 -6526
rect 9119 -6556 9151 -6554
rect 9119 -6686 9151 -6684
rect 9119 -6714 9121 -6686
rect 9121 -6714 9149 -6686
rect 9149 -6714 9151 -6686
rect 9119 -6716 9151 -6714
rect 9119 -6846 9151 -6844
rect 9119 -6874 9121 -6846
rect 9121 -6874 9149 -6846
rect 9149 -6874 9151 -6846
rect 9119 -6876 9151 -6874
rect 9119 -7006 9151 -7004
rect 9119 -7034 9121 -7006
rect 9121 -7034 9149 -7006
rect 9149 -7034 9151 -7006
rect 9119 -7036 9151 -7034
rect 9119 -7166 9151 -7164
rect 9119 -7194 9121 -7166
rect 9121 -7194 9149 -7166
rect 9149 -7194 9151 -7166
rect 9119 -7196 9151 -7194
rect 9119 -7326 9151 -7324
rect 9119 -7354 9121 -7326
rect 9121 -7354 9149 -7326
rect 9149 -7354 9151 -7326
rect 9119 -7356 9151 -7354
rect 9119 -7486 9151 -7484
rect 9119 -7514 9121 -7486
rect 9121 -7514 9149 -7486
rect 9149 -7514 9151 -7486
rect 9119 -7516 9151 -7514
rect 9119 -7646 9151 -7644
rect 9119 -7674 9121 -7646
rect 9121 -7674 9149 -7646
rect 9149 -7674 9151 -7646
rect 9119 -7676 9151 -7674
rect 9119 -7806 9151 -7804
rect 9119 -7834 9121 -7806
rect 9121 -7834 9149 -7806
rect 9149 -7834 9151 -7806
rect 9119 -7836 9151 -7834
rect 9119 -7966 9151 -7964
rect 9119 -7994 9121 -7966
rect 9121 -7994 9149 -7966
rect 9149 -7994 9151 -7966
rect 9119 -7996 9151 -7994
rect 9119 -8126 9151 -8124
rect 9119 -8154 9121 -8126
rect 9121 -8154 9149 -8126
rect 9149 -8154 9151 -8126
rect 9119 -8156 9151 -8154
rect 9119 -8286 9151 -8284
rect 9119 -8314 9121 -8286
rect 9121 -8314 9149 -8286
rect 9149 -8314 9151 -8286
rect 9119 -8316 9151 -8314
rect 9119 -8446 9151 -8444
rect 9119 -8474 9121 -8446
rect 9121 -8474 9149 -8446
rect 9149 -8474 9151 -8446
rect 9119 -8476 9151 -8474
rect 9119 -8606 9151 -8604
rect 9119 -8634 9121 -8606
rect 9121 -8634 9149 -8606
rect 9149 -8634 9151 -8606
rect 9119 -8636 9151 -8634
rect 9119 -8766 9151 -8764
rect 9119 -8794 9121 -8766
rect 9121 -8794 9149 -8766
rect 9149 -8794 9151 -8766
rect 9119 -8796 9151 -8794
rect 9119 -8926 9151 -8924
rect 9119 -8954 9121 -8926
rect 9121 -8954 9149 -8926
rect 9149 -8954 9151 -8926
rect 9119 -8956 9151 -8954
rect 9119 -9086 9151 -9084
rect 9119 -9114 9121 -9086
rect 9121 -9114 9149 -9086
rect 9149 -9114 9151 -9086
rect 9119 -9116 9151 -9114
rect 12852 -5886 12884 -5884
rect 12852 -5914 12854 -5886
rect 12854 -5914 12882 -5886
rect 12882 -5914 12884 -5886
rect 12852 -5916 12884 -5914
rect 12852 -6046 12884 -6044
rect 12852 -6074 12854 -6046
rect 12854 -6074 12882 -6046
rect 12882 -6074 12884 -6046
rect 12852 -6076 12884 -6074
rect 12852 -6206 12884 -6204
rect 12852 -6234 12854 -6206
rect 12854 -6234 12882 -6206
rect 12882 -6234 12884 -6206
rect 12852 -6236 12884 -6234
rect 12852 -6366 12884 -6364
rect 12852 -6394 12854 -6366
rect 12854 -6394 12882 -6366
rect 12882 -6394 12884 -6366
rect 12852 -6396 12884 -6394
rect 12852 -6526 12884 -6524
rect 12852 -6554 12854 -6526
rect 12854 -6554 12882 -6526
rect 12882 -6554 12884 -6526
rect 12852 -6556 12884 -6554
rect 12852 -6686 12884 -6684
rect 12852 -6714 12854 -6686
rect 12854 -6714 12882 -6686
rect 12882 -6714 12884 -6686
rect 12852 -6716 12884 -6714
rect 12852 -6846 12884 -6844
rect 12852 -6874 12854 -6846
rect 12854 -6874 12882 -6846
rect 12882 -6874 12884 -6846
rect 12852 -6876 12884 -6874
rect 12852 -7006 12884 -7004
rect 12852 -7034 12854 -7006
rect 12854 -7034 12882 -7006
rect 12882 -7034 12884 -7006
rect 12852 -7036 12884 -7034
rect 12852 -7166 12884 -7164
rect 12852 -7194 12854 -7166
rect 12854 -7194 12882 -7166
rect 12882 -7194 12884 -7166
rect 12852 -7196 12884 -7194
rect 12852 -7326 12884 -7324
rect 12852 -7354 12854 -7326
rect 12854 -7354 12882 -7326
rect 12882 -7354 12884 -7326
rect 12852 -7356 12884 -7354
rect 12852 -7486 12884 -7484
rect 12852 -7514 12854 -7486
rect 12854 -7514 12882 -7486
rect 12882 -7514 12884 -7486
rect 12852 -7516 12884 -7514
rect 12852 -7646 12884 -7644
rect 12852 -7674 12854 -7646
rect 12854 -7674 12882 -7646
rect 12882 -7674 12884 -7646
rect 12852 -7676 12884 -7674
rect 12852 -7806 12884 -7804
rect 12852 -7834 12854 -7806
rect 12854 -7834 12882 -7806
rect 12882 -7834 12884 -7806
rect 12852 -7836 12884 -7834
rect 15304 -5623 15336 -5621
rect 15304 -5651 15306 -5623
rect 15306 -5651 15334 -5623
rect 15334 -5651 15336 -5623
rect 15304 -5653 15336 -5651
rect 15464 -5623 15496 -5621
rect 15464 -5651 15466 -5623
rect 15466 -5651 15494 -5623
rect 15494 -5651 15496 -5623
rect 15464 -5653 15496 -5651
rect 15624 -5623 15656 -5621
rect 15624 -5651 15626 -5623
rect 15626 -5651 15654 -5623
rect 15654 -5651 15656 -5623
rect 15624 -5653 15656 -5651
rect 15784 -5623 15816 -5621
rect 15784 -5651 15786 -5623
rect 15786 -5651 15814 -5623
rect 15814 -5651 15816 -5623
rect 15784 -5653 15816 -5651
rect 15944 -5623 15976 -5621
rect 15944 -5651 15946 -5623
rect 15946 -5651 15974 -5623
rect 15974 -5651 15976 -5623
rect 15944 -5653 15976 -5651
rect 16104 -5623 16136 -5621
rect 16104 -5651 16106 -5623
rect 16106 -5651 16134 -5623
rect 16134 -5651 16136 -5623
rect 16104 -5653 16136 -5651
rect 16264 -5623 16296 -5621
rect 16264 -5651 16266 -5623
rect 16266 -5651 16294 -5623
rect 16294 -5651 16296 -5623
rect 16264 -5653 16296 -5651
rect 16424 -5623 16456 -5621
rect 16424 -5651 16426 -5623
rect 16426 -5651 16454 -5623
rect 16454 -5651 16456 -5623
rect 16424 -5653 16456 -5651
rect 16584 -5623 16616 -5621
rect 16584 -5651 16586 -5623
rect 16586 -5651 16614 -5623
rect 16614 -5651 16616 -5623
rect 16584 -5653 16616 -5651
rect 16744 -5623 16776 -5621
rect 16744 -5651 16746 -5623
rect 16746 -5651 16774 -5623
rect 16774 -5651 16776 -5623
rect 16744 -5653 16776 -5651
rect 16904 -5623 16936 -5621
rect 16904 -5651 16906 -5623
rect 16906 -5651 16934 -5623
rect 16934 -5651 16936 -5623
rect 16904 -5653 16936 -5651
rect 17064 -5623 17096 -5621
rect 17064 -5651 17066 -5623
rect 17066 -5651 17094 -5623
rect 17094 -5651 17096 -5623
rect 17064 -5653 17096 -5651
rect 17224 -5623 17256 -5621
rect 17224 -5651 17226 -5623
rect 17226 -5651 17254 -5623
rect 17254 -5651 17256 -5623
rect 17224 -5653 17256 -5651
rect 17384 -5623 17416 -5621
rect 17384 -5651 17386 -5623
rect 17386 -5651 17414 -5623
rect 17414 -5651 17416 -5623
rect 17384 -5653 17416 -5651
rect 17544 -5623 17576 -5621
rect 17544 -5651 17546 -5623
rect 17546 -5651 17574 -5623
rect 17574 -5651 17576 -5623
rect 17544 -5653 17576 -5651
rect 17704 -5623 17736 -5621
rect 17704 -5651 17706 -5623
rect 17706 -5651 17734 -5623
rect 17734 -5651 17736 -5623
rect 17704 -5653 17736 -5651
rect 17864 -5623 17896 -5621
rect 17864 -5651 17866 -5623
rect 17866 -5651 17894 -5623
rect 17894 -5651 17896 -5623
rect 17864 -5653 17896 -5651
rect 18024 -5623 18056 -5621
rect 18024 -5651 18026 -5623
rect 18026 -5651 18054 -5623
rect 18054 -5651 18056 -5623
rect 18024 -5653 18056 -5651
rect 18184 -5623 18216 -5621
rect 18184 -5651 18186 -5623
rect 18186 -5651 18214 -5623
rect 18214 -5651 18216 -5623
rect 18184 -5653 18216 -5651
rect 18344 -5623 18376 -5621
rect 18344 -5651 18346 -5623
rect 18346 -5651 18374 -5623
rect 18374 -5651 18376 -5623
rect 18344 -5653 18376 -5651
rect 18504 -5623 18536 -5621
rect 18504 -5651 18506 -5623
rect 18506 -5651 18534 -5623
rect 18534 -5651 18536 -5623
rect 18504 -5653 18536 -5651
rect 18664 -5623 18696 -5621
rect 18664 -5651 18666 -5623
rect 18666 -5651 18694 -5623
rect 18694 -5651 18696 -5623
rect 18664 -5653 18696 -5651
rect 15119 -5726 15151 -5724
rect 15119 -5754 15121 -5726
rect 15121 -5754 15149 -5726
rect 15149 -5754 15151 -5726
rect 15119 -5756 15151 -5754
rect 18852 -5726 18884 -5724
rect 18852 -5754 18854 -5726
rect 18854 -5754 18882 -5726
rect 18882 -5754 18884 -5726
rect 18852 -5756 18884 -5754
rect 15119 -5886 15151 -5884
rect 15119 -5914 15121 -5886
rect 15121 -5914 15149 -5886
rect 15149 -5914 15151 -5886
rect 15119 -5916 15151 -5914
rect 15119 -6046 15151 -6044
rect 15119 -6074 15121 -6046
rect 15121 -6074 15149 -6046
rect 15149 -6074 15151 -6046
rect 15119 -6076 15151 -6074
rect 15119 -6206 15151 -6204
rect 15119 -6234 15121 -6206
rect 15121 -6234 15149 -6206
rect 15149 -6234 15151 -6206
rect 15119 -6236 15151 -6234
rect 15119 -6366 15151 -6364
rect 15119 -6394 15121 -6366
rect 15121 -6394 15149 -6366
rect 15149 -6394 15151 -6366
rect 15119 -6396 15151 -6394
rect 15119 -6526 15151 -6524
rect 15119 -6554 15121 -6526
rect 15121 -6554 15149 -6526
rect 15149 -6554 15151 -6526
rect 15119 -6556 15151 -6554
rect 15119 -6686 15151 -6684
rect 15119 -6714 15121 -6686
rect 15121 -6714 15149 -6686
rect 15149 -6714 15151 -6686
rect 15119 -6716 15151 -6714
rect 15119 -6846 15151 -6844
rect 15119 -6874 15121 -6846
rect 15121 -6874 15149 -6846
rect 15149 -6874 15151 -6846
rect 15119 -6876 15151 -6874
rect 15119 -7006 15151 -7004
rect 15119 -7034 15121 -7006
rect 15121 -7034 15149 -7006
rect 15149 -7034 15151 -7006
rect 15119 -7036 15151 -7034
rect 15119 -7166 15151 -7164
rect 15119 -7194 15121 -7166
rect 15121 -7194 15149 -7166
rect 15149 -7194 15151 -7166
rect 15119 -7196 15151 -7194
rect 15119 -7326 15151 -7324
rect 15119 -7354 15121 -7326
rect 15121 -7354 15149 -7326
rect 15149 -7354 15151 -7326
rect 15119 -7356 15151 -7354
rect 15119 -7486 15151 -7484
rect 15119 -7514 15121 -7486
rect 15121 -7514 15149 -7486
rect 15149 -7514 15151 -7486
rect 15119 -7516 15151 -7514
rect 15119 -7646 15151 -7644
rect 15119 -7674 15121 -7646
rect 15121 -7674 15149 -7646
rect 15149 -7674 15151 -7646
rect 15119 -7676 15151 -7674
rect 12852 -7966 12884 -7964
rect 12852 -7994 12854 -7966
rect 12854 -7994 12882 -7966
rect 12882 -7994 12884 -7966
rect 12852 -7996 12884 -7994
rect 12852 -8126 12884 -8124
rect 12852 -8154 12854 -8126
rect 12854 -8154 12882 -8126
rect 12882 -8154 12884 -8126
rect 12852 -8156 12884 -8154
rect 12852 -8286 12884 -8284
rect 12852 -8314 12854 -8286
rect 12854 -8314 12882 -8286
rect 12882 -8314 12884 -8286
rect 12852 -8316 12884 -8314
rect 12852 -8446 12884 -8444
rect 12852 -8474 12854 -8446
rect 12854 -8474 12882 -8446
rect 12882 -8474 12884 -8446
rect 12852 -8476 12884 -8474
rect 12852 -8606 12884 -8604
rect 12852 -8634 12854 -8606
rect 12854 -8634 12882 -8606
rect 12882 -8634 12884 -8606
rect 12852 -8636 12884 -8634
rect 12852 -8766 12884 -8764
rect 12852 -8794 12854 -8766
rect 12854 -8794 12882 -8766
rect 12882 -8794 12884 -8766
rect 12852 -8796 12884 -8794
rect 12852 -8926 12884 -8924
rect 12852 -8954 12854 -8926
rect 12854 -8954 12882 -8926
rect 12882 -8954 12884 -8926
rect 12852 -8956 12884 -8954
rect 12852 -9086 12884 -9084
rect 12852 -9114 12854 -9086
rect 12854 -9114 12882 -9086
rect 12882 -9114 12884 -9086
rect 12852 -9116 12884 -9114
rect 9119 -9246 9151 -9244
rect 9119 -9274 9121 -9246
rect 9121 -9274 9149 -9246
rect 9149 -9274 9151 -9246
rect 9119 -9276 9151 -9274
rect 12852 -9246 12884 -9244
rect 12852 -9274 12854 -9246
rect 12854 -9274 12882 -9246
rect 12882 -9274 12884 -9246
rect 12852 -9276 12884 -9274
rect 9304 -9351 9336 -9349
rect 9304 -9379 9306 -9351
rect 9306 -9379 9334 -9351
rect 9334 -9379 9336 -9351
rect 9304 -9381 9336 -9379
rect 9464 -9351 9496 -9349
rect 9464 -9379 9466 -9351
rect 9466 -9379 9494 -9351
rect 9494 -9379 9496 -9351
rect 9464 -9381 9496 -9379
rect 9624 -9351 9656 -9349
rect 9624 -9379 9626 -9351
rect 9626 -9379 9654 -9351
rect 9654 -9379 9656 -9351
rect 9624 -9381 9656 -9379
rect 9784 -9351 9816 -9349
rect 9784 -9379 9786 -9351
rect 9786 -9379 9814 -9351
rect 9814 -9379 9816 -9351
rect 9784 -9381 9816 -9379
rect 9944 -9351 9976 -9349
rect 9944 -9379 9946 -9351
rect 9946 -9379 9974 -9351
rect 9974 -9379 9976 -9351
rect 9944 -9381 9976 -9379
rect 10104 -9351 10136 -9349
rect 10104 -9379 10106 -9351
rect 10106 -9379 10134 -9351
rect 10134 -9379 10136 -9351
rect 10104 -9381 10136 -9379
rect 10264 -9351 10296 -9349
rect 10264 -9379 10266 -9351
rect 10266 -9379 10294 -9351
rect 10294 -9379 10296 -9351
rect 10264 -9381 10296 -9379
rect 10424 -9351 10456 -9349
rect 10424 -9379 10426 -9351
rect 10426 -9379 10454 -9351
rect 10454 -9379 10456 -9351
rect 10424 -9381 10456 -9379
rect 10584 -9351 10616 -9349
rect 10584 -9379 10586 -9351
rect 10586 -9379 10614 -9351
rect 10614 -9379 10616 -9351
rect 10584 -9381 10616 -9379
rect 10744 -9351 10776 -9349
rect 10744 -9379 10746 -9351
rect 10746 -9379 10774 -9351
rect 10774 -9379 10776 -9351
rect 10744 -9381 10776 -9379
rect 10904 -9351 10936 -9349
rect 10904 -9379 10906 -9351
rect 10906 -9379 10934 -9351
rect 10934 -9379 10936 -9351
rect 10904 -9381 10936 -9379
rect 11064 -9351 11096 -9349
rect 11064 -9379 11066 -9351
rect 11066 -9379 11094 -9351
rect 11094 -9379 11096 -9351
rect 11064 -9381 11096 -9379
rect 11224 -9351 11256 -9349
rect 11224 -9379 11226 -9351
rect 11226 -9379 11254 -9351
rect 11254 -9379 11256 -9351
rect 11224 -9381 11256 -9379
rect 11384 -9351 11416 -9349
rect 11384 -9379 11386 -9351
rect 11386 -9379 11414 -9351
rect 11414 -9379 11416 -9351
rect 11384 -9381 11416 -9379
rect 11544 -9351 11576 -9349
rect 11544 -9379 11546 -9351
rect 11546 -9379 11574 -9351
rect 11574 -9379 11576 -9351
rect 11544 -9381 11576 -9379
rect 11704 -9351 11736 -9349
rect 11704 -9379 11706 -9351
rect 11706 -9379 11734 -9351
rect 11734 -9379 11736 -9351
rect 11704 -9381 11736 -9379
rect 11864 -9351 11896 -9349
rect 11864 -9379 11866 -9351
rect 11866 -9379 11894 -9351
rect 11894 -9379 11896 -9351
rect 11864 -9381 11896 -9379
rect 12024 -9351 12056 -9349
rect 12024 -9379 12026 -9351
rect 12026 -9379 12054 -9351
rect 12054 -9379 12056 -9351
rect 12024 -9381 12056 -9379
rect 12184 -9351 12216 -9349
rect 12184 -9379 12186 -9351
rect 12186 -9379 12214 -9351
rect 12214 -9379 12216 -9351
rect 12184 -9381 12216 -9379
rect 12344 -9351 12376 -9349
rect 12344 -9379 12346 -9351
rect 12346 -9379 12374 -9351
rect 12374 -9379 12376 -9351
rect 12344 -9381 12376 -9379
rect 12504 -9351 12536 -9349
rect 12504 -9379 12506 -9351
rect 12506 -9379 12534 -9351
rect 12534 -9379 12536 -9351
rect 12504 -9381 12536 -9379
rect 12664 -9351 12696 -9349
rect 12664 -9379 12666 -9351
rect 12666 -9379 12694 -9351
rect 12694 -9379 12696 -9351
rect 12664 -9381 12696 -9379
rect 15119 -7806 15151 -7804
rect 15119 -7834 15121 -7806
rect 15121 -7834 15149 -7806
rect 15149 -7834 15151 -7806
rect 15119 -7836 15151 -7834
rect 15119 -7966 15151 -7964
rect 15119 -7994 15121 -7966
rect 15121 -7994 15149 -7966
rect 15149 -7994 15151 -7966
rect 15119 -7996 15151 -7994
rect 15119 -8126 15151 -8124
rect 15119 -8154 15121 -8126
rect 15121 -8154 15149 -8126
rect 15149 -8154 15151 -8126
rect 15119 -8156 15151 -8154
rect 15119 -8286 15151 -8284
rect 15119 -8314 15121 -8286
rect 15121 -8314 15149 -8286
rect 15149 -8314 15151 -8286
rect 15119 -8316 15151 -8314
rect 15119 -8446 15151 -8444
rect 15119 -8474 15121 -8446
rect 15121 -8474 15149 -8446
rect 15149 -8474 15151 -8446
rect 15119 -8476 15151 -8474
rect 15119 -8606 15151 -8604
rect 15119 -8634 15121 -8606
rect 15121 -8634 15149 -8606
rect 15149 -8634 15151 -8606
rect 15119 -8636 15151 -8634
rect 15119 -8766 15151 -8764
rect 15119 -8794 15121 -8766
rect 15121 -8794 15149 -8766
rect 15149 -8794 15151 -8766
rect 15119 -8796 15151 -8794
rect 15119 -8926 15151 -8924
rect 15119 -8954 15121 -8926
rect 15121 -8954 15149 -8926
rect 15149 -8954 15151 -8926
rect 15119 -8956 15151 -8954
rect 15119 -9086 15151 -9084
rect 15119 -9114 15121 -9086
rect 15121 -9114 15149 -9086
rect 15149 -9114 15151 -9086
rect 15119 -9116 15151 -9114
rect 18852 -5886 18884 -5884
rect 18852 -5914 18854 -5886
rect 18854 -5914 18882 -5886
rect 18882 -5914 18884 -5886
rect 18852 -5916 18884 -5914
rect 18852 -6046 18884 -6044
rect 18852 -6074 18854 -6046
rect 18854 -6074 18882 -6046
rect 18882 -6074 18884 -6046
rect 18852 -6076 18884 -6074
rect 18852 -6206 18884 -6204
rect 18852 -6234 18854 -6206
rect 18854 -6234 18882 -6206
rect 18882 -6234 18884 -6206
rect 18852 -6236 18884 -6234
rect 18852 -6366 18884 -6364
rect 18852 -6394 18854 -6366
rect 18854 -6394 18882 -6366
rect 18882 -6394 18884 -6366
rect 18852 -6396 18884 -6394
rect 18852 -6526 18884 -6524
rect 18852 -6554 18854 -6526
rect 18854 -6554 18882 -6526
rect 18882 -6554 18884 -6526
rect 18852 -6556 18884 -6554
rect 18852 -6686 18884 -6684
rect 18852 -6714 18854 -6686
rect 18854 -6714 18882 -6686
rect 18882 -6714 18884 -6686
rect 18852 -6716 18884 -6714
rect 18852 -6846 18884 -6844
rect 18852 -6874 18854 -6846
rect 18854 -6874 18882 -6846
rect 18882 -6874 18884 -6846
rect 18852 -6876 18884 -6874
rect 18852 -7006 18884 -7004
rect 18852 -7034 18854 -7006
rect 18854 -7034 18882 -7006
rect 18882 -7034 18884 -7006
rect 18852 -7036 18884 -7034
rect 18852 -7166 18884 -7164
rect 18852 -7194 18854 -7166
rect 18854 -7194 18882 -7166
rect 18882 -7194 18884 -7166
rect 18852 -7196 18884 -7194
rect 18852 -7326 18884 -7324
rect 18852 -7354 18854 -7326
rect 18854 -7354 18882 -7326
rect 18882 -7354 18884 -7326
rect 18852 -7356 18884 -7354
rect 18852 -7486 18884 -7484
rect 18852 -7514 18854 -7486
rect 18854 -7514 18882 -7486
rect 18882 -7514 18884 -7486
rect 18852 -7516 18884 -7514
rect 18852 -7646 18884 -7644
rect 18852 -7674 18854 -7646
rect 18854 -7674 18882 -7646
rect 18882 -7674 18884 -7646
rect 18852 -7676 18884 -7674
rect 18852 -7806 18884 -7804
rect 18852 -7834 18854 -7806
rect 18854 -7834 18882 -7806
rect 18882 -7834 18884 -7806
rect 18852 -7836 18884 -7834
rect 18852 -7966 18884 -7964
rect 18852 -7994 18854 -7966
rect 18854 -7994 18882 -7966
rect 18882 -7994 18884 -7966
rect 18852 -7996 18884 -7994
rect 18852 -8126 18884 -8124
rect 18852 -8154 18854 -8126
rect 18854 -8154 18882 -8126
rect 18882 -8154 18884 -8126
rect 18852 -8156 18884 -8154
rect 18852 -8286 18884 -8284
rect 18852 -8314 18854 -8286
rect 18854 -8314 18882 -8286
rect 18882 -8314 18884 -8286
rect 18852 -8316 18884 -8314
rect 18852 -8446 18884 -8444
rect 18852 -8474 18854 -8446
rect 18854 -8474 18882 -8446
rect 18882 -8474 18884 -8446
rect 18852 -8476 18884 -8474
rect 18852 -8606 18884 -8604
rect 18852 -8634 18854 -8606
rect 18854 -8634 18882 -8606
rect 18882 -8634 18884 -8606
rect 18852 -8636 18884 -8634
rect 18852 -8766 18884 -8764
rect 18852 -8794 18854 -8766
rect 18854 -8794 18882 -8766
rect 18882 -8794 18884 -8766
rect 18852 -8796 18884 -8794
rect 18852 -8926 18884 -8924
rect 18852 -8954 18854 -8926
rect 18854 -8954 18882 -8926
rect 18882 -8954 18884 -8926
rect 18852 -8956 18884 -8954
rect 18852 -9086 18884 -9084
rect 18852 -9114 18854 -9086
rect 18854 -9114 18882 -9086
rect 18882 -9114 18884 -9086
rect 18852 -9116 18884 -9114
rect 15119 -9246 15151 -9244
rect 15119 -9274 15121 -9246
rect 15121 -9274 15149 -9246
rect 15149 -9274 15151 -9246
rect 15119 -9276 15151 -9274
rect 18852 -9246 18884 -9244
rect 18852 -9274 18854 -9246
rect 18854 -9274 18882 -9246
rect 18882 -9274 18884 -9246
rect 18852 -9276 18884 -9274
rect 15304 -9351 15336 -9349
rect 15304 -9379 15306 -9351
rect 15306 -9379 15334 -9351
rect 15334 -9379 15336 -9351
rect 15304 -9381 15336 -9379
rect 15464 -9351 15496 -9349
rect 15464 -9379 15466 -9351
rect 15466 -9379 15494 -9351
rect 15494 -9379 15496 -9351
rect 15464 -9381 15496 -9379
rect 15624 -9351 15656 -9349
rect 15624 -9379 15626 -9351
rect 15626 -9379 15654 -9351
rect 15654 -9379 15656 -9351
rect 15624 -9381 15656 -9379
rect 15784 -9351 15816 -9349
rect 15784 -9379 15786 -9351
rect 15786 -9379 15814 -9351
rect 15814 -9379 15816 -9351
rect 15784 -9381 15816 -9379
rect 15944 -9351 15976 -9349
rect 15944 -9379 15946 -9351
rect 15946 -9379 15974 -9351
rect 15974 -9379 15976 -9351
rect 15944 -9381 15976 -9379
rect 16104 -9351 16136 -9349
rect 16104 -9379 16106 -9351
rect 16106 -9379 16134 -9351
rect 16134 -9379 16136 -9351
rect 16104 -9381 16136 -9379
rect 16264 -9351 16296 -9349
rect 16264 -9379 16266 -9351
rect 16266 -9379 16294 -9351
rect 16294 -9379 16296 -9351
rect 16264 -9381 16296 -9379
rect 16424 -9351 16456 -9349
rect 16424 -9379 16426 -9351
rect 16426 -9379 16454 -9351
rect 16454 -9379 16456 -9351
rect 16424 -9381 16456 -9379
rect 16584 -9351 16616 -9349
rect 16584 -9379 16586 -9351
rect 16586 -9379 16614 -9351
rect 16614 -9379 16616 -9351
rect 16584 -9381 16616 -9379
rect 16744 -9351 16776 -9349
rect 16744 -9379 16746 -9351
rect 16746 -9379 16774 -9351
rect 16774 -9379 16776 -9351
rect 16744 -9381 16776 -9379
rect 16904 -9351 16936 -9349
rect 16904 -9379 16906 -9351
rect 16906 -9379 16934 -9351
rect 16934 -9379 16936 -9351
rect 16904 -9381 16936 -9379
rect 17064 -9351 17096 -9349
rect 17064 -9379 17066 -9351
rect 17066 -9379 17094 -9351
rect 17094 -9379 17096 -9351
rect 17064 -9381 17096 -9379
rect 17224 -9351 17256 -9349
rect 17224 -9379 17226 -9351
rect 17226 -9379 17254 -9351
rect 17254 -9379 17256 -9351
rect 17224 -9381 17256 -9379
rect 17384 -9351 17416 -9349
rect 17384 -9379 17386 -9351
rect 17386 -9379 17414 -9351
rect 17414 -9379 17416 -9351
rect 17384 -9381 17416 -9379
rect 17544 -9351 17576 -9349
rect 17544 -9379 17546 -9351
rect 17546 -9379 17574 -9351
rect 17574 -9379 17576 -9351
rect 17544 -9381 17576 -9379
rect 17704 -9351 17736 -9349
rect 17704 -9379 17706 -9351
rect 17706 -9379 17734 -9351
rect 17734 -9379 17736 -9351
rect 17704 -9381 17736 -9379
rect 17864 -9351 17896 -9349
rect 17864 -9379 17866 -9351
rect 17866 -9379 17894 -9351
rect 17894 -9379 17896 -9351
rect 17864 -9381 17896 -9379
rect 18024 -9351 18056 -9349
rect 18024 -9379 18026 -9351
rect 18026 -9379 18054 -9351
rect 18054 -9379 18056 -9351
rect 18024 -9381 18056 -9379
rect 18184 -9351 18216 -9349
rect 18184 -9379 18186 -9351
rect 18186 -9379 18214 -9351
rect 18214 -9379 18216 -9351
rect 18184 -9381 18216 -9379
rect 18344 -9351 18376 -9349
rect 18344 -9379 18346 -9351
rect 18346 -9379 18374 -9351
rect 18374 -9379 18376 -9351
rect 18344 -9381 18376 -9379
rect 18504 -9351 18536 -9349
rect 18504 -9379 18506 -9351
rect 18506 -9379 18534 -9351
rect 18534 -9379 18536 -9351
rect 18504 -9381 18536 -9379
rect 18664 -9351 18696 -9349
rect 18664 -9379 18666 -9351
rect 18666 -9379 18694 -9351
rect 18694 -9379 18696 -9351
rect 18664 -9381 18696 -9379
rect 21304 -5623 21336 -5621
rect 21304 -5651 21306 -5623
rect 21306 -5651 21334 -5623
rect 21334 -5651 21336 -5623
rect 21304 -5653 21336 -5651
rect 21464 -5623 21496 -5621
rect 21464 -5651 21466 -5623
rect 21466 -5651 21494 -5623
rect 21494 -5651 21496 -5623
rect 21464 -5653 21496 -5651
rect 21624 -5623 21656 -5621
rect 21624 -5651 21626 -5623
rect 21626 -5651 21654 -5623
rect 21654 -5651 21656 -5623
rect 21624 -5653 21656 -5651
rect 21784 -5623 21816 -5621
rect 21784 -5651 21786 -5623
rect 21786 -5651 21814 -5623
rect 21814 -5651 21816 -5623
rect 21784 -5653 21816 -5651
rect 21944 -5623 21976 -5621
rect 21944 -5651 21946 -5623
rect 21946 -5651 21974 -5623
rect 21974 -5651 21976 -5623
rect 21944 -5653 21976 -5651
rect 22104 -5623 22136 -5621
rect 22104 -5651 22106 -5623
rect 22106 -5651 22134 -5623
rect 22134 -5651 22136 -5623
rect 22104 -5653 22136 -5651
rect 22264 -5623 22296 -5621
rect 22264 -5651 22266 -5623
rect 22266 -5651 22294 -5623
rect 22294 -5651 22296 -5623
rect 22264 -5653 22296 -5651
rect 22424 -5623 22456 -5621
rect 22424 -5651 22426 -5623
rect 22426 -5651 22454 -5623
rect 22454 -5651 22456 -5623
rect 22424 -5653 22456 -5651
rect 22584 -5623 22616 -5621
rect 22584 -5651 22586 -5623
rect 22586 -5651 22614 -5623
rect 22614 -5651 22616 -5623
rect 22584 -5653 22616 -5651
rect 22744 -5623 22776 -5621
rect 22744 -5651 22746 -5623
rect 22746 -5651 22774 -5623
rect 22774 -5651 22776 -5623
rect 22744 -5653 22776 -5651
rect 22904 -5623 22936 -5621
rect 22904 -5651 22906 -5623
rect 22906 -5651 22934 -5623
rect 22934 -5651 22936 -5623
rect 22904 -5653 22936 -5651
rect 23064 -5623 23096 -5621
rect 23064 -5651 23066 -5623
rect 23066 -5651 23094 -5623
rect 23094 -5651 23096 -5623
rect 23064 -5653 23096 -5651
rect 23224 -5623 23256 -5621
rect 23224 -5651 23226 -5623
rect 23226 -5651 23254 -5623
rect 23254 -5651 23256 -5623
rect 23224 -5653 23256 -5651
rect 23384 -5623 23416 -5621
rect 23384 -5651 23386 -5623
rect 23386 -5651 23414 -5623
rect 23414 -5651 23416 -5623
rect 23384 -5653 23416 -5651
rect 23544 -5623 23576 -5621
rect 23544 -5651 23546 -5623
rect 23546 -5651 23574 -5623
rect 23574 -5651 23576 -5623
rect 23544 -5653 23576 -5651
rect 23704 -5623 23736 -5621
rect 23704 -5651 23706 -5623
rect 23706 -5651 23734 -5623
rect 23734 -5651 23736 -5623
rect 23704 -5653 23736 -5651
rect 23864 -5623 23896 -5621
rect 23864 -5651 23866 -5623
rect 23866 -5651 23894 -5623
rect 23894 -5651 23896 -5623
rect 23864 -5653 23896 -5651
rect 24024 -5623 24056 -5621
rect 24024 -5651 24026 -5623
rect 24026 -5651 24054 -5623
rect 24054 -5651 24056 -5623
rect 24024 -5653 24056 -5651
rect 24184 -5623 24216 -5621
rect 24184 -5651 24186 -5623
rect 24186 -5651 24214 -5623
rect 24214 -5651 24216 -5623
rect 24184 -5653 24216 -5651
rect 24344 -5623 24376 -5621
rect 24344 -5651 24346 -5623
rect 24346 -5651 24374 -5623
rect 24374 -5651 24376 -5623
rect 24344 -5653 24376 -5651
rect 24504 -5623 24536 -5621
rect 24504 -5651 24506 -5623
rect 24506 -5651 24534 -5623
rect 24534 -5651 24536 -5623
rect 24504 -5653 24536 -5651
rect 24664 -5623 24696 -5621
rect 24664 -5651 24666 -5623
rect 24666 -5651 24694 -5623
rect 24694 -5651 24696 -5623
rect 24664 -5653 24696 -5651
rect 21119 -5726 21151 -5724
rect 21119 -5754 21121 -5726
rect 21121 -5754 21149 -5726
rect 21149 -5754 21151 -5726
rect 21119 -5756 21151 -5754
rect 24852 -5726 24884 -5724
rect 24852 -5754 24854 -5726
rect 24854 -5754 24882 -5726
rect 24882 -5754 24884 -5726
rect 24852 -5756 24884 -5754
rect 21119 -5886 21151 -5884
rect 21119 -5914 21121 -5886
rect 21121 -5914 21149 -5886
rect 21149 -5914 21151 -5886
rect 21119 -5916 21151 -5914
rect 21119 -6046 21151 -6044
rect 21119 -6074 21121 -6046
rect 21121 -6074 21149 -6046
rect 21149 -6074 21151 -6046
rect 21119 -6076 21151 -6074
rect 21119 -6206 21151 -6204
rect 21119 -6234 21121 -6206
rect 21121 -6234 21149 -6206
rect 21149 -6234 21151 -6206
rect 21119 -6236 21151 -6234
rect 21119 -6366 21151 -6364
rect 21119 -6394 21121 -6366
rect 21121 -6394 21149 -6366
rect 21149 -6394 21151 -6366
rect 21119 -6396 21151 -6394
rect 21119 -6526 21151 -6524
rect 21119 -6554 21121 -6526
rect 21121 -6554 21149 -6526
rect 21149 -6554 21151 -6526
rect 21119 -6556 21151 -6554
rect 21119 -6686 21151 -6684
rect 21119 -6714 21121 -6686
rect 21121 -6714 21149 -6686
rect 21149 -6714 21151 -6686
rect 21119 -6716 21151 -6714
rect 21119 -6846 21151 -6844
rect 21119 -6874 21121 -6846
rect 21121 -6874 21149 -6846
rect 21149 -6874 21151 -6846
rect 21119 -6876 21151 -6874
rect 21119 -7006 21151 -7004
rect 21119 -7034 21121 -7006
rect 21121 -7034 21149 -7006
rect 21149 -7034 21151 -7006
rect 21119 -7036 21151 -7034
rect 21119 -7166 21151 -7164
rect 21119 -7194 21121 -7166
rect 21121 -7194 21149 -7166
rect 21149 -7194 21151 -7166
rect 21119 -7196 21151 -7194
rect 21119 -7326 21151 -7324
rect 21119 -7354 21121 -7326
rect 21121 -7354 21149 -7326
rect 21149 -7354 21151 -7326
rect 21119 -7356 21151 -7354
rect 21119 -7486 21151 -7484
rect 21119 -7514 21121 -7486
rect 21121 -7514 21149 -7486
rect 21149 -7514 21151 -7486
rect 21119 -7516 21151 -7514
rect 21119 -7646 21151 -7644
rect 21119 -7674 21121 -7646
rect 21121 -7674 21149 -7646
rect 21149 -7674 21151 -7646
rect 21119 -7676 21151 -7674
rect 21119 -7806 21151 -7804
rect 21119 -7834 21121 -7806
rect 21121 -7834 21149 -7806
rect 21149 -7834 21151 -7806
rect 21119 -7836 21151 -7834
rect 21119 -7966 21151 -7964
rect 21119 -7994 21121 -7966
rect 21121 -7994 21149 -7966
rect 21149 -7994 21151 -7966
rect 21119 -7996 21151 -7994
rect 21119 -8126 21151 -8124
rect 21119 -8154 21121 -8126
rect 21121 -8154 21149 -8126
rect 21149 -8154 21151 -8126
rect 21119 -8156 21151 -8154
rect 21119 -8286 21151 -8284
rect 21119 -8314 21121 -8286
rect 21121 -8314 21149 -8286
rect 21149 -8314 21151 -8286
rect 21119 -8316 21151 -8314
rect 21119 -8446 21151 -8444
rect 21119 -8474 21121 -8446
rect 21121 -8474 21149 -8446
rect 21149 -8474 21151 -8446
rect 21119 -8476 21151 -8474
rect 21119 -8606 21151 -8604
rect 21119 -8634 21121 -8606
rect 21121 -8634 21149 -8606
rect 21149 -8634 21151 -8606
rect 21119 -8636 21151 -8634
rect 21119 -8766 21151 -8764
rect 21119 -8794 21121 -8766
rect 21121 -8794 21149 -8766
rect 21149 -8794 21151 -8766
rect 21119 -8796 21151 -8794
rect 21119 -8926 21151 -8924
rect 21119 -8954 21121 -8926
rect 21121 -8954 21149 -8926
rect 21149 -8954 21151 -8926
rect 21119 -8956 21151 -8954
rect 21119 -9086 21151 -9084
rect 21119 -9114 21121 -9086
rect 21121 -9114 21149 -9086
rect 21149 -9114 21151 -9086
rect 21119 -9116 21151 -9114
rect 24852 -5886 24884 -5884
rect 24852 -5914 24854 -5886
rect 24854 -5914 24882 -5886
rect 24882 -5914 24884 -5886
rect 24852 -5916 24884 -5914
rect 24852 -6046 24884 -6044
rect 24852 -6074 24854 -6046
rect 24854 -6074 24882 -6046
rect 24882 -6074 24884 -6046
rect 24852 -6076 24884 -6074
rect 24852 -6206 24884 -6204
rect 24852 -6234 24854 -6206
rect 24854 -6234 24882 -6206
rect 24882 -6234 24884 -6206
rect 24852 -6236 24884 -6234
rect 24852 -6366 24884 -6364
rect 24852 -6394 24854 -6366
rect 24854 -6394 24882 -6366
rect 24882 -6394 24884 -6366
rect 24852 -6396 24884 -6394
rect 24852 -6526 24884 -6524
rect 24852 -6554 24854 -6526
rect 24854 -6554 24882 -6526
rect 24882 -6554 24884 -6526
rect 24852 -6556 24884 -6554
rect 24852 -6686 24884 -6684
rect 24852 -6714 24854 -6686
rect 24854 -6714 24882 -6686
rect 24882 -6714 24884 -6686
rect 24852 -6716 24884 -6714
rect 24852 -6846 24884 -6844
rect 24852 -6874 24854 -6846
rect 24854 -6874 24882 -6846
rect 24882 -6874 24884 -6846
rect 24852 -6876 24884 -6874
rect 24852 -7006 24884 -7004
rect 24852 -7034 24854 -7006
rect 24854 -7034 24882 -7006
rect 24882 -7034 24884 -7006
rect 24852 -7036 24884 -7034
rect 24852 -7166 24884 -7164
rect 24852 -7194 24854 -7166
rect 24854 -7194 24882 -7166
rect 24882 -7194 24884 -7166
rect 24852 -7196 24884 -7194
rect 24852 -7326 24884 -7324
rect 24852 -7354 24854 -7326
rect 24854 -7354 24882 -7326
rect 24882 -7354 24884 -7326
rect 24852 -7356 24884 -7354
rect 24852 -7486 24884 -7484
rect 24852 -7514 24854 -7486
rect 24854 -7514 24882 -7486
rect 24882 -7514 24884 -7486
rect 24852 -7516 24884 -7514
rect 24852 -7646 24884 -7644
rect 24852 -7674 24854 -7646
rect 24854 -7674 24882 -7646
rect 24882 -7674 24884 -7646
rect 24852 -7676 24884 -7674
rect 24852 -7806 24884 -7804
rect 24852 -7834 24854 -7806
rect 24854 -7834 24882 -7806
rect 24882 -7834 24884 -7806
rect 24852 -7836 24884 -7834
rect 24852 -7966 24884 -7964
rect 24852 -7994 24854 -7966
rect 24854 -7994 24882 -7966
rect 24882 -7994 24884 -7966
rect 24852 -7996 24884 -7994
rect 24852 -8126 24884 -8124
rect 24852 -8154 24854 -8126
rect 24854 -8154 24882 -8126
rect 24882 -8154 24884 -8126
rect 24852 -8156 24884 -8154
rect 24852 -8286 24884 -8284
rect 24852 -8314 24854 -8286
rect 24854 -8314 24882 -8286
rect 24882 -8314 24884 -8286
rect 24852 -8316 24884 -8314
rect 24852 -8446 24884 -8444
rect 24852 -8474 24854 -8446
rect 24854 -8474 24882 -8446
rect 24882 -8474 24884 -8446
rect 24852 -8476 24884 -8474
rect 24852 -8606 24884 -8604
rect 24852 -8634 24854 -8606
rect 24854 -8634 24882 -8606
rect 24882 -8634 24884 -8606
rect 24852 -8636 24884 -8634
rect 24852 -8766 24884 -8764
rect 24852 -8794 24854 -8766
rect 24854 -8794 24882 -8766
rect 24882 -8794 24884 -8766
rect 24852 -8796 24884 -8794
rect 24852 -8926 24884 -8924
rect 24852 -8954 24854 -8926
rect 24854 -8954 24882 -8926
rect 24882 -8954 24884 -8926
rect 24852 -8956 24884 -8954
rect 24852 -9086 24884 -9084
rect 24852 -9114 24854 -9086
rect 24854 -9114 24882 -9086
rect 24882 -9114 24884 -9086
rect 24852 -9116 24884 -9114
rect 21119 -9246 21151 -9244
rect 21119 -9274 21121 -9246
rect 21121 -9274 21149 -9246
rect 21149 -9274 21151 -9246
rect 21119 -9276 21151 -9274
rect 24852 -9246 24884 -9244
rect 24852 -9274 24854 -9246
rect 24854 -9274 24882 -9246
rect 24882 -9274 24884 -9246
rect 24852 -9276 24884 -9274
rect 21304 -9351 21336 -9349
rect 21304 -9379 21306 -9351
rect 21306 -9379 21334 -9351
rect 21334 -9379 21336 -9351
rect 21304 -9381 21336 -9379
rect 21464 -9351 21496 -9349
rect 21464 -9379 21466 -9351
rect 21466 -9379 21494 -9351
rect 21494 -9379 21496 -9351
rect 21464 -9381 21496 -9379
rect 21624 -9351 21656 -9349
rect 21624 -9379 21626 -9351
rect 21626 -9379 21654 -9351
rect 21654 -9379 21656 -9351
rect 21624 -9381 21656 -9379
rect 21784 -9351 21816 -9349
rect 21784 -9379 21786 -9351
rect 21786 -9379 21814 -9351
rect 21814 -9379 21816 -9351
rect 21784 -9381 21816 -9379
rect 21944 -9351 21976 -9349
rect 21944 -9379 21946 -9351
rect 21946 -9379 21974 -9351
rect 21974 -9379 21976 -9351
rect 21944 -9381 21976 -9379
rect 22104 -9351 22136 -9349
rect 22104 -9379 22106 -9351
rect 22106 -9379 22134 -9351
rect 22134 -9379 22136 -9351
rect 22104 -9381 22136 -9379
rect 22264 -9351 22296 -9349
rect 22264 -9379 22266 -9351
rect 22266 -9379 22294 -9351
rect 22294 -9379 22296 -9351
rect 22264 -9381 22296 -9379
rect 22424 -9351 22456 -9349
rect 22424 -9379 22426 -9351
rect 22426 -9379 22454 -9351
rect 22454 -9379 22456 -9351
rect 22424 -9381 22456 -9379
rect 22584 -9351 22616 -9349
rect 22584 -9379 22586 -9351
rect 22586 -9379 22614 -9351
rect 22614 -9379 22616 -9351
rect 22584 -9381 22616 -9379
rect 22744 -9351 22776 -9349
rect 22744 -9379 22746 -9351
rect 22746 -9379 22774 -9351
rect 22774 -9379 22776 -9351
rect 22744 -9381 22776 -9379
rect 22904 -9351 22936 -9349
rect 22904 -9379 22906 -9351
rect 22906 -9379 22934 -9351
rect 22934 -9379 22936 -9351
rect 22904 -9381 22936 -9379
rect 23064 -9351 23096 -9349
rect 23064 -9379 23066 -9351
rect 23066 -9379 23094 -9351
rect 23094 -9379 23096 -9351
rect 23064 -9381 23096 -9379
rect 23224 -9351 23256 -9349
rect 23224 -9379 23226 -9351
rect 23226 -9379 23254 -9351
rect 23254 -9379 23256 -9351
rect 23224 -9381 23256 -9379
rect 23384 -9351 23416 -9349
rect 23384 -9379 23386 -9351
rect 23386 -9379 23414 -9351
rect 23414 -9379 23416 -9351
rect 23384 -9381 23416 -9379
rect 23544 -9351 23576 -9349
rect 23544 -9379 23546 -9351
rect 23546 -9379 23574 -9351
rect 23574 -9379 23576 -9351
rect 23544 -9381 23576 -9379
rect 23704 -9351 23736 -9349
rect 23704 -9379 23706 -9351
rect 23706 -9379 23734 -9351
rect 23734 -9379 23736 -9351
rect 23704 -9381 23736 -9379
rect 23864 -9351 23896 -9349
rect 23864 -9379 23866 -9351
rect 23866 -9379 23894 -9351
rect 23894 -9379 23896 -9351
rect 23864 -9381 23896 -9379
rect 24024 -9351 24056 -9349
rect 24024 -9379 24026 -9351
rect 24026 -9379 24054 -9351
rect 24054 -9379 24056 -9351
rect 24024 -9381 24056 -9379
rect 24184 -9351 24216 -9349
rect 24184 -9379 24186 -9351
rect 24186 -9379 24214 -9351
rect 24214 -9379 24216 -9351
rect 24184 -9381 24216 -9379
rect 24344 -9351 24376 -9349
rect 24344 -9379 24346 -9351
rect 24346 -9379 24374 -9351
rect 24374 -9379 24376 -9351
rect 24344 -9381 24376 -9379
rect 24504 -9351 24536 -9349
rect 24504 -9379 24506 -9351
rect 24506 -9379 24534 -9351
rect 24534 -9379 24536 -9351
rect 24504 -9381 24536 -9379
rect 24664 -9351 24696 -9349
rect 24664 -9379 24666 -9351
rect 24666 -9379 24694 -9351
rect 24694 -9379 24696 -9351
rect 24664 -9381 24696 -9379
rect 9304 -11623 9336 -11621
rect 9304 -11651 9306 -11623
rect 9306 -11651 9334 -11623
rect 9334 -11651 9336 -11623
rect 9304 -11653 9336 -11651
rect 9464 -11623 9496 -11621
rect 9464 -11651 9466 -11623
rect 9466 -11651 9494 -11623
rect 9494 -11651 9496 -11623
rect 9464 -11653 9496 -11651
rect 9624 -11623 9656 -11621
rect 9624 -11651 9626 -11623
rect 9626 -11651 9654 -11623
rect 9654 -11651 9656 -11623
rect 9624 -11653 9656 -11651
rect 9784 -11623 9816 -11621
rect 9784 -11651 9786 -11623
rect 9786 -11651 9814 -11623
rect 9814 -11651 9816 -11623
rect 9784 -11653 9816 -11651
rect 9944 -11623 9976 -11621
rect 9944 -11651 9946 -11623
rect 9946 -11651 9974 -11623
rect 9974 -11651 9976 -11623
rect 9944 -11653 9976 -11651
rect 10104 -11623 10136 -11621
rect 10104 -11651 10106 -11623
rect 10106 -11651 10134 -11623
rect 10134 -11651 10136 -11623
rect 10104 -11653 10136 -11651
rect 10264 -11623 10296 -11621
rect 10264 -11651 10266 -11623
rect 10266 -11651 10294 -11623
rect 10294 -11651 10296 -11623
rect 10264 -11653 10296 -11651
rect 10424 -11623 10456 -11621
rect 10424 -11651 10426 -11623
rect 10426 -11651 10454 -11623
rect 10454 -11651 10456 -11623
rect 10424 -11653 10456 -11651
rect 10584 -11623 10616 -11621
rect 10584 -11651 10586 -11623
rect 10586 -11651 10614 -11623
rect 10614 -11651 10616 -11623
rect 10584 -11653 10616 -11651
rect 10744 -11623 10776 -11621
rect 10744 -11651 10746 -11623
rect 10746 -11651 10774 -11623
rect 10774 -11651 10776 -11623
rect 10744 -11653 10776 -11651
rect 10904 -11623 10936 -11621
rect 10904 -11651 10906 -11623
rect 10906 -11651 10934 -11623
rect 10934 -11651 10936 -11623
rect 10904 -11653 10936 -11651
rect 11064 -11623 11096 -11621
rect 11064 -11651 11066 -11623
rect 11066 -11651 11094 -11623
rect 11094 -11651 11096 -11623
rect 11064 -11653 11096 -11651
rect 11224 -11623 11256 -11621
rect 11224 -11651 11226 -11623
rect 11226 -11651 11254 -11623
rect 11254 -11651 11256 -11623
rect 11224 -11653 11256 -11651
rect 11384 -11623 11416 -11621
rect 11384 -11651 11386 -11623
rect 11386 -11651 11414 -11623
rect 11414 -11651 11416 -11623
rect 11384 -11653 11416 -11651
rect 11544 -11623 11576 -11621
rect 11544 -11651 11546 -11623
rect 11546 -11651 11574 -11623
rect 11574 -11651 11576 -11623
rect 11544 -11653 11576 -11651
rect 11704 -11623 11736 -11621
rect 11704 -11651 11706 -11623
rect 11706 -11651 11734 -11623
rect 11734 -11651 11736 -11623
rect 11704 -11653 11736 -11651
rect 11864 -11623 11896 -11621
rect 11864 -11651 11866 -11623
rect 11866 -11651 11894 -11623
rect 11894 -11651 11896 -11623
rect 11864 -11653 11896 -11651
rect 12024 -11623 12056 -11621
rect 12024 -11651 12026 -11623
rect 12026 -11651 12054 -11623
rect 12054 -11651 12056 -11623
rect 12024 -11653 12056 -11651
rect 12184 -11623 12216 -11621
rect 12184 -11651 12186 -11623
rect 12186 -11651 12214 -11623
rect 12214 -11651 12216 -11623
rect 12184 -11653 12216 -11651
rect 12344 -11623 12376 -11621
rect 12344 -11651 12346 -11623
rect 12346 -11651 12374 -11623
rect 12374 -11651 12376 -11623
rect 12344 -11653 12376 -11651
rect 12504 -11623 12536 -11621
rect 12504 -11651 12506 -11623
rect 12506 -11651 12534 -11623
rect 12534 -11651 12536 -11623
rect 12504 -11653 12536 -11651
rect 12664 -11623 12696 -11621
rect 12664 -11651 12666 -11623
rect 12666 -11651 12694 -11623
rect 12694 -11651 12696 -11623
rect 12664 -11653 12696 -11651
rect 9119 -11726 9151 -11724
rect 9119 -11754 9121 -11726
rect 9121 -11754 9149 -11726
rect 9149 -11754 9151 -11726
rect 9119 -11756 9151 -11754
rect 12852 -11726 12884 -11724
rect 12852 -11754 12854 -11726
rect 12854 -11754 12882 -11726
rect 12882 -11754 12884 -11726
rect 12852 -11756 12884 -11754
rect 9119 -11886 9151 -11884
rect 9119 -11914 9121 -11886
rect 9121 -11914 9149 -11886
rect 9149 -11914 9151 -11886
rect 9119 -11916 9151 -11914
rect 9119 -12046 9151 -12044
rect 9119 -12074 9121 -12046
rect 9121 -12074 9149 -12046
rect 9149 -12074 9151 -12046
rect 9119 -12076 9151 -12074
rect 9119 -12206 9151 -12204
rect 9119 -12234 9121 -12206
rect 9121 -12234 9149 -12206
rect 9149 -12234 9151 -12206
rect 9119 -12236 9151 -12234
rect 9119 -12366 9151 -12364
rect 9119 -12394 9121 -12366
rect 9121 -12394 9149 -12366
rect 9149 -12394 9151 -12366
rect 9119 -12396 9151 -12394
rect 9119 -12526 9151 -12524
rect 9119 -12554 9121 -12526
rect 9121 -12554 9149 -12526
rect 9149 -12554 9151 -12526
rect 9119 -12556 9151 -12554
rect 9119 -12686 9151 -12684
rect 9119 -12714 9121 -12686
rect 9121 -12714 9149 -12686
rect 9149 -12714 9151 -12686
rect 9119 -12716 9151 -12714
rect 9119 -12846 9151 -12844
rect 9119 -12874 9121 -12846
rect 9121 -12874 9149 -12846
rect 9149 -12874 9151 -12846
rect 9119 -12876 9151 -12874
rect 6852 -13006 6884 -13004
rect 6852 -13034 6854 -13006
rect 6854 -13034 6882 -13006
rect 6882 -13034 6884 -13006
rect 6852 -13036 6884 -13034
rect 6852 -13166 6884 -13164
rect 6852 -13194 6854 -13166
rect 6854 -13194 6882 -13166
rect 6882 -13194 6884 -13166
rect 6852 -13196 6884 -13194
rect 6852 -13326 6884 -13324
rect 6852 -13354 6854 -13326
rect 6854 -13354 6882 -13326
rect 6882 -13354 6884 -13326
rect 6852 -13356 6884 -13354
rect 6852 -13486 6884 -13484
rect 6852 -13514 6854 -13486
rect 6854 -13514 6882 -13486
rect 6882 -13514 6884 -13486
rect 6852 -13516 6884 -13514
rect 6852 -13646 6884 -13644
rect 6852 -13674 6854 -13646
rect 6854 -13674 6882 -13646
rect 6882 -13674 6884 -13646
rect 6852 -13676 6884 -13674
rect 6852 -13806 6884 -13804
rect 6852 -13834 6854 -13806
rect 6854 -13834 6882 -13806
rect 6882 -13834 6884 -13806
rect 6852 -13836 6884 -13834
rect 6852 -13966 6884 -13964
rect 6852 -13994 6854 -13966
rect 6854 -13994 6882 -13966
rect 6882 -13994 6884 -13966
rect 6852 -13996 6884 -13994
rect 6852 -14126 6884 -14124
rect 6852 -14154 6854 -14126
rect 6854 -14154 6882 -14126
rect 6882 -14154 6884 -14126
rect 6852 -14156 6884 -14154
rect 6852 -14286 6884 -14284
rect 6852 -14314 6854 -14286
rect 6854 -14314 6882 -14286
rect 6882 -14314 6884 -14286
rect 6852 -14316 6884 -14314
rect 6852 -14446 6884 -14444
rect 6852 -14474 6854 -14446
rect 6854 -14474 6882 -14446
rect 6882 -14474 6884 -14446
rect 6852 -14476 6884 -14474
rect 6852 -14606 6884 -14604
rect 6852 -14634 6854 -14606
rect 6854 -14634 6882 -14606
rect 6882 -14634 6884 -14606
rect 6852 -14636 6884 -14634
rect 6852 -14766 6884 -14764
rect 6852 -14794 6854 -14766
rect 6854 -14794 6882 -14766
rect 6882 -14794 6884 -14766
rect 6852 -14796 6884 -14794
rect 6852 -14926 6884 -14924
rect 6852 -14954 6854 -14926
rect 6854 -14954 6882 -14926
rect 6882 -14954 6884 -14926
rect 6852 -14956 6884 -14954
rect 6852 -15086 6884 -15084
rect 6852 -15114 6854 -15086
rect 6854 -15114 6882 -15086
rect 6882 -15114 6884 -15086
rect 6852 -15116 6884 -15114
rect 3119 -15246 3151 -15244
rect 3119 -15274 3121 -15246
rect 3121 -15274 3149 -15246
rect 3149 -15274 3151 -15246
rect 3119 -15276 3151 -15274
rect 6852 -15246 6884 -15244
rect 6852 -15274 6854 -15246
rect 6854 -15274 6882 -15246
rect 6882 -15274 6884 -15246
rect 6852 -15276 6884 -15274
rect 3304 -15351 3336 -15349
rect 3304 -15379 3306 -15351
rect 3306 -15379 3334 -15351
rect 3334 -15379 3336 -15351
rect 3304 -15381 3336 -15379
rect 3464 -15351 3496 -15349
rect 3464 -15379 3466 -15351
rect 3466 -15379 3494 -15351
rect 3494 -15379 3496 -15351
rect 3464 -15381 3496 -15379
rect 3624 -15351 3656 -15349
rect 3624 -15379 3626 -15351
rect 3626 -15379 3654 -15351
rect 3654 -15379 3656 -15351
rect 3624 -15381 3656 -15379
rect 3784 -15351 3816 -15349
rect 3784 -15379 3786 -15351
rect 3786 -15379 3814 -15351
rect 3814 -15379 3816 -15351
rect 3784 -15381 3816 -15379
rect 3944 -15351 3976 -15349
rect 3944 -15379 3946 -15351
rect 3946 -15379 3974 -15351
rect 3974 -15379 3976 -15351
rect 3944 -15381 3976 -15379
rect 4104 -15351 4136 -15349
rect 4104 -15379 4106 -15351
rect 4106 -15379 4134 -15351
rect 4134 -15379 4136 -15351
rect 4104 -15381 4136 -15379
rect 4264 -15351 4296 -15349
rect 4264 -15379 4266 -15351
rect 4266 -15379 4294 -15351
rect 4294 -15379 4296 -15351
rect 4264 -15381 4296 -15379
rect 4424 -15351 4456 -15349
rect 4424 -15379 4426 -15351
rect 4426 -15379 4454 -15351
rect 4454 -15379 4456 -15351
rect 4424 -15381 4456 -15379
rect 4584 -15351 4616 -15349
rect 4584 -15379 4586 -15351
rect 4586 -15379 4614 -15351
rect 4614 -15379 4616 -15351
rect 4584 -15381 4616 -15379
rect 4744 -15351 4776 -15349
rect 4744 -15379 4746 -15351
rect 4746 -15379 4774 -15351
rect 4774 -15379 4776 -15351
rect 4744 -15381 4776 -15379
rect 4904 -15351 4936 -15349
rect 4904 -15379 4906 -15351
rect 4906 -15379 4934 -15351
rect 4934 -15379 4936 -15351
rect 4904 -15381 4936 -15379
rect 5064 -15351 5096 -15349
rect 5064 -15379 5066 -15351
rect 5066 -15379 5094 -15351
rect 5094 -15379 5096 -15351
rect 5064 -15381 5096 -15379
rect 5224 -15351 5256 -15349
rect 5224 -15379 5226 -15351
rect 5226 -15379 5254 -15351
rect 5254 -15379 5256 -15351
rect 5224 -15381 5256 -15379
rect 5384 -15351 5416 -15349
rect 5384 -15379 5386 -15351
rect 5386 -15379 5414 -15351
rect 5414 -15379 5416 -15351
rect 5384 -15381 5416 -15379
rect 5544 -15351 5576 -15349
rect 5544 -15379 5546 -15351
rect 5546 -15379 5574 -15351
rect 5574 -15379 5576 -15351
rect 5544 -15381 5576 -15379
rect 5704 -15351 5736 -15349
rect 5704 -15379 5706 -15351
rect 5706 -15379 5734 -15351
rect 5734 -15379 5736 -15351
rect 5704 -15381 5736 -15379
rect 5864 -15351 5896 -15349
rect 5864 -15379 5866 -15351
rect 5866 -15379 5894 -15351
rect 5894 -15379 5896 -15351
rect 5864 -15381 5896 -15379
rect 6024 -15351 6056 -15349
rect 6024 -15379 6026 -15351
rect 6026 -15379 6054 -15351
rect 6054 -15379 6056 -15351
rect 6024 -15381 6056 -15379
rect 6184 -15351 6216 -15349
rect 6184 -15379 6186 -15351
rect 6186 -15379 6214 -15351
rect 6214 -15379 6216 -15351
rect 6184 -15381 6216 -15379
rect 6344 -15351 6376 -15349
rect 6344 -15379 6346 -15351
rect 6346 -15379 6374 -15351
rect 6374 -15379 6376 -15351
rect 6344 -15381 6376 -15379
rect 6504 -15351 6536 -15349
rect 6504 -15379 6506 -15351
rect 6506 -15379 6534 -15351
rect 6534 -15379 6536 -15351
rect 6504 -15381 6536 -15379
rect 6664 -15351 6696 -15349
rect 6664 -15379 6666 -15351
rect 6666 -15379 6694 -15351
rect 6694 -15379 6696 -15351
rect 6664 -15381 6696 -15379
rect 9119 -13006 9151 -13004
rect 9119 -13034 9121 -13006
rect 9121 -13034 9149 -13006
rect 9149 -13034 9151 -13006
rect 9119 -13036 9151 -13034
rect 9119 -13166 9151 -13164
rect 9119 -13194 9121 -13166
rect 9121 -13194 9149 -13166
rect 9149 -13194 9151 -13166
rect 9119 -13196 9151 -13194
rect 9119 -13326 9151 -13324
rect 9119 -13354 9121 -13326
rect 9121 -13354 9149 -13326
rect 9149 -13354 9151 -13326
rect 9119 -13356 9151 -13354
rect 9119 -13486 9151 -13484
rect 9119 -13514 9121 -13486
rect 9121 -13514 9149 -13486
rect 9149 -13514 9151 -13486
rect 9119 -13516 9151 -13514
rect 9119 -13646 9151 -13644
rect 9119 -13674 9121 -13646
rect 9121 -13674 9149 -13646
rect 9149 -13674 9151 -13646
rect 9119 -13676 9151 -13674
rect 9119 -13806 9151 -13804
rect 9119 -13834 9121 -13806
rect 9121 -13834 9149 -13806
rect 9149 -13834 9151 -13806
rect 9119 -13836 9151 -13834
rect 9119 -13966 9151 -13964
rect 9119 -13994 9121 -13966
rect 9121 -13994 9149 -13966
rect 9149 -13994 9151 -13966
rect 9119 -13996 9151 -13994
rect 9119 -14126 9151 -14124
rect 9119 -14154 9121 -14126
rect 9121 -14154 9149 -14126
rect 9149 -14154 9151 -14126
rect 9119 -14156 9151 -14154
rect 9119 -14286 9151 -14284
rect 9119 -14314 9121 -14286
rect 9121 -14314 9149 -14286
rect 9149 -14314 9151 -14286
rect 9119 -14316 9151 -14314
rect 9119 -14446 9151 -14444
rect 9119 -14474 9121 -14446
rect 9121 -14474 9149 -14446
rect 9149 -14474 9151 -14446
rect 9119 -14476 9151 -14474
rect 9119 -14606 9151 -14604
rect 9119 -14634 9121 -14606
rect 9121 -14634 9149 -14606
rect 9149 -14634 9151 -14606
rect 9119 -14636 9151 -14634
rect 9119 -14766 9151 -14764
rect 9119 -14794 9121 -14766
rect 9121 -14794 9149 -14766
rect 9149 -14794 9151 -14766
rect 9119 -14796 9151 -14794
rect 9119 -14926 9151 -14924
rect 9119 -14954 9121 -14926
rect 9121 -14954 9149 -14926
rect 9149 -14954 9151 -14926
rect 9119 -14956 9151 -14954
rect 9119 -15086 9151 -15084
rect 9119 -15114 9121 -15086
rect 9121 -15114 9149 -15086
rect 9149 -15114 9151 -15086
rect 9119 -15116 9151 -15114
rect 12852 -11886 12884 -11884
rect 12852 -11914 12854 -11886
rect 12854 -11914 12882 -11886
rect 12882 -11914 12884 -11886
rect 12852 -11916 12884 -11914
rect 12852 -12046 12884 -12044
rect 12852 -12074 12854 -12046
rect 12854 -12074 12882 -12046
rect 12882 -12074 12884 -12046
rect 12852 -12076 12884 -12074
rect 12852 -12206 12884 -12204
rect 12852 -12234 12854 -12206
rect 12854 -12234 12882 -12206
rect 12882 -12234 12884 -12206
rect 12852 -12236 12884 -12234
rect 12852 -12366 12884 -12364
rect 12852 -12394 12854 -12366
rect 12854 -12394 12882 -12366
rect 12882 -12394 12884 -12366
rect 12852 -12396 12884 -12394
rect 12852 -12526 12884 -12524
rect 12852 -12554 12854 -12526
rect 12854 -12554 12882 -12526
rect 12882 -12554 12884 -12526
rect 12852 -12556 12884 -12554
rect 12852 -12686 12884 -12684
rect 12852 -12714 12854 -12686
rect 12854 -12714 12882 -12686
rect 12882 -12714 12884 -12686
rect 12852 -12716 12884 -12714
rect 12852 -12846 12884 -12844
rect 12852 -12874 12854 -12846
rect 12854 -12874 12882 -12846
rect 12882 -12874 12884 -12846
rect 12852 -12876 12884 -12874
rect 15304 -11623 15336 -11621
rect 15304 -11651 15306 -11623
rect 15306 -11651 15334 -11623
rect 15334 -11651 15336 -11623
rect 15304 -11653 15336 -11651
rect 15464 -11623 15496 -11621
rect 15464 -11651 15466 -11623
rect 15466 -11651 15494 -11623
rect 15494 -11651 15496 -11623
rect 15464 -11653 15496 -11651
rect 15624 -11623 15656 -11621
rect 15624 -11651 15626 -11623
rect 15626 -11651 15654 -11623
rect 15654 -11651 15656 -11623
rect 15624 -11653 15656 -11651
rect 15784 -11623 15816 -11621
rect 15784 -11651 15786 -11623
rect 15786 -11651 15814 -11623
rect 15814 -11651 15816 -11623
rect 15784 -11653 15816 -11651
rect 15944 -11623 15976 -11621
rect 15944 -11651 15946 -11623
rect 15946 -11651 15974 -11623
rect 15974 -11651 15976 -11623
rect 15944 -11653 15976 -11651
rect 16104 -11623 16136 -11621
rect 16104 -11651 16106 -11623
rect 16106 -11651 16134 -11623
rect 16134 -11651 16136 -11623
rect 16104 -11653 16136 -11651
rect 16264 -11623 16296 -11621
rect 16264 -11651 16266 -11623
rect 16266 -11651 16294 -11623
rect 16294 -11651 16296 -11623
rect 16264 -11653 16296 -11651
rect 16424 -11623 16456 -11621
rect 16424 -11651 16426 -11623
rect 16426 -11651 16454 -11623
rect 16454 -11651 16456 -11623
rect 16424 -11653 16456 -11651
rect 16584 -11623 16616 -11621
rect 16584 -11651 16586 -11623
rect 16586 -11651 16614 -11623
rect 16614 -11651 16616 -11623
rect 16584 -11653 16616 -11651
rect 16744 -11623 16776 -11621
rect 16744 -11651 16746 -11623
rect 16746 -11651 16774 -11623
rect 16774 -11651 16776 -11623
rect 16744 -11653 16776 -11651
rect 16904 -11623 16936 -11621
rect 16904 -11651 16906 -11623
rect 16906 -11651 16934 -11623
rect 16934 -11651 16936 -11623
rect 16904 -11653 16936 -11651
rect 17064 -11623 17096 -11621
rect 17064 -11651 17066 -11623
rect 17066 -11651 17094 -11623
rect 17094 -11651 17096 -11623
rect 17064 -11653 17096 -11651
rect 17224 -11623 17256 -11621
rect 17224 -11651 17226 -11623
rect 17226 -11651 17254 -11623
rect 17254 -11651 17256 -11623
rect 17224 -11653 17256 -11651
rect 17384 -11623 17416 -11621
rect 17384 -11651 17386 -11623
rect 17386 -11651 17414 -11623
rect 17414 -11651 17416 -11623
rect 17384 -11653 17416 -11651
rect 17544 -11623 17576 -11621
rect 17544 -11651 17546 -11623
rect 17546 -11651 17574 -11623
rect 17574 -11651 17576 -11623
rect 17544 -11653 17576 -11651
rect 17704 -11623 17736 -11621
rect 17704 -11651 17706 -11623
rect 17706 -11651 17734 -11623
rect 17734 -11651 17736 -11623
rect 17704 -11653 17736 -11651
rect 17864 -11623 17896 -11621
rect 17864 -11651 17866 -11623
rect 17866 -11651 17894 -11623
rect 17894 -11651 17896 -11623
rect 17864 -11653 17896 -11651
rect 18024 -11623 18056 -11621
rect 18024 -11651 18026 -11623
rect 18026 -11651 18054 -11623
rect 18054 -11651 18056 -11623
rect 18024 -11653 18056 -11651
rect 18184 -11623 18216 -11621
rect 18184 -11651 18186 -11623
rect 18186 -11651 18214 -11623
rect 18214 -11651 18216 -11623
rect 18184 -11653 18216 -11651
rect 18344 -11623 18376 -11621
rect 18344 -11651 18346 -11623
rect 18346 -11651 18374 -11623
rect 18374 -11651 18376 -11623
rect 18344 -11653 18376 -11651
rect 18504 -11623 18536 -11621
rect 18504 -11651 18506 -11623
rect 18506 -11651 18534 -11623
rect 18534 -11651 18536 -11623
rect 18504 -11653 18536 -11651
rect 18664 -11623 18696 -11621
rect 18664 -11651 18666 -11623
rect 18666 -11651 18694 -11623
rect 18694 -11651 18696 -11623
rect 18664 -11653 18696 -11651
rect 15119 -11726 15151 -11724
rect 15119 -11754 15121 -11726
rect 15121 -11754 15149 -11726
rect 15149 -11754 15151 -11726
rect 15119 -11756 15151 -11754
rect 18852 -11726 18884 -11724
rect 18852 -11754 18854 -11726
rect 18854 -11754 18882 -11726
rect 18882 -11754 18884 -11726
rect 18852 -11756 18884 -11754
rect 15119 -11886 15151 -11884
rect 15119 -11914 15121 -11886
rect 15121 -11914 15149 -11886
rect 15149 -11914 15151 -11886
rect 15119 -11916 15151 -11914
rect 15119 -12046 15151 -12044
rect 15119 -12074 15121 -12046
rect 15121 -12074 15149 -12046
rect 15149 -12074 15151 -12046
rect 15119 -12076 15151 -12074
rect 15119 -12206 15151 -12204
rect 15119 -12234 15121 -12206
rect 15121 -12234 15149 -12206
rect 15149 -12234 15151 -12206
rect 15119 -12236 15151 -12234
rect 15119 -12366 15151 -12364
rect 15119 -12394 15121 -12366
rect 15121 -12394 15149 -12366
rect 15149 -12394 15151 -12366
rect 15119 -12396 15151 -12394
rect 15119 -12526 15151 -12524
rect 15119 -12554 15121 -12526
rect 15121 -12554 15149 -12526
rect 15149 -12554 15151 -12526
rect 15119 -12556 15151 -12554
rect 15119 -12686 15151 -12684
rect 15119 -12714 15121 -12686
rect 15121 -12714 15149 -12686
rect 15149 -12714 15151 -12686
rect 15119 -12716 15151 -12714
rect 15119 -12846 15151 -12844
rect 15119 -12874 15121 -12846
rect 15121 -12874 15149 -12846
rect 15149 -12874 15151 -12846
rect 15119 -12876 15151 -12874
rect 12852 -13006 12884 -13004
rect 12852 -13034 12854 -13006
rect 12854 -13034 12882 -13006
rect 12882 -13034 12884 -13006
rect 12852 -13036 12884 -13034
rect 12852 -13166 12884 -13164
rect 12852 -13194 12854 -13166
rect 12854 -13194 12882 -13166
rect 12882 -13194 12884 -13166
rect 12852 -13196 12884 -13194
rect 12852 -13326 12884 -13324
rect 12852 -13354 12854 -13326
rect 12854 -13354 12882 -13326
rect 12882 -13354 12884 -13326
rect 12852 -13356 12884 -13354
rect 12852 -13486 12884 -13484
rect 12852 -13514 12854 -13486
rect 12854 -13514 12882 -13486
rect 12882 -13514 12884 -13486
rect 12852 -13516 12884 -13514
rect 12852 -13646 12884 -13644
rect 12852 -13674 12854 -13646
rect 12854 -13674 12882 -13646
rect 12882 -13674 12884 -13646
rect 12852 -13676 12884 -13674
rect 12852 -13806 12884 -13804
rect 12852 -13834 12854 -13806
rect 12854 -13834 12882 -13806
rect 12882 -13834 12884 -13806
rect 12852 -13836 12884 -13834
rect 12852 -13966 12884 -13964
rect 12852 -13994 12854 -13966
rect 12854 -13994 12882 -13966
rect 12882 -13994 12884 -13966
rect 12852 -13996 12884 -13994
rect 12852 -14126 12884 -14124
rect 12852 -14154 12854 -14126
rect 12854 -14154 12882 -14126
rect 12882 -14154 12884 -14126
rect 12852 -14156 12884 -14154
rect 12852 -14286 12884 -14284
rect 12852 -14314 12854 -14286
rect 12854 -14314 12882 -14286
rect 12882 -14314 12884 -14286
rect 12852 -14316 12884 -14314
rect 12852 -14446 12884 -14444
rect 12852 -14474 12854 -14446
rect 12854 -14474 12882 -14446
rect 12882 -14474 12884 -14446
rect 12852 -14476 12884 -14474
rect 12852 -14606 12884 -14604
rect 12852 -14634 12854 -14606
rect 12854 -14634 12882 -14606
rect 12882 -14634 12884 -14606
rect 12852 -14636 12884 -14634
rect 12852 -14766 12884 -14764
rect 12852 -14794 12854 -14766
rect 12854 -14794 12882 -14766
rect 12882 -14794 12884 -14766
rect 12852 -14796 12884 -14794
rect 12852 -14926 12884 -14924
rect 12852 -14954 12854 -14926
rect 12854 -14954 12882 -14926
rect 12882 -14954 12884 -14926
rect 12852 -14956 12884 -14954
rect 12852 -15086 12884 -15084
rect 12852 -15114 12854 -15086
rect 12854 -15114 12882 -15086
rect 12882 -15114 12884 -15086
rect 12852 -15116 12884 -15114
rect 9119 -15246 9151 -15244
rect 9119 -15274 9121 -15246
rect 9121 -15274 9149 -15246
rect 9149 -15274 9151 -15246
rect 9119 -15276 9151 -15274
rect 12852 -15246 12884 -15244
rect 12852 -15274 12854 -15246
rect 12854 -15274 12882 -15246
rect 12882 -15274 12884 -15246
rect 12852 -15276 12884 -15274
rect 9304 -15351 9336 -15349
rect 9304 -15379 9306 -15351
rect 9306 -15379 9334 -15351
rect 9334 -15379 9336 -15351
rect 9304 -15381 9336 -15379
rect 9464 -15351 9496 -15349
rect 9464 -15379 9466 -15351
rect 9466 -15379 9494 -15351
rect 9494 -15379 9496 -15351
rect 9464 -15381 9496 -15379
rect 9624 -15351 9656 -15349
rect 9624 -15379 9626 -15351
rect 9626 -15379 9654 -15351
rect 9654 -15379 9656 -15351
rect 9624 -15381 9656 -15379
rect 9784 -15351 9816 -15349
rect 9784 -15379 9786 -15351
rect 9786 -15379 9814 -15351
rect 9814 -15379 9816 -15351
rect 9784 -15381 9816 -15379
rect 9944 -15351 9976 -15349
rect 9944 -15379 9946 -15351
rect 9946 -15379 9974 -15351
rect 9974 -15379 9976 -15351
rect 9944 -15381 9976 -15379
rect 10104 -15351 10136 -15349
rect 10104 -15379 10106 -15351
rect 10106 -15379 10134 -15351
rect 10134 -15379 10136 -15351
rect 10104 -15381 10136 -15379
rect 10264 -15351 10296 -15349
rect 10264 -15379 10266 -15351
rect 10266 -15379 10294 -15351
rect 10294 -15379 10296 -15351
rect 10264 -15381 10296 -15379
rect 10424 -15351 10456 -15349
rect 10424 -15379 10426 -15351
rect 10426 -15379 10454 -15351
rect 10454 -15379 10456 -15351
rect 10424 -15381 10456 -15379
rect 10584 -15351 10616 -15349
rect 10584 -15379 10586 -15351
rect 10586 -15379 10614 -15351
rect 10614 -15379 10616 -15351
rect 10584 -15381 10616 -15379
rect 10744 -15351 10776 -15349
rect 10744 -15379 10746 -15351
rect 10746 -15379 10774 -15351
rect 10774 -15379 10776 -15351
rect 10744 -15381 10776 -15379
rect 10904 -15351 10936 -15349
rect 10904 -15379 10906 -15351
rect 10906 -15379 10934 -15351
rect 10934 -15379 10936 -15351
rect 10904 -15381 10936 -15379
rect 11064 -15351 11096 -15349
rect 11064 -15379 11066 -15351
rect 11066 -15379 11094 -15351
rect 11094 -15379 11096 -15351
rect 11064 -15381 11096 -15379
rect 11224 -15351 11256 -15349
rect 11224 -15379 11226 -15351
rect 11226 -15379 11254 -15351
rect 11254 -15379 11256 -15351
rect 11224 -15381 11256 -15379
rect 11384 -15351 11416 -15349
rect 11384 -15379 11386 -15351
rect 11386 -15379 11414 -15351
rect 11414 -15379 11416 -15351
rect 11384 -15381 11416 -15379
rect 11544 -15351 11576 -15349
rect 11544 -15379 11546 -15351
rect 11546 -15379 11574 -15351
rect 11574 -15379 11576 -15351
rect 11544 -15381 11576 -15379
rect 11704 -15351 11736 -15349
rect 11704 -15379 11706 -15351
rect 11706 -15379 11734 -15351
rect 11734 -15379 11736 -15351
rect 11704 -15381 11736 -15379
rect 11864 -15351 11896 -15349
rect 11864 -15379 11866 -15351
rect 11866 -15379 11894 -15351
rect 11894 -15379 11896 -15351
rect 11864 -15381 11896 -15379
rect 12024 -15351 12056 -15349
rect 12024 -15379 12026 -15351
rect 12026 -15379 12054 -15351
rect 12054 -15379 12056 -15351
rect 12024 -15381 12056 -15379
rect 12184 -15351 12216 -15349
rect 12184 -15379 12186 -15351
rect 12186 -15379 12214 -15351
rect 12214 -15379 12216 -15351
rect 12184 -15381 12216 -15379
rect 12344 -15351 12376 -15349
rect 12344 -15379 12346 -15351
rect 12346 -15379 12374 -15351
rect 12374 -15379 12376 -15351
rect 12344 -15381 12376 -15379
rect 12504 -15351 12536 -15349
rect 12504 -15379 12506 -15351
rect 12506 -15379 12534 -15351
rect 12534 -15379 12536 -15351
rect 12504 -15381 12536 -15379
rect 12664 -15351 12696 -15349
rect 12664 -15379 12666 -15351
rect 12666 -15379 12694 -15351
rect 12694 -15379 12696 -15351
rect 12664 -15381 12696 -15379
rect 15119 -13006 15151 -13004
rect 15119 -13034 15121 -13006
rect 15121 -13034 15149 -13006
rect 15149 -13034 15151 -13006
rect 15119 -13036 15151 -13034
rect 15119 -13166 15151 -13164
rect 15119 -13194 15121 -13166
rect 15121 -13194 15149 -13166
rect 15149 -13194 15151 -13166
rect 15119 -13196 15151 -13194
rect 15119 -13326 15151 -13324
rect 15119 -13354 15121 -13326
rect 15121 -13354 15149 -13326
rect 15149 -13354 15151 -13326
rect 15119 -13356 15151 -13354
rect 15119 -13486 15151 -13484
rect 15119 -13514 15121 -13486
rect 15121 -13514 15149 -13486
rect 15149 -13514 15151 -13486
rect 15119 -13516 15151 -13514
rect 15119 -13646 15151 -13644
rect 15119 -13674 15121 -13646
rect 15121 -13674 15149 -13646
rect 15149 -13674 15151 -13646
rect 15119 -13676 15151 -13674
rect 15119 -13806 15151 -13804
rect 15119 -13834 15121 -13806
rect 15121 -13834 15149 -13806
rect 15149 -13834 15151 -13806
rect 15119 -13836 15151 -13834
rect 15119 -13966 15151 -13964
rect 15119 -13994 15121 -13966
rect 15121 -13994 15149 -13966
rect 15149 -13994 15151 -13966
rect 15119 -13996 15151 -13994
rect 15119 -14126 15151 -14124
rect 15119 -14154 15121 -14126
rect 15121 -14154 15149 -14126
rect 15149 -14154 15151 -14126
rect 15119 -14156 15151 -14154
rect 15119 -14286 15151 -14284
rect 15119 -14314 15121 -14286
rect 15121 -14314 15149 -14286
rect 15149 -14314 15151 -14286
rect 15119 -14316 15151 -14314
rect 15119 -14446 15151 -14444
rect 15119 -14474 15121 -14446
rect 15121 -14474 15149 -14446
rect 15149 -14474 15151 -14446
rect 15119 -14476 15151 -14474
rect 15119 -14606 15151 -14604
rect 15119 -14634 15121 -14606
rect 15121 -14634 15149 -14606
rect 15149 -14634 15151 -14606
rect 15119 -14636 15151 -14634
rect 15119 -14766 15151 -14764
rect 15119 -14794 15121 -14766
rect 15121 -14794 15149 -14766
rect 15149 -14794 15151 -14766
rect 15119 -14796 15151 -14794
rect 15119 -14926 15151 -14924
rect 15119 -14954 15121 -14926
rect 15121 -14954 15149 -14926
rect 15149 -14954 15151 -14926
rect 15119 -14956 15151 -14954
rect 15119 -15086 15151 -15084
rect 15119 -15114 15121 -15086
rect 15121 -15114 15149 -15086
rect 15149 -15114 15151 -15086
rect 15119 -15116 15151 -15114
rect 18852 -11886 18884 -11884
rect 18852 -11914 18854 -11886
rect 18854 -11914 18882 -11886
rect 18882 -11914 18884 -11886
rect 18852 -11916 18884 -11914
rect 18852 -12046 18884 -12044
rect 18852 -12074 18854 -12046
rect 18854 -12074 18882 -12046
rect 18882 -12074 18884 -12046
rect 18852 -12076 18884 -12074
rect 18852 -12206 18884 -12204
rect 18852 -12234 18854 -12206
rect 18854 -12234 18882 -12206
rect 18882 -12234 18884 -12206
rect 18852 -12236 18884 -12234
rect 18852 -12366 18884 -12364
rect 18852 -12394 18854 -12366
rect 18854 -12394 18882 -12366
rect 18882 -12394 18884 -12366
rect 18852 -12396 18884 -12394
rect 18852 -12526 18884 -12524
rect 18852 -12554 18854 -12526
rect 18854 -12554 18882 -12526
rect 18882 -12554 18884 -12526
rect 18852 -12556 18884 -12554
rect 18852 -12686 18884 -12684
rect 18852 -12714 18854 -12686
rect 18854 -12714 18882 -12686
rect 18882 -12714 18884 -12686
rect 18852 -12716 18884 -12714
rect 18852 -12846 18884 -12844
rect 18852 -12874 18854 -12846
rect 18854 -12874 18882 -12846
rect 18882 -12874 18884 -12846
rect 18852 -12876 18884 -12874
rect 18852 -13006 18884 -13004
rect 18852 -13034 18854 -13006
rect 18854 -13034 18882 -13006
rect 18882 -13034 18884 -13006
rect 18852 -13036 18884 -13034
rect 18852 -13166 18884 -13164
rect 18852 -13194 18854 -13166
rect 18854 -13194 18882 -13166
rect 18882 -13194 18884 -13166
rect 18852 -13196 18884 -13194
rect 18852 -13326 18884 -13324
rect 18852 -13354 18854 -13326
rect 18854 -13354 18882 -13326
rect 18882 -13354 18884 -13326
rect 18852 -13356 18884 -13354
rect 18852 -13486 18884 -13484
rect 18852 -13514 18854 -13486
rect 18854 -13514 18882 -13486
rect 18882 -13514 18884 -13486
rect 18852 -13516 18884 -13514
rect 18852 -13646 18884 -13644
rect 18852 -13674 18854 -13646
rect 18854 -13674 18882 -13646
rect 18882 -13674 18884 -13646
rect 18852 -13676 18884 -13674
rect 18852 -13806 18884 -13804
rect 18852 -13834 18854 -13806
rect 18854 -13834 18882 -13806
rect 18882 -13834 18884 -13806
rect 18852 -13836 18884 -13834
rect 18852 -13966 18884 -13964
rect 18852 -13994 18854 -13966
rect 18854 -13994 18882 -13966
rect 18882 -13994 18884 -13966
rect 18852 -13996 18884 -13994
rect 18852 -14126 18884 -14124
rect 18852 -14154 18854 -14126
rect 18854 -14154 18882 -14126
rect 18882 -14154 18884 -14126
rect 18852 -14156 18884 -14154
rect 18852 -14286 18884 -14284
rect 18852 -14314 18854 -14286
rect 18854 -14314 18882 -14286
rect 18882 -14314 18884 -14286
rect 18852 -14316 18884 -14314
rect 18852 -14446 18884 -14444
rect 18852 -14474 18854 -14446
rect 18854 -14474 18882 -14446
rect 18882 -14474 18884 -14446
rect 18852 -14476 18884 -14474
rect 18852 -14606 18884 -14604
rect 18852 -14634 18854 -14606
rect 18854 -14634 18882 -14606
rect 18882 -14634 18884 -14606
rect 18852 -14636 18884 -14634
rect 18852 -14766 18884 -14764
rect 18852 -14794 18854 -14766
rect 18854 -14794 18882 -14766
rect 18882 -14794 18884 -14766
rect 18852 -14796 18884 -14794
rect 18852 -14926 18884 -14924
rect 18852 -14954 18854 -14926
rect 18854 -14954 18882 -14926
rect 18882 -14954 18884 -14926
rect 18852 -14956 18884 -14954
rect 18852 -15086 18884 -15084
rect 18852 -15114 18854 -15086
rect 18854 -15114 18882 -15086
rect 18882 -15114 18884 -15086
rect 18852 -15116 18884 -15114
rect 15119 -15246 15151 -15244
rect 15119 -15274 15121 -15246
rect 15121 -15274 15149 -15246
rect 15149 -15274 15151 -15246
rect 15119 -15276 15151 -15274
rect 18852 -15246 18884 -15244
rect 18852 -15274 18854 -15246
rect 18854 -15274 18882 -15246
rect 18882 -15274 18884 -15246
rect 18852 -15276 18884 -15274
rect 15304 -15351 15336 -15349
rect 15304 -15379 15306 -15351
rect 15306 -15379 15334 -15351
rect 15334 -15379 15336 -15351
rect 15304 -15381 15336 -15379
rect 15464 -15351 15496 -15349
rect 15464 -15379 15466 -15351
rect 15466 -15379 15494 -15351
rect 15494 -15379 15496 -15351
rect 15464 -15381 15496 -15379
rect 15624 -15351 15656 -15349
rect 15624 -15379 15626 -15351
rect 15626 -15379 15654 -15351
rect 15654 -15379 15656 -15351
rect 15624 -15381 15656 -15379
rect 15784 -15351 15816 -15349
rect 15784 -15379 15786 -15351
rect 15786 -15379 15814 -15351
rect 15814 -15379 15816 -15351
rect 15784 -15381 15816 -15379
rect 15944 -15351 15976 -15349
rect 15944 -15379 15946 -15351
rect 15946 -15379 15974 -15351
rect 15974 -15379 15976 -15351
rect 15944 -15381 15976 -15379
rect 16104 -15351 16136 -15349
rect 16104 -15379 16106 -15351
rect 16106 -15379 16134 -15351
rect 16134 -15379 16136 -15351
rect 16104 -15381 16136 -15379
rect 16264 -15351 16296 -15349
rect 16264 -15379 16266 -15351
rect 16266 -15379 16294 -15351
rect 16294 -15379 16296 -15351
rect 16264 -15381 16296 -15379
rect 16424 -15351 16456 -15349
rect 16424 -15379 16426 -15351
rect 16426 -15379 16454 -15351
rect 16454 -15379 16456 -15351
rect 16424 -15381 16456 -15379
rect 16584 -15351 16616 -15349
rect 16584 -15379 16586 -15351
rect 16586 -15379 16614 -15351
rect 16614 -15379 16616 -15351
rect 16584 -15381 16616 -15379
rect 16744 -15351 16776 -15349
rect 16744 -15379 16746 -15351
rect 16746 -15379 16774 -15351
rect 16774 -15379 16776 -15351
rect 16744 -15381 16776 -15379
rect 16904 -15351 16936 -15349
rect 16904 -15379 16906 -15351
rect 16906 -15379 16934 -15351
rect 16934 -15379 16936 -15351
rect 16904 -15381 16936 -15379
rect 17064 -15351 17096 -15349
rect 17064 -15379 17066 -15351
rect 17066 -15379 17094 -15351
rect 17094 -15379 17096 -15351
rect 17064 -15381 17096 -15379
rect 17224 -15351 17256 -15349
rect 17224 -15379 17226 -15351
rect 17226 -15379 17254 -15351
rect 17254 -15379 17256 -15351
rect 17224 -15381 17256 -15379
rect 17384 -15351 17416 -15349
rect 17384 -15379 17386 -15351
rect 17386 -15379 17414 -15351
rect 17414 -15379 17416 -15351
rect 17384 -15381 17416 -15379
rect 17544 -15351 17576 -15349
rect 17544 -15379 17546 -15351
rect 17546 -15379 17574 -15351
rect 17574 -15379 17576 -15351
rect 17544 -15381 17576 -15379
rect 17704 -15351 17736 -15349
rect 17704 -15379 17706 -15351
rect 17706 -15379 17734 -15351
rect 17734 -15379 17736 -15351
rect 17704 -15381 17736 -15379
rect 17864 -15351 17896 -15349
rect 17864 -15379 17866 -15351
rect 17866 -15379 17894 -15351
rect 17894 -15379 17896 -15351
rect 17864 -15381 17896 -15379
rect 18024 -15351 18056 -15349
rect 18024 -15379 18026 -15351
rect 18026 -15379 18054 -15351
rect 18054 -15379 18056 -15351
rect 18024 -15381 18056 -15379
rect 18184 -15351 18216 -15349
rect 18184 -15379 18186 -15351
rect 18186 -15379 18214 -15351
rect 18214 -15379 18216 -15351
rect 18184 -15381 18216 -15379
rect 18344 -15351 18376 -15349
rect 18344 -15379 18346 -15351
rect 18346 -15379 18374 -15351
rect 18374 -15379 18376 -15351
rect 18344 -15381 18376 -15379
rect 18504 -15351 18536 -15349
rect 18504 -15379 18506 -15351
rect 18506 -15379 18534 -15351
rect 18534 -15379 18536 -15351
rect 18504 -15381 18536 -15379
rect 18664 -15351 18696 -15349
rect 18664 -15379 18666 -15351
rect 18666 -15379 18694 -15351
rect 18694 -15379 18696 -15351
rect 18664 -15381 18696 -15379
rect 21304 -11623 21336 -11621
rect 21304 -11651 21306 -11623
rect 21306 -11651 21334 -11623
rect 21334 -11651 21336 -11623
rect 21304 -11653 21336 -11651
rect 21464 -11623 21496 -11621
rect 21464 -11651 21466 -11623
rect 21466 -11651 21494 -11623
rect 21494 -11651 21496 -11623
rect 21464 -11653 21496 -11651
rect 21624 -11623 21656 -11621
rect 21624 -11651 21626 -11623
rect 21626 -11651 21654 -11623
rect 21654 -11651 21656 -11623
rect 21624 -11653 21656 -11651
rect 21784 -11623 21816 -11621
rect 21784 -11651 21786 -11623
rect 21786 -11651 21814 -11623
rect 21814 -11651 21816 -11623
rect 21784 -11653 21816 -11651
rect 21944 -11623 21976 -11621
rect 21944 -11651 21946 -11623
rect 21946 -11651 21974 -11623
rect 21974 -11651 21976 -11623
rect 21944 -11653 21976 -11651
rect 22104 -11623 22136 -11621
rect 22104 -11651 22106 -11623
rect 22106 -11651 22134 -11623
rect 22134 -11651 22136 -11623
rect 22104 -11653 22136 -11651
rect 22264 -11623 22296 -11621
rect 22264 -11651 22266 -11623
rect 22266 -11651 22294 -11623
rect 22294 -11651 22296 -11623
rect 22264 -11653 22296 -11651
rect 22424 -11623 22456 -11621
rect 22424 -11651 22426 -11623
rect 22426 -11651 22454 -11623
rect 22454 -11651 22456 -11623
rect 22424 -11653 22456 -11651
rect 22584 -11623 22616 -11621
rect 22584 -11651 22586 -11623
rect 22586 -11651 22614 -11623
rect 22614 -11651 22616 -11623
rect 22584 -11653 22616 -11651
rect 22744 -11623 22776 -11621
rect 22744 -11651 22746 -11623
rect 22746 -11651 22774 -11623
rect 22774 -11651 22776 -11623
rect 22744 -11653 22776 -11651
rect 22904 -11623 22936 -11621
rect 22904 -11651 22906 -11623
rect 22906 -11651 22934 -11623
rect 22934 -11651 22936 -11623
rect 22904 -11653 22936 -11651
rect 23064 -11623 23096 -11621
rect 23064 -11651 23066 -11623
rect 23066 -11651 23094 -11623
rect 23094 -11651 23096 -11623
rect 23064 -11653 23096 -11651
rect 23224 -11623 23256 -11621
rect 23224 -11651 23226 -11623
rect 23226 -11651 23254 -11623
rect 23254 -11651 23256 -11623
rect 23224 -11653 23256 -11651
rect 23384 -11623 23416 -11621
rect 23384 -11651 23386 -11623
rect 23386 -11651 23414 -11623
rect 23414 -11651 23416 -11623
rect 23384 -11653 23416 -11651
rect 23544 -11623 23576 -11621
rect 23544 -11651 23546 -11623
rect 23546 -11651 23574 -11623
rect 23574 -11651 23576 -11623
rect 23544 -11653 23576 -11651
rect 23704 -11623 23736 -11621
rect 23704 -11651 23706 -11623
rect 23706 -11651 23734 -11623
rect 23734 -11651 23736 -11623
rect 23704 -11653 23736 -11651
rect 23864 -11623 23896 -11621
rect 23864 -11651 23866 -11623
rect 23866 -11651 23894 -11623
rect 23894 -11651 23896 -11623
rect 23864 -11653 23896 -11651
rect 24024 -11623 24056 -11621
rect 24024 -11651 24026 -11623
rect 24026 -11651 24054 -11623
rect 24054 -11651 24056 -11623
rect 24024 -11653 24056 -11651
rect 24184 -11623 24216 -11621
rect 24184 -11651 24186 -11623
rect 24186 -11651 24214 -11623
rect 24214 -11651 24216 -11623
rect 24184 -11653 24216 -11651
rect 24344 -11623 24376 -11621
rect 24344 -11651 24346 -11623
rect 24346 -11651 24374 -11623
rect 24374 -11651 24376 -11623
rect 24344 -11653 24376 -11651
rect 24504 -11623 24536 -11621
rect 24504 -11651 24506 -11623
rect 24506 -11651 24534 -11623
rect 24534 -11651 24536 -11623
rect 24504 -11653 24536 -11651
rect 24664 -11623 24696 -11621
rect 24664 -11651 24666 -11623
rect 24666 -11651 24694 -11623
rect 24694 -11651 24696 -11623
rect 24664 -11653 24696 -11651
rect 21119 -11726 21151 -11724
rect 21119 -11754 21121 -11726
rect 21121 -11754 21149 -11726
rect 21149 -11754 21151 -11726
rect 21119 -11756 21151 -11754
rect 24852 -11726 24884 -11724
rect 24852 -11754 24854 -11726
rect 24854 -11754 24882 -11726
rect 24882 -11754 24884 -11726
rect 24852 -11756 24884 -11754
rect 21119 -11886 21151 -11884
rect 21119 -11914 21121 -11886
rect 21121 -11914 21149 -11886
rect 21149 -11914 21151 -11886
rect 21119 -11916 21151 -11914
rect 21119 -12046 21151 -12044
rect 21119 -12074 21121 -12046
rect 21121 -12074 21149 -12046
rect 21149 -12074 21151 -12046
rect 21119 -12076 21151 -12074
rect 21119 -12206 21151 -12204
rect 21119 -12234 21121 -12206
rect 21121 -12234 21149 -12206
rect 21149 -12234 21151 -12206
rect 21119 -12236 21151 -12234
rect 21119 -12366 21151 -12364
rect 21119 -12394 21121 -12366
rect 21121 -12394 21149 -12366
rect 21149 -12394 21151 -12366
rect 21119 -12396 21151 -12394
rect 21119 -12526 21151 -12524
rect 21119 -12554 21121 -12526
rect 21121 -12554 21149 -12526
rect 21149 -12554 21151 -12526
rect 21119 -12556 21151 -12554
rect 21119 -12686 21151 -12684
rect 21119 -12714 21121 -12686
rect 21121 -12714 21149 -12686
rect 21149 -12714 21151 -12686
rect 21119 -12716 21151 -12714
rect 21119 -12846 21151 -12844
rect 21119 -12874 21121 -12846
rect 21121 -12874 21149 -12846
rect 21149 -12874 21151 -12846
rect 21119 -12876 21151 -12874
rect 21119 -13006 21151 -13004
rect 21119 -13034 21121 -13006
rect 21121 -13034 21149 -13006
rect 21149 -13034 21151 -13006
rect 21119 -13036 21151 -13034
rect 21119 -13166 21151 -13164
rect 21119 -13194 21121 -13166
rect 21121 -13194 21149 -13166
rect 21149 -13194 21151 -13166
rect 21119 -13196 21151 -13194
rect 21119 -13326 21151 -13324
rect 21119 -13354 21121 -13326
rect 21121 -13354 21149 -13326
rect 21149 -13354 21151 -13326
rect 21119 -13356 21151 -13354
rect 21119 -13486 21151 -13484
rect 21119 -13514 21121 -13486
rect 21121 -13514 21149 -13486
rect 21149 -13514 21151 -13486
rect 21119 -13516 21151 -13514
rect 21119 -13646 21151 -13644
rect 21119 -13674 21121 -13646
rect 21121 -13674 21149 -13646
rect 21149 -13674 21151 -13646
rect 21119 -13676 21151 -13674
rect 21119 -13806 21151 -13804
rect 21119 -13834 21121 -13806
rect 21121 -13834 21149 -13806
rect 21149 -13834 21151 -13806
rect 21119 -13836 21151 -13834
rect 21119 -13966 21151 -13964
rect 21119 -13994 21121 -13966
rect 21121 -13994 21149 -13966
rect 21149 -13994 21151 -13966
rect 21119 -13996 21151 -13994
rect 21119 -14126 21151 -14124
rect 21119 -14154 21121 -14126
rect 21121 -14154 21149 -14126
rect 21149 -14154 21151 -14126
rect 21119 -14156 21151 -14154
rect 21119 -14286 21151 -14284
rect 21119 -14314 21121 -14286
rect 21121 -14314 21149 -14286
rect 21149 -14314 21151 -14286
rect 21119 -14316 21151 -14314
rect 21119 -14446 21151 -14444
rect 21119 -14474 21121 -14446
rect 21121 -14474 21149 -14446
rect 21149 -14474 21151 -14446
rect 21119 -14476 21151 -14474
rect 21119 -14606 21151 -14604
rect 21119 -14634 21121 -14606
rect 21121 -14634 21149 -14606
rect 21149 -14634 21151 -14606
rect 21119 -14636 21151 -14634
rect 21119 -14766 21151 -14764
rect 21119 -14794 21121 -14766
rect 21121 -14794 21149 -14766
rect 21149 -14794 21151 -14766
rect 21119 -14796 21151 -14794
rect 21119 -14926 21151 -14924
rect 21119 -14954 21121 -14926
rect 21121 -14954 21149 -14926
rect 21149 -14954 21151 -14926
rect 21119 -14956 21151 -14954
rect 21119 -15086 21151 -15084
rect 21119 -15114 21121 -15086
rect 21121 -15114 21149 -15086
rect 21149 -15114 21151 -15086
rect 21119 -15116 21151 -15114
rect 24852 -11886 24884 -11884
rect 24852 -11914 24854 -11886
rect 24854 -11914 24882 -11886
rect 24882 -11914 24884 -11886
rect 24852 -11916 24884 -11914
rect 24852 -12046 24884 -12044
rect 24852 -12074 24854 -12046
rect 24854 -12074 24882 -12046
rect 24882 -12074 24884 -12046
rect 24852 -12076 24884 -12074
rect 24852 -12206 24884 -12204
rect 24852 -12234 24854 -12206
rect 24854 -12234 24882 -12206
rect 24882 -12234 24884 -12206
rect 24852 -12236 24884 -12234
rect 24852 -12366 24884 -12364
rect 24852 -12394 24854 -12366
rect 24854 -12394 24882 -12366
rect 24882 -12394 24884 -12366
rect 24852 -12396 24884 -12394
rect 24852 -12526 24884 -12524
rect 24852 -12554 24854 -12526
rect 24854 -12554 24882 -12526
rect 24882 -12554 24884 -12526
rect 24852 -12556 24884 -12554
rect 24852 -12686 24884 -12684
rect 24852 -12714 24854 -12686
rect 24854 -12714 24882 -12686
rect 24882 -12714 24884 -12686
rect 24852 -12716 24884 -12714
rect 24852 -12846 24884 -12844
rect 24852 -12874 24854 -12846
rect 24854 -12874 24882 -12846
rect 24882 -12874 24884 -12846
rect 24852 -12876 24884 -12874
rect 24852 -13006 24884 -13004
rect 24852 -13034 24854 -13006
rect 24854 -13034 24882 -13006
rect 24882 -13034 24884 -13006
rect 24852 -13036 24884 -13034
rect 24852 -13166 24884 -13164
rect 24852 -13194 24854 -13166
rect 24854 -13194 24882 -13166
rect 24882 -13194 24884 -13166
rect 24852 -13196 24884 -13194
rect 24852 -13326 24884 -13324
rect 24852 -13354 24854 -13326
rect 24854 -13354 24882 -13326
rect 24882 -13354 24884 -13326
rect 24852 -13356 24884 -13354
rect 24852 -13486 24884 -13484
rect 24852 -13514 24854 -13486
rect 24854 -13514 24882 -13486
rect 24882 -13514 24884 -13486
rect 24852 -13516 24884 -13514
rect 24852 -13646 24884 -13644
rect 24852 -13674 24854 -13646
rect 24854 -13674 24882 -13646
rect 24882 -13674 24884 -13646
rect 24852 -13676 24884 -13674
rect 24852 -13806 24884 -13804
rect 24852 -13834 24854 -13806
rect 24854 -13834 24882 -13806
rect 24882 -13834 24884 -13806
rect 24852 -13836 24884 -13834
rect 24852 -13966 24884 -13964
rect 24852 -13994 24854 -13966
rect 24854 -13994 24882 -13966
rect 24882 -13994 24884 -13966
rect 24852 -13996 24884 -13994
rect 24852 -14126 24884 -14124
rect 24852 -14154 24854 -14126
rect 24854 -14154 24882 -14126
rect 24882 -14154 24884 -14126
rect 24852 -14156 24884 -14154
rect 24852 -14286 24884 -14284
rect 24852 -14314 24854 -14286
rect 24854 -14314 24882 -14286
rect 24882 -14314 24884 -14286
rect 24852 -14316 24884 -14314
rect 24852 -14446 24884 -14444
rect 24852 -14474 24854 -14446
rect 24854 -14474 24882 -14446
rect 24882 -14474 24884 -14446
rect 24852 -14476 24884 -14474
rect 24852 -14606 24884 -14604
rect 24852 -14634 24854 -14606
rect 24854 -14634 24882 -14606
rect 24882 -14634 24884 -14606
rect 24852 -14636 24884 -14634
rect 24852 -14766 24884 -14764
rect 24852 -14794 24854 -14766
rect 24854 -14794 24882 -14766
rect 24882 -14794 24884 -14766
rect 24852 -14796 24884 -14794
rect 24852 -14926 24884 -14924
rect 24852 -14954 24854 -14926
rect 24854 -14954 24882 -14926
rect 24882 -14954 24884 -14926
rect 24852 -14956 24884 -14954
rect 24852 -15086 24884 -15084
rect 24852 -15114 24854 -15086
rect 24854 -15114 24882 -15086
rect 24882 -15114 24884 -15086
rect 24852 -15116 24884 -15114
rect 21119 -15246 21151 -15244
rect 21119 -15274 21121 -15246
rect 21121 -15274 21149 -15246
rect 21149 -15274 21151 -15246
rect 21119 -15276 21151 -15274
rect 24852 -15246 24884 -15244
rect 24852 -15274 24854 -15246
rect 24854 -15274 24882 -15246
rect 24882 -15274 24884 -15246
rect 24852 -15276 24884 -15274
rect 21304 -15351 21336 -15349
rect 21304 -15379 21306 -15351
rect 21306 -15379 21334 -15351
rect 21334 -15379 21336 -15351
rect 21304 -15381 21336 -15379
rect 21464 -15351 21496 -15349
rect 21464 -15379 21466 -15351
rect 21466 -15379 21494 -15351
rect 21494 -15379 21496 -15351
rect 21464 -15381 21496 -15379
rect 21624 -15351 21656 -15349
rect 21624 -15379 21626 -15351
rect 21626 -15379 21654 -15351
rect 21654 -15379 21656 -15351
rect 21624 -15381 21656 -15379
rect 21784 -15351 21816 -15349
rect 21784 -15379 21786 -15351
rect 21786 -15379 21814 -15351
rect 21814 -15379 21816 -15351
rect 21784 -15381 21816 -15379
rect 21944 -15351 21976 -15349
rect 21944 -15379 21946 -15351
rect 21946 -15379 21974 -15351
rect 21974 -15379 21976 -15351
rect 21944 -15381 21976 -15379
rect 22104 -15351 22136 -15349
rect 22104 -15379 22106 -15351
rect 22106 -15379 22134 -15351
rect 22134 -15379 22136 -15351
rect 22104 -15381 22136 -15379
rect 22264 -15351 22296 -15349
rect 22264 -15379 22266 -15351
rect 22266 -15379 22294 -15351
rect 22294 -15379 22296 -15351
rect 22264 -15381 22296 -15379
rect 22424 -15351 22456 -15349
rect 22424 -15379 22426 -15351
rect 22426 -15379 22454 -15351
rect 22454 -15379 22456 -15351
rect 22424 -15381 22456 -15379
rect 22584 -15351 22616 -15349
rect 22584 -15379 22586 -15351
rect 22586 -15379 22614 -15351
rect 22614 -15379 22616 -15351
rect 22584 -15381 22616 -15379
rect 22744 -15351 22776 -15349
rect 22744 -15379 22746 -15351
rect 22746 -15379 22774 -15351
rect 22774 -15379 22776 -15351
rect 22744 -15381 22776 -15379
rect 22904 -15351 22936 -15349
rect 22904 -15379 22906 -15351
rect 22906 -15379 22934 -15351
rect 22934 -15379 22936 -15351
rect 22904 -15381 22936 -15379
rect 23064 -15351 23096 -15349
rect 23064 -15379 23066 -15351
rect 23066 -15379 23094 -15351
rect 23094 -15379 23096 -15351
rect 23064 -15381 23096 -15379
rect 23224 -15351 23256 -15349
rect 23224 -15379 23226 -15351
rect 23226 -15379 23254 -15351
rect 23254 -15379 23256 -15351
rect 23224 -15381 23256 -15379
rect 23384 -15351 23416 -15349
rect 23384 -15379 23386 -15351
rect 23386 -15379 23414 -15351
rect 23414 -15379 23416 -15351
rect 23384 -15381 23416 -15379
rect 23544 -15351 23576 -15349
rect 23544 -15379 23546 -15351
rect 23546 -15379 23574 -15351
rect 23574 -15379 23576 -15351
rect 23544 -15381 23576 -15379
rect 23704 -15351 23736 -15349
rect 23704 -15379 23706 -15351
rect 23706 -15379 23734 -15351
rect 23734 -15379 23736 -15351
rect 23704 -15381 23736 -15379
rect 23864 -15351 23896 -15349
rect 23864 -15379 23866 -15351
rect 23866 -15379 23894 -15351
rect 23894 -15379 23896 -15351
rect 23864 -15381 23896 -15379
rect 24024 -15351 24056 -15349
rect 24024 -15379 24026 -15351
rect 24026 -15379 24054 -15351
rect 24054 -15379 24056 -15351
rect 24024 -15381 24056 -15379
rect 24184 -15351 24216 -15349
rect 24184 -15379 24186 -15351
rect 24186 -15379 24214 -15351
rect 24214 -15379 24216 -15351
rect 24184 -15381 24216 -15379
rect 24344 -15351 24376 -15349
rect 24344 -15379 24346 -15351
rect 24346 -15379 24374 -15351
rect 24374 -15379 24376 -15351
rect 24344 -15381 24376 -15379
rect 24504 -15351 24536 -15349
rect 24504 -15379 24506 -15351
rect 24506 -15379 24534 -15351
rect 24534 -15379 24536 -15351
rect 24504 -15381 24536 -15379
rect 24664 -15351 24696 -15349
rect 24664 -15379 24666 -15351
rect 24666 -15379 24694 -15351
rect 24694 -15379 24696 -15351
rect 24664 -15381 24696 -15379
<< metal4 >>
rect 11750 -2770 12450 -2750
rect 11065 -2800 12450 -2770
rect 11750 -2850 12450 -2800
rect 5500 -4550 6600 -3950
rect 5500 -5500 6150 -4550
rect 12350 -5150 12450 -2850
rect 9000 -5500 11100 -5150
rect 12350 -5250 13550 -5150
rect 13450 -5350 13550 -5250
rect 13450 -5450 19350 -5350
rect 3000 -5578 7000 -5500
rect 3000 -5681 3261 -5578
rect 3000 -5799 3076 -5681
rect 3194 -5696 3261 -5681
rect 3379 -5696 3421 -5578
rect 3539 -5696 3581 -5578
rect 3699 -5696 3741 -5578
rect 3859 -5696 3901 -5578
rect 4019 -5696 4061 -5578
rect 4179 -5696 4221 -5578
rect 4339 -5696 4381 -5578
rect 4499 -5696 4541 -5578
rect 4659 -5696 4701 -5578
rect 4819 -5696 4861 -5578
rect 4979 -5696 5021 -5578
rect 5139 -5696 5181 -5578
rect 5299 -5696 5341 -5578
rect 5459 -5696 5501 -5578
rect 5619 -5696 5661 -5578
rect 5779 -5696 5821 -5578
rect 5939 -5696 5981 -5578
rect 6099 -5696 6141 -5578
rect 6259 -5696 6301 -5578
rect 6419 -5696 6461 -5578
rect 6579 -5696 6621 -5578
rect 6739 -5681 7000 -5578
rect 6739 -5696 6809 -5681
rect 3194 -5770 6809 -5696
rect 3194 -5799 3270 -5770
rect 3000 -5841 3270 -5799
rect 3000 -5959 3076 -5841
rect 3194 -5959 3270 -5841
rect 3000 -6001 3270 -5959
rect 3000 -6119 3076 -6001
rect 3194 -6119 3270 -6001
rect 3000 -6161 3270 -6119
rect 3000 -6279 3076 -6161
rect 3194 -6279 3270 -6161
rect 3000 -6321 3270 -6279
rect 3000 -6439 3076 -6321
rect 3194 -6439 3270 -6321
rect 3000 -6481 3270 -6439
rect 3000 -6599 3076 -6481
rect 3194 -6599 3270 -6481
rect 3000 -6641 3270 -6599
rect 3000 -6759 3076 -6641
rect 3194 -6759 3270 -6641
rect 3000 -6801 3270 -6759
rect 3000 -6919 3076 -6801
rect 3194 -6919 3270 -6801
rect 3000 -6961 3270 -6919
rect 3000 -7079 3076 -6961
rect 3194 -7079 3270 -6961
rect 3000 -7121 3270 -7079
rect 3000 -7239 3076 -7121
rect 3194 -7239 3270 -7121
rect 3000 -7281 3270 -7239
rect 3000 -7399 3076 -7281
rect 3194 -7399 3270 -7281
rect 3000 -7441 3270 -7399
rect 3000 -7559 3076 -7441
rect 3194 -7559 3270 -7441
rect 3000 -7601 3270 -7559
rect 3000 -7719 3076 -7601
rect 3194 -7719 3270 -7601
rect 3000 -7761 3270 -7719
rect 3000 -7879 3076 -7761
rect 3194 -7879 3270 -7761
rect 3000 -7921 3270 -7879
rect 3000 -8039 3076 -7921
rect 3194 -8039 3270 -7921
rect 3000 -8081 3270 -8039
rect 3000 -8199 3076 -8081
rect 3194 -8199 3270 -8081
rect 3000 -8241 3270 -8199
rect 3000 -8359 3076 -8241
rect 3194 -8359 3270 -8241
rect 3000 -8401 3270 -8359
rect 3000 -8519 3076 -8401
rect 3194 -8519 3270 -8401
rect 3000 -8561 3270 -8519
rect 3000 -8679 3076 -8561
rect 3194 -8679 3270 -8561
rect 3000 -8721 3270 -8679
rect 3000 -8839 3076 -8721
rect 3194 -8839 3270 -8721
rect 3000 -8881 3270 -8839
rect 3000 -8999 3076 -8881
rect 3194 -8999 3270 -8881
rect 3000 -9041 3270 -8999
rect 3000 -9159 3076 -9041
rect 3194 -9159 3270 -9041
rect 3000 -9201 3270 -9159
rect 3000 -9319 3076 -9201
rect 3194 -9230 3270 -9201
rect 6730 -5799 6809 -5770
rect 6927 -5799 7000 -5681
rect 6730 -5841 7000 -5799
rect 6730 -5959 6809 -5841
rect 6927 -5959 7000 -5841
rect 6730 -6001 7000 -5959
rect 6730 -6119 6809 -6001
rect 6927 -6119 7000 -6001
rect 6730 -6161 7000 -6119
rect 6730 -6279 6809 -6161
rect 6927 -6279 7000 -6161
rect 6730 -6321 7000 -6279
rect 6730 -6439 6809 -6321
rect 6927 -6439 7000 -6321
rect 6730 -6481 7000 -6439
rect 6730 -6599 6809 -6481
rect 6927 -6599 7000 -6481
rect 6730 -6641 7000 -6599
rect 6730 -6759 6809 -6641
rect 6927 -6759 7000 -6641
rect 6730 -6801 7000 -6759
rect 6730 -6919 6809 -6801
rect 6927 -6919 7000 -6801
rect 6730 -6961 7000 -6919
rect 6730 -7079 6809 -6961
rect 6927 -7079 7000 -6961
rect 6730 -7121 7000 -7079
rect 6730 -7239 6809 -7121
rect 6927 -7239 7000 -7121
rect 6730 -7281 7000 -7239
rect 6730 -7399 6809 -7281
rect 6927 -7399 7000 -7281
rect 6730 -7441 7000 -7399
rect 6730 -7559 6809 -7441
rect 6927 -7559 7000 -7441
rect 6730 -7601 7000 -7559
rect 6730 -7719 6809 -7601
rect 6927 -7719 7000 -7601
rect 6730 -7761 7000 -7719
rect 6730 -7879 6809 -7761
rect 6927 -7879 7000 -7761
rect 6730 -7921 7000 -7879
rect 6730 -8039 6809 -7921
rect 6927 -8039 7000 -7921
rect 6730 -8081 7000 -8039
rect 6730 -8199 6809 -8081
rect 6927 -8199 7000 -8081
rect 6730 -8241 7000 -8199
rect 6730 -8359 6809 -8241
rect 6927 -8359 7000 -8241
rect 6730 -8401 7000 -8359
rect 6730 -8519 6809 -8401
rect 6927 -8519 7000 -8401
rect 6730 -8561 7000 -8519
rect 6730 -8679 6809 -8561
rect 6927 -8679 7000 -8561
rect 6730 -8721 7000 -8679
rect 6730 -8839 6809 -8721
rect 6927 -8839 7000 -8721
rect 6730 -8881 7000 -8839
rect 6730 -8999 6809 -8881
rect 6927 -8999 7000 -8881
rect 6730 -9041 7000 -8999
rect 6730 -9159 6809 -9041
rect 6927 -9159 7000 -9041
rect 6730 -9201 7000 -9159
rect 6730 -9230 6809 -9201
rect 3194 -9306 6809 -9230
rect 3194 -9319 3261 -9306
rect 3000 -9424 3261 -9319
rect 3379 -9424 3421 -9306
rect 3539 -9424 3581 -9306
rect 3699 -9424 3741 -9306
rect 3859 -9424 3901 -9306
rect 4019 -9424 4061 -9306
rect 4179 -9424 4221 -9306
rect 4339 -9424 4381 -9306
rect 4499 -9424 4541 -9306
rect 4659 -9424 4701 -9306
rect 4819 -9424 4861 -9306
rect 4979 -9424 5021 -9306
rect 5139 -9424 5181 -9306
rect 5299 -9424 5341 -9306
rect 5459 -9424 5501 -9306
rect 5619 -9424 5661 -9306
rect 5779 -9424 5821 -9306
rect 5939 -9424 5981 -9306
rect 6099 -9424 6141 -9306
rect 6259 -9424 6301 -9306
rect 6419 -9424 6461 -9306
rect 6579 -9424 6621 -9306
rect 6739 -9319 6809 -9306
rect 6927 -9319 7000 -9201
rect 6739 -9424 7000 -9319
rect 3000 -9500 7000 -9424
rect 9000 -5578 13000 -5500
rect 9000 -5681 9261 -5578
rect 9000 -5799 9076 -5681
rect 9194 -5696 9261 -5681
rect 9379 -5696 9421 -5578
rect 9539 -5696 9581 -5578
rect 9699 -5696 9741 -5578
rect 9859 -5696 9901 -5578
rect 10019 -5696 10061 -5578
rect 10179 -5696 10221 -5578
rect 10339 -5696 10381 -5578
rect 10499 -5696 10541 -5578
rect 10659 -5696 10701 -5578
rect 10819 -5696 10861 -5578
rect 10979 -5696 11021 -5578
rect 11139 -5696 11181 -5578
rect 11299 -5696 11341 -5578
rect 11459 -5696 11501 -5578
rect 11619 -5696 11661 -5578
rect 11779 -5696 11821 -5578
rect 11939 -5696 11981 -5578
rect 12099 -5696 12141 -5578
rect 12259 -5696 12301 -5578
rect 12419 -5696 12461 -5578
rect 12579 -5696 12621 -5578
rect 12739 -5681 13000 -5578
rect 12739 -5696 12809 -5681
rect 9194 -5770 12809 -5696
rect 9194 -5799 9270 -5770
rect 9000 -5841 9270 -5799
rect 9000 -5959 9076 -5841
rect 9194 -5959 9270 -5841
rect 9000 -6001 9270 -5959
rect 9000 -6119 9076 -6001
rect 9194 -6119 9270 -6001
rect 9000 -6161 9270 -6119
rect 9000 -6279 9076 -6161
rect 9194 -6279 9270 -6161
rect 9000 -6321 9270 -6279
rect 9000 -6439 9076 -6321
rect 9194 -6439 9270 -6321
rect 9000 -6481 9270 -6439
rect 9000 -6599 9076 -6481
rect 9194 -6599 9270 -6481
rect 9000 -6641 9270 -6599
rect 9000 -6759 9076 -6641
rect 9194 -6759 9270 -6641
rect 9000 -6801 9270 -6759
rect 9000 -6919 9076 -6801
rect 9194 -6919 9270 -6801
rect 9000 -6961 9270 -6919
rect 9000 -7079 9076 -6961
rect 9194 -7079 9270 -6961
rect 9000 -7121 9270 -7079
rect 9000 -7239 9076 -7121
rect 9194 -7239 9270 -7121
rect 9000 -7281 9270 -7239
rect 9000 -7399 9076 -7281
rect 9194 -7399 9270 -7281
rect 9000 -7441 9270 -7399
rect 9000 -7559 9076 -7441
rect 9194 -7559 9270 -7441
rect 9000 -7601 9270 -7559
rect 9000 -7719 9076 -7601
rect 9194 -7719 9270 -7601
rect 9000 -7761 9270 -7719
rect 9000 -7879 9076 -7761
rect 9194 -7879 9270 -7761
rect 9000 -7921 9270 -7879
rect 9000 -8039 9076 -7921
rect 9194 -8039 9270 -7921
rect 9000 -8081 9270 -8039
rect 9000 -8199 9076 -8081
rect 9194 -8199 9270 -8081
rect 9000 -8241 9270 -8199
rect 9000 -8359 9076 -8241
rect 9194 -8359 9270 -8241
rect 9000 -8401 9270 -8359
rect 9000 -8519 9076 -8401
rect 9194 -8519 9270 -8401
rect 9000 -8561 9270 -8519
rect 9000 -8679 9076 -8561
rect 9194 -8679 9270 -8561
rect 9000 -8721 9270 -8679
rect 9000 -8839 9076 -8721
rect 9194 -8839 9270 -8721
rect 9000 -8881 9270 -8839
rect 9000 -8999 9076 -8881
rect 9194 -8999 9270 -8881
rect 9000 -9041 9270 -8999
rect 9000 -9159 9076 -9041
rect 9194 -9159 9270 -9041
rect 9000 -9201 9270 -9159
rect 9000 -9319 9076 -9201
rect 9194 -9230 9270 -9201
rect 12730 -5799 12809 -5770
rect 12927 -5799 13000 -5681
rect 12730 -5841 13000 -5799
rect 12730 -5959 12809 -5841
rect 12927 -5959 13000 -5841
rect 12730 -6001 13000 -5959
rect 12730 -6119 12809 -6001
rect 12927 -6119 13000 -6001
rect 12730 -6161 13000 -6119
rect 12730 -6279 12809 -6161
rect 12927 -6279 13000 -6161
rect 12730 -6321 13000 -6279
rect 12730 -6439 12809 -6321
rect 12927 -6439 13000 -6321
rect 12730 -6481 13000 -6439
rect 12730 -6599 12809 -6481
rect 12927 -6599 13000 -6481
rect 12730 -6641 13000 -6599
rect 12730 -6759 12809 -6641
rect 12927 -6759 13000 -6641
rect 12730 -6801 13000 -6759
rect 12730 -6919 12809 -6801
rect 12927 -6919 13000 -6801
rect 12730 -6961 13000 -6919
rect 12730 -7079 12809 -6961
rect 12927 -7079 13000 -6961
rect 12730 -7121 13000 -7079
rect 12730 -7239 12809 -7121
rect 12927 -7239 13000 -7121
rect 12730 -7281 13000 -7239
rect 12730 -7399 12809 -7281
rect 12927 -7399 13000 -7281
rect 12730 -7441 13000 -7399
rect 12730 -7559 12809 -7441
rect 12927 -7559 13000 -7441
rect 12730 -7601 13000 -7559
rect 12730 -7719 12809 -7601
rect 12927 -7719 13000 -7601
rect 12730 -7761 13000 -7719
rect 12730 -7879 12809 -7761
rect 12927 -7879 13000 -7761
rect 12730 -7921 13000 -7879
rect 12730 -8039 12809 -7921
rect 12927 -8039 13000 -7921
rect 12730 -8081 13000 -8039
rect 12730 -8199 12809 -8081
rect 12927 -8199 13000 -8081
rect 12730 -8241 13000 -8199
rect 12730 -8359 12809 -8241
rect 12927 -8359 13000 -8241
rect 12730 -8401 13000 -8359
rect 12730 -8519 12809 -8401
rect 12927 -8519 13000 -8401
rect 12730 -8561 13000 -8519
rect 12730 -8679 12809 -8561
rect 12927 -8679 13000 -8561
rect 12730 -8721 13000 -8679
rect 12730 -8839 12809 -8721
rect 12927 -8839 13000 -8721
rect 12730 -8881 13000 -8839
rect 12730 -8999 12809 -8881
rect 12927 -8999 13000 -8881
rect 12730 -9041 13000 -8999
rect 12730 -9159 12809 -9041
rect 12927 -9159 13000 -9041
rect 12730 -9201 13000 -9159
rect 12730 -9230 12809 -9201
rect 9194 -9306 12809 -9230
rect 9194 -9319 9261 -9306
rect 9000 -9424 9261 -9319
rect 9379 -9424 9421 -9306
rect 9539 -9424 9581 -9306
rect 9699 -9424 9741 -9306
rect 9859 -9424 9901 -9306
rect 10019 -9424 10061 -9306
rect 10179 -9424 10221 -9306
rect 10339 -9424 10381 -9306
rect 10499 -9424 10541 -9306
rect 10659 -9424 10701 -9306
rect 10819 -9424 10861 -9306
rect 10979 -9424 11021 -9306
rect 11139 -9424 11181 -9306
rect 11299 -9424 11341 -9306
rect 11459 -9424 11501 -9306
rect 11619 -9424 11661 -9306
rect 11779 -9424 11821 -9306
rect 11939 -9424 11981 -9306
rect 12099 -9424 12141 -9306
rect 12259 -9424 12301 -9306
rect 12419 -9424 12461 -9306
rect 12579 -9424 12621 -9306
rect 12739 -9319 12809 -9306
rect 12927 -9319 13000 -9201
rect 12739 -9424 13000 -9319
rect 9000 -9500 13000 -9424
rect 15000 -5578 19000 -5500
rect 15000 -5681 15261 -5578
rect 15000 -5799 15076 -5681
rect 15194 -5696 15261 -5681
rect 15379 -5696 15421 -5578
rect 15539 -5696 15581 -5578
rect 15699 -5696 15741 -5578
rect 15859 -5696 15901 -5578
rect 16019 -5696 16061 -5578
rect 16179 -5696 16221 -5578
rect 16339 -5696 16381 -5578
rect 16499 -5696 16541 -5578
rect 16659 -5696 16701 -5578
rect 16819 -5696 16861 -5578
rect 16979 -5696 17021 -5578
rect 17139 -5696 17181 -5578
rect 17299 -5696 17341 -5578
rect 17459 -5696 17501 -5578
rect 17619 -5696 17661 -5578
rect 17779 -5696 17821 -5578
rect 17939 -5696 17981 -5578
rect 18099 -5696 18141 -5578
rect 18259 -5696 18301 -5578
rect 18419 -5696 18461 -5578
rect 18579 -5696 18621 -5578
rect 18739 -5681 19000 -5578
rect 18739 -5696 18809 -5681
rect 15194 -5770 18809 -5696
rect 15194 -5799 15270 -5770
rect 15000 -5841 15270 -5799
rect 15000 -5959 15076 -5841
rect 15194 -5959 15270 -5841
rect 15000 -6001 15270 -5959
rect 15000 -6119 15076 -6001
rect 15194 -6119 15270 -6001
rect 15000 -6161 15270 -6119
rect 15000 -6279 15076 -6161
rect 15194 -6279 15270 -6161
rect 15000 -6321 15270 -6279
rect 15000 -6439 15076 -6321
rect 15194 -6439 15270 -6321
rect 15000 -6481 15270 -6439
rect 15000 -6599 15076 -6481
rect 15194 -6599 15270 -6481
rect 15000 -6641 15270 -6599
rect 15000 -6759 15076 -6641
rect 15194 -6759 15270 -6641
rect 15000 -6801 15270 -6759
rect 15000 -6919 15076 -6801
rect 15194 -6919 15270 -6801
rect 15000 -6961 15270 -6919
rect 15000 -7079 15076 -6961
rect 15194 -7079 15270 -6961
rect 15000 -7121 15270 -7079
rect 15000 -7239 15076 -7121
rect 15194 -7239 15270 -7121
rect 15000 -7281 15270 -7239
rect 15000 -7399 15076 -7281
rect 15194 -7399 15270 -7281
rect 15000 -7441 15270 -7399
rect 15000 -7559 15076 -7441
rect 15194 -7559 15270 -7441
rect 15000 -7601 15270 -7559
rect 15000 -7719 15076 -7601
rect 15194 -7719 15270 -7601
rect 15000 -7761 15270 -7719
rect 15000 -7879 15076 -7761
rect 15194 -7879 15270 -7761
rect 15000 -7921 15270 -7879
rect 15000 -8039 15076 -7921
rect 15194 -8039 15270 -7921
rect 15000 -8081 15270 -8039
rect 15000 -8199 15076 -8081
rect 15194 -8199 15270 -8081
rect 15000 -8241 15270 -8199
rect 15000 -8359 15076 -8241
rect 15194 -8359 15270 -8241
rect 15000 -8401 15270 -8359
rect 15000 -8519 15076 -8401
rect 15194 -8519 15270 -8401
rect 15000 -8561 15270 -8519
rect 15000 -8679 15076 -8561
rect 15194 -8679 15270 -8561
rect 15000 -8721 15270 -8679
rect 15000 -8839 15076 -8721
rect 15194 -8839 15270 -8721
rect 15000 -8881 15270 -8839
rect 15000 -8999 15076 -8881
rect 15194 -8999 15270 -8881
rect 15000 -9041 15270 -8999
rect 15000 -9159 15076 -9041
rect 15194 -9159 15270 -9041
rect 15000 -9201 15270 -9159
rect 15000 -9319 15076 -9201
rect 15194 -9230 15270 -9201
rect 18730 -5799 18809 -5770
rect 18927 -5799 19000 -5681
rect 19250 -5650 19350 -5450
rect 21000 -5578 25000 -5500
rect 21000 -5650 21261 -5578
rect 19250 -5681 21261 -5650
rect 19250 -5750 21076 -5681
rect 21194 -5696 21261 -5681
rect 21379 -5696 21421 -5578
rect 21539 -5696 21581 -5578
rect 21699 -5696 21741 -5578
rect 21859 -5696 21901 -5578
rect 22019 -5696 22061 -5578
rect 22179 -5696 22221 -5578
rect 22339 -5696 22381 -5578
rect 22499 -5696 22541 -5578
rect 22659 -5696 22701 -5578
rect 22819 -5696 22861 -5578
rect 22979 -5696 23021 -5578
rect 23139 -5696 23181 -5578
rect 23299 -5696 23341 -5578
rect 23459 -5696 23501 -5578
rect 23619 -5696 23661 -5578
rect 23779 -5696 23821 -5578
rect 23939 -5696 23981 -5578
rect 24099 -5696 24141 -5578
rect 24259 -5696 24301 -5578
rect 24419 -5696 24461 -5578
rect 24579 -5696 24621 -5578
rect 24739 -5681 25000 -5578
rect 24739 -5696 24809 -5681
rect 18730 -5841 19000 -5799
rect 18730 -5959 18809 -5841
rect 18927 -5959 19000 -5841
rect 18730 -6001 19000 -5959
rect 18730 -6119 18809 -6001
rect 18927 -6119 19000 -6001
rect 18730 -6161 19000 -6119
rect 18730 -6279 18809 -6161
rect 18927 -6279 19000 -6161
rect 18730 -6321 19000 -6279
rect 18730 -6439 18809 -6321
rect 18927 -6439 19000 -6321
rect 18730 -6481 19000 -6439
rect 18730 -6599 18809 -6481
rect 18927 -6599 19000 -6481
rect 18730 -6641 19000 -6599
rect 18730 -6759 18809 -6641
rect 18927 -6759 19000 -6641
rect 18730 -6801 19000 -6759
rect 18730 -6919 18809 -6801
rect 18927 -6919 19000 -6801
rect 18730 -6961 19000 -6919
rect 18730 -7079 18809 -6961
rect 18927 -7079 19000 -6961
rect 18730 -7121 19000 -7079
rect 18730 -7239 18809 -7121
rect 18927 -7239 19000 -7121
rect 18730 -7281 19000 -7239
rect 18730 -7399 18809 -7281
rect 18927 -7399 19000 -7281
rect 18730 -7441 19000 -7399
rect 18730 -7559 18809 -7441
rect 18927 -7559 19000 -7441
rect 18730 -7601 19000 -7559
rect 18730 -7719 18809 -7601
rect 18927 -7719 19000 -7601
rect 18730 -7761 19000 -7719
rect 18730 -7879 18809 -7761
rect 18927 -7879 19000 -7761
rect 18730 -7921 19000 -7879
rect 18730 -8039 18809 -7921
rect 18927 -8039 19000 -7921
rect 18730 -8081 19000 -8039
rect 18730 -8199 18809 -8081
rect 18927 -8199 19000 -8081
rect 18730 -8241 19000 -8199
rect 18730 -8359 18809 -8241
rect 18927 -8359 19000 -8241
rect 18730 -8401 19000 -8359
rect 18730 -8519 18809 -8401
rect 18927 -8519 19000 -8401
rect 18730 -8561 19000 -8519
rect 18730 -8679 18809 -8561
rect 18927 -8679 19000 -8561
rect 18730 -8721 19000 -8679
rect 18730 -8839 18809 -8721
rect 18927 -8839 19000 -8721
rect 18730 -8881 19000 -8839
rect 18730 -8999 18809 -8881
rect 18927 -8999 19000 -8881
rect 18730 -9041 19000 -8999
rect 18730 -9159 18809 -9041
rect 18927 -9159 19000 -9041
rect 18730 -9201 19000 -9159
rect 18730 -9230 18809 -9201
rect 15194 -9306 18809 -9230
rect 15194 -9319 15261 -9306
rect 15000 -9424 15261 -9319
rect 15379 -9424 15421 -9306
rect 15539 -9424 15581 -9306
rect 15699 -9424 15741 -9306
rect 15859 -9424 15901 -9306
rect 16019 -9424 16061 -9306
rect 16179 -9424 16221 -9306
rect 16339 -9424 16381 -9306
rect 16499 -9424 16541 -9306
rect 16659 -9424 16701 -9306
rect 16819 -9424 16861 -9306
rect 16979 -9424 17021 -9306
rect 17139 -9424 17181 -9306
rect 17299 -9424 17341 -9306
rect 17459 -9424 17501 -9306
rect 17619 -9424 17661 -9306
rect 17779 -9424 17821 -9306
rect 17939 -9424 17981 -9306
rect 18099 -9424 18141 -9306
rect 18259 -9424 18301 -9306
rect 18419 -9424 18461 -9306
rect 18579 -9424 18621 -9306
rect 18739 -9319 18809 -9306
rect 18927 -9319 19000 -9201
rect 18739 -9424 19000 -9319
rect 15000 -9500 19000 -9424
rect 21000 -5799 21076 -5750
rect 21194 -5770 24809 -5696
rect 21194 -5799 21270 -5770
rect 21000 -5841 21270 -5799
rect 21000 -5959 21076 -5841
rect 21194 -5959 21270 -5841
rect 21000 -6001 21270 -5959
rect 21000 -6119 21076 -6001
rect 21194 -6119 21270 -6001
rect 21000 -6161 21270 -6119
rect 21000 -6279 21076 -6161
rect 21194 -6279 21270 -6161
rect 21000 -6321 21270 -6279
rect 21000 -6439 21076 -6321
rect 21194 -6439 21270 -6321
rect 21000 -6481 21270 -6439
rect 21000 -6599 21076 -6481
rect 21194 -6599 21270 -6481
rect 21000 -6641 21270 -6599
rect 21000 -6759 21076 -6641
rect 21194 -6759 21270 -6641
rect 21000 -6801 21270 -6759
rect 21000 -6919 21076 -6801
rect 21194 -6919 21270 -6801
rect 21000 -6961 21270 -6919
rect 21000 -7079 21076 -6961
rect 21194 -7079 21270 -6961
rect 21000 -7121 21270 -7079
rect 21000 -7239 21076 -7121
rect 21194 -7239 21270 -7121
rect 21000 -7281 21270 -7239
rect 21000 -7399 21076 -7281
rect 21194 -7399 21270 -7281
rect 21000 -7441 21270 -7399
rect 21000 -7559 21076 -7441
rect 21194 -7559 21270 -7441
rect 21000 -7601 21270 -7559
rect 21000 -7719 21076 -7601
rect 21194 -7719 21270 -7601
rect 21000 -7761 21270 -7719
rect 21000 -7879 21076 -7761
rect 21194 -7879 21270 -7761
rect 21000 -7921 21270 -7879
rect 21000 -8039 21076 -7921
rect 21194 -8039 21270 -7921
rect 21000 -8081 21270 -8039
rect 21000 -8199 21076 -8081
rect 21194 -8199 21270 -8081
rect 21000 -8241 21270 -8199
rect 21000 -8359 21076 -8241
rect 21194 -8359 21270 -8241
rect 21000 -8401 21270 -8359
rect 21000 -8519 21076 -8401
rect 21194 -8519 21270 -8401
rect 21000 -8561 21270 -8519
rect 21000 -8679 21076 -8561
rect 21194 -8679 21270 -8561
rect 21000 -8721 21270 -8679
rect 21000 -8839 21076 -8721
rect 21194 -8839 21270 -8721
rect 21000 -8881 21270 -8839
rect 21000 -8999 21076 -8881
rect 21194 -8999 21270 -8881
rect 21000 -9041 21270 -8999
rect 21000 -9159 21076 -9041
rect 21194 -9159 21270 -9041
rect 21000 -9201 21270 -9159
rect 21000 -9319 21076 -9201
rect 21194 -9230 21270 -9201
rect 24730 -5799 24809 -5770
rect 24927 -5799 25000 -5681
rect 24730 -5841 25000 -5799
rect 24730 -5959 24809 -5841
rect 24927 -5959 25000 -5841
rect 24730 -6001 25000 -5959
rect 24730 -6119 24809 -6001
rect 24927 -6119 25000 -6001
rect 24730 -6161 25000 -6119
rect 24730 -6279 24809 -6161
rect 24927 -6279 25000 -6161
rect 24730 -6321 25000 -6279
rect 24730 -6439 24809 -6321
rect 24927 -6439 25000 -6321
rect 24730 -6481 25000 -6439
rect 24730 -6599 24809 -6481
rect 24927 -6599 25000 -6481
rect 24730 -6641 25000 -6599
rect 24730 -6759 24809 -6641
rect 24927 -6759 25000 -6641
rect 24730 -6801 25000 -6759
rect 24730 -6919 24809 -6801
rect 24927 -6919 25000 -6801
rect 24730 -6961 25000 -6919
rect 24730 -7079 24809 -6961
rect 24927 -7079 25000 -6961
rect 24730 -7121 25000 -7079
rect 24730 -7239 24809 -7121
rect 24927 -7239 25000 -7121
rect 24730 -7281 25000 -7239
rect 24730 -7399 24809 -7281
rect 24927 -7399 25000 -7281
rect 24730 -7441 25000 -7399
rect 24730 -7559 24809 -7441
rect 24927 -7559 25000 -7441
rect 24730 -7601 25000 -7559
rect 24730 -7719 24809 -7601
rect 24927 -7719 25000 -7601
rect 24730 -7761 25000 -7719
rect 24730 -7879 24809 -7761
rect 24927 -7879 25000 -7761
rect 24730 -7921 25000 -7879
rect 24730 -8039 24809 -7921
rect 24927 -8039 25000 -7921
rect 24730 -8081 25000 -8039
rect 24730 -8199 24809 -8081
rect 24927 -8199 25000 -8081
rect 24730 -8241 25000 -8199
rect 24730 -8359 24809 -8241
rect 24927 -8359 25000 -8241
rect 24730 -8401 25000 -8359
rect 24730 -8519 24809 -8401
rect 24927 -8519 25000 -8401
rect 24730 -8561 25000 -8519
rect 24730 -8679 24809 -8561
rect 24927 -8679 25000 -8561
rect 24730 -8721 25000 -8679
rect 24730 -8839 24809 -8721
rect 24927 -8839 25000 -8721
rect 24730 -8881 25000 -8839
rect 24730 -8999 24809 -8881
rect 24927 -8999 25000 -8881
rect 24730 -9041 25000 -8999
rect 24730 -9159 24809 -9041
rect 24927 -9159 25000 -9041
rect 24730 -9201 25000 -9159
rect 24730 -9230 24809 -9201
rect 21194 -9306 24809 -9230
rect 21194 -9319 21261 -9306
rect 21000 -9424 21261 -9319
rect 21379 -9424 21421 -9306
rect 21539 -9424 21581 -9306
rect 21699 -9424 21741 -9306
rect 21859 -9424 21901 -9306
rect 22019 -9424 22061 -9306
rect 22179 -9424 22221 -9306
rect 22339 -9424 22381 -9306
rect 22499 -9424 22541 -9306
rect 22659 -9424 22701 -9306
rect 22819 -9424 22861 -9306
rect 22979 -9424 23021 -9306
rect 23139 -9424 23181 -9306
rect 23299 -9424 23341 -9306
rect 23459 -9424 23501 -9306
rect 23619 -9424 23661 -9306
rect 23779 -9424 23821 -9306
rect 23939 -9424 23981 -9306
rect 24099 -9424 24141 -9306
rect 24259 -9424 24301 -9306
rect 24419 -9424 24461 -9306
rect 24579 -9424 24621 -9306
rect 24739 -9319 24809 -9306
rect 24927 -9319 25000 -9201
rect 24739 -9424 25000 -9319
rect 21000 -9500 25000 -9424
rect 3050 -9800 3150 -9550
rect 3250 -9800 3350 -9550
rect 3050 -9850 3350 -9800
rect 3450 -9600 3700 -9550
rect 3850 -9600 4100 -9550
rect 3450 -9650 3750 -9600
rect 3450 -9850 3550 -9650
rect 3650 -9850 3750 -9650
rect 3100 -9900 3300 -9850
rect 3450 -9900 3750 -9850
rect 3850 -9650 4150 -9600
rect 3850 -9850 3950 -9650
rect 4050 -9850 4150 -9650
rect 9050 -9800 9150 -9550
rect 9250 -9800 9350 -9550
rect 9450 -9650 9750 -9550
rect 9850 -9650 10150 -9550
rect 9450 -9700 9550 -9650
rect 9850 -9700 9950 -9650
rect 9450 -9750 9700 -9700
rect 9850 -9750 10100 -9700
rect 9500 -9800 9750 -9750
rect 9900 -9800 10150 -9750
rect 9050 -9850 9350 -9800
rect 9650 -9850 9750 -9800
rect 10050 -9850 10150 -9800
rect 15050 -9800 15150 -9550
rect 15250 -9800 15350 -9550
rect 15450 -9650 15750 -9550
rect 15050 -9850 15350 -9800
rect 15550 -9850 15650 -9650
rect 15950 -9700 16050 -9600
rect 15850 -9800 16150 -9700
rect 21050 -9800 21150 -9550
rect 21250 -9800 21350 -9550
rect 21500 -9600 21700 -9550
rect 3850 -9900 4150 -9850
rect 9100 -9900 9300 -9850
rect 3150 -9950 3250 -9900
rect 3450 -9950 3700 -9900
rect 3850 -9950 4100 -9900
rect 9150 -9950 9250 -9900
rect 9450 -9950 9750 -9850
rect 9850 -9950 10150 -9850
rect 15100 -9900 15300 -9850
rect 15150 -9950 15250 -9900
rect 15450 -9950 15750 -9850
rect 15950 -9900 16050 -9800
rect 21050 -9850 21350 -9800
rect 21450 -9650 21750 -9600
rect 21450 -9850 21550 -9650
rect 21650 -9850 21750 -9650
rect 21950 -9700 22050 -9600
rect 21850 -9800 22150 -9700
rect 21100 -9900 21300 -9850
rect 21450 -9900 21750 -9850
rect 21950 -9900 22050 -9800
rect 21150 -9950 21250 -9900
rect 21500 -9950 21700 -9900
rect 9050 -11000 9350 -10950
rect 3050 -11150 3350 -11050
rect 9050 -11150 9350 -11050
rect 3050 -11200 3150 -11150
rect 9050 -11200 9150 -11150
rect 3050 -11250 3300 -11200
rect 9050 -11250 9300 -11200
rect 3100 -11300 3350 -11250
rect 9100 -11300 9350 -11250
rect 3250 -11350 3350 -11300
rect 9250 -11350 9350 -11300
rect 15050 -11300 15150 -11050
rect 15250 -11300 15350 -11050
rect 15050 -11350 15350 -11300
rect 15450 -11100 15700 -11050
rect 15450 -11150 15750 -11100
rect 15450 -11250 15550 -11150
rect 15650 -11250 15750 -11150
rect 15850 -11150 16150 -11050
rect 16250 -11150 16550 -11050
rect 15850 -11200 15950 -11150
rect 16250 -11200 16350 -11150
rect 15450 -11350 15700 -11250
rect 15850 -11300 16100 -11200
rect 16250 -11300 16500 -11200
rect 21050 -11300 21150 -11050
rect 21250 -11300 21350 -11050
rect 21450 -11150 21750 -11050
rect 15850 -11350 15950 -11300
rect 3050 -11450 3350 -11350
rect 9050 -11450 9350 -11350
rect 15100 -11400 15300 -11350
rect 15150 -11450 15250 -11400
rect 15450 -11450 15550 -11350
rect 15650 -11450 15750 -11350
rect 15850 -11450 16150 -11350
rect 16250 -11450 16350 -11300
rect 21050 -11350 21350 -11300
rect 21550 -11350 21650 -11150
rect 21850 -11300 22150 -11200
rect 21100 -11400 21300 -11350
rect 21150 -11450 21250 -11400
rect 21450 -11450 21750 -11350
rect 3000 -11578 7000 -11500
rect 3000 -11681 3261 -11578
rect 3000 -11799 3076 -11681
rect 3194 -11696 3261 -11681
rect 3379 -11696 3421 -11578
rect 3539 -11696 3581 -11578
rect 3699 -11696 3741 -11578
rect 3859 -11696 3901 -11578
rect 4019 -11696 4061 -11578
rect 4179 -11696 4221 -11578
rect 4339 -11696 4381 -11578
rect 4499 -11696 4541 -11578
rect 4659 -11696 4701 -11578
rect 4819 -11696 4861 -11578
rect 4979 -11696 5021 -11578
rect 5139 -11696 5181 -11578
rect 5299 -11696 5341 -11578
rect 5459 -11696 5501 -11578
rect 5619 -11696 5661 -11578
rect 5779 -11696 5821 -11578
rect 5939 -11696 5981 -11578
rect 6099 -11696 6141 -11578
rect 6259 -11696 6301 -11578
rect 6419 -11696 6461 -11578
rect 6579 -11696 6621 -11578
rect 6739 -11681 7000 -11578
rect 6739 -11696 6809 -11681
rect 3194 -11770 6809 -11696
rect 3194 -11799 3270 -11770
rect 3000 -11841 3270 -11799
rect 3000 -11959 3076 -11841
rect 3194 -11959 3270 -11841
rect 3000 -12001 3270 -11959
rect 3000 -12119 3076 -12001
rect 3194 -12119 3270 -12001
rect 3000 -12161 3270 -12119
rect 3000 -12279 3076 -12161
rect 3194 -12279 3270 -12161
rect 3000 -12321 3270 -12279
rect 3000 -12439 3076 -12321
rect 3194 -12439 3270 -12321
rect 3000 -12481 3270 -12439
rect 3000 -12599 3076 -12481
rect 3194 -12599 3270 -12481
rect 3000 -12641 3270 -12599
rect 3000 -12759 3076 -12641
rect 3194 -12759 3270 -12641
rect 3000 -12801 3270 -12759
rect 3000 -12919 3076 -12801
rect 3194 -12919 3270 -12801
rect 3000 -12961 3270 -12919
rect 3000 -13079 3076 -12961
rect 3194 -13079 3270 -12961
rect 3000 -13121 3270 -13079
rect 3000 -13239 3076 -13121
rect 3194 -13239 3270 -13121
rect 3000 -13281 3270 -13239
rect 3000 -13399 3076 -13281
rect 3194 -13399 3270 -13281
rect 3000 -13441 3270 -13399
rect 3000 -13559 3076 -13441
rect 3194 -13559 3270 -13441
rect 3000 -13601 3270 -13559
rect 3000 -13719 3076 -13601
rect 3194 -13719 3270 -13601
rect 3000 -13761 3270 -13719
rect 3000 -13879 3076 -13761
rect 3194 -13879 3270 -13761
rect 3000 -13921 3270 -13879
rect 3000 -14039 3076 -13921
rect 3194 -14039 3270 -13921
rect 3000 -14081 3270 -14039
rect 3000 -14199 3076 -14081
rect 3194 -14199 3270 -14081
rect 3000 -14241 3270 -14199
rect 3000 -14359 3076 -14241
rect 3194 -14359 3270 -14241
rect 3000 -14401 3270 -14359
rect 3000 -14519 3076 -14401
rect 3194 -14519 3270 -14401
rect 3000 -14561 3270 -14519
rect 3000 -14679 3076 -14561
rect 3194 -14679 3270 -14561
rect 3000 -14721 3270 -14679
rect 3000 -14839 3076 -14721
rect 3194 -14839 3270 -14721
rect 3000 -14881 3270 -14839
rect 3000 -14999 3076 -14881
rect 3194 -14999 3270 -14881
rect 3000 -15041 3270 -14999
rect 3000 -15159 3076 -15041
rect 3194 -15159 3270 -15041
rect 3000 -15201 3270 -15159
rect 3000 -15319 3076 -15201
rect 3194 -15230 3270 -15201
rect 6730 -11799 6809 -11770
rect 6927 -11799 7000 -11681
rect 6730 -11841 7000 -11799
rect 6730 -11959 6809 -11841
rect 6927 -11959 7000 -11841
rect 6730 -12001 7000 -11959
rect 6730 -12119 6809 -12001
rect 6927 -12119 7000 -12001
rect 6730 -12161 7000 -12119
rect 6730 -12279 6809 -12161
rect 6927 -12279 7000 -12161
rect 6730 -12321 7000 -12279
rect 6730 -12439 6809 -12321
rect 6927 -12439 7000 -12321
rect 6730 -12481 7000 -12439
rect 6730 -12599 6809 -12481
rect 6927 -12599 7000 -12481
rect 6730 -12641 7000 -12599
rect 6730 -12759 6809 -12641
rect 6927 -12759 7000 -12641
rect 6730 -12801 7000 -12759
rect 6730 -12919 6809 -12801
rect 6927 -12919 7000 -12801
rect 6730 -12961 7000 -12919
rect 6730 -13079 6809 -12961
rect 6927 -13079 7000 -12961
rect 6730 -13121 7000 -13079
rect 6730 -13239 6809 -13121
rect 6927 -13239 7000 -13121
rect 6730 -13281 7000 -13239
rect 6730 -13399 6809 -13281
rect 6927 -13399 7000 -13281
rect 6730 -13441 7000 -13399
rect 6730 -13559 6809 -13441
rect 6927 -13559 7000 -13441
rect 6730 -13601 7000 -13559
rect 6730 -13719 6809 -13601
rect 6927 -13719 7000 -13601
rect 6730 -13761 7000 -13719
rect 6730 -13879 6809 -13761
rect 6927 -13879 7000 -13761
rect 6730 -13921 7000 -13879
rect 6730 -14039 6809 -13921
rect 6927 -14039 7000 -13921
rect 6730 -14081 7000 -14039
rect 6730 -14199 6809 -14081
rect 6927 -14199 7000 -14081
rect 6730 -14241 7000 -14199
rect 6730 -14359 6809 -14241
rect 6927 -14359 7000 -14241
rect 6730 -14401 7000 -14359
rect 6730 -14519 6809 -14401
rect 6927 -14519 7000 -14401
rect 6730 -14561 7000 -14519
rect 6730 -14679 6809 -14561
rect 6927 -14679 7000 -14561
rect 6730 -14721 7000 -14679
rect 6730 -14839 6809 -14721
rect 6927 -14839 7000 -14721
rect 6730 -14881 7000 -14839
rect 6730 -14999 6809 -14881
rect 6927 -14999 7000 -14881
rect 6730 -15041 7000 -14999
rect 6730 -15159 6809 -15041
rect 6927 -15159 7000 -15041
rect 6730 -15201 7000 -15159
rect 6730 -15230 6809 -15201
rect 3194 -15306 6809 -15230
rect 3194 -15319 3261 -15306
rect 3000 -15424 3261 -15319
rect 3379 -15424 3421 -15306
rect 3539 -15424 3581 -15306
rect 3699 -15424 3741 -15306
rect 3859 -15424 3901 -15306
rect 4019 -15424 4061 -15306
rect 4179 -15424 4221 -15306
rect 4339 -15424 4381 -15306
rect 4499 -15424 4541 -15306
rect 4659 -15424 4701 -15306
rect 4819 -15424 4861 -15306
rect 4979 -15424 5021 -15306
rect 5139 -15424 5181 -15306
rect 5299 -15424 5341 -15306
rect 5459 -15424 5501 -15306
rect 5619 -15424 5661 -15306
rect 5779 -15424 5821 -15306
rect 5939 -15424 5981 -15306
rect 6099 -15424 6141 -15306
rect 6259 -15424 6301 -15306
rect 6419 -15424 6461 -15306
rect 6579 -15424 6621 -15306
rect 6739 -15319 6809 -15306
rect 6927 -15319 7000 -15201
rect 6739 -15424 7000 -15319
rect 3000 -15500 7000 -15424
rect 9000 -11578 13000 -11500
rect 9000 -11681 9261 -11578
rect 9000 -11799 9076 -11681
rect 9194 -11696 9261 -11681
rect 9379 -11696 9421 -11578
rect 9539 -11696 9581 -11578
rect 9699 -11696 9741 -11578
rect 9859 -11696 9901 -11578
rect 10019 -11696 10061 -11578
rect 10179 -11696 10221 -11578
rect 10339 -11696 10381 -11578
rect 10499 -11696 10541 -11578
rect 10659 -11696 10701 -11578
rect 10819 -11696 10861 -11578
rect 10979 -11696 11021 -11578
rect 11139 -11696 11181 -11578
rect 11299 -11696 11341 -11578
rect 11459 -11696 11501 -11578
rect 11619 -11696 11661 -11578
rect 11779 -11696 11821 -11578
rect 11939 -11696 11981 -11578
rect 12099 -11696 12141 -11578
rect 12259 -11696 12301 -11578
rect 12419 -11696 12461 -11578
rect 12579 -11696 12621 -11578
rect 12739 -11681 13000 -11578
rect 12739 -11696 12809 -11681
rect 9194 -11770 12809 -11696
rect 9194 -11799 9270 -11770
rect 9000 -11841 9270 -11799
rect 9000 -11959 9076 -11841
rect 9194 -11959 9270 -11841
rect 9000 -12001 9270 -11959
rect 9000 -12119 9076 -12001
rect 9194 -12119 9270 -12001
rect 9000 -12161 9270 -12119
rect 9000 -12279 9076 -12161
rect 9194 -12279 9270 -12161
rect 9000 -12321 9270 -12279
rect 9000 -12439 9076 -12321
rect 9194 -12439 9270 -12321
rect 9000 -12481 9270 -12439
rect 9000 -12599 9076 -12481
rect 9194 -12599 9270 -12481
rect 9000 -12641 9270 -12599
rect 9000 -12759 9076 -12641
rect 9194 -12759 9270 -12641
rect 9000 -12801 9270 -12759
rect 9000 -12919 9076 -12801
rect 9194 -12919 9270 -12801
rect 9000 -12961 9270 -12919
rect 9000 -13079 9076 -12961
rect 9194 -13079 9270 -12961
rect 9000 -13121 9270 -13079
rect 9000 -13239 9076 -13121
rect 9194 -13239 9270 -13121
rect 9000 -13281 9270 -13239
rect 9000 -13399 9076 -13281
rect 9194 -13399 9270 -13281
rect 9000 -13441 9270 -13399
rect 9000 -13559 9076 -13441
rect 9194 -13559 9270 -13441
rect 9000 -13601 9270 -13559
rect 9000 -13719 9076 -13601
rect 9194 -13719 9270 -13601
rect 9000 -13761 9270 -13719
rect 9000 -13879 9076 -13761
rect 9194 -13879 9270 -13761
rect 9000 -13921 9270 -13879
rect 9000 -14039 9076 -13921
rect 9194 -14039 9270 -13921
rect 9000 -14081 9270 -14039
rect 9000 -14199 9076 -14081
rect 9194 -14199 9270 -14081
rect 9000 -14241 9270 -14199
rect 9000 -14359 9076 -14241
rect 9194 -14359 9270 -14241
rect 9000 -14401 9270 -14359
rect 9000 -14519 9076 -14401
rect 9194 -14519 9270 -14401
rect 9000 -14561 9270 -14519
rect 9000 -14679 9076 -14561
rect 9194 -14679 9270 -14561
rect 9000 -14721 9270 -14679
rect 9000 -14839 9076 -14721
rect 9194 -14839 9270 -14721
rect 9000 -14881 9270 -14839
rect 9000 -14999 9076 -14881
rect 9194 -14999 9270 -14881
rect 9000 -15041 9270 -14999
rect 9000 -15159 9076 -15041
rect 9194 -15159 9270 -15041
rect 9000 -15201 9270 -15159
rect 9000 -15319 9076 -15201
rect 9194 -15230 9270 -15201
rect 12730 -11799 12809 -11770
rect 12927 -11799 13000 -11681
rect 12730 -11841 13000 -11799
rect 12730 -11959 12809 -11841
rect 12927 -11959 13000 -11841
rect 12730 -12001 13000 -11959
rect 12730 -12119 12809 -12001
rect 12927 -12119 13000 -12001
rect 12730 -12161 13000 -12119
rect 12730 -12279 12809 -12161
rect 12927 -12279 13000 -12161
rect 12730 -12321 13000 -12279
rect 12730 -12439 12809 -12321
rect 12927 -12439 13000 -12321
rect 12730 -12481 13000 -12439
rect 12730 -12599 12809 -12481
rect 12927 -12599 13000 -12481
rect 12730 -12641 13000 -12599
rect 12730 -12759 12809 -12641
rect 12927 -12759 13000 -12641
rect 12730 -12801 13000 -12759
rect 12730 -12919 12809 -12801
rect 12927 -12919 13000 -12801
rect 12730 -12961 13000 -12919
rect 12730 -13079 12809 -12961
rect 12927 -13079 13000 -12961
rect 12730 -13121 13000 -13079
rect 12730 -13239 12809 -13121
rect 12927 -13239 13000 -13121
rect 12730 -13281 13000 -13239
rect 12730 -13399 12809 -13281
rect 12927 -13399 13000 -13281
rect 12730 -13441 13000 -13399
rect 12730 -13559 12809 -13441
rect 12927 -13559 13000 -13441
rect 12730 -13601 13000 -13559
rect 12730 -13719 12809 -13601
rect 12927 -13719 13000 -13601
rect 12730 -13761 13000 -13719
rect 12730 -13879 12809 -13761
rect 12927 -13879 13000 -13761
rect 12730 -13921 13000 -13879
rect 12730 -14039 12809 -13921
rect 12927 -14039 13000 -13921
rect 12730 -14081 13000 -14039
rect 12730 -14199 12809 -14081
rect 12927 -14199 13000 -14081
rect 12730 -14241 13000 -14199
rect 12730 -14359 12809 -14241
rect 12927 -14359 13000 -14241
rect 12730 -14401 13000 -14359
rect 12730 -14519 12809 -14401
rect 12927 -14519 13000 -14401
rect 12730 -14561 13000 -14519
rect 12730 -14679 12809 -14561
rect 12927 -14679 13000 -14561
rect 12730 -14721 13000 -14679
rect 12730 -14839 12809 -14721
rect 12927 -14839 13000 -14721
rect 12730 -14881 13000 -14839
rect 12730 -14999 12809 -14881
rect 12927 -14999 13000 -14881
rect 12730 -15041 13000 -14999
rect 12730 -15159 12809 -15041
rect 12927 -15159 13000 -15041
rect 12730 -15201 13000 -15159
rect 12730 -15230 12809 -15201
rect 9194 -15306 12809 -15230
rect 9194 -15319 9261 -15306
rect 9000 -15424 9261 -15319
rect 9379 -15424 9421 -15306
rect 9539 -15424 9581 -15306
rect 9699 -15424 9741 -15306
rect 9859 -15424 9901 -15306
rect 10019 -15424 10061 -15306
rect 10179 -15424 10221 -15306
rect 10339 -15424 10381 -15306
rect 10499 -15424 10541 -15306
rect 10659 -15424 10701 -15306
rect 10819 -15424 10861 -15306
rect 10979 -15424 11021 -15306
rect 11139 -15424 11181 -15306
rect 11299 -15424 11341 -15306
rect 11459 -15424 11501 -15306
rect 11619 -15424 11661 -15306
rect 11779 -15424 11821 -15306
rect 11939 -15424 11981 -15306
rect 12099 -15424 12141 -15306
rect 12259 -15424 12301 -15306
rect 12419 -15424 12461 -15306
rect 12579 -15424 12621 -15306
rect 12739 -15319 12809 -15306
rect 12927 -15319 13000 -15201
rect 12739 -15424 13000 -15319
rect 9000 -15500 13000 -15424
rect 15000 -11578 19000 -11500
rect 15000 -11681 15261 -11578
rect 15000 -11799 15076 -11681
rect 15194 -11696 15261 -11681
rect 15379 -11696 15421 -11578
rect 15539 -11696 15581 -11578
rect 15699 -11696 15741 -11578
rect 15859 -11696 15901 -11578
rect 16019 -11696 16061 -11578
rect 16179 -11696 16221 -11578
rect 16339 -11696 16381 -11578
rect 16499 -11696 16541 -11578
rect 16659 -11696 16701 -11578
rect 16819 -11696 16861 -11578
rect 16979 -11696 17021 -11578
rect 17139 -11696 17181 -11578
rect 17299 -11696 17341 -11578
rect 17459 -11696 17501 -11578
rect 17619 -11696 17661 -11578
rect 17779 -11696 17821 -11578
rect 17939 -11696 17981 -11578
rect 18099 -11696 18141 -11578
rect 18259 -11696 18301 -11578
rect 18419 -11696 18461 -11578
rect 18579 -11696 18621 -11578
rect 18739 -11681 19000 -11578
rect 18739 -11696 18809 -11681
rect 15194 -11770 18809 -11696
rect 15194 -11799 15270 -11770
rect 15000 -11841 15270 -11799
rect 15000 -11959 15076 -11841
rect 15194 -11959 15270 -11841
rect 15000 -12001 15270 -11959
rect 15000 -12119 15076 -12001
rect 15194 -12119 15270 -12001
rect 15000 -12161 15270 -12119
rect 15000 -12279 15076 -12161
rect 15194 -12279 15270 -12161
rect 15000 -12321 15270 -12279
rect 15000 -12439 15076 -12321
rect 15194 -12439 15270 -12321
rect 15000 -12481 15270 -12439
rect 15000 -12599 15076 -12481
rect 15194 -12599 15270 -12481
rect 15000 -12641 15270 -12599
rect 15000 -12759 15076 -12641
rect 15194 -12759 15270 -12641
rect 15000 -12801 15270 -12759
rect 15000 -12919 15076 -12801
rect 15194 -12919 15270 -12801
rect 15000 -12961 15270 -12919
rect 15000 -13079 15076 -12961
rect 15194 -13079 15270 -12961
rect 15000 -13121 15270 -13079
rect 15000 -13239 15076 -13121
rect 15194 -13239 15270 -13121
rect 15000 -13281 15270 -13239
rect 15000 -13399 15076 -13281
rect 15194 -13399 15270 -13281
rect 15000 -13441 15270 -13399
rect 15000 -13559 15076 -13441
rect 15194 -13559 15270 -13441
rect 15000 -13601 15270 -13559
rect 15000 -13719 15076 -13601
rect 15194 -13719 15270 -13601
rect 15000 -13761 15270 -13719
rect 15000 -13879 15076 -13761
rect 15194 -13879 15270 -13761
rect 15000 -13921 15270 -13879
rect 15000 -14039 15076 -13921
rect 15194 -14039 15270 -13921
rect 15000 -14081 15270 -14039
rect 15000 -14199 15076 -14081
rect 15194 -14199 15270 -14081
rect 15000 -14241 15270 -14199
rect 15000 -14359 15076 -14241
rect 15194 -14359 15270 -14241
rect 15000 -14401 15270 -14359
rect 15000 -14519 15076 -14401
rect 15194 -14519 15270 -14401
rect 15000 -14561 15270 -14519
rect 15000 -14679 15076 -14561
rect 15194 -14679 15270 -14561
rect 15000 -14721 15270 -14679
rect 15000 -14839 15076 -14721
rect 15194 -14839 15270 -14721
rect 15000 -14881 15270 -14839
rect 15000 -14999 15076 -14881
rect 15194 -14999 15270 -14881
rect 15000 -15041 15270 -14999
rect 15000 -15159 15076 -15041
rect 15194 -15159 15270 -15041
rect 15000 -15201 15270 -15159
rect 15000 -15319 15076 -15201
rect 15194 -15230 15270 -15201
rect 18730 -11799 18809 -11770
rect 18927 -11799 19000 -11681
rect 18730 -11841 19000 -11799
rect 18730 -11959 18809 -11841
rect 18927 -11959 19000 -11841
rect 18730 -12001 19000 -11959
rect 18730 -12119 18809 -12001
rect 18927 -12119 19000 -12001
rect 18730 -12161 19000 -12119
rect 18730 -12279 18809 -12161
rect 18927 -12279 19000 -12161
rect 18730 -12321 19000 -12279
rect 18730 -12439 18809 -12321
rect 18927 -12439 19000 -12321
rect 18730 -12481 19000 -12439
rect 18730 -12599 18809 -12481
rect 18927 -12599 19000 -12481
rect 18730 -12641 19000 -12599
rect 18730 -12759 18809 -12641
rect 18927 -12759 19000 -12641
rect 18730 -12801 19000 -12759
rect 18730 -12919 18809 -12801
rect 18927 -12919 19000 -12801
rect 18730 -12961 19000 -12919
rect 18730 -13079 18809 -12961
rect 18927 -13079 19000 -12961
rect 18730 -13121 19000 -13079
rect 18730 -13239 18809 -13121
rect 18927 -13239 19000 -13121
rect 18730 -13281 19000 -13239
rect 18730 -13399 18809 -13281
rect 18927 -13399 19000 -13281
rect 18730 -13441 19000 -13399
rect 18730 -13559 18809 -13441
rect 18927 -13559 19000 -13441
rect 18730 -13601 19000 -13559
rect 18730 -13719 18809 -13601
rect 18927 -13719 19000 -13601
rect 18730 -13761 19000 -13719
rect 18730 -13879 18809 -13761
rect 18927 -13879 19000 -13761
rect 18730 -13921 19000 -13879
rect 18730 -14039 18809 -13921
rect 18927 -14039 19000 -13921
rect 18730 -14081 19000 -14039
rect 18730 -14199 18809 -14081
rect 18927 -14199 19000 -14081
rect 18730 -14241 19000 -14199
rect 18730 -14359 18809 -14241
rect 18927 -14359 19000 -14241
rect 18730 -14401 19000 -14359
rect 18730 -14519 18809 -14401
rect 18927 -14519 19000 -14401
rect 18730 -14561 19000 -14519
rect 18730 -14679 18809 -14561
rect 18927 -14679 19000 -14561
rect 18730 -14721 19000 -14679
rect 18730 -14839 18809 -14721
rect 18927 -14839 19000 -14721
rect 18730 -14881 19000 -14839
rect 18730 -14999 18809 -14881
rect 18927 -14999 19000 -14881
rect 18730 -15041 19000 -14999
rect 18730 -15159 18809 -15041
rect 18927 -15159 19000 -15041
rect 18730 -15201 19000 -15159
rect 18730 -15230 18809 -15201
rect 15194 -15306 18809 -15230
rect 15194 -15319 15261 -15306
rect 15000 -15424 15261 -15319
rect 15379 -15424 15421 -15306
rect 15539 -15424 15581 -15306
rect 15699 -15424 15741 -15306
rect 15859 -15424 15901 -15306
rect 16019 -15424 16061 -15306
rect 16179 -15424 16221 -15306
rect 16339 -15424 16381 -15306
rect 16499 -15424 16541 -15306
rect 16659 -15424 16701 -15306
rect 16819 -15424 16861 -15306
rect 16979 -15424 17021 -15306
rect 17139 -15424 17181 -15306
rect 17299 -15424 17341 -15306
rect 17459 -15424 17501 -15306
rect 17619 -15424 17661 -15306
rect 17779 -15424 17821 -15306
rect 17939 -15424 17981 -15306
rect 18099 -15424 18141 -15306
rect 18259 -15424 18301 -15306
rect 18419 -15424 18461 -15306
rect 18579 -15424 18621 -15306
rect 18739 -15319 18809 -15306
rect 18927 -15319 19000 -15201
rect 18739 -15424 19000 -15319
rect 15000 -15500 19000 -15424
rect 21000 -11578 25000 -11500
rect 21000 -11681 21261 -11578
rect 21000 -11799 21076 -11681
rect 21194 -11696 21261 -11681
rect 21379 -11696 21421 -11578
rect 21539 -11696 21581 -11578
rect 21699 -11696 21741 -11578
rect 21859 -11696 21901 -11578
rect 22019 -11696 22061 -11578
rect 22179 -11696 22221 -11578
rect 22339 -11696 22381 -11578
rect 22499 -11696 22541 -11578
rect 22659 -11696 22701 -11578
rect 22819 -11696 22861 -11578
rect 22979 -11696 23021 -11578
rect 23139 -11696 23181 -11578
rect 23299 -11696 23341 -11578
rect 23459 -11696 23501 -11578
rect 23619 -11696 23661 -11578
rect 23779 -11696 23821 -11578
rect 23939 -11696 23981 -11578
rect 24099 -11696 24141 -11578
rect 24259 -11696 24301 -11578
rect 24419 -11696 24461 -11578
rect 24579 -11696 24621 -11578
rect 24739 -11681 25000 -11578
rect 24739 -11696 24809 -11681
rect 21194 -11770 24809 -11696
rect 21194 -11799 21270 -11770
rect 21000 -11841 21270 -11799
rect 21000 -11959 21076 -11841
rect 21194 -11959 21270 -11841
rect 21000 -12001 21270 -11959
rect 21000 -12119 21076 -12001
rect 21194 -12119 21270 -12001
rect 21000 -12161 21270 -12119
rect 21000 -12279 21076 -12161
rect 21194 -12279 21270 -12161
rect 21000 -12321 21270 -12279
rect 21000 -12439 21076 -12321
rect 21194 -12439 21270 -12321
rect 21000 -12481 21270 -12439
rect 21000 -12599 21076 -12481
rect 21194 -12599 21270 -12481
rect 21000 -12641 21270 -12599
rect 21000 -12759 21076 -12641
rect 21194 -12759 21270 -12641
rect 21000 -12801 21270 -12759
rect 21000 -12919 21076 -12801
rect 21194 -12919 21270 -12801
rect 21000 -12961 21270 -12919
rect 21000 -13079 21076 -12961
rect 21194 -13079 21270 -12961
rect 21000 -13121 21270 -13079
rect 21000 -13239 21076 -13121
rect 21194 -13239 21270 -13121
rect 21000 -13281 21270 -13239
rect 21000 -13399 21076 -13281
rect 21194 -13399 21270 -13281
rect 21000 -13441 21270 -13399
rect 21000 -13559 21076 -13441
rect 21194 -13559 21270 -13441
rect 21000 -13601 21270 -13559
rect 21000 -13719 21076 -13601
rect 21194 -13719 21270 -13601
rect 21000 -13761 21270 -13719
rect 21000 -13879 21076 -13761
rect 21194 -13879 21270 -13761
rect 21000 -13921 21270 -13879
rect 21000 -14039 21076 -13921
rect 21194 -14039 21270 -13921
rect 21000 -14081 21270 -14039
rect 21000 -14199 21076 -14081
rect 21194 -14199 21270 -14081
rect 21000 -14241 21270 -14199
rect 21000 -14359 21076 -14241
rect 21194 -14359 21270 -14241
rect 21000 -14401 21270 -14359
rect 21000 -14519 21076 -14401
rect 21194 -14519 21270 -14401
rect 21000 -14561 21270 -14519
rect 21000 -14679 21076 -14561
rect 21194 -14679 21270 -14561
rect 21000 -14721 21270 -14679
rect 21000 -14839 21076 -14721
rect 21194 -14839 21270 -14721
rect 21000 -14881 21270 -14839
rect 21000 -14999 21076 -14881
rect 21194 -14999 21270 -14881
rect 21000 -15041 21270 -14999
rect 21000 -15159 21076 -15041
rect 21194 -15159 21270 -15041
rect 21000 -15201 21270 -15159
rect 21000 -15319 21076 -15201
rect 21194 -15230 21270 -15201
rect 24730 -11799 24809 -11770
rect 24927 -11799 25000 -11681
rect 24730 -11841 25000 -11799
rect 24730 -11959 24809 -11841
rect 24927 -11959 25000 -11841
rect 24730 -12001 25000 -11959
rect 24730 -12119 24809 -12001
rect 24927 -12119 25000 -12001
rect 24730 -12161 25000 -12119
rect 24730 -12279 24809 -12161
rect 24927 -12279 25000 -12161
rect 24730 -12321 25000 -12279
rect 24730 -12439 24809 -12321
rect 24927 -12439 25000 -12321
rect 24730 -12481 25000 -12439
rect 24730 -12599 24809 -12481
rect 24927 -12599 25000 -12481
rect 24730 -12641 25000 -12599
rect 24730 -12759 24809 -12641
rect 24927 -12759 25000 -12641
rect 24730 -12801 25000 -12759
rect 24730 -12919 24809 -12801
rect 24927 -12919 25000 -12801
rect 24730 -12961 25000 -12919
rect 24730 -13079 24809 -12961
rect 24927 -13079 25000 -12961
rect 24730 -13121 25000 -13079
rect 24730 -13239 24809 -13121
rect 24927 -13239 25000 -13121
rect 24730 -13281 25000 -13239
rect 24730 -13399 24809 -13281
rect 24927 -13399 25000 -13281
rect 24730 -13441 25000 -13399
rect 24730 -13559 24809 -13441
rect 24927 -13559 25000 -13441
rect 24730 -13601 25000 -13559
rect 24730 -13719 24809 -13601
rect 24927 -13719 25000 -13601
rect 24730 -13761 25000 -13719
rect 24730 -13879 24809 -13761
rect 24927 -13879 25000 -13761
rect 24730 -13921 25000 -13879
rect 24730 -14039 24809 -13921
rect 24927 -14039 25000 -13921
rect 24730 -14081 25000 -14039
rect 24730 -14199 24809 -14081
rect 24927 -14199 25000 -14081
rect 24730 -14241 25000 -14199
rect 24730 -14359 24809 -14241
rect 24927 -14359 25000 -14241
rect 24730 -14401 25000 -14359
rect 24730 -14519 24809 -14401
rect 24927 -14519 25000 -14401
rect 24730 -14561 25000 -14519
rect 24730 -14679 24809 -14561
rect 24927 -14679 25000 -14561
rect 24730 -14721 25000 -14679
rect 24730 -14839 24809 -14721
rect 24927 -14839 25000 -14721
rect 24730 -14881 25000 -14839
rect 24730 -14999 24809 -14881
rect 24927 -14999 25000 -14881
rect 24730 -15041 25000 -14999
rect 24730 -15159 24809 -15041
rect 24927 -15159 25000 -15041
rect 24730 -15201 25000 -15159
rect 24730 -15230 24809 -15201
rect 21194 -15306 24809 -15230
rect 21194 -15319 21261 -15306
rect 21000 -15424 21261 -15319
rect 21379 -15424 21421 -15306
rect 21539 -15424 21581 -15306
rect 21699 -15424 21741 -15306
rect 21859 -15424 21901 -15306
rect 22019 -15424 22061 -15306
rect 22179 -15424 22221 -15306
rect 22339 -15424 22381 -15306
rect 22499 -15424 22541 -15306
rect 22659 -15424 22701 -15306
rect 22819 -15424 22861 -15306
rect 22979 -15424 23021 -15306
rect 23139 -15424 23181 -15306
rect 23299 -15424 23341 -15306
rect 23459 -15424 23501 -15306
rect 23619 -15424 23661 -15306
rect 23779 -15424 23821 -15306
rect 23939 -15424 23981 -15306
rect 24099 -15424 24141 -15306
rect 24259 -15424 24301 -15306
rect 24419 -15424 24461 -15306
rect 24579 -15424 24621 -15306
rect 24739 -15319 24809 -15306
rect 24927 -15319 25000 -15201
rect 24739 -15424 25000 -15319
rect 21000 -15500 25000 -15424
<< via4 >>
rect 3261 -5621 3379 -5578
rect 3261 -5653 3304 -5621
rect 3304 -5653 3336 -5621
rect 3336 -5653 3379 -5621
rect 3076 -5724 3194 -5681
rect 3261 -5696 3379 -5653
rect 3421 -5621 3539 -5578
rect 3421 -5653 3464 -5621
rect 3464 -5653 3496 -5621
rect 3496 -5653 3539 -5621
rect 3421 -5696 3539 -5653
rect 3581 -5621 3699 -5578
rect 3581 -5653 3624 -5621
rect 3624 -5653 3656 -5621
rect 3656 -5653 3699 -5621
rect 3581 -5696 3699 -5653
rect 3741 -5621 3859 -5578
rect 3741 -5653 3784 -5621
rect 3784 -5653 3816 -5621
rect 3816 -5653 3859 -5621
rect 3741 -5696 3859 -5653
rect 3901 -5621 4019 -5578
rect 3901 -5653 3944 -5621
rect 3944 -5653 3976 -5621
rect 3976 -5653 4019 -5621
rect 3901 -5696 4019 -5653
rect 4061 -5621 4179 -5578
rect 4061 -5653 4104 -5621
rect 4104 -5653 4136 -5621
rect 4136 -5653 4179 -5621
rect 4061 -5696 4179 -5653
rect 4221 -5621 4339 -5578
rect 4221 -5653 4264 -5621
rect 4264 -5653 4296 -5621
rect 4296 -5653 4339 -5621
rect 4221 -5696 4339 -5653
rect 4381 -5621 4499 -5578
rect 4381 -5653 4424 -5621
rect 4424 -5653 4456 -5621
rect 4456 -5653 4499 -5621
rect 4381 -5696 4499 -5653
rect 4541 -5621 4659 -5578
rect 4541 -5653 4584 -5621
rect 4584 -5653 4616 -5621
rect 4616 -5653 4659 -5621
rect 4541 -5696 4659 -5653
rect 4701 -5621 4819 -5578
rect 4701 -5653 4744 -5621
rect 4744 -5653 4776 -5621
rect 4776 -5653 4819 -5621
rect 4701 -5696 4819 -5653
rect 4861 -5621 4979 -5578
rect 4861 -5653 4904 -5621
rect 4904 -5653 4936 -5621
rect 4936 -5653 4979 -5621
rect 4861 -5696 4979 -5653
rect 5021 -5621 5139 -5578
rect 5021 -5653 5064 -5621
rect 5064 -5653 5096 -5621
rect 5096 -5653 5139 -5621
rect 5021 -5696 5139 -5653
rect 5181 -5621 5299 -5578
rect 5181 -5653 5224 -5621
rect 5224 -5653 5256 -5621
rect 5256 -5653 5299 -5621
rect 5181 -5696 5299 -5653
rect 5341 -5621 5459 -5578
rect 5341 -5653 5384 -5621
rect 5384 -5653 5416 -5621
rect 5416 -5653 5459 -5621
rect 5341 -5696 5459 -5653
rect 5501 -5621 5619 -5578
rect 5501 -5653 5544 -5621
rect 5544 -5653 5576 -5621
rect 5576 -5653 5619 -5621
rect 5501 -5696 5619 -5653
rect 5661 -5621 5779 -5578
rect 5661 -5653 5704 -5621
rect 5704 -5653 5736 -5621
rect 5736 -5653 5779 -5621
rect 5661 -5696 5779 -5653
rect 5821 -5621 5939 -5578
rect 5821 -5653 5864 -5621
rect 5864 -5653 5896 -5621
rect 5896 -5653 5939 -5621
rect 5821 -5696 5939 -5653
rect 5981 -5621 6099 -5578
rect 5981 -5653 6024 -5621
rect 6024 -5653 6056 -5621
rect 6056 -5653 6099 -5621
rect 5981 -5696 6099 -5653
rect 6141 -5621 6259 -5578
rect 6141 -5653 6184 -5621
rect 6184 -5653 6216 -5621
rect 6216 -5653 6259 -5621
rect 6141 -5696 6259 -5653
rect 6301 -5621 6419 -5578
rect 6301 -5653 6344 -5621
rect 6344 -5653 6376 -5621
rect 6376 -5653 6419 -5621
rect 6301 -5696 6419 -5653
rect 6461 -5621 6579 -5578
rect 6461 -5653 6504 -5621
rect 6504 -5653 6536 -5621
rect 6536 -5653 6579 -5621
rect 6461 -5696 6579 -5653
rect 6621 -5621 6739 -5578
rect 6621 -5653 6664 -5621
rect 6664 -5653 6696 -5621
rect 6696 -5653 6739 -5621
rect 6621 -5696 6739 -5653
rect 3076 -5756 3119 -5724
rect 3119 -5756 3151 -5724
rect 3151 -5756 3194 -5724
rect 3076 -5799 3194 -5756
rect 6809 -5724 6927 -5681
rect 6809 -5756 6852 -5724
rect 6852 -5756 6884 -5724
rect 6884 -5756 6927 -5724
rect 3076 -5884 3194 -5841
rect 3076 -5916 3119 -5884
rect 3119 -5916 3151 -5884
rect 3151 -5916 3194 -5884
rect 3076 -5959 3194 -5916
rect 3076 -6044 3194 -6001
rect 3076 -6076 3119 -6044
rect 3119 -6076 3151 -6044
rect 3151 -6076 3194 -6044
rect 3076 -6119 3194 -6076
rect 3076 -6204 3194 -6161
rect 3076 -6236 3119 -6204
rect 3119 -6236 3151 -6204
rect 3151 -6236 3194 -6204
rect 3076 -6279 3194 -6236
rect 3076 -6364 3194 -6321
rect 3076 -6396 3119 -6364
rect 3119 -6396 3151 -6364
rect 3151 -6396 3194 -6364
rect 3076 -6439 3194 -6396
rect 3076 -6524 3194 -6481
rect 3076 -6556 3119 -6524
rect 3119 -6556 3151 -6524
rect 3151 -6556 3194 -6524
rect 3076 -6599 3194 -6556
rect 3076 -6684 3194 -6641
rect 3076 -6716 3119 -6684
rect 3119 -6716 3151 -6684
rect 3151 -6716 3194 -6684
rect 3076 -6759 3194 -6716
rect 3076 -6844 3194 -6801
rect 3076 -6876 3119 -6844
rect 3119 -6876 3151 -6844
rect 3151 -6876 3194 -6844
rect 3076 -6919 3194 -6876
rect 3076 -7004 3194 -6961
rect 3076 -7036 3119 -7004
rect 3119 -7036 3151 -7004
rect 3151 -7036 3194 -7004
rect 3076 -7079 3194 -7036
rect 3076 -7164 3194 -7121
rect 3076 -7196 3119 -7164
rect 3119 -7196 3151 -7164
rect 3151 -7196 3194 -7164
rect 3076 -7239 3194 -7196
rect 3076 -7324 3194 -7281
rect 3076 -7356 3119 -7324
rect 3119 -7356 3151 -7324
rect 3151 -7356 3194 -7324
rect 3076 -7399 3194 -7356
rect 3076 -7484 3194 -7441
rect 3076 -7516 3119 -7484
rect 3119 -7516 3151 -7484
rect 3151 -7516 3194 -7484
rect 3076 -7559 3194 -7516
rect 3076 -7644 3194 -7601
rect 3076 -7676 3119 -7644
rect 3119 -7676 3151 -7644
rect 3151 -7676 3194 -7644
rect 3076 -7719 3194 -7676
rect 3076 -7804 3194 -7761
rect 3076 -7836 3119 -7804
rect 3119 -7836 3151 -7804
rect 3151 -7836 3194 -7804
rect 3076 -7879 3194 -7836
rect 3076 -7964 3194 -7921
rect 3076 -7996 3119 -7964
rect 3119 -7996 3151 -7964
rect 3151 -7996 3194 -7964
rect 3076 -8039 3194 -7996
rect 3076 -8124 3194 -8081
rect 3076 -8156 3119 -8124
rect 3119 -8156 3151 -8124
rect 3151 -8156 3194 -8124
rect 3076 -8199 3194 -8156
rect 3076 -8284 3194 -8241
rect 3076 -8316 3119 -8284
rect 3119 -8316 3151 -8284
rect 3151 -8316 3194 -8284
rect 3076 -8359 3194 -8316
rect 3076 -8444 3194 -8401
rect 3076 -8476 3119 -8444
rect 3119 -8476 3151 -8444
rect 3151 -8476 3194 -8444
rect 3076 -8519 3194 -8476
rect 3076 -8604 3194 -8561
rect 3076 -8636 3119 -8604
rect 3119 -8636 3151 -8604
rect 3151 -8636 3194 -8604
rect 3076 -8679 3194 -8636
rect 3076 -8764 3194 -8721
rect 3076 -8796 3119 -8764
rect 3119 -8796 3151 -8764
rect 3151 -8796 3194 -8764
rect 3076 -8839 3194 -8796
rect 3076 -8924 3194 -8881
rect 3076 -8956 3119 -8924
rect 3119 -8956 3151 -8924
rect 3151 -8956 3194 -8924
rect 3076 -8999 3194 -8956
rect 3076 -9084 3194 -9041
rect 3076 -9116 3119 -9084
rect 3119 -9116 3151 -9084
rect 3151 -9116 3194 -9084
rect 3076 -9159 3194 -9116
rect 3076 -9244 3194 -9201
rect 6809 -5799 6927 -5756
rect 6809 -5884 6927 -5841
rect 6809 -5916 6852 -5884
rect 6852 -5916 6884 -5884
rect 6884 -5916 6927 -5884
rect 6809 -5959 6927 -5916
rect 6809 -6044 6927 -6001
rect 6809 -6076 6852 -6044
rect 6852 -6076 6884 -6044
rect 6884 -6076 6927 -6044
rect 6809 -6119 6927 -6076
rect 6809 -6204 6927 -6161
rect 6809 -6236 6852 -6204
rect 6852 -6236 6884 -6204
rect 6884 -6236 6927 -6204
rect 6809 -6279 6927 -6236
rect 6809 -6364 6927 -6321
rect 6809 -6396 6852 -6364
rect 6852 -6396 6884 -6364
rect 6884 -6396 6927 -6364
rect 6809 -6439 6927 -6396
rect 6809 -6524 6927 -6481
rect 6809 -6556 6852 -6524
rect 6852 -6556 6884 -6524
rect 6884 -6556 6927 -6524
rect 6809 -6599 6927 -6556
rect 6809 -6684 6927 -6641
rect 6809 -6716 6852 -6684
rect 6852 -6716 6884 -6684
rect 6884 -6716 6927 -6684
rect 6809 -6759 6927 -6716
rect 6809 -6844 6927 -6801
rect 6809 -6876 6852 -6844
rect 6852 -6876 6884 -6844
rect 6884 -6876 6927 -6844
rect 6809 -6919 6927 -6876
rect 6809 -7004 6927 -6961
rect 6809 -7036 6852 -7004
rect 6852 -7036 6884 -7004
rect 6884 -7036 6927 -7004
rect 6809 -7079 6927 -7036
rect 6809 -7164 6927 -7121
rect 6809 -7196 6852 -7164
rect 6852 -7196 6884 -7164
rect 6884 -7196 6927 -7164
rect 6809 -7239 6927 -7196
rect 6809 -7324 6927 -7281
rect 6809 -7356 6852 -7324
rect 6852 -7356 6884 -7324
rect 6884 -7356 6927 -7324
rect 6809 -7399 6927 -7356
rect 6809 -7484 6927 -7441
rect 6809 -7516 6852 -7484
rect 6852 -7516 6884 -7484
rect 6884 -7516 6927 -7484
rect 6809 -7559 6927 -7516
rect 6809 -7644 6927 -7601
rect 6809 -7676 6852 -7644
rect 6852 -7676 6884 -7644
rect 6884 -7676 6927 -7644
rect 6809 -7719 6927 -7676
rect 6809 -7804 6927 -7761
rect 6809 -7836 6852 -7804
rect 6852 -7836 6884 -7804
rect 6884 -7836 6927 -7804
rect 6809 -7879 6927 -7836
rect 6809 -7964 6927 -7921
rect 6809 -7996 6852 -7964
rect 6852 -7996 6884 -7964
rect 6884 -7996 6927 -7964
rect 6809 -8039 6927 -7996
rect 6809 -8124 6927 -8081
rect 6809 -8156 6852 -8124
rect 6852 -8156 6884 -8124
rect 6884 -8156 6927 -8124
rect 6809 -8199 6927 -8156
rect 6809 -8284 6927 -8241
rect 6809 -8316 6852 -8284
rect 6852 -8316 6884 -8284
rect 6884 -8316 6927 -8284
rect 6809 -8359 6927 -8316
rect 6809 -8444 6927 -8401
rect 6809 -8476 6852 -8444
rect 6852 -8476 6884 -8444
rect 6884 -8476 6927 -8444
rect 6809 -8519 6927 -8476
rect 6809 -8604 6927 -8561
rect 6809 -8636 6852 -8604
rect 6852 -8636 6884 -8604
rect 6884 -8636 6927 -8604
rect 6809 -8679 6927 -8636
rect 6809 -8764 6927 -8721
rect 6809 -8796 6852 -8764
rect 6852 -8796 6884 -8764
rect 6884 -8796 6927 -8764
rect 6809 -8839 6927 -8796
rect 6809 -8924 6927 -8881
rect 6809 -8956 6852 -8924
rect 6852 -8956 6884 -8924
rect 6884 -8956 6927 -8924
rect 6809 -8999 6927 -8956
rect 6809 -9084 6927 -9041
rect 6809 -9116 6852 -9084
rect 6852 -9116 6884 -9084
rect 6884 -9116 6927 -9084
rect 6809 -9159 6927 -9116
rect 3076 -9276 3119 -9244
rect 3119 -9276 3151 -9244
rect 3151 -9276 3194 -9244
rect 3076 -9319 3194 -9276
rect 6809 -9244 6927 -9201
rect 6809 -9276 6852 -9244
rect 6852 -9276 6884 -9244
rect 6884 -9276 6927 -9244
rect 3261 -9349 3379 -9306
rect 3261 -9381 3304 -9349
rect 3304 -9381 3336 -9349
rect 3336 -9381 3379 -9349
rect 3261 -9424 3379 -9381
rect 3421 -9349 3539 -9306
rect 3421 -9381 3464 -9349
rect 3464 -9381 3496 -9349
rect 3496 -9381 3539 -9349
rect 3421 -9424 3539 -9381
rect 3581 -9349 3699 -9306
rect 3581 -9381 3624 -9349
rect 3624 -9381 3656 -9349
rect 3656 -9381 3699 -9349
rect 3581 -9424 3699 -9381
rect 3741 -9349 3859 -9306
rect 3741 -9381 3784 -9349
rect 3784 -9381 3816 -9349
rect 3816 -9381 3859 -9349
rect 3741 -9424 3859 -9381
rect 3901 -9349 4019 -9306
rect 3901 -9381 3944 -9349
rect 3944 -9381 3976 -9349
rect 3976 -9381 4019 -9349
rect 3901 -9424 4019 -9381
rect 4061 -9349 4179 -9306
rect 4061 -9381 4104 -9349
rect 4104 -9381 4136 -9349
rect 4136 -9381 4179 -9349
rect 4061 -9424 4179 -9381
rect 4221 -9349 4339 -9306
rect 4221 -9381 4264 -9349
rect 4264 -9381 4296 -9349
rect 4296 -9381 4339 -9349
rect 4221 -9424 4339 -9381
rect 4381 -9349 4499 -9306
rect 4381 -9381 4424 -9349
rect 4424 -9381 4456 -9349
rect 4456 -9381 4499 -9349
rect 4381 -9424 4499 -9381
rect 4541 -9349 4659 -9306
rect 4541 -9381 4584 -9349
rect 4584 -9381 4616 -9349
rect 4616 -9381 4659 -9349
rect 4541 -9424 4659 -9381
rect 4701 -9349 4819 -9306
rect 4701 -9381 4744 -9349
rect 4744 -9381 4776 -9349
rect 4776 -9381 4819 -9349
rect 4701 -9424 4819 -9381
rect 4861 -9349 4979 -9306
rect 4861 -9381 4904 -9349
rect 4904 -9381 4936 -9349
rect 4936 -9381 4979 -9349
rect 4861 -9424 4979 -9381
rect 5021 -9349 5139 -9306
rect 5021 -9381 5064 -9349
rect 5064 -9381 5096 -9349
rect 5096 -9381 5139 -9349
rect 5021 -9424 5139 -9381
rect 5181 -9349 5299 -9306
rect 5181 -9381 5224 -9349
rect 5224 -9381 5256 -9349
rect 5256 -9381 5299 -9349
rect 5181 -9424 5299 -9381
rect 5341 -9349 5459 -9306
rect 5341 -9381 5384 -9349
rect 5384 -9381 5416 -9349
rect 5416 -9381 5459 -9349
rect 5341 -9424 5459 -9381
rect 5501 -9349 5619 -9306
rect 5501 -9381 5544 -9349
rect 5544 -9381 5576 -9349
rect 5576 -9381 5619 -9349
rect 5501 -9424 5619 -9381
rect 5661 -9349 5779 -9306
rect 5661 -9381 5704 -9349
rect 5704 -9381 5736 -9349
rect 5736 -9381 5779 -9349
rect 5661 -9424 5779 -9381
rect 5821 -9349 5939 -9306
rect 5821 -9381 5864 -9349
rect 5864 -9381 5896 -9349
rect 5896 -9381 5939 -9349
rect 5821 -9424 5939 -9381
rect 5981 -9349 6099 -9306
rect 5981 -9381 6024 -9349
rect 6024 -9381 6056 -9349
rect 6056 -9381 6099 -9349
rect 5981 -9424 6099 -9381
rect 6141 -9349 6259 -9306
rect 6141 -9381 6184 -9349
rect 6184 -9381 6216 -9349
rect 6216 -9381 6259 -9349
rect 6141 -9424 6259 -9381
rect 6301 -9349 6419 -9306
rect 6301 -9381 6344 -9349
rect 6344 -9381 6376 -9349
rect 6376 -9381 6419 -9349
rect 6301 -9424 6419 -9381
rect 6461 -9349 6579 -9306
rect 6461 -9381 6504 -9349
rect 6504 -9381 6536 -9349
rect 6536 -9381 6579 -9349
rect 6461 -9424 6579 -9381
rect 6621 -9349 6739 -9306
rect 6809 -9319 6927 -9276
rect 6621 -9381 6664 -9349
rect 6664 -9381 6696 -9349
rect 6696 -9381 6739 -9349
rect 6621 -9424 6739 -9381
rect 9261 -5621 9379 -5578
rect 9261 -5653 9304 -5621
rect 9304 -5653 9336 -5621
rect 9336 -5653 9379 -5621
rect 9076 -5724 9194 -5681
rect 9261 -5696 9379 -5653
rect 9421 -5621 9539 -5578
rect 9421 -5653 9464 -5621
rect 9464 -5653 9496 -5621
rect 9496 -5653 9539 -5621
rect 9421 -5696 9539 -5653
rect 9581 -5621 9699 -5578
rect 9581 -5653 9624 -5621
rect 9624 -5653 9656 -5621
rect 9656 -5653 9699 -5621
rect 9581 -5696 9699 -5653
rect 9741 -5621 9859 -5578
rect 9741 -5653 9784 -5621
rect 9784 -5653 9816 -5621
rect 9816 -5653 9859 -5621
rect 9741 -5696 9859 -5653
rect 9901 -5621 10019 -5578
rect 9901 -5653 9944 -5621
rect 9944 -5653 9976 -5621
rect 9976 -5653 10019 -5621
rect 9901 -5696 10019 -5653
rect 10061 -5621 10179 -5578
rect 10061 -5653 10104 -5621
rect 10104 -5653 10136 -5621
rect 10136 -5653 10179 -5621
rect 10061 -5696 10179 -5653
rect 10221 -5621 10339 -5578
rect 10221 -5653 10264 -5621
rect 10264 -5653 10296 -5621
rect 10296 -5653 10339 -5621
rect 10221 -5696 10339 -5653
rect 10381 -5621 10499 -5578
rect 10381 -5653 10424 -5621
rect 10424 -5653 10456 -5621
rect 10456 -5653 10499 -5621
rect 10381 -5696 10499 -5653
rect 10541 -5621 10659 -5578
rect 10541 -5653 10584 -5621
rect 10584 -5653 10616 -5621
rect 10616 -5653 10659 -5621
rect 10541 -5696 10659 -5653
rect 10701 -5621 10819 -5578
rect 10701 -5653 10744 -5621
rect 10744 -5653 10776 -5621
rect 10776 -5653 10819 -5621
rect 10701 -5696 10819 -5653
rect 10861 -5621 10979 -5578
rect 10861 -5653 10904 -5621
rect 10904 -5653 10936 -5621
rect 10936 -5653 10979 -5621
rect 10861 -5696 10979 -5653
rect 11021 -5621 11139 -5578
rect 11021 -5653 11064 -5621
rect 11064 -5653 11096 -5621
rect 11096 -5653 11139 -5621
rect 11021 -5696 11139 -5653
rect 11181 -5621 11299 -5578
rect 11181 -5653 11224 -5621
rect 11224 -5653 11256 -5621
rect 11256 -5653 11299 -5621
rect 11181 -5696 11299 -5653
rect 11341 -5621 11459 -5578
rect 11341 -5653 11384 -5621
rect 11384 -5653 11416 -5621
rect 11416 -5653 11459 -5621
rect 11341 -5696 11459 -5653
rect 11501 -5621 11619 -5578
rect 11501 -5653 11544 -5621
rect 11544 -5653 11576 -5621
rect 11576 -5653 11619 -5621
rect 11501 -5696 11619 -5653
rect 11661 -5621 11779 -5578
rect 11661 -5653 11704 -5621
rect 11704 -5653 11736 -5621
rect 11736 -5653 11779 -5621
rect 11661 -5696 11779 -5653
rect 11821 -5621 11939 -5578
rect 11821 -5653 11864 -5621
rect 11864 -5653 11896 -5621
rect 11896 -5653 11939 -5621
rect 11821 -5696 11939 -5653
rect 11981 -5621 12099 -5578
rect 11981 -5653 12024 -5621
rect 12024 -5653 12056 -5621
rect 12056 -5653 12099 -5621
rect 11981 -5696 12099 -5653
rect 12141 -5621 12259 -5578
rect 12141 -5653 12184 -5621
rect 12184 -5653 12216 -5621
rect 12216 -5653 12259 -5621
rect 12141 -5696 12259 -5653
rect 12301 -5621 12419 -5578
rect 12301 -5653 12344 -5621
rect 12344 -5653 12376 -5621
rect 12376 -5653 12419 -5621
rect 12301 -5696 12419 -5653
rect 12461 -5621 12579 -5578
rect 12461 -5653 12504 -5621
rect 12504 -5653 12536 -5621
rect 12536 -5653 12579 -5621
rect 12461 -5696 12579 -5653
rect 12621 -5621 12739 -5578
rect 12621 -5653 12664 -5621
rect 12664 -5653 12696 -5621
rect 12696 -5653 12739 -5621
rect 12621 -5696 12739 -5653
rect 9076 -5756 9119 -5724
rect 9119 -5756 9151 -5724
rect 9151 -5756 9194 -5724
rect 9076 -5799 9194 -5756
rect 12809 -5724 12927 -5681
rect 12809 -5756 12852 -5724
rect 12852 -5756 12884 -5724
rect 12884 -5756 12927 -5724
rect 9076 -5884 9194 -5841
rect 9076 -5916 9119 -5884
rect 9119 -5916 9151 -5884
rect 9151 -5916 9194 -5884
rect 9076 -5959 9194 -5916
rect 9076 -6044 9194 -6001
rect 9076 -6076 9119 -6044
rect 9119 -6076 9151 -6044
rect 9151 -6076 9194 -6044
rect 9076 -6119 9194 -6076
rect 9076 -6204 9194 -6161
rect 9076 -6236 9119 -6204
rect 9119 -6236 9151 -6204
rect 9151 -6236 9194 -6204
rect 9076 -6279 9194 -6236
rect 9076 -6364 9194 -6321
rect 9076 -6396 9119 -6364
rect 9119 -6396 9151 -6364
rect 9151 -6396 9194 -6364
rect 9076 -6439 9194 -6396
rect 9076 -6524 9194 -6481
rect 9076 -6556 9119 -6524
rect 9119 -6556 9151 -6524
rect 9151 -6556 9194 -6524
rect 9076 -6599 9194 -6556
rect 9076 -6684 9194 -6641
rect 9076 -6716 9119 -6684
rect 9119 -6716 9151 -6684
rect 9151 -6716 9194 -6684
rect 9076 -6759 9194 -6716
rect 9076 -6844 9194 -6801
rect 9076 -6876 9119 -6844
rect 9119 -6876 9151 -6844
rect 9151 -6876 9194 -6844
rect 9076 -6919 9194 -6876
rect 9076 -7004 9194 -6961
rect 9076 -7036 9119 -7004
rect 9119 -7036 9151 -7004
rect 9151 -7036 9194 -7004
rect 9076 -7079 9194 -7036
rect 9076 -7164 9194 -7121
rect 9076 -7196 9119 -7164
rect 9119 -7196 9151 -7164
rect 9151 -7196 9194 -7164
rect 9076 -7239 9194 -7196
rect 9076 -7324 9194 -7281
rect 9076 -7356 9119 -7324
rect 9119 -7356 9151 -7324
rect 9151 -7356 9194 -7324
rect 9076 -7399 9194 -7356
rect 9076 -7484 9194 -7441
rect 9076 -7516 9119 -7484
rect 9119 -7516 9151 -7484
rect 9151 -7516 9194 -7484
rect 9076 -7559 9194 -7516
rect 9076 -7644 9194 -7601
rect 9076 -7676 9119 -7644
rect 9119 -7676 9151 -7644
rect 9151 -7676 9194 -7644
rect 9076 -7719 9194 -7676
rect 9076 -7804 9194 -7761
rect 9076 -7836 9119 -7804
rect 9119 -7836 9151 -7804
rect 9151 -7836 9194 -7804
rect 9076 -7879 9194 -7836
rect 9076 -7964 9194 -7921
rect 9076 -7996 9119 -7964
rect 9119 -7996 9151 -7964
rect 9151 -7996 9194 -7964
rect 9076 -8039 9194 -7996
rect 9076 -8124 9194 -8081
rect 9076 -8156 9119 -8124
rect 9119 -8156 9151 -8124
rect 9151 -8156 9194 -8124
rect 9076 -8199 9194 -8156
rect 9076 -8284 9194 -8241
rect 9076 -8316 9119 -8284
rect 9119 -8316 9151 -8284
rect 9151 -8316 9194 -8284
rect 9076 -8359 9194 -8316
rect 9076 -8444 9194 -8401
rect 9076 -8476 9119 -8444
rect 9119 -8476 9151 -8444
rect 9151 -8476 9194 -8444
rect 9076 -8519 9194 -8476
rect 9076 -8604 9194 -8561
rect 9076 -8636 9119 -8604
rect 9119 -8636 9151 -8604
rect 9151 -8636 9194 -8604
rect 9076 -8679 9194 -8636
rect 9076 -8764 9194 -8721
rect 9076 -8796 9119 -8764
rect 9119 -8796 9151 -8764
rect 9151 -8796 9194 -8764
rect 9076 -8839 9194 -8796
rect 9076 -8924 9194 -8881
rect 9076 -8956 9119 -8924
rect 9119 -8956 9151 -8924
rect 9151 -8956 9194 -8924
rect 9076 -8999 9194 -8956
rect 9076 -9084 9194 -9041
rect 9076 -9116 9119 -9084
rect 9119 -9116 9151 -9084
rect 9151 -9116 9194 -9084
rect 9076 -9159 9194 -9116
rect 9076 -9244 9194 -9201
rect 12809 -5799 12927 -5756
rect 12809 -5884 12927 -5841
rect 12809 -5916 12852 -5884
rect 12852 -5916 12884 -5884
rect 12884 -5916 12927 -5884
rect 12809 -5959 12927 -5916
rect 12809 -6044 12927 -6001
rect 12809 -6076 12852 -6044
rect 12852 -6076 12884 -6044
rect 12884 -6076 12927 -6044
rect 12809 -6119 12927 -6076
rect 12809 -6204 12927 -6161
rect 12809 -6236 12852 -6204
rect 12852 -6236 12884 -6204
rect 12884 -6236 12927 -6204
rect 12809 -6279 12927 -6236
rect 12809 -6364 12927 -6321
rect 12809 -6396 12852 -6364
rect 12852 -6396 12884 -6364
rect 12884 -6396 12927 -6364
rect 12809 -6439 12927 -6396
rect 12809 -6524 12927 -6481
rect 12809 -6556 12852 -6524
rect 12852 -6556 12884 -6524
rect 12884 -6556 12927 -6524
rect 12809 -6599 12927 -6556
rect 12809 -6684 12927 -6641
rect 12809 -6716 12852 -6684
rect 12852 -6716 12884 -6684
rect 12884 -6716 12927 -6684
rect 12809 -6759 12927 -6716
rect 12809 -6844 12927 -6801
rect 12809 -6876 12852 -6844
rect 12852 -6876 12884 -6844
rect 12884 -6876 12927 -6844
rect 12809 -6919 12927 -6876
rect 12809 -7004 12927 -6961
rect 12809 -7036 12852 -7004
rect 12852 -7036 12884 -7004
rect 12884 -7036 12927 -7004
rect 12809 -7079 12927 -7036
rect 12809 -7164 12927 -7121
rect 12809 -7196 12852 -7164
rect 12852 -7196 12884 -7164
rect 12884 -7196 12927 -7164
rect 12809 -7239 12927 -7196
rect 12809 -7324 12927 -7281
rect 12809 -7356 12852 -7324
rect 12852 -7356 12884 -7324
rect 12884 -7356 12927 -7324
rect 12809 -7399 12927 -7356
rect 12809 -7484 12927 -7441
rect 12809 -7516 12852 -7484
rect 12852 -7516 12884 -7484
rect 12884 -7516 12927 -7484
rect 12809 -7559 12927 -7516
rect 12809 -7644 12927 -7601
rect 12809 -7676 12852 -7644
rect 12852 -7676 12884 -7644
rect 12884 -7676 12927 -7644
rect 12809 -7719 12927 -7676
rect 12809 -7804 12927 -7761
rect 12809 -7836 12852 -7804
rect 12852 -7836 12884 -7804
rect 12884 -7836 12927 -7804
rect 12809 -7879 12927 -7836
rect 12809 -7964 12927 -7921
rect 12809 -7996 12852 -7964
rect 12852 -7996 12884 -7964
rect 12884 -7996 12927 -7964
rect 12809 -8039 12927 -7996
rect 12809 -8124 12927 -8081
rect 12809 -8156 12852 -8124
rect 12852 -8156 12884 -8124
rect 12884 -8156 12927 -8124
rect 12809 -8199 12927 -8156
rect 12809 -8284 12927 -8241
rect 12809 -8316 12852 -8284
rect 12852 -8316 12884 -8284
rect 12884 -8316 12927 -8284
rect 12809 -8359 12927 -8316
rect 12809 -8444 12927 -8401
rect 12809 -8476 12852 -8444
rect 12852 -8476 12884 -8444
rect 12884 -8476 12927 -8444
rect 12809 -8519 12927 -8476
rect 12809 -8604 12927 -8561
rect 12809 -8636 12852 -8604
rect 12852 -8636 12884 -8604
rect 12884 -8636 12927 -8604
rect 12809 -8679 12927 -8636
rect 12809 -8764 12927 -8721
rect 12809 -8796 12852 -8764
rect 12852 -8796 12884 -8764
rect 12884 -8796 12927 -8764
rect 12809 -8839 12927 -8796
rect 12809 -8924 12927 -8881
rect 12809 -8956 12852 -8924
rect 12852 -8956 12884 -8924
rect 12884 -8956 12927 -8924
rect 12809 -8999 12927 -8956
rect 12809 -9084 12927 -9041
rect 12809 -9116 12852 -9084
rect 12852 -9116 12884 -9084
rect 12884 -9116 12927 -9084
rect 12809 -9159 12927 -9116
rect 9076 -9276 9119 -9244
rect 9119 -9276 9151 -9244
rect 9151 -9276 9194 -9244
rect 9076 -9319 9194 -9276
rect 12809 -9244 12927 -9201
rect 12809 -9276 12852 -9244
rect 12852 -9276 12884 -9244
rect 12884 -9276 12927 -9244
rect 9261 -9349 9379 -9306
rect 9261 -9381 9304 -9349
rect 9304 -9381 9336 -9349
rect 9336 -9381 9379 -9349
rect 9261 -9424 9379 -9381
rect 9421 -9349 9539 -9306
rect 9421 -9381 9464 -9349
rect 9464 -9381 9496 -9349
rect 9496 -9381 9539 -9349
rect 9421 -9424 9539 -9381
rect 9581 -9349 9699 -9306
rect 9581 -9381 9624 -9349
rect 9624 -9381 9656 -9349
rect 9656 -9381 9699 -9349
rect 9581 -9424 9699 -9381
rect 9741 -9349 9859 -9306
rect 9741 -9381 9784 -9349
rect 9784 -9381 9816 -9349
rect 9816 -9381 9859 -9349
rect 9741 -9424 9859 -9381
rect 9901 -9349 10019 -9306
rect 9901 -9381 9944 -9349
rect 9944 -9381 9976 -9349
rect 9976 -9381 10019 -9349
rect 9901 -9424 10019 -9381
rect 10061 -9349 10179 -9306
rect 10061 -9381 10104 -9349
rect 10104 -9381 10136 -9349
rect 10136 -9381 10179 -9349
rect 10061 -9424 10179 -9381
rect 10221 -9349 10339 -9306
rect 10221 -9381 10264 -9349
rect 10264 -9381 10296 -9349
rect 10296 -9381 10339 -9349
rect 10221 -9424 10339 -9381
rect 10381 -9349 10499 -9306
rect 10381 -9381 10424 -9349
rect 10424 -9381 10456 -9349
rect 10456 -9381 10499 -9349
rect 10381 -9424 10499 -9381
rect 10541 -9349 10659 -9306
rect 10541 -9381 10584 -9349
rect 10584 -9381 10616 -9349
rect 10616 -9381 10659 -9349
rect 10541 -9424 10659 -9381
rect 10701 -9349 10819 -9306
rect 10701 -9381 10744 -9349
rect 10744 -9381 10776 -9349
rect 10776 -9381 10819 -9349
rect 10701 -9424 10819 -9381
rect 10861 -9349 10979 -9306
rect 10861 -9381 10904 -9349
rect 10904 -9381 10936 -9349
rect 10936 -9381 10979 -9349
rect 10861 -9424 10979 -9381
rect 11021 -9349 11139 -9306
rect 11021 -9381 11064 -9349
rect 11064 -9381 11096 -9349
rect 11096 -9381 11139 -9349
rect 11021 -9424 11139 -9381
rect 11181 -9349 11299 -9306
rect 11181 -9381 11224 -9349
rect 11224 -9381 11256 -9349
rect 11256 -9381 11299 -9349
rect 11181 -9424 11299 -9381
rect 11341 -9349 11459 -9306
rect 11341 -9381 11384 -9349
rect 11384 -9381 11416 -9349
rect 11416 -9381 11459 -9349
rect 11341 -9424 11459 -9381
rect 11501 -9349 11619 -9306
rect 11501 -9381 11544 -9349
rect 11544 -9381 11576 -9349
rect 11576 -9381 11619 -9349
rect 11501 -9424 11619 -9381
rect 11661 -9349 11779 -9306
rect 11661 -9381 11704 -9349
rect 11704 -9381 11736 -9349
rect 11736 -9381 11779 -9349
rect 11661 -9424 11779 -9381
rect 11821 -9349 11939 -9306
rect 11821 -9381 11864 -9349
rect 11864 -9381 11896 -9349
rect 11896 -9381 11939 -9349
rect 11821 -9424 11939 -9381
rect 11981 -9349 12099 -9306
rect 11981 -9381 12024 -9349
rect 12024 -9381 12056 -9349
rect 12056 -9381 12099 -9349
rect 11981 -9424 12099 -9381
rect 12141 -9349 12259 -9306
rect 12141 -9381 12184 -9349
rect 12184 -9381 12216 -9349
rect 12216 -9381 12259 -9349
rect 12141 -9424 12259 -9381
rect 12301 -9349 12419 -9306
rect 12301 -9381 12344 -9349
rect 12344 -9381 12376 -9349
rect 12376 -9381 12419 -9349
rect 12301 -9424 12419 -9381
rect 12461 -9349 12579 -9306
rect 12461 -9381 12504 -9349
rect 12504 -9381 12536 -9349
rect 12536 -9381 12579 -9349
rect 12461 -9424 12579 -9381
rect 12621 -9349 12739 -9306
rect 12809 -9319 12927 -9276
rect 12621 -9381 12664 -9349
rect 12664 -9381 12696 -9349
rect 12696 -9381 12739 -9349
rect 12621 -9424 12739 -9381
rect 15261 -5621 15379 -5578
rect 15261 -5653 15304 -5621
rect 15304 -5653 15336 -5621
rect 15336 -5653 15379 -5621
rect 15076 -5724 15194 -5681
rect 15261 -5696 15379 -5653
rect 15421 -5621 15539 -5578
rect 15421 -5653 15464 -5621
rect 15464 -5653 15496 -5621
rect 15496 -5653 15539 -5621
rect 15421 -5696 15539 -5653
rect 15581 -5621 15699 -5578
rect 15581 -5653 15624 -5621
rect 15624 -5653 15656 -5621
rect 15656 -5653 15699 -5621
rect 15581 -5696 15699 -5653
rect 15741 -5621 15859 -5578
rect 15741 -5653 15784 -5621
rect 15784 -5653 15816 -5621
rect 15816 -5653 15859 -5621
rect 15741 -5696 15859 -5653
rect 15901 -5621 16019 -5578
rect 15901 -5653 15944 -5621
rect 15944 -5653 15976 -5621
rect 15976 -5653 16019 -5621
rect 15901 -5696 16019 -5653
rect 16061 -5621 16179 -5578
rect 16061 -5653 16104 -5621
rect 16104 -5653 16136 -5621
rect 16136 -5653 16179 -5621
rect 16061 -5696 16179 -5653
rect 16221 -5621 16339 -5578
rect 16221 -5653 16264 -5621
rect 16264 -5653 16296 -5621
rect 16296 -5653 16339 -5621
rect 16221 -5696 16339 -5653
rect 16381 -5621 16499 -5578
rect 16381 -5653 16424 -5621
rect 16424 -5653 16456 -5621
rect 16456 -5653 16499 -5621
rect 16381 -5696 16499 -5653
rect 16541 -5621 16659 -5578
rect 16541 -5653 16584 -5621
rect 16584 -5653 16616 -5621
rect 16616 -5653 16659 -5621
rect 16541 -5696 16659 -5653
rect 16701 -5621 16819 -5578
rect 16701 -5653 16744 -5621
rect 16744 -5653 16776 -5621
rect 16776 -5653 16819 -5621
rect 16701 -5696 16819 -5653
rect 16861 -5621 16979 -5578
rect 16861 -5653 16904 -5621
rect 16904 -5653 16936 -5621
rect 16936 -5653 16979 -5621
rect 16861 -5696 16979 -5653
rect 17021 -5621 17139 -5578
rect 17021 -5653 17064 -5621
rect 17064 -5653 17096 -5621
rect 17096 -5653 17139 -5621
rect 17021 -5696 17139 -5653
rect 17181 -5621 17299 -5578
rect 17181 -5653 17224 -5621
rect 17224 -5653 17256 -5621
rect 17256 -5653 17299 -5621
rect 17181 -5696 17299 -5653
rect 17341 -5621 17459 -5578
rect 17341 -5653 17384 -5621
rect 17384 -5653 17416 -5621
rect 17416 -5653 17459 -5621
rect 17341 -5696 17459 -5653
rect 17501 -5621 17619 -5578
rect 17501 -5653 17544 -5621
rect 17544 -5653 17576 -5621
rect 17576 -5653 17619 -5621
rect 17501 -5696 17619 -5653
rect 17661 -5621 17779 -5578
rect 17661 -5653 17704 -5621
rect 17704 -5653 17736 -5621
rect 17736 -5653 17779 -5621
rect 17661 -5696 17779 -5653
rect 17821 -5621 17939 -5578
rect 17821 -5653 17864 -5621
rect 17864 -5653 17896 -5621
rect 17896 -5653 17939 -5621
rect 17821 -5696 17939 -5653
rect 17981 -5621 18099 -5578
rect 17981 -5653 18024 -5621
rect 18024 -5653 18056 -5621
rect 18056 -5653 18099 -5621
rect 17981 -5696 18099 -5653
rect 18141 -5621 18259 -5578
rect 18141 -5653 18184 -5621
rect 18184 -5653 18216 -5621
rect 18216 -5653 18259 -5621
rect 18141 -5696 18259 -5653
rect 18301 -5621 18419 -5578
rect 18301 -5653 18344 -5621
rect 18344 -5653 18376 -5621
rect 18376 -5653 18419 -5621
rect 18301 -5696 18419 -5653
rect 18461 -5621 18579 -5578
rect 18461 -5653 18504 -5621
rect 18504 -5653 18536 -5621
rect 18536 -5653 18579 -5621
rect 18461 -5696 18579 -5653
rect 18621 -5621 18739 -5578
rect 18621 -5653 18664 -5621
rect 18664 -5653 18696 -5621
rect 18696 -5653 18739 -5621
rect 18621 -5696 18739 -5653
rect 15076 -5756 15119 -5724
rect 15119 -5756 15151 -5724
rect 15151 -5756 15194 -5724
rect 15076 -5799 15194 -5756
rect 18809 -5724 18927 -5681
rect 18809 -5756 18852 -5724
rect 18852 -5756 18884 -5724
rect 18884 -5756 18927 -5724
rect 15076 -5884 15194 -5841
rect 15076 -5916 15119 -5884
rect 15119 -5916 15151 -5884
rect 15151 -5916 15194 -5884
rect 15076 -5959 15194 -5916
rect 15076 -6044 15194 -6001
rect 15076 -6076 15119 -6044
rect 15119 -6076 15151 -6044
rect 15151 -6076 15194 -6044
rect 15076 -6119 15194 -6076
rect 15076 -6204 15194 -6161
rect 15076 -6236 15119 -6204
rect 15119 -6236 15151 -6204
rect 15151 -6236 15194 -6204
rect 15076 -6279 15194 -6236
rect 15076 -6364 15194 -6321
rect 15076 -6396 15119 -6364
rect 15119 -6396 15151 -6364
rect 15151 -6396 15194 -6364
rect 15076 -6439 15194 -6396
rect 15076 -6524 15194 -6481
rect 15076 -6556 15119 -6524
rect 15119 -6556 15151 -6524
rect 15151 -6556 15194 -6524
rect 15076 -6599 15194 -6556
rect 15076 -6684 15194 -6641
rect 15076 -6716 15119 -6684
rect 15119 -6716 15151 -6684
rect 15151 -6716 15194 -6684
rect 15076 -6759 15194 -6716
rect 15076 -6844 15194 -6801
rect 15076 -6876 15119 -6844
rect 15119 -6876 15151 -6844
rect 15151 -6876 15194 -6844
rect 15076 -6919 15194 -6876
rect 15076 -7004 15194 -6961
rect 15076 -7036 15119 -7004
rect 15119 -7036 15151 -7004
rect 15151 -7036 15194 -7004
rect 15076 -7079 15194 -7036
rect 15076 -7164 15194 -7121
rect 15076 -7196 15119 -7164
rect 15119 -7196 15151 -7164
rect 15151 -7196 15194 -7164
rect 15076 -7239 15194 -7196
rect 15076 -7324 15194 -7281
rect 15076 -7356 15119 -7324
rect 15119 -7356 15151 -7324
rect 15151 -7356 15194 -7324
rect 15076 -7399 15194 -7356
rect 15076 -7484 15194 -7441
rect 15076 -7516 15119 -7484
rect 15119 -7516 15151 -7484
rect 15151 -7516 15194 -7484
rect 15076 -7559 15194 -7516
rect 15076 -7644 15194 -7601
rect 15076 -7676 15119 -7644
rect 15119 -7676 15151 -7644
rect 15151 -7676 15194 -7644
rect 15076 -7719 15194 -7676
rect 15076 -7804 15194 -7761
rect 15076 -7836 15119 -7804
rect 15119 -7836 15151 -7804
rect 15151 -7836 15194 -7804
rect 15076 -7879 15194 -7836
rect 15076 -7964 15194 -7921
rect 15076 -7996 15119 -7964
rect 15119 -7996 15151 -7964
rect 15151 -7996 15194 -7964
rect 15076 -8039 15194 -7996
rect 15076 -8124 15194 -8081
rect 15076 -8156 15119 -8124
rect 15119 -8156 15151 -8124
rect 15151 -8156 15194 -8124
rect 15076 -8199 15194 -8156
rect 15076 -8284 15194 -8241
rect 15076 -8316 15119 -8284
rect 15119 -8316 15151 -8284
rect 15151 -8316 15194 -8284
rect 15076 -8359 15194 -8316
rect 15076 -8444 15194 -8401
rect 15076 -8476 15119 -8444
rect 15119 -8476 15151 -8444
rect 15151 -8476 15194 -8444
rect 15076 -8519 15194 -8476
rect 15076 -8604 15194 -8561
rect 15076 -8636 15119 -8604
rect 15119 -8636 15151 -8604
rect 15151 -8636 15194 -8604
rect 15076 -8679 15194 -8636
rect 15076 -8764 15194 -8721
rect 15076 -8796 15119 -8764
rect 15119 -8796 15151 -8764
rect 15151 -8796 15194 -8764
rect 15076 -8839 15194 -8796
rect 15076 -8924 15194 -8881
rect 15076 -8956 15119 -8924
rect 15119 -8956 15151 -8924
rect 15151 -8956 15194 -8924
rect 15076 -8999 15194 -8956
rect 15076 -9084 15194 -9041
rect 15076 -9116 15119 -9084
rect 15119 -9116 15151 -9084
rect 15151 -9116 15194 -9084
rect 15076 -9159 15194 -9116
rect 15076 -9244 15194 -9201
rect 18809 -5799 18927 -5756
rect 21261 -5621 21379 -5578
rect 21261 -5653 21304 -5621
rect 21304 -5653 21336 -5621
rect 21336 -5653 21379 -5621
rect 21076 -5724 21194 -5681
rect 21261 -5696 21379 -5653
rect 21421 -5621 21539 -5578
rect 21421 -5653 21464 -5621
rect 21464 -5653 21496 -5621
rect 21496 -5653 21539 -5621
rect 21421 -5696 21539 -5653
rect 21581 -5621 21699 -5578
rect 21581 -5653 21624 -5621
rect 21624 -5653 21656 -5621
rect 21656 -5653 21699 -5621
rect 21581 -5696 21699 -5653
rect 21741 -5621 21859 -5578
rect 21741 -5653 21784 -5621
rect 21784 -5653 21816 -5621
rect 21816 -5653 21859 -5621
rect 21741 -5696 21859 -5653
rect 21901 -5621 22019 -5578
rect 21901 -5653 21944 -5621
rect 21944 -5653 21976 -5621
rect 21976 -5653 22019 -5621
rect 21901 -5696 22019 -5653
rect 22061 -5621 22179 -5578
rect 22061 -5653 22104 -5621
rect 22104 -5653 22136 -5621
rect 22136 -5653 22179 -5621
rect 22061 -5696 22179 -5653
rect 22221 -5621 22339 -5578
rect 22221 -5653 22264 -5621
rect 22264 -5653 22296 -5621
rect 22296 -5653 22339 -5621
rect 22221 -5696 22339 -5653
rect 22381 -5621 22499 -5578
rect 22381 -5653 22424 -5621
rect 22424 -5653 22456 -5621
rect 22456 -5653 22499 -5621
rect 22381 -5696 22499 -5653
rect 22541 -5621 22659 -5578
rect 22541 -5653 22584 -5621
rect 22584 -5653 22616 -5621
rect 22616 -5653 22659 -5621
rect 22541 -5696 22659 -5653
rect 22701 -5621 22819 -5578
rect 22701 -5653 22744 -5621
rect 22744 -5653 22776 -5621
rect 22776 -5653 22819 -5621
rect 22701 -5696 22819 -5653
rect 22861 -5621 22979 -5578
rect 22861 -5653 22904 -5621
rect 22904 -5653 22936 -5621
rect 22936 -5653 22979 -5621
rect 22861 -5696 22979 -5653
rect 23021 -5621 23139 -5578
rect 23021 -5653 23064 -5621
rect 23064 -5653 23096 -5621
rect 23096 -5653 23139 -5621
rect 23021 -5696 23139 -5653
rect 23181 -5621 23299 -5578
rect 23181 -5653 23224 -5621
rect 23224 -5653 23256 -5621
rect 23256 -5653 23299 -5621
rect 23181 -5696 23299 -5653
rect 23341 -5621 23459 -5578
rect 23341 -5653 23384 -5621
rect 23384 -5653 23416 -5621
rect 23416 -5653 23459 -5621
rect 23341 -5696 23459 -5653
rect 23501 -5621 23619 -5578
rect 23501 -5653 23544 -5621
rect 23544 -5653 23576 -5621
rect 23576 -5653 23619 -5621
rect 23501 -5696 23619 -5653
rect 23661 -5621 23779 -5578
rect 23661 -5653 23704 -5621
rect 23704 -5653 23736 -5621
rect 23736 -5653 23779 -5621
rect 23661 -5696 23779 -5653
rect 23821 -5621 23939 -5578
rect 23821 -5653 23864 -5621
rect 23864 -5653 23896 -5621
rect 23896 -5653 23939 -5621
rect 23821 -5696 23939 -5653
rect 23981 -5621 24099 -5578
rect 23981 -5653 24024 -5621
rect 24024 -5653 24056 -5621
rect 24056 -5653 24099 -5621
rect 23981 -5696 24099 -5653
rect 24141 -5621 24259 -5578
rect 24141 -5653 24184 -5621
rect 24184 -5653 24216 -5621
rect 24216 -5653 24259 -5621
rect 24141 -5696 24259 -5653
rect 24301 -5621 24419 -5578
rect 24301 -5653 24344 -5621
rect 24344 -5653 24376 -5621
rect 24376 -5653 24419 -5621
rect 24301 -5696 24419 -5653
rect 24461 -5621 24579 -5578
rect 24461 -5653 24504 -5621
rect 24504 -5653 24536 -5621
rect 24536 -5653 24579 -5621
rect 24461 -5696 24579 -5653
rect 24621 -5621 24739 -5578
rect 24621 -5653 24664 -5621
rect 24664 -5653 24696 -5621
rect 24696 -5653 24739 -5621
rect 24621 -5696 24739 -5653
rect 18809 -5884 18927 -5841
rect 18809 -5916 18852 -5884
rect 18852 -5916 18884 -5884
rect 18884 -5916 18927 -5884
rect 18809 -5959 18927 -5916
rect 18809 -6044 18927 -6001
rect 18809 -6076 18852 -6044
rect 18852 -6076 18884 -6044
rect 18884 -6076 18927 -6044
rect 18809 -6119 18927 -6076
rect 18809 -6204 18927 -6161
rect 18809 -6236 18852 -6204
rect 18852 -6236 18884 -6204
rect 18884 -6236 18927 -6204
rect 18809 -6279 18927 -6236
rect 18809 -6364 18927 -6321
rect 18809 -6396 18852 -6364
rect 18852 -6396 18884 -6364
rect 18884 -6396 18927 -6364
rect 18809 -6439 18927 -6396
rect 18809 -6524 18927 -6481
rect 18809 -6556 18852 -6524
rect 18852 -6556 18884 -6524
rect 18884 -6556 18927 -6524
rect 18809 -6599 18927 -6556
rect 18809 -6684 18927 -6641
rect 18809 -6716 18852 -6684
rect 18852 -6716 18884 -6684
rect 18884 -6716 18927 -6684
rect 18809 -6759 18927 -6716
rect 18809 -6844 18927 -6801
rect 18809 -6876 18852 -6844
rect 18852 -6876 18884 -6844
rect 18884 -6876 18927 -6844
rect 18809 -6919 18927 -6876
rect 18809 -7004 18927 -6961
rect 18809 -7036 18852 -7004
rect 18852 -7036 18884 -7004
rect 18884 -7036 18927 -7004
rect 18809 -7079 18927 -7036
rect 18809 -7164 18927 -7121
rect 18809 -7196 18852 -7164
rect 18852 -7196 18884 -7164
rect 18884 -7196 18927 -7164
rect 18809 -7239 18927 -7196
rect 18809 -7324 18927 -7281
rect 18809 -7356 18852 -7324
rect 18852 -7356 18884 -7324
rect 18884 -7356 18927 -7324
rect 18809 -7399 18927 -7356
rect 18809 -7484 18927 -7441
rect 18809 -7516 18852 -7484
rect 18852 -7516 18884 -7484
rect 18884 -7516 18927 -7484
rect 18809 -7559 18927 -7516
rect 18809 -7644 18927 -7601
rect 18809 -7676 18852 -7644
rect 18852 -7676 18884 -7644
rect 18884 -7676 18927 -7644
rect 18809 -7719 18927 -7676
rect 18809 -7804 18927 -7761
rect 18809 -7836 18852 -7804
rect 18852 -7836 18884 -7804
rect 18884 -7836 18927 -7804
rect 18809 -7879 18927 -7836
rect 18809 -7964 18927 -7921
rect 18809 -7996 18852 -7964
rect 18852 -7996 18884 -7964
rect 18884 -7996 18927 -7964
rect 18809 -8039 18927 -7996
rect 18809 -8124 18927 -8081
rect 18809 -8156 18852 -8124
rect 18852 -8156 18884 -8124
rect 18884 -8156 18927 -8124
rect 18809 -8199 18927 -8156
rect 18809 -8284 18927 -8241
rect 18809 -8316 18852 -8284
rect 18852 -8316 18884 -8284
rect 18884 -8316 18927 -8284
rect 18809 -8359 18927 -8316
rect 18809 -8444 18927 -8401
rect 18809 -8476 18852 -8444
rect 18852 -8476 18884 -8444
rect 18884 -8476 18927 -8444
rect 18809 -8519 18927 -8476
rect 18809 -8604 18927 -8561
rect 18809 -8636 18852 -8604
rect 18852 -8636 18884 -8604
rect 18884 -8636 18927 -8604
rect 18809 -8679 18927 -8636
rect 18809 -8764 18927 -8721
rect 18809 -8796 18852 -8764
rect 18852 -8796 18884 -8764
rect 18884 -8796 18927 -8764
rect 18809 -8839 18927 -8796
rect 18809 -8924 18927 -8881
rect 18809 -8956 18852 -8924
rect 18852 -8956 18884 -8924
rect 18884 -8956 18927 -8924
rect 18809 -8999 18927 -8956
rect 18809 -9084 18927 -9041
rect 18809 -9116 18852 -9084
rect 18852 -9116 18884 -9084
rect 18884 -9116 18927 -9084
rect 18809 -9159 18927 -9116
rect 15076 -9276 15119 -9244
rect 15119 -9276 15151 -9244
rect 15151 -9276 15194 -9244
rect 15076 -9319 15194 -9276
rect 18809 -9244 18927 -9201
rect 18809 -9276 18852 -9244
rect 18852 -9276 18884 -9244
rect 18884 -9276 18927 -9244
rect 15261 -9349 15379 -9306
rect 15261 -9381 15304 -9349
rect 15304 -9381 15336 -9349
rect 15336 -9381 15379 -9349
rect 15261 -9424 15379 -9381
rect 15421 -9349 15539 -9306
rect 15421 -9381 15464 -9349
rect 15464 -9381 15496 -9349
rect 15496 -9381 15539 -9349
rect 15421 -9424 15539 -9381
rect 15581 -9349 15699 -9306
rect 15581 -9381 15624 -9349
rect 15624 -9381 15656 -9349
rect 15656 -9381 15699 -9349
rect 15581 -9424 15699 -9381
rect 15741 -9349 15859 -9306
rect 15741 -9381 15784 -9349
rect 15784 -9381 15816 -9349
rect 15816 -9381 15859 -9349
rect 15741 -9424 15859 -9381
rect 15901 -9349 16019 -9306
rect 15901 -9381 15944 -9349
rect 15944 -9381 15976 -9349
rect 15976 -9381 16019 -9349
rect 15901 -9424 16019 -9381
rect 16061 -9349 16179 -9306
rect 16061 -9381 16104 -9349
rect 16104 -9381 16136 -9349
rect 16136 -9381 16179 -9349
rect 16061 -9424 16179 -9381
rect 16221 -9349 16339 -9306
rect 16221 -9381 16264 -9349
rect 16264 -9381 16296 -9349
rect 16296 -9381 16339 -9349
rect 16221 -9424 16339 -9381
rect 16381 -9349 16499 -9306
rect 16381 -9381 16424 -9349
rect 16424 -9381 16456 -9349
rect 16456 -9381 16499 -9349
rect 16381 -9424 16499 -9381
rect 16541 -9349 16659 -9306
rect 16541 -9381 16584 -9349
rect 16584 -9381 16616 -9349
rect 16616 -9381 16659 -9349
rect 16541 -9424 16659 -9381
rect 16701 -9349 16819 -9306
rect 16701 -9381 16744 -9349
rect 16744 -9381 16776 -9349
rect 16776 -9381 16819 -9349
rect 16701 -9424 16819 -9381
rect 16861 -9349 16979 -9306
rect 16861 -9381 16904 -9349
rect 16904 -9381 16936 -9349
rect 16936 -9381 16979 -9349
rect 16861 -9424 16979 -9381
rect 17021 -9349 17139 -9306
rect 17021 -9381 17064 -9349
rect 17064 -9381 17096 -9349
rect 17096 -9381 17139 -9349
rect 17021 -9424 17139 -9381
rect 17181 -9349 17299 -9306
rect 17181 -9381 17224 -9349
rect 17224 -9381 17256 -9349
rect 17256 -9381 17299 -9349
rect 17181 -9424 17299 -9381
rect 17341 -9349 17459 -9306
rect 17341 -9381 17384 -9349
rect 17384 -9381 17416 -9349
rect 17416 -9381 17459 -9349
rect 17341 -9424 17459 -9381
rect 17501 -9349 17619 -9306
rect 17501 -9381 17544 -9349
rect 17544 -9381 17576 -9349
rect 17576 -9381 17619 -9349
rect 17501 -9424 17619 -9381
rect 17661 -9349 17779 -9306
rect 17661 -9381 17704 -9349
rect 17704 -9381 17736 -9349
rect 17736 -9381 17779 -9349
rect 17661 -9424 17779 -9381
rect 17821 -9349 17939 -9306
rect 17821 -9381 17864 -9349
rect 17864 -9381 17896 -9349
rect 17896 -9381 17939 -9349
rect 17821 -9424 17939 -9381
rect 17981 -9349 18099 -9306
rect 17981 -9381 18024 -9349
rect 18024 -9381 18056 -9349
rect 18056 -9381 18099 -9349
rect 17981 -9424 18099 -9381
rect 18141 -9349 18259 -9306
rect 18141 -9381 18184 -9349
rect 18184 -9381 18216 -9349
rect 18216 -9381 18259 -9349
rect 18141 -9424 18259 -9381
rect 18301 -9349 18419 -9306
rect 18301 -9381 18344 -9349
rect 18344 -9381 18376 -9349
rect 18376 -9381 18419 -9349
rect 18301 -9424 18419 -9381
rect 18461 -9349 18579 -9306
rect 18461 -9381 18504 -9349
rect 18504 -9381 18536 -9349
rect 18536 -9381 18579 -9349
rect 18461 -9424 18579 -9381
rect 18621 -9349 18739 -9306
rect 18809 -9319 18927 -9276
rect 18621 -9381 18664 -9349
rect 18664 -9381 18696 -9349
rect 18696 -9381 18739 -9349
rect 18621 -9424 18739 -9381
rect 21076 -5756 21119 -5724
rect 21119 -5756 21151 -5724
rect 21151 -5756 21194 -5724
rect 21076 -5799 21194 -5756
rect 24809 -5724 24927 -5681
rect 24809 -5756 24852 -5724
rect 24852 -5756 24884 -5724
rect 24884 -5756 24927 -5724
rect 21076 -5884 21194 -5841
rect 21076 -5916 21119 -5884
rect 21119 -5916 21151 -5884
rect 21151 -5916 21194 -5884
rect 21076 -5959 21194 -5916
rect 21076 -6044 21194 -6001
rect 21076 -6076 21119 -6044
rect 21119 -6076 21151 -6044
rect 21151 -6076 21194 -6044
rect 21076 -6119 21194 -6076
rect 21076 -6204 21194 -6161
rect 21076 -6236 21119 -6204
rect 21119 -6236 21151 -6204
rect 21151 -6236 21194 -6204
rect 21076 -6279 21194 -6236
rect 21076 -6364 21194 -6321
rect 21076 -6396 21119 -6364
rect 21119 -6396 21151 -6364
rect 21151 -6396 21194 -6364
rect 21076 -6439 21194 -6396
rect 21076 -6524 21194 -6481
rect 21076 -6556 21119 -6524
rect 21119 -6556 21151 -6524
rect 21151 -6556 21194 -6524
rect 21076 -6599 21194 -6556
rect 21076 -6684 21194 -6641
rect 21076 -6716 21119 -6684
rect 21119 -6716 21151 -6684
rect 21151 -6716 21194 -6684
rect 21076 -6759 21194 -6716
rect 21076 -6844 21194 -6801
rect 21076 -6876 21119 -6844
rect 21119 -6876 21151 -6844
rect 21151 -6876 21194 -6844
rect 21076 -6919 21194 -6876
rect 21076 -7004 21194 -6961
rect 21076 -7036 21119 -7004
rect 21119 -7036 21151 -7004
rect 21151 -7036 21194 -7004
rect 21076 -7079 21194 -7036
rect 21076 -7164 21194 -7121
rect 21076 -7196 21119 -7164
rect 21119 -7196 21151 -7164
rect 21151 -7196 21194 -7164
rect 21076 -7239 21194 -7196
rect 21076 -7324 21194 -7281
rect 21076 -7356 21119 -7324
rect 21119 -7356 21151 -7324
rect 21151 -7356 21194 -7324
rect 21076 -7399 21194 -7356
rect 21076 -7484 21194 -7441
rect 21076 -7516 21119 -7484
rect 21119 -7516 21151 -7484
rect 21151 -7516 21194 -7484
rect 21076 -7559 21194 -7516
rect 21076 -7644 21194 -7601
rect 21076 -7676 21119 -7644
rect 21119 -7676 21151 -7644
rect 21151 -7676 21194 -7644
rect 21076 -7719 21194 -7676
rect 21076 -7804 21194 -7761
rect 21076 -7836 21119 -7804
rect 21119 -7836 21151 -7804
rect 21151 -7836 21194 -7804
rect 21076 -7879 21194 -7836
rect 21076 -7964 21194 -7921
rect 21076 -7996 21119 -7964
rect 21119 -7996 21151 -7964
rect 21151 -7996 21194 -7964
rect 21076 -8039 21194 -7996
rect 21076 -8124 21194 -8081
rect 21076 -8156 21119 -8124
rect 21119 -8156 21151 -8124
rect 21151 -8156 21194 -8124
rect 21076 -8199 21194 -8156
rect 21076 -8284 21194 -8241
rect 21076 -8316 21119 -8284
rect 21119 -8316 21151 -8284
rect 21151 -8316 21194 -8284
rect 21076 -8359 21194 -8316
rect 21076 -8444 21194 -8401
rect 21076 -8476 21119 -8444
rect 21119 -8476 21151 -8444
rect 21151 -8476 21194 -8444
rect 21076 -8519 21194 -8476
rect 21076 -8604 21194 -8561
rect 21076 -8636 21119 -8604
rect 21119 -8636 21151 -8604
rect 21151 -8636 21194 -8604
rect 21076 -8679 21194 -8636
rect 21076 -8764 21194 -8721
rect 21076 -8796 21119 -8764
rect 21119 -8796 21151 -8764
rect 21151 -8796 21194 -8764
rect 21076 -8839 21194 -8796
rect 21076 -8924 21194 -8881
rect 21076 -8956 21119 -8924
rect 21119 -8956 21151 -8924
rect 21151 -8956 21194 -8924
rect 21076 -8999 21194 -8956
rect 21076 -9084 21194 -9041
rect 21076 -9116 21119 -9084
rect 21119 -9116 21151 -9084
rect 21151 -9116 21194 -9084
rect 21076 -9159 21194 -9116
rect 21076 -9244 21194 -9201
rect 24809 -5799 24927 -5756
rect 24809 -5884 24927 -5841
rect 24809 -5916 24852 -5884
rect 24852 -5916 24884 -5884
rect 24884 -5916 24927 -5884
rect 24809 -5959 24927 -5916
rect 24809 -6044 24927 -6001
rect 24809 -6076 24852 -6044
rect 24852 -6076 24884 -6044
rect 24884 -6076 24927 -6044
rect 24809 -6119 24927 -6076
rect 24809 -6204 24927 -6161
rect 24809 -6236 24852 -6204
rect 24852 -6236 24884 -6204
rect 24884 -6236 24927 -6204
rect 24809 -6279 24927 -6236
rect 24809 -6364 24927 -6321
rect 24809 -6396 24852 -6364
rect 24852 -6396 24884 -6364
rect 24884 -6396 24927 -6364
rect 24809 -6439 24927 -6396
rect 24809 -6524 24927 -6481
rect 24809 -6556 24852 -6524
rect 24852 -6556 24884 -6524
rect 24884 -6556 24927 -6524
rect 24809 -6599 24927 -6556
rect 24809 -6684 24927 -6641
rect 24809 -6716 24852 -6684
rect 24852 -6716 24884 -6684
rect 24884 -6716 24927 -6684
rect 24809 -6759 24927 -6716
rect 24809 -6844 24927 -6801
rect 24809 -6876 24852 -6844
rect 24852 -6876 24884 -6844
rect 24884 -6876 24927 -6844
rect 24809 -6919 24927 -6876
rect 24809 -7004 24927 -6961
rect 24809 -7036 24852 -7004
rect 24852 -7036 24884 -7004
rect 24884 -7036 24927 -7004
rect 24809 -7079 24927 -7036
rect 24809 -7164 24927 -7121
rect 24809 -7196 24852 -7164
rect 24852 -7196 24884 -7164
rect 24884 -7196 24927 -7164
rect 24809 -7239 24927 -7196
rect 24809 -7324 24927 -7281
rect 24809 -7356 24852 -7324
rect 24852 -7356 24884 -7324
rect 24884 -7356 24927 -7324
rect 24809 -7399 24927 -7356
rect 24809 -7484 24927 -7441
rect 24809 -7516 24852 -7484
rect 24852 -7516 24884 -7484
rect 24884 -7516 24927 -7484
rect 24809 -7559 24927 -7516
rect 24809 -7644 24927 -7601
rect 24809 -7676 24852 -7644
rect 24852 -7676 24884 -7644
rect 24884 -7676 24927 -7644
rect 24809 -7719 24927 -7676
rect 24809 -7804 24927 -7761
rect 24809 -7836 24852 -7804
rect 24852 -7836 24884 -7804
rect 24884 -7836 24927 -7804
rect 24809 -7879 24927 -7836
rect 24809 -7964 24927 -7921
rect 24809 -7996 24852 -7964
rect 24852 -7996 24884 -7964
rect 24884 -7996 24927 -7964
rect 24809 -8039 24927 -7996
rect 24809 -8124 24927 -8081
rect 24809 -8156 24852 -8124
rect 24852 -8156 24884 -8124
rect 24884 -8156 24927 -8124
rect 24809 -8199 24927 -8156
rect 24809 -8284 24927 -8241
rect 24809 -8316 24852 -8284
rect 24852 -8316 24884 -8284
rect 24884 -8316 24927 -8284
rect 24809 -8359 24927 -8316
rect 24809 -8444 24927 -8401
rect 24809 -8476 24852 -8444
rect 24852 -8476 24884 -8444
rect 24884 -8476 24927 -8444
rect 24809 -8519 24927 -8476
rect 24809 -8604 24927 -8561
rect 24809 -8636 24852 -8604
rect 24852 -8636 24884 -8604
rect 24884 -8636 24927 -8604
rect 24809 -8679 24927 -8636
rect 24809 -8764 24927 -8721
rect 24809 -8796 24852 -8764
rect 24852 -8796 24884 -8764
rect 24884 -8796 24927 -8764
rect 24809 -8839 24927 -8796
rect 24809 -8924 24927 -8881
rect 24809 -8956 24852 -8924
rect 24852 -8956 24884 -8924
rect 24884 -8956 24927 -8924
rect 24809 -8999 24927 -8956
rect 24809 -9084 24927 -9041
rect 24809 -9116 24852 -9084
rect 24852 -9116 24884 -9084
rect 24884 -9116 24927 -9084
rect 24809 -9159 24927 -9116
rect 21076 -9276 21119 -9244
rect 21119 -9276 21151 -9244
rect 21151 -9276 21194 -9244
rect 21076 -9319 21194 -9276
rect 24809 -9244 24927 -9201
rect 24809 -9276 24852 -9244
rect 24852 -9276 24884 -9244
rect 24884 -9276 24927 -9244
rect 21261 -9349 21379 -9306
rect 21261 -9381 21304 -9349
rect 21304 -9381 21336 -9349
rect 21336 -9381 21379 -9349
rect 21261 -9424 21379 -9381
rect 21421 -9349 21539 -9306
rect 21421 -9381 21464 -9349
rect 21464 -9381 21496 -9349
rect 21496 -9381 21539 -9349
rect 21421 -9424 21539 -9381
rect 21581 -9349 21699 -9306
rect 21581 -9381 21624 -9349
rect 21624 -9381 21656 -9349
rect 21656 -9381 21699 -9349
rect 21581 -9424 21699 -9381
rect 21741 -9349 21859 -9306
rect 21741 -9381 21784 -9349
rect 21784 -9381 21816 -9349
rect 21816 -9381 21859 -9349
rect 21741 -9424 21859 -9381
rect 21901 -9349 22019 -9306
rect 21901 -9381 21944 -9349
rect 21944 -9381 21976 -9349
rect 21976 -9381 22019 -9349
rect 21901 -9424 22019 -9381
rect 22061 -9349 22179 -9306
rect 22061 -9381 22104 -9349
rect 22104 -9381 22136 -9349
rect 22136 -9381 22179 -9349
rect 22061 -9424 22179 -9381
rect 22221 -9349 22339 -9306
rect 22221 -9381 22264 -9349
rect 22264 -9381 22296 -9349
rect 22296 -9381 22339 -9349
rect 22221 -9424 22339 -9381
rect 22381 -9349 22499 -9306
rect 22381 -9381 22424 -9349
rect 22424 -9381 22456 -9349
rect 22456 -9381 22499 -9349
rect 22381 -9424 22499 -9381
rect 22541 -9349 22659 -9306
rect 22541 -9381 22584 -9349
rect 22584 -9381 22616 -9349
rect 22616 -9381 22659 -9349
rect 22541 -9424 22659 -9381
rect 22701 -9349 22819 -9306
rect 22701 -9381 22744 -9349
rect 22744 -9381 22776 -9349
rect 22776 -9381 22819 -9349
rect 22701 -9424 22819 -9381
rect 22861 -9349 22979 -9306
rect 22861 -9381 22904 -9349
rect 22904 -9381 22936 -9349
rect 22936 -9381 22979 -9349
rect 22861 -9424 22979 -9381
rect 23021 -9349 23139 -9306
rect 23021 -9381 23064 -9349
rect 23064 -9381 23096 -9349
rect 23096 -9381 23139 -9349
rect 23021 -9424 23139 -9381
rect 23181 -9349 23299 -9306
rect 23181 -9381 23224 -9349
rect 23224 -9381 23256 -9349
rect 23256 -9381 23299 -9349
rect 23181 -9424 23299 -9381
rect 23341 -9349 23459 -9306
rect 23341 -9381 23384 -9349
rect 23384 -9381 23416 -9349
rect 23416 -9381 23459 -9349
rect 23341 -9424 23459 -9381
rect 23501 -9349 23619 -9306
rect 23501 -9381 23544 -9349
rect 23544 -9381 23576 -9349
rect 23576 -9381 23619 -9349
rect 23501 -9424 23619 -9381
rect 23661 -9349 23779 -9306
rect 23661 -9381 23704 -9349
rect 23704 -9381 23736 -9349
rect 23736 -9381 23779 -9349
rect 23661 -9424 23779 -9381
rect 23821 -9349 23939 -9306
rect 23821 -9381 23864 -9349
rect 23864 -9381 23896 -9349
rect 23896 -9381 23939 -9349
rect 23821 -9424 23939 -9381
rect 23981 -9349 24099 -9306
rect 23981 -9381 24024 -9349
rect 24024 -9381 24056 -9349
rect 24056 -9381 24099 -9349
rect 23981 -9424 24099 -9381
rect 24141 -9349 24259 -9306
rect 24141 -9381 24184 -9349
rect 24184 -9381 24216 -9349
rect 24216 -9381 24259 -9349
rect 24141 -9424 24259 -9381
rect 24301 -9349 24419 -9306
rect 24301 -9381 24344 -9349
rect 24344 -9381 24376 -9349
rect 24376 -9381 24419 -9349
rect 24301 -9424 24419 -9381
rect 24461 -9349 24579 -9306
rect 24461 -9381 24504 -9349
rect 24504 -9381 24536 -9349
rect 24536 -9381 24579 -9349
rect 24461 -9424 24579 -9381
rect 24621 -9349 24739 -9306
rect 24809 -9319 24927 -9276
rect 24621 -9381 24664 -9349
rect 24664 -9381 24696 -9349
rect 24696 -9381 24739 -9349
rect 24621 -9424 24739 -9381
rect 3261 -11621 3379 -11578
rect 3261 -11653 3304 -11621
rect 3304 -11653 3336 -11621
rect 3336 -11653 3379 -11621
rect 3076 -11724 3194 -11681
rect 3261 -11696 3379 -11653
rect 3421 -11621 3539 -11578
rect 3421 -11653 3464 -11621
rect 3464 -11653 3496 -11621
rect 3496 -11653 3539 -11621
rect 3421 -11696 3539 -11653
rect 3581 -11621 3699 -11578
rect 3581 -11653 3624 -11621
rect 3624 -11653 3656 -11621
rect 3656 -11653 3699 -11621
rect 3581 -11696 3699 -11653
rect 3741 -11621 3859 -11578
rect 3741 -11653 3784 -11621
rect 3784 -11653 3816 -11621
rect 3816 -11653 3859 -11621
rect 3741 -11696 3859 -11653
rect 3901 -11621 4019 -11578
rect 3901 -11653 3944 -11621
rect 3944 -11653 3976 -11621
rect 3976 -11653 4019 -11621
rect 3901 -11696 4019 -11653
rect 4061 -11621 4179 -11578
rect 4061 -11653 4104 -11621
rect 4104 -11653 4136 -11621
rect 4136 -11653 4179 -11621
rect 4061 -11696 4179 -11653
rect 4221 -11621 4339 -11578
rect 4221 -11653 4264 -11621
rect 4264 -11653 4296 -11621
rect 4296 -11653 4339 -11621
rect 4221 -11696 4339 -11653
rect 4381 -11621 4499 -11578
rect 4381 -11653 4424 -11621
rect 4424 -11653 4456 -11621
rect 4456 -11653 4499 -11621
rect 4381 -11696 4499 -11653
rect 4541 -11621 4659 -11578
rect 4541 -11653 4584 -11621
rect 4584 -11653 4616 -11621
rect 4616 -11653 4659 -11621
rect 4541 -11696 4659 -11653
rect 4701 -11621 4819 -11578
rect 4701 -11653 4744 -11621
rect 4744 -11653 4776 -11621
rect 4776 -11653 4819 -11621
rect 4701 -11696 4819 -11653
rect 4861 -11621 4979 -11578
rect 4861 -11653 4904 -11621
rect 4904 -11653 4936 -11621
rect 4936 -11653 4979 -11621
rect 4861 -11696 4979 -11653
rect 5021 -11621 5139 -11578
rect 5021 -11653 5064 -11621
rect 5064 -11653 5096 -11621
rect 5096 -11653 5139 -11621
rect 5021 -11696 5139 -11653
rect 5181 -11621 5299 -11578
rect 5181 -11653 5224 -11621
rect 5224 -11653 5256 -11621
rect 5256 -11653 5299 -11621
rect 5181 -11696 5299 -11653
rect 5341 -11621 5459 -11578
rect 5341 -11653 5384 -11621
rect 5384 -11653 5416 -11621
rect 5416 -11653 5459 -11621
rect 5341 -11696 5459 -11653
rect 5501 -11621 5619 -11578
rect 5501 -11653 5544 -11621
rect 5544 -11653 5576 -11621
rect 5576 -11653 5619 -11621
rect 5501 -11696 5619 -11653
rect 5661 -11621 5779 -11578
rect 5661 -11653 5704 -11621
rect 5704 -11653 5736 -11621
rect 5736 -11653 5779 -11621
rect 5661 -11696 5779 -11653
rect 5821 -11621 5939 -11578
rect 5821 -11653 5864 -11621
rect 5864 -11653 5896 -11621
rect 5896 -11653 5939 -11621
rect 5821 -11696 5939 -11653
rect 5981 -11621 6099 -11578
rect 5981 -11653 6024 -11621
rect 6024 -11653 6056 -11621
rect 6056 -11653 6099 -11621
rect 5981 -11696 6099 -11653
rect 6141 -11621 6259 -11578
rect 6141 -11653 6184 -11621
rect 6184 -11653 6216 -11621
rect 6216 -11653 6259 -11621
rect 6141 -11696 6259 -11653
rect 6301 -11621 6419 -11578
rect 6301 -11653 6344 -11621
rect 6344 -11653 6376 -11621
rect 6376 -11653 6419 -11621
rect 6301 -11696 6419 -11653
rect 6461 -11621 6579 -11578
rect 6461 -11653 6504 -11621
rect 6504 -11653 6536 -11621
rect 6536 -11653 6579 -11621
rect 6461 -11696 6579 -11653
rect 6621 -11621 6739 -11578
rect 6621 -11653 6664 -11621
rect 6664 -11653 6696 -11621
rect 6696 -11653 6739 -11621
rect 6621 -11696 6739 -11653
rect 3076 -11756 3119 -11724
rect 3119 -11756 3151 -11724
rect 3151 -11756 3194 -11724
rect 3076 -11799 3194 -11756
rect 6809 -11724 6927 -11681
rect 6809 -11756 6852 -11724
rect 6852 -11756 6884 -11724
rect 6884 -11756 6927 -11724
rect 3076 -11884 3194 -11841
rect 3076 -11916 3119 -11884
rect 3119 -11916 3151 -11884
rect 3151 -11916 3194 -11884
rect 3076 -11959 3194 -11916
rect 3076 -12044 3194 -12001
rect 3076 -12076 3119 -12044
rect 3119 -12076 3151 -12044
rect 3151 -12076 3194 -12044
rect 3076 -12119 3194 -12076
rect 3076 -12204 3194 -12161
rect 3076 -12236 3119 -12204
rect 3119 -12236 3151 -12204
rect 3151 -12236 3194 -12204
rect 3076 -12279 3194 -12236
rect 3076 -12364 3194 -12321
rect 3076 -12396 3119 -12364
rect 3119 -12396 3151 -12364
rect 3151 -12396 3194 -12364
rect 3076 -12439 3194 -12396
rect 3076 -12524 3194 -12481
rect 3076 -12556 3119 -12524
rect 3119 -12556 3151 -12524
rect 3151 -12556 3194 -12524
rect 3076 -12599 3194 -12556
rect 3076 -12684 3194 -12641
rect 3076 -12716 3119 -12684
rect 3119 -12716 3151 -12684
rect 3151 -12716 3194 -12684
rect 3076 -12759 3194 -12716
rect 3076 -12844 3194 -12801
rect 3076 -12876 3119 -12844
rect 3119 -12876 3151 -12844
rect 3151 -12876 3194 -12844
rect 3076 -12919 3194 -12876
rect 3076 -13004 3194 -12961
rect 3076 -13036 3119 -13004
rect 3119 -13036 3151 -13004
rect 3151 -13036 3194 -13004
rect 3076 -13079 3194 -13036
rect 3076 -13164 3194 -13121
rect 3076 -13196 3119 -13164
rect 3119 -13196 3151 -13164
rect 3151 -13196 3194 -13164
rect 3076 -13239 3194 -13196
rect 3076 -13324 3194 -13281
rect 3076 -13356 3119 -13324
rect 3119 -13356 3151 -13324
rect 3151 -13356 3194 -13324
rect 3076 -13399 3194 -13356
rect 3076 -13484 3194 -13441
rect 3076 -13516 3119 -13484
rect 3119 -13516 3151 -13484
rect 3151 -13516 3194 -13484
rect 3076 -13559 3194 -13516
rect 3076 -13644 3194 -13601
rect 3076 -13676 3119 -13644
rect 3119 -13676 3151 -13644
rect 3151 -13676 3194 -13644
rect 3076 -13719 3194 -13676
rect 3076 -13804 3194 -13761
rect 3076 -13836 3119 -13804
rect 3119 -13836 3151 -13804
rect 3151 -13836 3194 -13804
rect 3076 -13879 3194 -13836
rect 3076 -13964 3194 -13921
rect 3076 -13996 3119 -13964
rect 3119 -13996 3151 -13964
rect 3151 -13996 3194 -13964
rect 3076 -14039 3194 -13996
rect 3076 -14124 3194 -14081
rect 3076 -14156 3119 -14124
rect 3119 -14156 3151 -14124
rect 3151 -14156 3194 -14124
rect 3076 -14199 3194 -14156
rect 3076 -14284 3194 -14241
rect 3076 -14316 3119 -14284
rect 3119 -14316 3151 -14284
rect 3151 -14316 3194 -14284
rect 3076 -14359 3194 -14316
rect 3076 -14444 3194 -14401
rect 3076 -14476 3119 -14444
rect 3119 -14476 3151 -14444
rect 3151 -14476 3194 -14444
rect 3076 -14519 3194 -14476
rect 3076 -14604 3194 -14561
rect 3076 -14636 3119 -14604
rect 3119 -14636 3151 -14604
rect 3151 -14636 3194 -14604
rect 3076 -14679 3194 -14636
rect 3076 -14764 3194 -14721
rect 3076 -14796 3119 -14764
rect 3119 -14796 3151 -14764
rect 3151 -14796 3194 -14764
rect 3076 -14839 3194 -14796
rect 3076 -14924 3194 -14881
rect 3076 -14956 3119 -14924
rect 3119 -14956 3151 -14924
rect 3151 -14956 3194 -14924
rect 3076 -14999 3194 -14956
rect 3076 -15084 3194 -15041
rect 3076 -15116 3119 -15084
rect 3119 -15116 3151 -15084
rect 3151 -15116 3194 -15084
rect 3076 -15159 3194 -15116
rect 3076 -15244 3194 -15201
rect 6809 -11799 6927 -11756
rect 6809 -11884 6927 -11841
rect 6809 -11916 6852 -11884
rect 6852 -11916 6884 -11884
rect 6884 -11916 6927 -11884
rect 6809 -11959 6927 -11916
rect 6809 -12044 6927 -12001
rect 6809 -12076 6852 -12044
rect 6852 -12076 6884 -12044
rect 6884 -12076 6927 -12044
rect 6809 -12119 6927 -12076
rect 6809 -12204 6927 -12161
rect 6809 -12236 6852 -12204
rect 6852 -12236 6884 -12204
rect 6884 -12236 6927 -12204
rect 6809 -12279 6927 -12236
rect 6809 -12364 6927 -12321
rect 6809 -12396 6852 -12364
rect 6852 -12396 6884 -12364
rect 6884 -12396 6927 -12364
rect 6809 -12439 6927 -12396
rect 6809 -12524 6927 -12481
rect 6809 -12556 6852 -12524
rect 6852 -12556 6884 -12524
rect 6884 -12556 6927 -12524
rect 6809 -12599 6927 -12556
rect 6809 -12684 6927 -12641
rect 6809 -12716 6852 -12684
rect 6852 -12716 6884 -12684
rect 6884 -12716 6927 -12684
rect 6809 -12759 6927 -12716
rect 6809 -12844 6927 -12801
rect 6809 -12876 6852 -12844
rect 6852 -12876 6884 -12844
rect 6884 -12876 6927 -12844
rect 6809 -12919 6927 -12876
rect 6809 -13004 6927 -12961
rect 6809 -13036 6852 -13004
rect 6852 -13036 6884 -13004
rect 6884 -13036 6927 -13004
rect 6809 -13079 6927 -13036
rect 6809 -13164 6927 -13121
rect 6809 -13196 6852 -13164
rect 6852 -13196 6884 -13164
rect 6884 -13196 6927 -13164
rect 6809 -13239 6927 -13196
rect 6809 -13324 6927 -13281
rect 6809 -13356 6852 -13324
rect 6852 -13356 6884 -13324
rect 6884 -13356 6927 -13324
rect 6809 -13399 6927 -13356
rect 6809 -13484 6927 -13441
rect 6809 -13516 6852 -13484
rect 6852 -13516 6884 -13484
rect 6884 -13516 6927 -13484
rect 6809 -13559 6927 -13516
rect 6809 -13644 6927 -13601
rect 6809 -13676 6852 -13644
rect 6852 -13676 6884 -13644
rect 6884 -13676 6927 -13644
rect 6809 -13719 6927 -13676
rect 6809 -13804 6927 -13761
rect 6809 -13836 6852 -13804
rect 6852 -13836 6884 -13804
rect 6884 -13836 6927 -13804
rect 6809 -13879 6927 -13836
rect 6809 -13964 6927 -13921
rect 6809 -13996 6852 -13964
rect 6852 -13996 6884 -13964
rect 6884 -13996 6927 -13964
rect 6809 -14039 6927 -13996
rect 6809 -14124 6927 -14081
rect 6809 -14156 6852 -14124
rect 6852 -14156 6884 -14124
rect 6884 -14156 6927 -14124
rect 6809 -14199 6927 -14156
rect 6809 -14284 6927 -14241
rect 6809 -14316 6852 -14284
rect 6852 -14316 6884 -14284
rect 6884 -14316 6927 -14284
rect 6809 -14359 6927 -14316
rect 6809 -14444 6927 -14401
rect 6809 -14476 6852 -14444
rect 6852 -14476 6884 -14444
rect 6884 -14476 6927 -14444
rect 6809 -14519 6927 -14476
rect 6809 -14604 6927 -14561
rect 6809 -14636 6852 -14604
rect 6852 -14636 6884 -14604
rect 6884 -14636 6927 -14604
rect 6809 -14679 6927 -14636
rect 6809 -14764 6927 -14721
rect 6809 -14796 6852 -14764
rect 6852 -14796 6884 -14764
rect 6884 -14796 6927 -14764
rect 6809 -14839 6927 -14796
rect 6809 -14924 6927 -14881
rect 6809 -14956 6852 -14924
rect 6852 -14956 6884 -14924
rect 6884 -14956 6927 -14924
rect 6809 -14999 6927 -14956
rect 6809 -15084 6927 -15041
rect 6809 -15116 6852 -15084
rect 6852 -15116 6884 -15084
rect 6884 -15116 6927 -15084
rect 6809 -15159 6927 -15116
rect 3076 -15276 3119 -15244
rect 3119 -15276 3151 -15244
rect 3151 -15276 3194 -15244
rect 3076 -15319 3194 -15276
rect 6809 -15244 6927 -15201
rect 6809 -15276 6852 -15244
rect 6852 -15276 6884 -15244
rect 6884 -15276 6927 -15244
rect 3261 -15349 3379 -15306
rect 3261 -15381 3304 -15349
rect 3304 -15381 3336 -15349
rect 3336 -15381 3379 -15349
rect 3261 -15424 3379 -15381
rect 3421 -15349 3539 -15306
rect 3421 -15381 3464 -15349
rect 3464 -15381 3496 -15349
rect 3496 -15381 3539 -15349
rect 3421 -15424 3539 -15381
rect 3581 -15349 3699 -15306
rect 3581 -15381 3624 -15349
rect 3624 -15381 3656 -15349
rect 3656 -15381 3699 -15349
rect 3581 -15424 3699 -15381
rect 3741 -15349 3859 -15306
rect 3741 -15381 3784 -15349
rect 3784 -15381 3816 -15349
rect 3816 -15381 3859 -15349
rect 3741 -15424 3859 -15381
rect 3901 -15349 4019 -15306
rect 3901 -15381 3944 -15349
rect 3944 -15381 3976 -15349
rect 3976 -15381 4019 -15349
rect 3901 -15424 4019 -15381
rect 4061 -15349 4179 -15306
rect 4061 -15381 4104 -15349
rect 4104 -15381 4136 -15349
rect 4136 -15381 4179 -15349
rect 4061 -15424 4179 -15381
rect 4221 -15349 4339 -15306
rect 4221 -15381 4264 -15349
rect 4264 -15381 4296 -15349
rect 4296 -15381 4339 -15349
rect 4221 -15424 4339 -15381
rect 4381 -15349 4499 -15306
rect 4381 -15381 4424 -15349
rect 4424 -15381 4456 -15349
rect 4456 -15381 4499 -15349
rect 4381 -15424 4499 -15381
rect 4541 -15349 4659 -15306
rect 4541 -15381 4584 -15349
rect 4584 -15381 4616 -15349
rect 4616 -15381 4659 -15349
rect 4541 -15424 4659 -15381
rect 4701 -15349 4819 -15306
rect 4701 -15381 4744 -15349
rect 4744 -15381 4776 -15349
rect 4776 -15381 4819 -15349
rect 4701 -15424 4819 -15381
rect 4861 -15349 4979 -15306
rect 4861 -15381 4904 -15349
rect 4904 -15381 4936 -15349
rect 4936 -15381 4979 -15349
rect 4861 -15424 4979 -15381
rect 5021 -15349 5139 -15306
rect 5021 -15381 5064 -15349
rect 5064 -15381 5096 -15349
rect 5096 -15381 5139 -15349
rect 5021 -15424 5139 -15381
rect 5181 -15349 5299 -15306
rect 5181 -15381 5224 -15349
rect 5224 -15381 5256 -15349
rect 5256 -15381 5299 -15349
rect 5181 -15424 5299 -15381
rect 5341 -15349 5459 -15306
rect 5341 -15381 5384 -15349
rect 5384 -15381 5416 -15349
rect 5416 -15381 5459 -15349
rect 5341 -15424 5459 -15381
rect 5501 -15349 5619 -15306
rect 5501 -15381 5544 -15349
rect 5544 -15381 5576 -15349
rect 5576 -15381 5619 -15349
rect 5501 -15424 5619 -15381
rect 5661 -15349 5779 -15306
rect 5661 -15381 5704 -15349
rect 5704 -15381 5736 -15349
rect 5736 -15381 5779 -15349
rect 5661 -15424 5779 -15381
rect 5821 -15349 5939 -15306
rect 5821 -15381 5864 -15349
rect 5864 -15381 5896 -15349
rect 5896 -15381 5939 -15349
rect 5821 -15424 5939 -15381
rect 5981 -15349 6099 -15306
rect 5981 -15381 6024 -15349
rect 6024 -15381 6056 -15349
rect 6056 -15381 6099 -15349
rect 5981 -15424 6099 -15381
rect 6141 -15349 6259 -15306
rect 6141 -15381 6184 -15349
rect 6184 -15381 6216 -15349
rect 6216 -15381 6259 -15349
rect 6141 -15424 6259 -15381
rect 6301 -15349 6419 -15306
rect 6301 -15381 6344 -15349
rect 6344 -15381 6376 -15349
rect 6376 -15381 6419 -15349
rect 6301 -15424 6419 -15381
rect 6461 -15349 6579 -15306
rect 6461 -15381 6504 -15349
rect 6504 -15381 6536 -15349
rect 6536 -15381 6579 -15349
rect 6461 -15424 6579 -15381
rect 6621 -15349 6739 -15306
rect 6809 -15319 6927 -15276
rect 6621 -15381 6664 -15349
rect 6664 -15381 6696 -15349
rect 6696 -15381 6739 -15349
rect 6621 -15424 6739 -15381
rect 9261 -11621 9379 -11578
rect 9261 -11653 9304 -11621
rect 9304 -11653 9336 -11621
rect 9336 -11653 9379 -11621
rect 9076 -11724 9194 -11681
rect 9261 -11696 9379 -11653
rect 9421 -11621 9539 -11578
rect 9421 -11653 9464 -11621
rect 9464 -11653 9496 -11621
rect 9496 -11653 9539 -11621
rect 9421 -11696 9539 -11653
rect 9581 -11621 9699 -11578
rect 9581 -11653 9624 -11621
rect 9624 -11653 9656 -11621
rect 9656 -11653 9699 -11621
rect 9581 -11696 9699 -11653
rect 9741 -11621 9859 -11578
rect 9741 -11653 9784 -11621
rect 9784 -11653 9816 -11621
rect 9816 -11653 9859 -11621
rect 9741 -11696 9859 -11653
rect 9901 -11621 10019 -11578
rect 9901 -11653 9944 -11621
rect 9944 -11653 9976 -11621
rect 9976 -11653 10019 -11621
rect 9901 -11696 10019 -11653
rect 10061 -11621 10179 -11578
rect 10061 -11653 10104 -11621
rect 10104 -11653 10136 -11621
rect 10136 -11653 10179 -11621
rect 10061 -11696 10179 -11653
rect 10221 -11621 10339 -11578
rect 10221 -11653 10264 -11621
rect 10264 -11653 10296 -11621
rect 10296 -11653 10339 -11621
rect 10221 -11696 10339 -11653
rect 10381 -11621 10499 -11578
rect 10381 -11653 10424 -11621
rect 10424 -11653 10456 -11621
rect 10456 -11653 10499 -11621
rect 10381 -11696 10499 -11653
rect 10541 -11621 10659 -11578
rect 10541 -11653 10584 -11621
rect 10584 -11653 10616 -11621
rect 10616 -11653 10659 -11621
rect 10541 -11696 10659 -11653
rect 10701 -11621 10819 -11578
rect 10701 -11653 10744 -11621
rect 10744 -11653 10776 -11621
rect 10776 -11653 10819 -11621
rect 10701 -11696 10819 -11653
rect 10861 -11621 10979 -11578
rect 10861 -11653 10904 -11621
rect 10904 -11653 10936 -11621
rect 10936 -11653 10979 -11621
rect 10861 -11696 10979 -11653
rect 11021 -11621 11139 -11578
rect 11021 -11653 11064 -11621
rect 11064 -11653 11096 -11621
rect 11096 -11653 11139 -11621
rect 11021 -11696 11139 -11653
rect 11181 -11621 11299 -11578
rect 11181 -11653 11224 -11621
rect 11224 -11653 11256 -11621
rect 11256 -11653 11299 -11621
rect 11181 -11696 11299 -11653
rect 11341 -11621 11459 -11578
rect 11341 -11653 11384 -11621
rect 11384 -11653 11416 -11621
rect 11416 -11653 11459 -11621
rect 11341 -11696 11459 -11653
rect 11501 -11621 11619 -11578
rect 11501 -11653 11544 -11621
rect 11544 -11653 11576 -11621
rect 11576 -11653 11619 -11621
rect 11501 -11696 11619 -11653
rect 11661 -11621 11779 -11578
rect 11661 -11653 11704 -11621
rect 11704 -11653 11736 -11621
rect 11736 -11653 11779 -11621
rect 11661 -11696 11779 -11653
rect 11821 -11621 11939 -11578
rect 11821 -11653 11864 -11621
rect 11864 -11653 11896 -11621
rect 11896 -11653 11939 -11621
rect 11821 -11696 11939 -11653
rect 11981 -11621 12099 -11578
rect 11981 -11653 12024 -11621
rect 12024 -11653 12056 -11621
rect 12056 -11653 12099 -11621
rect 11981 -11696 12099 -11653
rect 12141 -11621 12259 -11578
rect 12141 -11653 12184 -11621
rect 12184 -11653 12216 -11621
rect 12216 -11653 12259 -11621
rect 12141 -11696 12259 -11653
rect 12301 -11621 12419 -11578
rect 12301 -11653 12344 -11621
rect 12344 -11653 12376 -11621
rect 12376 -11653 12419 -11621
rect 12301 -11696 12419 -11653
rect 12461 -11621 12579 -11578
rect 12461 -11653 12504 -11621
rect 12504 -11653 12536 -11621
rect 12536 -11653 12579 -11621
rect 12461 -11696 12579 -11653
rect 12621 -11621 12739 -11578
rect 12621 -11653 12664 -11621
rect 12664 -11653 12696 -11621
rect 12696 -11653 12739 -11621
rect 12621 -11696 12739 -11653
rect 9076 -11756 9119 -11724
rect 9119 -11756 9151 -11724
rect 9151 -11756 9194 -11724
rect 9076 -11799 9194 -11756
rect 12809 -11724 12927 -11681
rect 12809 -11756 12852 -11724
rect 12852 -11756 12884 -11724
rect 12884 -11756 12927 -11724
rect 9076 -11884 9194 -11841
rect 9076 -11916 9119 -11884
rect 9119 -11916 9151 -11884
rect 9151 -11916 9194 -11884
rect 9076 -11959 9194 -11916
rect 9076 -12044 9194 -12001
rect 9076 -12076 9119 -12044
rect 9119 -12076 9151 -12044
rect 9151 -12076 9194 -12044
rect 9076 -12119 9194 -12076
rect 9076 -12204 9194 -12161
rect 9076 -12236 9119 -12204
rect 9119 -12236 9151 -12204
rect 9151 -12236 9194 -12204
rect 9076 -12279 9194 -12236
rect 9076 -12364 9194 -12321
rect 9076 -12396 9119 -12364
rect 9119 -12396 9151 -12364
rect 9151 -12396 9194 -12364
rect 9076 -12439 9194 -12396
rect 9076 -12524 9194 -12481
rect 9076 -12556 9119 -12524
rect 9119 -12556 9151 -12524
rect 9151 -12556 9194 -12524
rect 9076 -12599 9194 -12556
rect 9076 -12684 9194 -12641
rect 9076 -12716 9119 -12684
rect 9119 -12716 9151 -12684
rect 9151 -12716 9194 -12684
rect 9076 -12759 9194 -12716
rect 9076 -12844 9194 -12801
rect 9076 -12876 9119 -12844
rect 9119 -12876 9151 -12844
rect 9151 -12876 9194 -12844
rect 9076 -12919 9194 -12876
rect 9076 -13004 9194 -12961
rect 9076 -13036 9119 -13004
rect 9119 -13036 9151 -13004
rect 9151 -13036 9194 -13004
rect 9076 -13079 9194 -13036
rect 9076 -13164 9194 -13121
rect 9076 -13196 9119 -13164
rect 9119 -13196 9151 -13164
rect 9151 -13196 9194 -13164
rect 9076 -13239 9194 -13196
rect 9076 -13324 9194 -13281
rect 9076 -13356 9119 -13324
rect 9119 -13356 9151 -13324
rect 9151 -13356 9194 -13324
rect 9076 -13399 9194 -13356
rect 9076 -13484 9194 -13441
rect 9076 -13516 9119 -13484
rect 9119 -13516 9151 -13484
rect 9151 -13516 9194 -13484
rect 9076 -13559 9194 -13516
rect 9076 -13644 9194 -13601
rect 9076 -13676 9119 -13644
rect 9119 -13676 9151 -13644
rect 9151 -13676 9194 -13644
rect 9076 -13719 9194 -13676
rect 9076 -13804 9194 -13761
rect 9076 -13836 9119 -13804
rect 9119 -13836 9151 -13804
rect 9151 -13836 9194 -13804
rect 9076 -13879 9194 -13836
rect 9076 -13964 9194 -13921
rect 9076 -13996 9119 -13964
rect 9119 -13996 9151 -13964
rect 9151 -13996 9194 -13964
rect 9076 -14039 9194 -13996
rect 9076 -14124 9194 -14081
rect 9076 -14156 9119 -14124
rect 9119 -14156 9151 -14124
rect 9151 -14156 9194 -14124
rect 9076 -14199 9194 -14156
rect 9076 -14284 9194 -14241
rect 9076 -14316 9119 -14284
rect 9119 -14316 9151 -14284
rect 9151 -14316 9194 -14284
rect 9076 -14359 9194 -14316
rect 9076 -14444 9194 -14401
rect 9076 -14476 9119 -14444
rect 9119 -14476 9151 -14444
rect 9151 -14476 9194 -14444
rect 9076 -14519 9194 -14476
rect 9076 -14604 9194 -14561
rect 9076 -14636 9119 -14604
rect 9119 -14636 9151 -14604
rect 9151 -14636 9194 -14604
rect 9076 -14679 9194 -14636
rect 9076 -14764 9194 -14721
rect 9076 -14796 9119 -14764
rect 9119 -14796 9151 -14764
rect 9151 -14796 9194 -14764
rect 9076 -14839 9194 -14796
rect 9076 -14924 9194 -14881
rect 9076 -14956 9119 -14924
rect 9119 -14956 9151 -14924
rect 9151 -14956 9194 -14924
rect 9076 -14999 9194 -14956
rect 9076 -15084 9194 -15041
rect 9076 -15116 9119 -15084
rect 9119 -15116 9151 -15084
rect 9151 -15116 9194 -15084
rect 9076 -15159 9194 -15116
rect 9076 -15244 9194 -15201
rect 12809 -11799 12927 -11756
rect 12809 -11884 12927 -11841
rect 12809 -11916 12852 -11884
rect 12852 -11916 12884 -11884
rect 12884 -11916 12927 -11884
rect 12809 -11959 12927 -11916
rect 12809 -12044 12927 -12001
rect 12809 -12076 12852 -12044
rect 12852 -12076 12884 -12044
rect 12884 -12076 12927 -12044
rect 12809 -12119 12927 -12076
rect 12809 -12204 12927 -12161
rect 12809 -12236 12852 -12204
rect 12852 -12236 12884 -12204
rect 12884 -12236 12927 -12204
rect 12809 -12279 12927 -12236
rect 12809 -12364 12927 -12321
rect 12809 -12396 12852 -12364
rect 12852 -12396 12884 -12364
rect 12884 -12396 12927 -12364
rect 12809 -12439 12927 -12396
rect 12809 -12524 12927 -12481
rect 12809 -12556 12852 -12524
rect 12852 -12556 12884 -12524
rect 12884 -12556 12927 -12524
rect 12809 -12599 12927 -12556
rect 12809 -12684 12927 -12641
rect 12809 -12716 12852 -12684
rect 12852 -12716 12884 -12684
rect 12884 -12716 12927 -12684
rect 12809 -12759 12927 -12716
rect 12809 -12844 12927 -12801
rect 12809 -12876 12852 -12844
rect 12852 -12876 12884 -12844
rect 12884 -12876 12927 -12844
rect 12809 -12919 12927 -12876
rect 12809 -13004 12927 -12961
rect 12809 -13036 12852 -13004
rect 12852 -13036 12884 -13004
rect 12884 -13036 12927 -13004
rect 12809 -13079 12927 -13036
rect 12809 -13164 12927 -13121
rect 12809 -13196 12852 -13164
rect 12852 -13196 12884 -13164
rect 12884 -13196 12927 -13164
rect 12809 -13239 12927 -13196
rect 12809 -13324 12927 -13281
rect 12809 -13356 12852 -13324
rect 12852 -13356 12884 -13324
rect 12884 -13356 12927 -13324
rect 12809 -13399 12927 -13356
rect 12809 -13484 12927 -13441
rect 12809 -13516 12852 -13484
rect 12852 -13516 12884 -13484
rect 12884 -13516 12927 -13484
rect 12809 -13559 12927 -13516
rect 12809 -13644 12927 -13601
rect 12809 -13676 12852 -13644
rect 12852 -13676 12884 -13644
rect 12884 -13676 12927 -13644
rect 12809 -13719 12927 -13676
rect 12809 -13804 12927 -13761
rect 12809 -13836 12852 -13804
rect 12852 -13836 12884 -13804
rect 12884 -13836 12927 -13804
rect 12809 -13879 12927 -13836
rect 12809 -13964 12927 -13921
rect 12809 -13996 12852 -13964
rect 12852 -13996 12884 -13964
rect 12884 -13996 12927 -13964
rect 12809 -14039 12927 -13996
rect 12809 -14124 12927 -14081
rect 12809 -14156 12852 -14124
rect 12852 -14156 12884 -14124
rect 12884 -14156 12927 -14124
rect 12809 -14199 12927 -14156
rect 12809 -14284 12927 -14241
rect 12809 -14316 12852 -14284
rect 12852 -14316 12884 -14284
rect 12884 -14316 12927 -14284
rect 12809 -14359 12927 -14316
rect 12809 -14444 12927 -14401
rect 12809 -14476 12852 -14444
rect 12852 -14476 12884 -14444
rect 12884 -14476 12927 -14444
rect 12809 -14519 12927 -14476
rect 12809 -14604 12927 -14561
rect 12809 -14636 12852 -14604
rect 12852 -14636 12884 -14604
rect 12884 -14636 12927 -14604
rect 12809 -14679 12927 -14636
rect 12809 -14764 12927 -14721
rect 12809 -14796 12852 -14764
rect 12852 -14796 12884 -14764
rect 12884 -14796 12927 -14764
rect 12809 -14839 12927 -14796
rect 12809 -14924 12927 -14881
rect 12809 -14956 12852 -14924
rect 12852 -14956 12884 -14924
rect 12884 -14956 12927 -14924
rect 12809 -14999 12927 -14956
rect 12809 -15084 12927 -15041
rect 12809 -15116 12852 -15084
rect 12852 -15116 12884 -15084
rect 12884 -15116 12927 -15084
rect 12809 -15159 12927 -15116
rect 9076 -15276 9119 -15244
rect 9119 -15276 9151 -15244
rect 9151 -15276 9194 -15244
rect 9076 -15319 9194 -15276
rect 12809 -15244 12927 -15201
rect 12809 -15276 12852 -15244
rect 12852 -15276 12884 -15244
rect 12884 -15276 12927 -15244
rect 9261 -15349 9379 -15306
rect 9261 -15381 9304 -15349
rect 9304 -15381 9336 -15349
rect 9336 -15381 9379 -15349
rect 9261 -15424 9379 -15381
rect 9421 -15349 9539 -15306
rect 9421 -15381 9464 -15349
rect 9464 -15381 9496 -15349
rect 9496 -15381 9539 -15349
rect 9421 -15424 9539 -15381
rect 9581 -15349 9699 -15306
rect 9581 -15381 9624 -15349
rect 9624 -15381 9656 -15349
rect 9656 -15381 9699 -15349
rect 9581 -15424 9699 -15381
rect 9741 -15349 9859 -15306
rect 9741 -15381 9784 -15349
rect 9784 -15381 9816 -15349
rect 9816 -15381 9859 -15349
rect 9741 -15424 9859 -15381
rect 9901 -15349 10019 -15306
rect 9901 -15381 9944 -15349
rect 9944 -15381 9976 -15349
rect 9976 -15381 10019 -15349
rect 9901 -15424 10019 -15381
rect 10061 -15349 10179 -15306
rect 10061 -15381 10104 -15349
rect 10104 -15381 10136 -15349
rect 10136 -15381 10179 -15349
rect 10061 -15424 10179 -15381
rect 10221 -15349 10339 -15306
rect 10221 -15381 10264 -15349
rect 10264 -15381 10296 -15349
rect 10296 -15381 10339 -15349
rect 10221 -15424 10339 -15381
rect 10381 -15349 10499 -15306
rect 10381 -15381 10424 -15349
rect 10424 -15381 10456 -15349
rect 10456 -15381 10499 -15349
rect 10381 -15424 10499 -15381
rect 10541 -15349 10659 -15306
rect 10541 -15381 10584 -15349
rect 10584 -15381 10616 -15349
rect 10616 -15381 10659 -15349
rect 10541 -15424 10659 -15381
rect 10701 -15349 10819 -15306
rect 10701 -15381 10744 -15349
rect 10744 -15381 10776 -15349
rect 10776 -15381 10819 -15349
rect 10701 -15424 10819 -15381
rect 10861 -15349 10979 -15306
rect 10861 -15381 10904 -15349
rect 10904 -15381 10936 -15349
rect 10936 -15381 10979 -15349
rect 10861 -15424 10979 -15381
rect 11021 -15349 11139 -15306
rect 11021 -15381 11064 -15349
rect 11064 -15381 11096 -15349
rect 11096 -15381 11139 -15349
rect 11021 -15424 11139 -15381
rect 11181 -15349 11299 -15306
rect 11181 -15381 11224 -15349
rect 11224 -15381 11256 -15349
rect 11256 -15381 11299 -15349
rect 11181 -15424 11299 -15381
rect 11341 -15349 11459 -15306
rect 11341 -15381 11384 -15349
rect 11384 -15381 11416 -15349
rect 11416 -15381 11459 -15349
rect 11341 -15424 11459 -15381
rect 11501 -15349 11619 -15306
rect 11501 -15381 11544 -15349
rect 11544 -15381 11576 -15349
rect 11576 -15381 11619 -15349
rect 11501 -15424 11619 -15381
rect 11661 -15349 11779 -15306
rect 11661 -15381 11704 -15349
rect 11704 -15381 11736 -15349
rect 11736 -15381 11779 -15349
rect 11661 -15424 11779 -15381
rect 11821 -15349 11939 -15306
rect 11821 -15381 11864 -15349
rect 11864 -15381 11896 -15349
rect 11896 -15381 11939 -15349
rect 11821 -15424 11939 -15381
rect 11981 -15349 12099 -15306
rect 11981 -15381 12024 -15349
rect 12024 -15381 12056 -15349
rect 12056 -15381 12099 -15349
rect 11981 -15424 12099 -15381
rect 12141 -15349 12259 -15306
rect 12141 -15381 12184 -15349
rect 12184 -15381 12216 -15349
rect 12216 -15381 12259 -15349
rect 12141 -15424 12259 -15381
rect 12301 -15349 12419 -15306
rect 12301 -15381 12344 -15349
rect 12344 -15381 12376 -15349
rect 12376 -15381 12419 -15349
rect 12301 -15424 12419 -15381
rect 12461 -15349 12579 -15306
rect 12461 -15381 12504 -15349
rect 12504 -15381 12536 -15349
rect 12536 -15381 12579 -15349
rect 12461 -15424 12579 -15381
rect 12621 -15349 12739 -15306
rect 12809 -15319 12927 -15276
rect 12621 -15381 12664 -15349
rect 12664 -15381 12696 -15349
rect 12696 -15381 12739 -15349
rect 12621 -15424 12739 -15381
rect 15261 -11621 15379 -11578
rect 15261 -11653 15304 -11621
rect 15304 -11653 15336 -11621
rect 15336 -11653 15379 -11621
rect 15076 -11724 15194 -11681
rect 15261 -11696 15379 -11653
rect 15421 -11621 15539 -11578
rect 15421 -11653 15464 -11621
rect 15464 -11653 15496 -11621
rect 15496 -11653 15539 -11621
rect 15421 -11696 15539 -11653
rect 15581 -11621 15699 -11578
rect 15581 -11653 15624 -11621
rect 15624 -11653 15656 -11621
rect 15656 -11653 15699 -11621
rect 15581 -11696 15699 -11653
rect 15741 -11621 15859 -11578
rect 15741 -11653 15784 -11621
rect 15784 -11653 15816 -11621
rect 15816 -11653 15859 -11621
rect 15741 -11696 15859 -11653
rect 15901 -11621 16019 -11578
rect 15901 -11653 15944 -11621
rect 15944 -11653 15976 -11621
rect 15976 -11653 16019 -11621
rect 15901 -11696 16019 -11653
rect 16061 -11621 16179 -11578
rect 16061 -11653 16104 -11621
rect 16104 -11653 16136 -11621
rect 16136 -11653 16179 -11621
rect 16061 -11696 16179 -11653
rect 16221 -11621 16339 -11578
rect 16221 -11653 16264 -11621
rect 16264 -11653 16296 -11621
rect 16296 -11653 16339 -11621
rect 16221 -11696 16339 -11653
rect 16381 -11621 16499 -11578
rect 16381 -11653 16424 -11621
rect 16424 -11653 16456 -11621
rect 16456 -11653 16499 -11621
rect 16381 -11696 16499 -11653
rect 16541 -11621 16659 -11578
rect 16541 -11653 16584 -11621
rect 16584 -11653 16616 -11621
rect 16616 -11653 16659 -11621
rect 16541 -11696 16659 -11653
rect 16701 -11621 16819 -11578
rect 16701 -11653 16744 -11621
rect 16744 -11653 16776 -11621
rect 16776 -11653 16819 -11621
rect 16701 -11696 16819 -11653
rect 16861 -11621 16979 -11578
rect 16861 -11653 16904 -11621
rect 16904 -11653 16936 -11621
rect 16936 -11653 16979 -11621
rect 16861 -11696 16979 -11653
rect 17021 -11621 17139 -11578
rect 17021 -11653 17064 -11621
rect 17064 -11653 17096 -11621
rect 17096 -11653 17139 -11621
rect 17021 -11696 17139 -11653
rect 17181 -11621 17299 -11578
rect 17181 -11653 17224 -11621
rect 17224 -11653 17256 -11621
rect 17256 -11653 17299 -11621
rect 17181 -11696 17299 -11653
rect 17341 -11621 17459 -11578
rect 17341 -11653 17384 -11621
rect 17384 -11653 17416 -11621
rect 17416 -11653 17459 -11621
rect 17341 -11696 17459 -11653
rect 17501 -11621 17619 -11578
rect 17501 -11653 17544 -11621
rect 17544 -11653 17576 -11621
rect 17576 -11653 17619 -11621
rect 17501 -11696 17619 -11653
rect 17661 -11621 17779 -11578
rect 17661 -11653 17704 -11621
rect 17704 -11653 17736 -11621
rect 17736 -11653 17779 -11621
rect 17661 -11696 17779 -11653
rect 17821 -11621 17939 -11578
rect 17821 -11653 17864 -11621
rect 17864 -11653 17896 -11621
rect 17896 -11653 17939 -11621
rect 17821 -11696 17939 -11653
rect 17981 -11621 18099 -11578
rect 17981 -11653 18024 -11621
rect 18024 -11653 18056 -11621
rect 18056 -11653 18099 -11621
rect 17981 -11696 18099 -11653
rect 18141 -11621 18259 -11578
rect 18141 -11653 18184 -11621
rect 18184 -11653 18216 -11621
rect 18216 -11653 18259 -11621
rect 18141 -11696 18259 -11653
rect 18301 -11621 18419 -11578
rect 18301 -11653 18344 -11621
rect 18344 -11653 18376 -11621
rect 18376 -11653 18419 -11621
rect 18301 -11696 18419 -11653
rect 18461 -11621 18579 -11578
rect 18461 -11653 18504 -11621
rect 18504 -11653 18536 -11621
rect 18536 -11653 18579 -11621
rect 18461 -11696 18579 -11653
rect 18621 -11621 18739 -11578
rect 18621 -11653 18664 -11621
rect 18664 -11653 18696 -11621
rect 18696 -11653 18739 -11621
rect 18621 -11696 18739 -11653
rect 15076 -11756 15119 -11724
rect 15119 -11756 15151 -11724
rect 15151 -11756 15194 -11724
rect 15076 -11799 15194 -11756
rect 18809 -11724 18927 -11681
rect 18809 -11756 18852 -11724
rect 18852 -11756 18884 -11724
rect 18884 -11756 18927 -11724
rect 15076 -11884 15194 -11841
rect 15076 -11916 15119 -11884
rect 15119 -11916 15151 -11884
rect 15151 -11916 15194 -11884
rect 15076 -11959 15194 -11916
rect 15076 -12044 15194 -12001
rect 15076 -12076 15119 -12044
rect 15119 -12076 15151 -12044
rect 15151 -12076 15194 -12044
rect 15076 -12119 15194 -12076
rect 15076 -12204 15194 -12161
rect 15076 -12236 15119 -12204
rect 15119 -12236 15151 -12204
rect 15151 -12236 15194 -12204
rect 15076 -12279 15194 -12236
rect 15076 -12364 15194 -12321
rect 15076 -12396 15119 -12364
rect 15119 -12396 15151 -12364
rect 15151 -12396 15194 -12364
rect 15076 -12439 15194 -12396
rect 15076 -12524 15194 -12481
rect 15076 -12556 15119 -12524
rect 15119 -12556 15151 -12524
rect 15151 -12556 15194 -12524
rect 15076 -12599 15194 -12556
rect 15076 -12684 15194 -12641
rect 15076 -12716 15119 -12684
rect 15119 -12716 15151 -12684
rect 15151 -12716 15194 -12684
rect 15076 -12759 15194 -12716
rect 15076 -12844 15194 -12801
rect 15076 -12876 15119 -12844
rect 15119 -12876 15151 -12844
rect 15151 -12876 15194 -12844
rect 15076 -12919 15194 -12876
rect 15076 -13004 15194 -12961
rect 15076 -13036 15119 -13004
rect 15119 -13036 15151 -13004
rect 15151 -13036 15194 -13004
rect 15076 -13079 15194 -13036
rect 15076 -13164 15194 -13121
rect 15076 -13196 15119 -13164
rect 15119 -13196 15151 -13164
rect 15151 -13196 15194 -13164
rect 15076 -13239 15194 -13196
rect 15076 -13324 15194 -13281
rect 15076 -13356 15119 -13324
rect 15119 -13356 15151 -13324
rect 15151 -13356 15194 -13324
rect 15076 -13399 15194 -13356
rect 15076 -13484 15194 -13441
rect 15076 -13516 15119 -13484
rect 15119 -13516 15151 -13484
rect 15151 -13516 15194 -13484
rect 15076 -13559 15194 -13516
rect 15076 -13644 15194 -13601
rect 15076 -13676 15119 -13644
rect 15119 -13676 15151 -13644
rect 15151 -13676 15194 -13644
rect 15076 -13719 15194 -13676
rect 15076 -13804 15194 -13761
rect 15076 -13836 15119 -13804
rect 15119 -13836 15151 -13804
rect 15151 -13836 15194 -13804
rect 15076 -13879 15194 -13836
rect 15076 -13964 15194 -13921
rect 15076 -13996 15119 -13964
rect 15119 -13996 15151 -13964
rect 15151 -13996 15194 -13964
rect 15076 -14039 15194 -13996
rect 15076 -14124 15194 -14081
rect 15076 -14156 15119 -14124
rect 15119 -14156 15151 -14124
rect 15151 -14156 15194 -14124
rect 15076 -14199 15194 -14156
rect 15076 -14284 15194 -14241
rect 15076 -14316 15119 -14284
rect 15119 -14316 15151 -14284
rect 15151 -14316 15194 -14284
rect 15076 -14359 15194 -14316
rect 15076 -14444 15194 -14401
rect 15076 -14476 15119 -14444
rect 15119 -14476 15151 -14444
rect 15151 -14476 15194 -14444
rect 15076 -14519 15194 -14476
rect 15076 -14604 15194 -14561
rect 15076 -14636 15119 -14604
rect 15119 -14636 15151 -14604
rect 15151 -14636 15194 -14604
rect 15076 -14679 15194 -14636
rect 15076 -14764 15194 -14721
rect 15076 -14796 15119 -14764
rect 15119 -14796 15151 -14764
rect 15151 -14796 15194 -14764
rect 15076 -14839 15194 -14796
rect 15076 -14924 15194 -14881
rect 15076 -14956 15119 -14924
rect 15119 -14956 15151 -14924
rect 15151 -14956 15194 -14924
rect 15076 -14999 15194 -14956
rect 15076 -15084 15194 -15041
rect 15076 -15116 15119 -15084
rect 15119 -15116 15151 -15084
rect 15151 -15116 15194 -15084
rect 15076 -15159 15194 -15116
rect 15076 -15244 15194 -15201
rect 18809 -11799 18927 -11756
rect 18809 -11884 18927 -11841
rect 18809 -11916 18852 -11884
rect 18852 -11916 18884 -11884
rect 18884 -11916 18927 -11884
rect 18809 -11959 18927 -11916
rect 18809 -12044 18927 -12001
rect 18809 -12076 18852 -12044
rect 18852 -12076 18884 -12044
rect 18884 -12076 18927 -12044
rect 18809 -12119 18927 -12076
rect 18809 -12204 18927 -12161
rect 18809 -12236 18852 -12204
rect 18852 -12236 18884 -12204
rect 18884 -12236 18927 -12204
rect 18809 -12279 18927 -12236
rect 18809 -12364 18927 -12321
rect 18809 -12396 18852 -12364
rect 18852 -12396 18884 -12364
rect 18884 -12396 18927 -12364
rect 18809 -12439 18927 -12396
rect 18809 -12524 18927 -12481
rect 18809 -12556 18852 -12524
rect 18852 -12556 18884 -12524
rect 18884 -12556 18927 -12524
rect 18809 -12599 18927 -12556
rect 18809 -12684 18927 -12641
rect 18809 -12716 18852 -12684
rect 18852 -12716 18884 -12684
rect 18884 -12716 18927 -12684
rect 18809 -12759 18927 -12716
rect 18809 -12844 18927 -12801
rect 18809 -12876 18852 -12844
rect 18852 -12876 18884 -12844
rect 18884 -12876 18927 -12844
rect 18809 -12919 18927 -12876
rect 18809 -13004 18927 -12961
rect 18809 -13036 18852 -13004
rect 18852 -13036 18884 -13004
rect 18884 -13036 18927 -13004
rect 18809 -13079 18927 -13036
rect 18809 -13164 18927 -13121
rect 18809 -13196 18852 -13164
rect 18852 -13196 18884 -13164
rect 18884 -13196 18927 -13164
rect 18809 -13239 18927 -13196
rect 18809 -13324 18927 -13281
rect 18809 -13356 18852 -13324
rect 18852 -13356 18884 -13324
rect 18884 -13356 18927 -13324
rect 18809 -13399 18927 -13356
rect 18809 -13484 18927 -13441
rect 18809 -13516 18852 -13484
rect 18852 -13516 18884 -13484
rect 18884 -13516 18927 -13484
rect 18809 -13559 18927 -13516
rect 18809 -13644 18927 -13601
rect 18809 -13676 18852 -13644
rect 18852 -13676 18884 -13644
rect 18884 -13676 18927 -13644
rect 18809 -13719 18927 -13676
rect 18809 -13804 18927 -13761
rect 18809 -13836 18852 -13804
rect 18852 -13836 18884 -13804
rect 18884 -13836 18927 -13804
rect 18809 -13879 18927 -13836
rect 18809 -13964 18927 -13921
rect 18809 -13996 18852 -13964
rect 18852 -13996 18884 -13964
rect 18884 -13996 18927 -13964
rect 18809 -14039 18927 -13996
rect 18809 -14124 18927 -14081
rect 18809 -14156 18852 -14124
rect 18852 -14156 18884 -14124
rect 18884 -14156 18927 -14124
rect 18809 -14199 18927 -14156
rect 18809 -14284 18927 -14241
rect 18809 -14316 18852 -14284
rect 18852 -14316 18884 -14284
rect 18884 -14316 18927 -14284
rect 18809 -14359 18927 -14316
rect 18809 -14444 18927 -14401
rect 18809 -14476 18852 -14444
rect 18852 -14476 18884 -14444
rect 18884 -14476 18927 -14444
rect 18809 -14519 18927 -14476
rect 18809 -14604 18927 -14561
rect 18809 -14636 18852 -14604
rect 18852 -14636 18884 -14604
rect 18884 -14636 18927 -14604
rect 18809 -14679 18927 -14636
rect 18809 -14764 18927 -14721
rect 18809 -14796 18852 -14764
rect 18852 -14796 18884 -14764
rect 18884 -14796 18927 -14764
rect 18809 -14839 18927 -14796
rect 18809 -14924 18927 -14881
rect 18809 -14956 18852 -14924
rect 18852 -14956 18884 -14924
rect 18884 -14956 18927 -14924
rect 18809 -14999 18927 -14956
rect 18809 -15084 18927 -15041
rect 18809 -15116 18852 -15084
rect 18852 -15116 18884 -15084
rect 18884 -15116 18927 -15084
rect 18809 -15159 18927 -15116
rect 15076 -15276 15119 -15244
rect 15119 -15276 15151 -15244
rect 15151 -15276 15194 -15244
rect 15076 -15319 15194 -15276
rect 18809 -15244 18927 -15201
rect 18809 -15276 18852 -15244
rect 18852 -15276 18884 -15244
rect 18884 -15276 18927 -15244
rect 15261 -15349 15379 -15306
rect 15261 -15381 15304 -15349
rect 15304 -15381 15336 -15349
rect 15336 -15381 15379 -15349
rect 15261 -15424 15379 -15381
rect 15421 -15349 15539 -15306
rect 15421 -15381 15464 -15349
rect 15464 -15381 15496 -15349
rect 15496 -15381 15539 -15349
rect 15421 -15424 15539 -15381
rect 15581 -15349 15699 -15306
rect 15581 -15381 15624 -15349
rect 15624 -15381 15656 -15349
rect 15656 -15381 15699 -15349
rect 15581 -15424 15699 -15381
rect 15741 -15349 15859 -15306
rect 15741 -15381 15784 -15349
rect 15784 -15381 15816 -15349
rect 15816 -15381 15859 -15349
rect 15741 -15424 15859 -15381
rect 15901 -15349 16019 -15306
rect 15901 -15381 15944 -15349
rect 15944 -15381 15976 -15349
rect 15976 -15381 16019 -15349
rect 15901 -15424 16019 -15381
rect 16061 -15349 16179 -15306
rect 16061 -15381 16104 -15349
rect 16104 -15381 16136 -15349
rect 16136 -15381 16179 -15349
rect 16061 -15424 16179 -15381
rect 16221 -15349 16339 -15306
rect 16221 -15381 16264 -15349
rect 16264 -15381 16296 -15349
rect 16296 -15381 16339 -15349
rect 16221 -15424 16339 -15381
rect 16381 -15349 16499 -15306
rect 16381 -15381 16424 -15349
rect 16424 -15381 16456 -15349
rect 16456 -15381 16499 -15349
rect 16381 -15424 16499 -15381
rect 16541 -15349 16659 -15306
rect 16541 -15381 16584 -15349
rect 16584 -15381 16616 -15349
rect 16616 -15381 16659 -15349
rect 16541 -15424 16659 -15381
rect 16701 -15349 16819 -15306
rect 16701 -15381 16744 -15349
rect 16744 -15381 16776 -15349
rect 16776 -15381 16819 -15349
rect 16701 -15424 16819 -15381
rect 16861 -15349 16979 -15306
rect 16861 -15381 16904 -15349
rect 16904 -15381 16936 -15349
rect 16936 -15381 16979 -15349
rect 16861 -15424 16979 -15381
rect 17021 -15349 17139 -15306
rect 17021 -15381 17064 -15349
rect 17064 -15381 17096 -15349
rect 17096 -15381 17139 -15349
rect 17021 -15424 17139 -15381
rect 17181 -15349 17299 -15306
rect 17181 -15381 17224 -15349
rect 17224 -15381 17256 -15349
rect 17256 -15381 17299 -15349
rect 17181 -15424 17299 -15381
rect 17341 -15349 17459 -15306
rect 17341 -15381 17384 -15349
rect 17384 -15381 17416 -15349
rect 17416 -15381 17459 -15349
rect 17341 -15424 17459 -15381
rect 17501 -15349 17619 -15306
rect 17501 -15381 17544 -15349
rect 17544 -15381 17576 -15349
rect 17576 -15381 17619 -15349
rect 17501 -15424 17619 -15381
rect 17661 -15349 17779 -15306
rect 17661 -15381 17704 -15349
rect 17704 -15381 17736 -15349
rect 17736 -15381 17779 -15349
rect 17661 -15424 17779 -15381
rect 17821 -15349 17939 -15306
rect 17821 -15381 17864 -15349
rect 17864 -15381 17896 -15349
rect 17896 -15381 17939 -15349
rect 17821 -15424 17939 -15381
rect 17981 -15349 18099 -15306
rect 17981 -15381 18024 -15349
rect 18024 -15381 18056 -15349
rect 18056 -15381 18099 -15349
rect 17981 -15424 18099 -15381
rect 18141 -15349 18259 -15306
rect 18141 -15381 18184 -15349
rect 18184 -15381 18216 -15349
rect 18216 -15381 18259 -15349
rect 18141 -15424 18259 -15381
rect 18301 -15349 18419 -15306
rect 18301 -15381 18344 -15349
rect 18344 -15381 18376 -15349
rect 18376 -15381 18419 -15349
rect 18301 -15424 18419 -15381
rect 18461 -15349 18579 -15306
rect 18461 -15381 18504 -15349
rect 18504 -15381 18536 -15349
rect 18536 -15381 18579 -15349
rect 18461 -15424 18579 -15381
rect 18621 -15349 18739 -15306
rect 18809 -15319 18927 -15276
rect 18621 -15381 18664 -15349
rect 18664 -15381 18696 -15349
rect 18696 -15381 18739 -15349
rect 18621 -15424 18739 -15381
rect 21261 -11621 21379 -11578
rect 21261 -11653 21304 -11621
rect 21304 -11653 21336 -11621
rect 21336 -11653 21379 -11621
rect 21076 -11724 21194 -11681
rect 21261 -11696 21379 -11653
rect 21421 -11621 21539 -11578
rect 21421 -11653 21464 -11621
rect 21464 -11653 21496 -11621
rect 21496 -11653 21539 -11621
rect 21421 -11696 21539 -11653
rect 21581 -11621 21699 -11578
rect 21581 -11653 21624 -11621
rect 21624 -11653 21656 -11621
rect 21656 -11653 21699 -11621
rect 21581 -11696 21699 -11653
rect 21741 -11621 21859 -11578
rect 21741 -11653 21784 -11621
rect 21784 -11653 21816 -11621
rect 21816 -11653 21859 -11621
rect 21741 -11696 21859 -11653
rect 21901 -11621 22019 -11578
rect 21901 -11653 21944 -11621
rect 21944 -11653 21976 -11621
rect 21976 -11653 22019 -11621
rect 21901 -11696 22019 -11653
rect 22061 -11621 22179 -11578
rect 22061 -11653 22104 -11621
rect 22104 -11653 22136 -11621
rect 22136 -11653 22179 -11621
rect 22061 -11696 22179 -11653
rect 22221 -11621 22339 -11578
rect 22221 -11653 22264 -11621
rect 22264 -11653 22296 -11621
rect 22296 -11653 22339 -11621
rect 22221 -11696 22339 -11653
rect 22381 -11621 22499 -11578
rect 22381 -11653 22424 -11621
rect 22424 -11653 22456 -11621
rect 22456 -11653 22499 -11621
rect 22381 -11696 22499 -11653
rect 22541 -11621 22659 -11578
rect 22541 -11653 22584 -11621
rect 22584 -11653 22616 -11621
rect 22616 -11653 22659 -11621
rect 22541 -11696 22659 -11653
rect 22701 -11621 22819 -11578
rect 22701 -11653 22744 -11621
rect 22744 -11653 22776 -11621
rect 22776 -11653 22819 -11621
rect 22701 -11696 22819 -11653
rect 22861 -11621 22979 -11578
rect 22861 -11653 22904 -11621
rect 22904 -11653 22936 -11621
rect 22936 -11653 22979 -11621
rect 22861 -11696 22979 -11653
rect 23021 -11621 23139 -11578
rect 23021 -11653 23064 -11621
rect 23064 -11653 23096 -11621
rect 23096 -11653 23139 -11621
rect 23021 -11696 23139 -11653
rect 23181 -11621 23299 -11578
rect 23181 -11653 23224 -11621
rect 23224 -11653 23256 -11621
rect 23256 -11653 23299 -11621
rect 23181 -11696 23299 -11653
rect 23341 -11621 23459 -11578
rect 23341 -11653 23384 -11621
rect 23384 -11653 23416 -11621
rect 23416 -11653 23459 -11621
rect 23341 -11696 23459 -11653
rect 23501 -11621 23619 -11578
rect 23501 -11653 23544 -11621
rect 23544 -11653 23576 -11621
rect 23576 -11653 23619 -11621
rect 23501 -11696 23619 -11653
rect 23661 -11621 23779 -11578
rect 23661 -11653 23704 -11621
rect 23704 -11653 23736 -11621
rect 23736 -11653 23779 -11621
rect 23661 -11696 23779 -11653
rect 23821 -11621 23939 -11578
rect 23821 -11653 23864 -11621
rect 23864 -11653 23896 -11621
rect 23896 -11653 23939 -11621
rect 23821 -11696 23939 -11653
rect 23981 -11621 24099 -11578
rect 23981 -11653 24024 -11621
rect 24024 -11653 24056 -11621
rect 24056 -11653 24099 -11621
rect 23981 -11696 24099 -11653
rect 24141 -11621 24259 -11578
rect 24141 -11653 24184 -11621
rect 24184 -11653 24216 -11621
rect 24216 -11653 24259 -11621
rect 24141 -11696 24259 -11653
rect 24301 -11621 24419 -11578
rect 24301 -11653 24344 -11621
rect 24344 -11653 24376 -11621
rect 24376 -11653 24419 -11621
rect 24301 -11696 24419 -11653
rect 24461 -11621 24579 -11578
rect 24461 -11653 24504 -11621
rect 24504 -11653 24536 -11621
rect 24536 -11653 24579 -11621
rect 24461 -11696 24579 -11653
rect 24621 -11621 24739 -11578
rect 24621 -11653 24664 -11621
rect 24664 -11653 24696 -11621
rect 24696 -11653 24739 -11621
rect 24621 -11696 24739 -11653
rect 21076 -11756 21119 -11724
rect 21119 -11756 21151 -11724
rect 21151 -11756 21194 -11724
rect 21076 -11799 21194 -11756
rect 24809 -11724 24927 -11681
rect 24809 -11756 24852 -11724
rect 24852 -11756 24884 -11724
rect 24884 -11756 24927 -11724
rect 21076 -11884 21194 -11841
rect 21076 -11916 21119 -11884
rect 21119 -11916 21151 -11884
rect 21151 -11916 21194 -11884
rect 21076 -11959 21194 -11916
rect 21076 -12044 21194 -12001
rect 21076 -12076 21119 -12044
rect 21119 -12076 21151 -12044
rect 21151 -12076 21194 -12044
rect 21076 -12119 21194 -12076
rect 21076 -12204 21194 -12161
rect 21076 -12236 21119 -12204
rect 21119 -12236 21151 -12204
rect 21151 -12236 21194 -12204
rect 21076 -12279 21194 -12236
rect 21076 -12364 21194 -12321
rect 21076 -12396 21119 -12364
rect 21119 -12396 21151 -12364
rect 21151 -12396 21194 -12364
rect 21076 -12439 21194 -12396
rect 21076 -12524 21194 -12481
rect 21076 -12556 21119 -12524
rect 21119 -12556 21151 -12524
rect 21151 -12556 21194 -12524
rect 21076 -12599 21194 -12556
rect 21076 -12684 21194 -12641
rect 21076 -12716 21119 -12684
rect 21119 -12716 21151 -12684
rect 21151 -12716 21194 -12684
rect 21076 -12759 21194 -12716
rect 21076 -12844 21194 -12801
rect 21076 -12876 21119 -12844
rect 21119 -12876 21151 -12844
rect 21151 -12876 21194 -12844
rect 21076 -12919 21194 -12876
rect 21076 -13004 21194 -12961
rect 21076 -13036 21119 -13004
rect 21119 -13036 21151 -13004
rect 21151 -13036 21194 -13004
rect 21076 -13079 21194 -13036
rect 21076 -13164 21194 -13121
rect 21076 -13196 21119 -13164
rect 21119 -13196 21151 -13164
rect 21151 -13196 21194 -13164
rect 21076 -13239 21194 -13196
rect 21076 -13324 21194 -13281
rect 21076 -13356 21119 -13324
rect 21119 -13356 21151 -13324
rect 21151 -13356 21194 -13324
rect 21076 -13399 21194 -13356
rect 21076 -13484 21194 -13441
rect 21076 -13516 21119 -13484
rect 21119 -13516 21151 -13484
rect 21151 -13516 21194 -13484
rect 21076 -13559 21194 -13516
rect 21076 -13644 21194 -13601
rect 21076 -13676 21119 -13644
rect 21119 -13676 21151 -13644
rect 21151 -13676 21194 -13644
rect 21076 -13719 21194 -13676
rect 21076 -13804 21194 -13761
rect 21076 -13836 21119 -13804
rect 21119 -13836 21151 -13804
rect 21151 -13836 21194 -13804
rect 21076 -13879 21194 -13836
rect 21076 -13964 21194 -13921
rect 21076 -13996 21119 -13964
rect 21119 -13996 21151 -13964
rect 21151 -13996 21194 -13964
rect 21076 -14039 21194 -13996
rect 21076 -14124 21194 -14081
rect 21076 -14156 21119 -14124
rect 21119 -14156 21151 -14124
rect 21151 -14156 21194 -14124
rect 21076 -14199 21194 -14156
rect 21076 -14284 21194 -14241
rect 21076 -14316 21119 -14284
rect 21119 -14316 21151 -14284
rect 21151 -14316 21194 -14284
rect 21076 -14359 21194 -14316
rect 21076 -14444 21194 -14401
rect 21076 -14476 21119 -14444
rect 21119 -14476 21151 -14444
rect 21151 -14476 21194 -14444
rect 21076 -14519 21194 -14476
rect 21076 -14604 21194 -14561
rect 21076 -14636 21119 -14604
rect 21119 -14636 21151 -14604
rect 21151 -14636 21194 -14604
rect 21076 -14679 21194 -14636
rect 21076 -14764 21194 -14721
rect 21076 -14796 21119 -14764
rect 21119 -14796 21151 -14764
rect 21151 -14796 21194 -14764
rect 21076 -14839 21194 -14796
rect 21076 -14924 21194 -14881
rect 21076 -14956 21119 -14924
rect 21119 -14956 21151 -14924
rect 21151 -14956 21194 -14924
rect 21076 -14999 21194 -14956
rect 21076 -15084 21194 -15041
rect 21076 -15116 21119 -15084
rect 21119 -15116 21151 -15084
rect 21151 -15116 21194 -15084
rect 21076 -15159 21194 -15116
rect 21076 -15244 21194 -15201
rect 24809 -11799 24927 -11756
rect 24809 -11884 24927 -11841
rect 24809 -11916 24852 -11884
rect 24852 -11916 24884 -11884
rect 24884 -11916 24927 -11884
rect 24809 -11959 24927 -11916
rect 24809 -12044 24927 -12001
rect 24809 -12076 24852 -12044
rect 24852 -12076 24884 -12044
rect 24884 -12076 24927 -12044
rect 24809 -12119 24927 -12076
rect 24809 -12204 24927 -12161
rect 24809 -12236 24852 -12204
rect 24852 -12236 24884 -12204
rect 24884 -12236 24927 -12204
rect 24809 -12279 24927 -12236
rect 24809 -12364 24927 -12321
rect 24809 -12396 24852 -12364
rect 24852 -12396 24884 -12364
rect 24884 -12396 24927 -12364
rect 24809 -12439 24927 -12396
rect 24809 -12524 24927 -12481
rect 24809 -12556 24852 -12524
rect 24852 -12556 24884 -12524
rect 24884 -12556 24927 -12524
rect 24809 -12599 24927 -12556
rect 24809 -12684 24927 -12641
rect 24809 -12716 24852 -12684
rect 24852 -12716 24884 -12684
rect 24884 -12716 24927 -12684
rect 24809 -12759 24927 -12716
rect 24809 -12844 24927 -12801
rect 24809 -12876 24852 -12844
rect 24852 -12876 24884 -12844
rect 24884 -12876 24927 -12844
rect 24809 -12919 24927 -12876
rect 24809 -13004 24927 -12961
rect 24809 -13036 24852 -13004
rect 24852 -13036 24884 -13004
rect 24884 -13036 24927 -13004
rect 24809 -13079 24927 -13036
rect 24809 -13164 24927 -13121
rect 24809 -13196 24852 -13164
rect 24852 -13196 24884 -13164
rect 24884 -13196 24927 -13164
rect 24809 -13239 24927 -13196
rect 24809 -13324 24927 -13281
rect 24809 -13356 24852 -13324
rect 24852 -13356 24884 -13324
rect 24884 -13356 24927 -13324
rect 24809 -13399 24927 -13356
rect 24809 -13484 24927 -13441
rect 24809 -13516 24852 -13484
rect 24852 -13516 24884 -13484
rect 24884 -13516 24927 -13484
rect 24809 -13559 24927 -13516
rect 24809 -13644 24927 -13601
rect 24809 -13676 24852 -13644
rect 24852 -13676 24884 -13644
rect 24884 -13676 24927 -13644
rect 24809 -13719 24927 -13676
rect 24809 -13804 24927 -13761
rect 24809 -13836 24852 -13804
rect 24852 -13836 24884 -13804
rect 24884 -13836 24927 -13804
rect 24809 -13879 24927 -13836
rect 24809 -13964 24927 -13921
rect 24809 -13996 24852 -13964
rect 24852 -13996 24884 -13964
rect 24884 -13996 24927 -13964
rect 24809 -14039 24927 -13996
rect 24809 -14124 24927 -14081
rect 24809 -14156 24852 -14124
rect 24852 -14156 24884 -14124
rect 24884 -14156 24927 -14124
rect 24809 -14199 24927 -14156
rect 24809 -14284 24927 -14241
rect 24809 -14316 24852 -14284
rect 24852 -14316 24884 -14284
rect 24884 -14316 24927 -14284
rect 24809 -14359 24927 -14316
rect 24809 -14444 24927 -14401
rect 24809 -14476 24852 -14444
rect 24852 -14476 24884 -14444
rect 24884 -14476 24927 -14444
rect 24809 -14519 24927 -14476
rect 24809 -14604 24927 -14561
rect 24809 -14636 24852 -14604
rect 24852 -14636 24884 -14604
rect 24884 -14636 24927 -14604
rect 24809 -14679 24927 -14636
rect 24809 -14764 24927 -14721
rect 24809 -14796 24852 -14764
rect 24852 -14796 24884 -14764
rect 24884 -14796 24927 -14764
rect 24809 -14839 24927 -14796
rect 24809 -14924 24927 -14881
rect 24809 -14956 24852 -14924
rect 24852 -14956 24884 -14924
rect 24884 -14956 24927 -14924
rect 24809 -14999 24927 -14956
rect 24809 -15084 24927 -15041
rect 24809 -15116 24852 -15084
rect 24852 -15116 24884 -15084
rect 24884 -15116 24927 -15084
rect 24809 -15159 24927 -15116
rect 21076 -15276 21119 -15244
rect 21119 -15276 21151 -15244
rect 21151 -15276 21194 -15244
rect 21076 -15319 21194 -15276
rect 24809 -15244 24927 -15201
rect 24809 -15276 24852 -15244
rect 24852 -15276 24884 -15244
rect 24884 -15276 24927 -15244
rect 21261 -15349 21379 -15306
rect 21261 -15381 21304 -15349
rect 21304 -15381 21336 -15349
rect 21336 -15381 21379 -15349
rect 21261 -15424 21379 -15381
rect 21421 -15349 21539 -15306
rect 21421 -15381 21464 -15349
rect 21464 -15381 21496 -15349
rect 21496 -15381 21539 -15349
rect 21421 -15424 21539 -15381
rect 21581 -15349 21699 -15306
rect 21581 -15381 21624 -15349
rect 21624 -15381 21656 -15349
rect 21656 -15381 21699 -15349
rect 21581 -15424 21699 -15381
rect 21741 -15349 21859 -15306
rect 21741 -15381 21784 -15349
rect 21784 -15381 21816 -15349
rect 21816 -15381 21859 -15349
rect 21741 -15424 21859 -15381
rect 21901 -15349 22019 -15306
rect 21901 -15381 21944 -15349
rect 21944 -15381 21976 -15349
rect 21976 -15381 22019 -15349
rect 21901 -15424 22019 -15381
rect 22061 -15349 22179 -15306
rect 22061 -15381 22104 -15349
rect 22104 -15381 22136 -15349
rect 22136 -15381 22179 -15349
rect 22061 -15424 22179 -15381
rect 22221 -15349 22339 -15306
rect 22221 -15381 22264 -15349
rect 22264 -15381 22296 -15349
rect 22296 -15381 22339 -15349
rect 22221 -15424 22339 -15381
rect 22381 -15349 22499 -15306
rect 22381 -15381 22424 -15349
rect 22424 -15381 22456 -15349
rect 22456 -15381 22499 -15349
rect 22381 -15424 22499 -15381
rect 22541 -15349 22659 -15306
rect 22541 -15381 22584 -15349
rect 22584 -15381 22616 -15349
rect 22616 -15381 22659 -15349
rect 22541 -15424 22659 -15381
rect 22701 -15349 22819 -15306
rect 22701 -15381 22744 -15349
rect 22744 -15381 22776 -15349
rect 22776 -15381 22819 -15349
rect 22701 -15424 22819 -15381
rect 22861 -15349 22979 -15306
rect 22861 -15381 22904 -15349
rect 22904 -15381 22936 -15349
rect 22936 -15381 22979 -15349
rect 22861 -15424 22979 -15381
rect 23021 -15349 23139 -15306
rect 23021 -15381 23064 -15349
rect 23064 -15381 23096 -15349
rect 23096 -15381 23139 -15349
rect 23021 -15424 23139 -15381
rect 23181 -15349 23299 -15306
rect 23181 -15381 23224 -15349
rect 23224 -15381 23256 -15349
rect 23256 -15381 23299 -15349
rect 23181 -15424 23299 -15381
rect 23341 -15349 23459 -15306
rect 23341 -15381 23384 -15349
rect 23384 -15381 23416 -15349
rect 23416 -15381 23459 -15349
rect 23341 -15424 23459 -15381
rect 23501 -15349 23619 -15306
rect 23501 -15381 23544 -15349
rect 23544 -15381 23576 -15349
rect 23576 -15381 23619 -15349
rect 23501 -15424 23619 -15381
rect 23661 -15349 23779 -15306
rect 23661 -15381 23704 -15349
rect 23704 -15381 23736 -15349
rect 23736 -15381 23779 -15349
rect 23661 -15424 23779 -15381
rect 23821 -15349 23939 -15306
rect 23821 -15381 23864 -15349
rect 23864 -15381 23896 -15349
rect 23896 -15381 23939 -15349
rect 23821 -15424 23939 -15381
rect 23981 -15349 24099 -15306
rect 23981 -15381 24024 -15349
rect 24024 -15381 24056 -15349
rect 24056 -15381 24099 -15349
rect 23981 -15424 24099 -15381
rect 24141 -15349 24259 -15306
rect 24141 -15381 24184 -15349
rect 24184 -15381 24216 -15349
rect 24216 -15381 24259 -15349
rect 24141 -15424 24259 -15381
rect 24301 -15349 24419 -15306
rect 24301 -15381 24344 -15349
rect 24344 -15381 24376 -15349
rect 24376 -15381 24419 -15349
rect 24301 -15424 24419 -15381
rect 24461 -15349 24579 -15306
rect 24461 -15381 24504 -15349
rect 24504 -15381 24536 -15349
rect 24536 -15381 24579 -15349
rect 24461 -15424 24579 -15381
rect 24621 -15349 24739 -15306
rect 24809 -15319 24927 -15276
rect 24621 -15381 24664 -15349
rect 24664 -15381 24696 -15349
rect 24696 -15381 24739 -15349
rect 24621 -15424 24739 -15381
<< metal5 >>
rect 3000 -5578 7000 -5500
rect 3000 -5681 3261 -5578
rect 3000 -5799 3076 -5681
rect 3194 -5696 3261 -5681
rect 3379 -5696 3421 -5578
rect 3539 -5696 3581 -5578
rect 3699 -5696 3741 -5578
rect 3859 -5696 3901 -5578
rect 4019 -5696 4061 -5578
rect 4179 -5696 4221 -5578
rect 4339 -5696 4381 -5578
rect 4499 -5696 4541 -5578
rect 4659 -5696 4701 -5578
rect 4819 -5696 4861 -5578
rect 4979 -5696 5021 -5578
rect 5139 -5696 5181 -5578
rect 5299 -5696 5341 -5578
rect 5459 -5696 5501 -5578
rect 5619 -5696 5661 -5578
rect 5779 -5696 5821 -5578
rect 5939 -5696 5981 -5578
rect 6099 -5696 6141 -5578
rect 6259 -5696 6301 -5578
rect 6419 -5696 6461 -5578
rect 6579 -5696 6621 -5578
rect 6739 -5681 7000 -5578
rect 6739 -5696 6809 -5681
rect 3194 -5799 6809 -5696
rect 6927 -5799 7000 -5681
rect 3000 -5841 7000 -5799
rect 3000 -5959 3076 -5841
rect 3194 -5959 6809 -5841
rect 6927 -5959 7000 -5841
rect 3000 -6001 7000 -5959
rect 3000 -6119 3076 -6001
rect 3194 -6119 6809 -6001
rect 6927 -6119 7000 -6001
rect 3000 -6161 7000 -6119
rect 3000 -6279 3076 -6161
rect 3194 -6279 6809 -6161
rect 6927 -6279 7000 -6161
rect 3000 -6321 7000 -6279
rect 3000 -6439 3076 -6321
rect 3194 -6439 6809 -6321
rect 6927 -6439 7000 -6321
rect 3000 -6481 7000 -6439
rect 3000 -6599 3076 -6481
rect 3194 -6599 6809 -6481
rect 6927 -6599 7000 -6481
rect 3000 -6641 7000 -6599
rect 3000 -6759 3076 -6641
rect 3194 -6759 6809 -6641
rect 6927 -6759 7000 -6641
rect 3000 -6801 7000 -6759
rect 3000 -6919 3076 -6801
rect 3194 -6919 6809 -6801
rect 6927 -6919 7000 -6801
rect 3000 -6961 7000 -6919
rect 3000 -7079 3076 -6961
rect 3194 -7079 6809 -6961
rect 6927 -7079 7000 -6961
rect 3000 -7121 7000 -7079
rect 3000 -7239 3076 -7121
rect 3194 -7239 6809 -7121
rect 6927 -7239 7000 -7121
rect 3000 -7281 7000 -7239
rect 3000 -7399 3076 -7281
rect 3194 -7399 6809 -7281
rect 6927 -7399 7000 -7281
rect 3000 -7441 7000 -7399
rect 3000 -7559 3076 -7441
rect 3194 -7559 6809 -7441
rect 6927 -7559 7000 -7441
rect 3000 -7601 7000 -7559
rect 3000 -7719 3076 -7601
rect 3194 -7719 6809 -7601
rect 6927 -7719 7000 -7601
rect 3000 -7761 7000 -7719
rect 3000 -7879 3076 -7761
rect 3194 -7879 6809 -7761
rect 6927 -7879 7000 -7761
rect 3000 -7921 7000 -7879
rect 3000 -8039 3076 -7921
rect 3194 -8039 6809 -7921
rect 6927 -8039 7000 -7921
rect 3000 -8081 7000 -8039
rect 3000 -8199 3076 -8081
rect 3194 -8199 6809 -8081
rect 6927 -8199 7000 -8081
rect 3000 -8241 7000 -8199
rect 3000 -8359 3076 -8241
rect 3194 -8359 6809 -8241
rect 6927 -8359 7000 -8241
rect 3000 -8401 7000 -8359
rect 3000 -8519 3076 -8401
rect 3194 -8519 6809 -8401
rect 6927 -8519 7000 -8401
rect 3000 -8561 7000 -8519
rect 3000 -8679 3076 -8561
rect 3194 -8679 6809 -8561
rect 6927 -8679 7000 -8561
rect 3000 -8721 7000 -8679
rect 3000 -8839 3076 -8721
rect 3194 -8839 6809 -8721
rect 6927 -8839 7000 -8721
rect 3000 -8881 7000 -8839
rect 3000 -8999 3076 -8881
rect 3194 -8999 6809 -8881
rect 6927 -8999 7000 -8881
rect 3000 -9041 7000 -8999
rect 3000 -9159 3076 -9041
rect 3194 -9159 6809 -9041
rect 6927 -9159 7000 -9041
rect 3000 -9201 7000 -9159
rect 3000 -9319 3076 -9201
rect 3194 -9306 6809 -9201
rect 3194 -9319 3261 -9306
rect 3000 -9424 3261 -9319
rect 3379 -9424 3421 -9306
rect 3539 -9424 3581 -9306
rect 3699 -9424 3741 -9306
rect 3859 -9424 3901 -9306
rect 4019 -9424 4061 -9306
rect 4179 -9424 4221 -9306
rect 4339 -9424 4381 -9306
rect 4499 -9424 4541 -9306
rect 4659 -9424 4701 -9306
rect 4819 -9424 4861 -9306
rect 4979 -9424 5021 -9306
rect 5139 -9424 5181 -9306
rect 5299 -9424 5341 -9306
rect 5459 -9424 5501 -9306
rect 5619 -9424 5661 -9306
rect 5779 -9424 5821 -9306
rect 5939 -9424 5981 -9306
rect 6099 -9424 6141 -9306
rect 6259 -9424 6301 -9306
rect 6419 -9424 6461 -9306
rect 6579 -9424 6621 -9306
rect 6739 -9319 6809 -9306
rect 6927 -9319 7000 -9201
rect 6739 -9424 7000 -9319
rect 3000 -9500 7000 -9424
rect 9000 -5578 13000 -5500
rect 9000 -5681 9261 -5578
rect 9000 -5799 9076 -5681
rect 9194 -5696 9261 -5681
rect 9379 -5696 9421 -5578
rect 9539 -5696 9581 -5578
rect 9699 -5696 9741 -5578
rect 9859 -5696 9901 -5578
rect 10019 -5696 10061 -5578
rect 10179 -5696 10221 -5578
rect 10339 -5696 10381 -5578
rect 10499 -5696 10541 -5578
rect 10659 -5696 10701 -5578
rect 10819 -5696 10861 -5578
rect 10979 -5696 11021 -5578
rect 11139 -5696 11181 -5578
rect 11299 -5696 11341 -5578
rect 11459 -5696 11501 -5578
rect 11619 -5696 11661 -5578
rect 11779 -5696 11821 -5578
rect 11939 -5696 11981 -5578
rect 12099 -5696 12141 -5578
rect 12259 -5696 12301 -5578
rect 12419 -5696 12461 -5578
rect 12579 -5696 12621 -5578
rect 12739 -5681 13000 -5578
rect 12739 -5696 12809 -5681
rect 9194 -5799 12809 -5696
rect 12927 -5799 13000 -5681
rect 9000 -5841 13000 -5799
rect 9000 -5959 9076 -5841
rect 9194 -5959 12809 -5841
rect 12927 -5959 13000 -5841
rect 9000 -6001 13000 -5959
rect 9000 -6119 9076 -6001
rect 9194 -6119 12809 -6001
rect 12927 -6119 13000 -6001
rect 9000 -6161 13000 -6119
rect 9000 -6279 9076 -6161
rect 9194 -6279 12809 -6161
rect 12927 -6279 13000 -6161
rect 9000 -6321 13000 -6279
rect 9000 -6439 9076 -6321
rect 9194 -6439 12809 -6321
rect 12927 -6439 13000 -6321
rect 9000 -6481 13000 -6439
rect 9000 -6599 9076 -6481
rect 9194 -6599 12809 -6481
rect 12927 -6599 13000 -6481
rect 9000 -6641 13000 -6599
rect 9000 -6759 9076 -6641
rect 9194 -6759 12809 -6641
rect 12927 -6759 13000 -6641
rect 9000 -6801 13000 -6759
rect 9000 -6919 9076 -6801
rect 9194 -6919 12809 -6801
rect 12927 -6919 13000 -6801
rect 9000 -6961 13000 -6919
rect 9000 -7079 9076 -6961
rect 9194 -7079 12809 -6961
rect 12927 -7079 13000 -6961
rect 9000 -7121 13000 -7079
rect 9000 -7239 9076 -7121
rect 9194 -7239 12809 -7121
rect 12927 -7239 13000 -7121
rect 9000 -7281 13000 -7239
rect 9000 -7399 9076 -7281
rect 9194 -7399 12809 -7281
rect 12927 -7399 13000 -7281
rect 9000 -7441 13000 -7399
rect 9000 -7559 9076 -7441
rect 9194 -7559 12809 -7441
rect 12927 -7559 13000 -7441
rect 9000 -7601 13000 -7559
rect 9000 -7719 9076 -7601
rect 9194 -7719 12809 -7601
rect 12927 -7719 13000 -7601
rect 9000 -7761 13000 -7719
rect 9000 -7879 9076 -7761
rect 9194 -7879 12809 -7761
rect 12927 -7879 13000 -7761
rect 9000 -7921 13000 -7879
rect 9000 -8039 9076 -7921
rect 9194 -8039 12809 -7921
rect 12927 -8039 13000 -7921
rect 9000 -8081 13000 -8039
rect 9000 -8199 9076 -8081
rect 9194 -8199 12809 -8081
rect 12927 -8199 13000 -8081
rect 9000 -8241 13000 -8199
rect 9000 -8359 9076 -8241
rect 9194 -8359 12809 -8241
rect 12927 -8359 13000 -8241
rect 9000 -8401 13000 -8359
rect 9000 -8519 9076 -8401
rect 9194 -8519 12809 -8401
rect 12927 -8519 13000 -8401
rect 9000 -8561 13000 -8519
rect 9000 -8679 9076 -8561
rect 9194 -8679 12809 -8561
rect 12927 -8679 13000 -8561
rect 9000 -8721 13000 -8679
rect 9000 -8839 9076 -8721
rect 9194 -8839 12809 -8721
rect 12927 -8839 13000 -8721
rect 9000 -8881 13000 -8839
rect 9000 -8999 9076 -8881
rect 9194 -8999 12809 -8881
rect 12927 -8999 13000 -8881
rect 9000 -9041 13000 -8999
rect 9000 -9159 9076 -9041
rect 9194 -9159 12809 -9041
rect 12927 -9159 13000 -9041
rect 9000 -9201 13000 -9159
rect 9000 -9319 9076 -9201
rect 9194 -9306 12809 -9201
rect 9194 -9319 9261 -9306
rect 9000 -9424 9261 -9319
rect 9379 -9424 9421 -9306
rect 9539 -9424 9581 -9306
rect 9699 -9424 9741 -9306
rect 9859 -9424 9901 -9306
rect 10019 -9424 10061 -9306
rect 10179 -9424 10221 -9306
rect 10339 -9424 10381 -9306
rect 10499 -9424 10541 -9306
rect 10659 -9424 10701 -9306
rect 10819 -9424 10861 -9306
rect 10979 -9424 11021 -9306
rect 11139 -9424 11181 -9306
rect 11299 -9424 11341 -9306
rect 11459 -9424 11501 -9306
rect 11619 -9424 11661 -9306
rect 11779 -9424 11821 -9306
rect 11939 -9424 11981 -9306
rect 12099 -9424 12141 -9306
rect 12259 -9424 12301 -9306
rect 12419 -9424 12461 -9306
rect 12579 -9424 12621 -9306
rect 12739 -9319 12809 -9306
rect 12927 -9319 13000 -9201
rect 12739 -9424 13000 -9319
rect 9000 -9500 13000 -9424
rect 15000 -5578 19000 -5500
rect 15000 -5681 15261 -5578
rect 15000 -5799 15076 -5681
rect 15194 -5696 15261 -5681
rect 15379 -5696 15421 -5578
rect 15539 -5696 15581 -5578
rect 15699 -5696 15741 -5578
rect 15859 -5696 15901 -5578
rect 16019 -5696 16061 -5578
rect 16179 -5696 16221 -5578
rect 16339 -5696 16381 -5578
rect 16499 -5696 16541 -5578
rect 16659 -5696 16701 -5578
rect 16819 -5696 16861 -5578
rect 16979 -5696 17021 -5578
rect 17139 -5696 17181 -5578
rect 17299 -5696 17341 -5578
rect 17459 -5696 17501 -5578
rect 17619 -5696 17661 -5578
rect 17779 -5696 17821 -5578
rect 17939 -5696 17981 -5578
rect 18099 -5696 18141 -5578
rect 18259 -5696 18301 -5578
rect 18419 -5696 18461 -5578
rect 18579 -5696 18621 -5578
rect 18739 -5681 19000 -5578
rect 18739 -5696 18809 -5681
rect 15194 -5799 18809 -5696
rect 18927 -5799 19000 -5681
rect 15000 -5841 19000 -5799
rect 15000 -5959 15076 -5841
rect 15194 -5959 18809 -5841
rect 18927 -5959 19000 -5841
rect 15000 -6001 19000 -5959
rect 15000 -6119 15076 -6001
rect 15194 -6119 18809 -6001
rect 18927 -6119 19000 -6001
rect 15000 -6161 19000 -6119
rect 15000 -6279 15076 -6161
rect 15194 -6279 18809 -6161
rect 18927 -6279 19000 -6161
rect 15000 -6321 19000 -6279
rect 15000 -6439 15076 -6321
rect 15194 -6439 18809 -6321
rect 18927 -6439 19000 -6321
rect 15000 -6481 19000 -6439
rect 15000 -6599 15076 -6481
rect 15194 -6599 18809 -6481
rect 18927 -6599 19000 -6481
rect 15000 -6641 19000 -6599
rect 15000 -6759 15076 -6641
rect 15194 -6759 18809 -6641
rect 18927 -6759 19000 -6641
rect 15000 -6801 19000 -6759
rect 15000 -6919 15076 -6801
rect 15194 -6919 18809 -6801
rect 18927 -6919 19000 -6801
rect 15000 -6961 19000 -6919
rect 15000 -7079 15076 -6961
rect 15194 -7079 18809 -6961
rect 18927 -7079 19000 -6961
rect 15000 -7121 19000 -7079
rect 15000 -7239 15076 -7121
rect 15194 -7239 18809 -7121
rect 18927 -7239 19000 -7121
rect 15000 -7281 19000 -7239
rect 15000 -7399 15076 -7281
rect 15194 -7399 18809 -7281
rect 18927 -7399 19000 -7281
rect 15000 -7441 19000 -7399
rect 15000 -7559 15076 -7441
rect 15194 -7559 18809 -7441
rect 18927 -7559 19000 -7441
rect 15000 -7601 19000 -7559
rect 15000 -7719 15076 -7601
rect 15194 -7719 18809 -7601
rect 18927 -7719 19000 -7601
rect 15000 -7761 19000 -7719
rect 15000 -7879 15076 -7761
rect 15194 -7879 18809 -7761
rect 18927 -7879 19000 -7761
rect 15000 -7921 19000 -7879
rect 15000 -8039 15076 -7921
rect 15194 -8039 18809 -7921
rect 18927 -8039 19000 -7921
rect 15000 -8081 19000 -8039
rect 15000 -8199 15076 -8081
rect 15194 -8199 18809 -8081
rect 18927 -8199 19000 -8081
rect 15000 -8241 19000 -8199
rect 15000 -8359 15076 -8241
rect 15194 -8359 18809 -8241
rect 18927 -8359 19000 -8241
rect 15000 -8401 19000 -8359
rect 15000 -8519 15076 -8401
rect 15194 -8519 18809 -8401
rect 18927 -8519 19000 -8401
rect 15000 -8561 19000 -8519
rect 15000 -8679 15076 -8561
rect 15194 -8679 18809 -8561
rect 18927 -8679 19000 -8561
rect 15000 -8721 19000 -8679
rect 15000 -8839 15076 -8721
rect 15194 -8839 18809 -8721
rect 18927 -8839 19000 -8721
rect 15000 -8881 19000 -8839
rect 15000 -8999 15076 -8881
rect 15194 -8999 18809 -8881
rect 18927 -8999 19000 -8881
rect 15000 -9041 19000 -8999
rect 15000 -9159 15076 -9041
rect 15194 -9159 18809 -9041
rect 18927 -9159 19000 -9041
rect 15000 -9201 19000 -9159
rect 15000 -9319 15076 -9201
rect 15194 -9306 18809 -9201
rect 15194 -9319 15261 -9306
rect 15000 -9424 15261 -9319
rect 15379 -9424 15421 -9306
rect 15539 -9424 15581 -9306
rect 15699 -9424 15741 -9306
rect 15859 -9424 15901 -9306
rect 16019 -9424 16061 -9306
rect 16179 -9424 16221 -9306
rect 16339 -9424 16381 -9306
rect 16499 -9424 16541 -9306
rect 16659 -9424 16701 -9306
rect 16819 -9424 16861 -9306
rect 16979 -9424 17021 -9306
rect 17139 -9424 17181 -9306
rect 17299 -9424 17341 -9306
rect 17459 -9424 17501 -9306
rect 17619 -9424 17661 -9306
rect 17779 -9424 17821 -9306
rect 17939 -9424 17981 -9306
rect 18099 -9424 18141 -9306
rect 18259 -9424 18301 -9306
rect 18419 -9424 18461 -9306
rect 18579 -9424 18621 -9306
rect 18739 -9319 18809 -9306
rect 18927 -9319 19000 -9201
rect 18739 -9424 19000 -9319
rect 15000 -9500 19000 -9424
rect 21000 -5578 25000 -5500
rect 21000 -5681 21261 -5578
rect 21000 -5799 21076 -5681
rect 21194 -5696 21261 -5681
rect 21379 -5696 21421 -5578
rect 21539 -5696 21581 -5578
rect 21699 -5696 21741 -5578
rect 21859 -5696 21901 -5578
rect 22019 -5696 22061 -5578
rect 22179 -5696 22221 -5578
rect 22339 -5696 22381 -5578
rect 22499 -5696 22541 -5578
rect 22659 -5696 22701 -5578
rect 22819 -5696 22861 -5578
rect 22979 -5696 23021 -5578
rect 23139 -5696 23181 -5578
rect 23299 -5696 23341 -5578
rect 23459 -5696 23501 -5578
rect 23619 -5696 23661 -5578
rect 23779 -5696 23821 -5578
rect 23939 -5696 23981 -5578
rect 24099 -5696 24141 -5578
rect 24259 -5696 24301 -5578
rect 24419 -5696 24461 -5578
rect 24579 -5696 24621 -5578
rect 24739 -5681 25000 -5578
rect 24739 -5696 24809 -5681
rect 21194 -5799 24809 -5696
rect 24927 -5799 25000 -5681
rect 21000 -5841 25000 -5799
rect 21000 -5959 21076 -5841
rect 21194 -5959 24809 -5841
rect 24927 -5959 25000 -5841
rect 21000 -6001 25000 -5959
rect 21000 -6119 21076 -6001
rect 21194 -6119 24809 -6001
rect 24927 -6119 25000 -6001
rect 21000 -6161 25000 -6119
rect 21000 -6279 21076 -6161
rect 21194 -6279 24809 -6161
rect 24927 -6279 25000 -6161
rect 21000 -6321 25000 -6279
rect 21000 -6439 21076 -6321
rect 21194 -6439 24809 -6321
rect 24927 -6439 25000 -6321
rect 21000 -6481 25000 -6439
rect 21000 -6599 21076 -6481
rect 21194 -6599 24809 -6481
rect 24927 -6599 25000 -6481
rect 21000 -6641 25000 -6599
rect 21000 -6759 21076 -6641
rect 21194 -6759 24809 -6641
rect 24927 -6759 25000 -6641
rect 21000 -6801 25000 -6759
rect 21000 -6919 21076 -6801
rect 21194 -6919 24809 -6801
rect 24927 -6919 25000 -6801
rect 21000 -6961 25000 -6919
rect 21000 -7079 21076 -6961
rect 21194 -7079 24809 -6961
rect 24927 -7079 25000 -6961
rect 21000 -7121 25000 -7079
rect 21000 -7239 21076 -7121
rect 21194 -7239 24809 -7121
rect 24927 -7239 25000 -7121
rect 21000 -7281 25000 -7239
rect 21000 -7399 21076 -7281
rect 21194 -7399 24809 -7281
rect 24927 -7399 25000 -7281
rect 21000 -7441 25000 -7399
rect 21000 -7559 21076 -7441
rect 21194 -7559 24809 -7441
rect 24927 -7559 25000 -7441
rect 21000 -7601 25000 -7559
rect 21000 -7719 21076 -7601
rect 21194 -7719 24809 -7601
rect 24927 -7719 25000 -7601
rect 21000 -7761 25000 -7719
rect 21000 -7879 21076 -7761
rect 21194 -7879 24809 -7761
rect 24927 -7879 25000 -7761
rect 21000 -7921 25000 -7879
rect 21000 -8039 21076 -7921
rect 21194 -8039 24809 -7921
rect 24927 -8039 25000 -7921
rect 21000 -8081 25000 -8039
rect 21000 -8199 21076 -8081
rect 21194 -8199 24809 -8081
rect 24927 -8199 25000 -8081
rect 21000 -8241 25000 -8199
rect 21000 -8359 21076 -8241
rect 21194 -8359 24809 -8241
rect 24927 -8359 25000 -8241
rect 21000 -8401 25000 -8359
rect 21000 -8519 21076 -8401
rect 21194 -8519 24809 -8401
rect 24927 -8519 25000 -8401
rect 21000 -8561 25000 -8519
rect 21000 -8679 21076 -8561
rect 21194 -8679 24809 -8561
rect 24927 -8679 25000 -8561
rect 21000 -8721 25000 -8679
rect 21000 -8839 21076 -8721
rect 21194 -8839 24809 -8721
rect 24927 -8839 25000 -8721
rect 21000 -8881 25000 -8839
rect 21000 -8999 21076 -8881
rect 21194 -8999 24809 -8881
rect 24927 -8999 25000 -8881
rect 21000 -9041 25000 -8999
rect 21000 -9159 21076 -9041
rect 21194 -9159 24809 -9041
rect 24927 -9159 25000 -9041
rect 21000 -9201 25000 -9159
rect 21000 -9319 21076 -9201
rect 21194 -9306 24809 -9201
rect 21194 -9319 21261 -9306
rect 21000 -9424 21261 -9319
rect 21379 -9424 21421 -9306
rect 21539 -9424 21581 -9306
rect 21699 -9424 21741 -9306
rect 21859 -9424 21901 -9306
rect 22019 -9424 22061 -9306
rect 22179 -9424 22221 -9306
rect 22339 -9424 22381 -9306
rect 22499 -9424 22541 -9306
rect 22659 -9424 22701 -9306
rect 22819 -9424 22861 -9306
rect 22979 -9424 23021 -9306
rect 23139 -9424 23181 -9306
rect 23299 -9424 23341 -9306
rect 23459 -9424 23501 -9306
rect 23619 -9424 23661 -9306
rect 23779 -9424 23821 -9306
rect 23939 -9424 23981 -9306
rect 24099 -9424 24141 -9306
rect 24259 -9424 24301 -9306
rect 24419 -9424 24461 -9306
rect 24579 -9424 24621 -9306
rect 24739 -9319 24809 -9306
rect 24927 -9319 25000 -9201
rect 24739 -9424 25000 -9319
rect 21000 -9500 25000 -9424
rect 3000 -11578 7000 -11500
rect 3000 -11681 3261 -11578
rect 3000 -11799 3076 -11681
rect 3194 -11696 3261 -11681
rect 3379 -11696 3421 -11578
rect 3539 -11696 3581 -11578
rect 3699 -11696 3741 -11578
rect 3859 -11696 3901 -11578
rect 4019 -11696 4061 -11578
rect 4179 -11696 4221 -11578
rect 4339 -11696 4381 -11578
rect 4499 -11696 4541 -11578
rect 4659 -11696 4701 -11578
rect 4819 -11696 4861 -11578
rect 4979 -11696 5021 -11578
rect 5139 -11696 5181 -11578
rect 5299 -11696 5341 -11578
rect 5459 -11696 5501 -11578
rect 5619 -11696 5661 -11578
rect 5779 -11696 5821 -11578
rect 5939 -11696 5981 -11578
rect 6099 -11696 6141 -11578
rect 6259 -11696 6301 -11578
rect 6419 -11696 6461 -11578
rect 6579 -11696 6621 -11578
rect 6739 -11681 7000 -11578
rect 6739 -11696 6809 -11681
rect 3194 -11799 6809 -11696
rect 6927 -11799 7000 -11681
rect 3000 -11841 7000 -11799
rect 3000 -11959 3076 -11841
rect 3194 -11959 6809 -11841
rect 6927 -11959 7000 -11841
rect 3000 -12001 7000 -11959
rect 3000 -12119 3076 -12001
rect 3194 -12119 6809 -12001
rect 6927 -12119 7000 -12001
rect 3000 -12161 7000 -12119
rect 3000 -12279 3076 -12161
rect 3194 -12279 6809 -12161
rect 6927 -12279 7000 -12161
rect 3000 -12321 7000 -12279
rect 3000 -12439 3076 -12321
rect 3194 -12439 6809 -12321
rect 6927 -12439 7000 -12321
rect 3000 -12481 7000 -12439
rect 3000 -12599 3076 -12481
rect 3194 -12599 6809 -12481
rect 6927 -12599 7000 -12481
rect 3000 -12641 7000 -12599
rect 3000 -12759 3076 -12641
rect 3194 -12759 6809 -12641
rect 6927 -12759 7000 -12641
rect 3000 -12801 7000 -12759
rect 3000 -12919 3076 -12801
rect 3194 -12919 6809 -12801
rect 6927 -12919 7000 -12801
rect 3000 -12961 7000 -12919
rect 3000 -13079 3076 -12961
rect 3194 -13079 6809 -12961
rect 6927 -13079 7000 -12961
rect 3000 -13121 7000 -13079
rect 3000 -13239 3076 -13121
rect 3194 -13239 6809 -13121
rect 6927 -13239 7000 -13121
rect 3000 -13281 7000 -13239
rect 3000 -13399 3076 -13281
rect 3194 -13399 6809 -13281
rect 6927 -13399 7000 -13281
rect 3000 -13441 7000 -13399
rect 3000 -13559 3076 -13441
rect 3194 -13559 6809 -13441
rect 6927 -13559 7000 -13441
rect 3000 -13601 7000 -13559
rect 3000 -13719 3076 -13601
rect 3194 -13719 6809 -13601
rect 6927 -13719 7000 -13601
rect 3000 -13761 7000 -13719
rect 3000 -13879 3076 -13761
rect 3194 -13879 6809 -13761
rect 6927 -13879 7000 -13761
rect 3000 -13921 7000 -13879
rect 3000 -14039 3076 -13921
rect 3194 -14039 6809 -13921
rect 6927 -14039 7000 -13921
rect 3000 -14081 7000 -14039
rect 3000 -14199 3076 -14081
rect 3194 -14199 6809 -14081
rect 6927 -14199 7000 -14081
rect 3000 -14241 7000 -14199
rect 3000 -14359 3076 -14241
rect 3194 -14359 6809 -14241
rect 6927 -14359 7000 -14241
rect 3000 -14401 7000 -14359
rect 3000 -14519 3076 -14401
rect 3194 -14519 6809 -14401
rect 6927 -14519 7000 -14401
rect 3000 -14561 7000 -14519
rect 3000 -14679 3076 -14561
rect 3194 -14679 6809 -14561
rect 6927 -14679 7000 -14561
rect 3000 -14721 7000 -14679
rect 3000 -14839 3076 -14721
rect 3194 -14839 6809 -14721
rect 6927 -14839 7000 -14721
rect 3000 -14881 7000 -14839
rect 3000 -14999 3076 -14881
rect 3194 -14999 6809 -14881
rect 6927 -14999 7000 -14881
rect 3000 -15041 7000 -14999
rect 3000 -15159 3076 -15041
rect 3194 -15159 6809 -15041
rect 6927 -15159 7000 -15041
rect 3000 -15201 7000 -15159
rect 3000 -15319 3076 -15201
rect 3194 -15306 6809 -15201
rect 3194 -15319 3261 -15306
rect 3000 -15424 3261 -15319
rect 3379 -15424 3421 -15306
rect 3539 -15424 3581 -15306
rect 3699 -15424 3741 -15306
rect 3859 -15424 3901 -15306
rect 4019 -15424 4061 -15306
rect 4179 -15424 4221 -15306
rect 4339 -15424 4381 -15306
rect 4499 -15424 4541 -15306
rect 4659 -15424 4701 -15306
rect 4819 -15424 4861 -15306
rect 4979 -15424 5021 -15306
rect 5139 -15424 5181 -15306
rect 5299 -15424 5341 -15306
rect 5459 -15424 5501 -15306
rect 5619 -15424 5661 -15306
rect 5779 -15424 5821 -15306
rect 5939 -15424 5981 -15306
rect 6099 -15424 6141 -15306
rect 6259 -15424 6301 -15306
rect 6419 -15424 6461 -15306
rect 6579 -15424 6621 -15306
rect 6739 -15319 6809 -15306
rect 6927 -15319 7000 -15201
rect 6739 -15424 7000 -15319
rect 3000 -15500 7000 -15424
rect 9000 -11578 13000 -11500
rect 9000 -11681 9261 -11578
rect 9000 -11799 9076 -11681
rect 9194 -11696 9261 -11681
rect 9379 -11696 9421 -11578
rect 9539 -11696 9581 -11578
rect 9699 -11696 9741 -11578
rect 9859 -11696 9901 -11578
rect 10019 -11696 10061 -11578
rect 10179 -11696 10221 -11578
rect 10339 -11696 10381 -11578
rect 10499 -11696 10541 -11578
rect 10659 -11696 10701 -11578
rect 10819 -11696 10861 -11578
rect 10979 -11696 11021 -11578
rect 11139 -11696 11181 -11578
rect 11299 -11696 11341 -11578
rect 11459 -11696 11501 -11578
rect 11619 -11696 11661 -11578
rect 11779 -11696 11821 -11578
rect 11939 -11696 11981 -11578
rect 12099 -11696 12141 -11578
rect 12259 -11696 12301 -11578
rect 12419 -11696 12461 -11578
rect 12579 -11696 12621 -11578
rect 12739 -11681 13000 -11578
rect 12739 -11696 12809 -11681
rect 9194 -11799 12809 -11696
rect 12927 -11799 13000 -11681
rect 9000 -11841 13000 -11799
rect 9000 -11959 9076 -11841
rect 9194 -11959 12809 -11841
rect 12927 -11959 13000 -11841
rect 9000 -12001 13000 -11959
rect 9000 -12119 9076 -12001
rect 9194 -12119 12809 -12001
rect 12927 -12119 13000 -12001
rect 9000 -12161 13000 -12119
rect 9000 -12279 9076 -12161
rect 9194 -12279 12809 -12161
rect 12927 -12279 13000 -12161
rect 9000 -12321 13000 -12279
rect 9000 -12439 9076 -12321
rect 9194 -12439 12809 -12321
rect 12927 -12439 13000 -12321
rect 9000 -12481 13000 -12439
rect 9000 -12599 9076 -12481
rect 9194 -12599 12809 -12481
rect 12927 -12599 13000 -12481
rect 9000 -12641 13000 -12599
rect 9000 -12759 9076 -12641
rect 9194 -12759 12809 -12641
rect 12927 -12759 13000 -12641
rect 9000 -12801 13000 -12759
rect 9000 -12919 9076 -12801
rect 9194 -12919 12809 -12801
rect 12927 -12919 13000 -12801
rect 9000 -12961 13000 -12919
rect 9000 -13079 9076 -12961
rect 9194 -13079 12809 -12961
rect 12927 -13079 13000 -12961
rect 9000 -13121 13000 -13079
rect 9000 -13239 9076 -13121
rect 9194 -13239 12809 -13121
rect 12927 -13239 13000 -13121
rect 9000 -13281 13000 -13239
rect 9000 -13399 9076 -13281
rect 9194 -13399 12809 -13281
rect 12927 -13399 13000 -13281
rect 9000 -13441 13000 -13399
rect 9000 -13559 9076 -13441
rect 9194 -13559 12809 -13441
rect 12927 -13559 13000 -13441
rect 9000 -13601 13000 -13559
rect 9000 -13719 9076 -13601
rect 9194 -13719 12809 -13601
rect 12927 -13719 13000 -13601
rect 9000 -13761 13000 -13719
rect 9000 -13879 9076 -13761
rect 9194 -13879 12809 -13761
rect 12927 -13879 13000 -13761
rect 9000 -13921 13000 -13879
rect 9000 -14039 9076 -13921
rect 9194 -14039 12809 -13921
rect 12927 -14039 13000 -13921
rect 9000 -14081 13000 -14039
rect 9000 -14199 9076 -14081
rect 9194 -14199 12809 -14081
rect 12927 -14199 13000 -14081
rect 9000 -14241 13000 -14199
rect 9000 -14359 9076 -14241
rect 9194 -14359 12809 -14241
rect 12927 -14359 13000 -14241
rect 9000 -14401 13000 -14359
rect 9000 -14519 9076 -14401
rect 9194 -14519 12809 -14401
rect 12927 -14519 13000 -14401
rect 9000 -14561 13000 -14519
rect 9000 -14679 9076 -14561
rect 9194 -14679 12809 -14561
rect 12927 -14679 13000 -14561
rect 9000 -14721 13000 -14679
rect 9000 -14839 9076 -14721
rect 9194 -14839 12809 -14721
rect 12927 -14839 13000 -14721
rect 9000 -14881 13000 -14839
rect 9000 -14999 9076 -14881
rect 9194 -14999 12809 -14881
rect 12927 -14999 13000 -14881
rect 9000 -15041 13000 -14999
rect 9000 -15159 9076 -15041
rect 9194 -15159 12809 -15041
rect 12927 -15159 13000 -15041
rect 9000 -15201 13000 -15159
rect 9000 -15319 9076 -15201
rect 9194 -15306 12809 -15201
rect 9194 -15319 9261 -15306
rect 9000 -15424 9261 -15319
rect 9379 -15424 9421 -15306
rect 9539 -15424 9581 -15306
rect 9699 -15424 9741 -15306
rect 9859 -15424 9901 -15306
rect 10019 -15424 10061 -15306
rect 10179 -15424 10221 -15306
rect 10339 -15424 10381 -15306
rect 10499 -15424 10541 -15306
rect 10659 -15424 10701 -15306
rect 10819 -15424 10861 -15306
rect 10979 -15424 11021 -15306
rect 11139 -15424 11181 -15306
rect 11299 -15424 11341 -15306
rect 11459 -15424 11501 -15306
rect 11619 -15424 11661 -15306
rect 11779 -15424 11821 -15306
rect 11939 -15424 11981 -15306
rect 12099 -15424 12141 -15306
rect 12259 -15424 12301 -15306
rect 12419 -15424 12461 -15306
rect 12579 -15424 12621 -15306
rect 12739 -15319 12809 -15306
rect 12927 -15319 13000 -15201
rect 12739 -15424 13000 -15319
rect 9000 -15500 13000 -15424
rect 15000 -11578 19000 -11500
rect 15000 -11681 15261 -11578
rect 15000 -11799 15076 -11681
rect 15194 -11696 15261 -11681
rect 15379 -11696 15421 -11578
rect 15539 -11696 15581 -11578
rect 15699 -11696 15741 -11578
rect 15859 -11696 15901 -11578
rect 16019 -11696 16061 -11578
rect 16179 -11696 16221 -11578
rect 16339 -11696 16381 -11578
rect 16499 -11696 16541 -11578
rect 16659 -11696 16701 -11578
rect 16819 -11696 16861 -11578
rect 16979 -11696 17021 -11578
rect 17139 -11696 17181 -11578
rect 17299 -11696 17341 -11578
rect 17459 -11696 17501 -11578
rect 17619 -11696 17661 -11578
rect 17779 -11696 17821 -11578
rect 17939 -11696 17981 -11578
rect 18099 -11696 18141 -11578
rect 18259 -11696 18301 -11578
rect 18419 -11696 18461 -11578
rect 18579 -11696 18621 -11578
rect 18739 -11681 19000 -11578
rect 18739 -11696 18809 -11681
rect 15194 -11799 18809 -11696
rect 18927 -11799 19000 -11681
rect 15000 -11841 19000 -11799
rect 15000 -11959 15076 -11841
rect 15194 -11959 18809 -11841
rect 18927 -11959 19000 -11841
rect 15000 -12001 19000 -11959
rect 15000 -12119 15076 -12001
rect 15194 -12119 18809 -12001
rect 18927 -12119 19000 -12001
rect 15000 -12161 19000 -12119
rect 15000 -12279 15076 -12161
rect 15194 -12279 18809 -12161
rect 18927 -12279 19000 -12161
rect 15000 -12321 19000 -12279
rect 15000 -12439 15076 -12321
rect 15194 -12439 18809 -12321
rect 18927 -12439 19000 -12321
rect 15000 -12481 19000 -12439
rect 15000 -12599 15076 -12481
rect 15194 -12599 18809 -12481
rect 18927 -12599 19000 -12481
rect 15000 -12641 19000 -12599
rect 15000 -12759 15076 -12641
rect 15194 -12759 18809 -12641
rect 18927 -12759 19000 -12641
rect 15000 -12801 19000 -12759
rect 15000 -12919 15076 -12801
rect 15194 -12919 18809 -12801
rect 18927 -12919 19000 -12801
rect 15000 -12961 19000 -12919
rect 15000 -13079 15076 -12961
rect 15194 -13079 18809 -12961
rect 18927 -13079 19000 -12961
rect 15000 -13121 19000 -13079
rect 15000 -13239 15076 -13121
rect 15194 -13239 18809 -13121
rect 18927 -13239 19000 -13121
rect 15000 -13281 19000 -13239
rect 15000 -13399 15076 -13281
rect 15194 -13399 18809 -13281
rect 18927 -13399 19000 -13281
rect 15000 -13441 19000 -13399
rect 15000 -13559 15076 -13441
rect 15194 -13559 18809 -13441
rect 18927 -13559 19000 -13441
rect 15000 -13601 19000 -13559
rect 15000 -13719 15076 -13601
rect 15194 -13719 18809 -13601
rect 18927 -13719 19000 -13601
rect 15000 -13761 19000 -13719
rect 15000 -13879 15076 -13761
rect 15194 -13879 18809 -13761
rect 18927 -13879 19000 -13761
rect 15000 -13921 19000 -13879
rect 15000 -14039 15076 -13921
rect 15194 -14039 18809 -13921
rect 18927 -14039 19000 -13921
rect 15000 -14081 19000 -14039
rect 15000 -14199 15076 -14081
rect 15194 -14199 18809 -14081
rect 18927 -14199 19000 -14081
rect 15000 -14241 19000 -14199
rect 15000 -14359 15076 -14241
rect 15194 -14359 18809 -14241
rect 18927 -14359 19000 -14241
rect 15000 -14401 19000 -14359
rect 15000 -14519 15076 -14401
rect 15194 -14519 18809 -14401
rect 18927 -14519 19000 -14401
rect 15000 -14561 19000 -14519
rect 15000 -14679 15076 -14561
rect 15194 -14679 18809 -14561
rect 18927 -14679 19000 -14561
rect 15000 -14721 19000 -14679
rect 15000 -14839 15076 -14721
rect 15194 -14839 18809 -14721
rect 18927 -14839 19000 -14721
rect 15000 -14881 19000 -14839
rect 15000 -14999 15076 -14881
rect 15194 -14999 18809 -14881
rect 18927 -14999 19000 -14881
rect 15000 -15041 19000 -14999
rect 15000 -15159 15076 -15041
rect 15194 -15159 18809 -15041
rect 18927 -15159 19000 -15041
rect 15000 -15201 19000 -15159
rect 15000 -15319 15076 -15201
rect 15194 -15306 18809 -15201
rect 15194 -15319 15261 -15306
rect 15000 -15424 15261 -15319
rect 15379 -15424 15421 -15306
rect 15539 -15424 15581 -15306
rect 15699 -15424 15741 -15306
rect 15859 -15424 15901 -15306
rect 16019 -15424 16061 -15306
rect 16179 -15424 16221 -15306
rect 16339 -15424 16381 -15306
rect 16499 -15424 16541 -15306
rect 16659 -15424 16701 -15306
rect 16819 -15424 16861 -15306
rect 16979 -15424 17021 -15306
rect 17139 -15424 17181 -15306
rect 17299 -15424 17341 -15306
rect 17459 -15424 17501 -15306
rect 17619 -15424 17661 -15306
rect 17779 -15424 17821 -15306
rect 17939 -15424 17981 -15306
rect 18099 -15424 18141 -15306
rect 18259 -15424 18301 -15306
rect 18419 -15424 18461 -15306
rect 18579 -15424 18621 -15306
rect 18739 -15319 18809 -15306
rect 18927 -15319 19000 -15201
rect 18739 -15424 19000 -15319
rect 15000 -15500 19000 -15424
rect 21000 -11578 25000 -11500
rect 21000 -11681 21261 -11578
rect 21000 -11799 21076 -11681
rect 21194 -11696 21261 -11681
rect 21379 -11696 21421 -11578
rect 21539 -11696 21581 -11578
rect 21699 -11696 21741 -11578
rect 21859 -11696 21901 -11578
rect 22019 -11696 22061 -11578
rect 22179 -11696 22221 -11578
rect 22339 -11696 22381 -11578
rect 22499 -11696 22541 -11578
rect 22659 -11696 22701 -11578
rect 22819 -11696 22861 -11578
rect 22979 -11696 23021 -11578
rect 23139 -11696 23181 -11578
rect 23299 -11696 23341 -11578
rect 23459 -11696 23501 -11578
rect 23619 -11696 23661 -11578
rect 23779 -11696 23821 -11578
rect 23939 -11696 23981 -11578
rect 24099 -11696 24141 -11578
rect 24259 -11696 24301 -11578
rect 24419 -11696 24461 -11578
rect 24579 -11696 24621 -11578
rect 24739 -11681 25000 -11578
rect 24739 -11696 24809 -11681
rect 21194 -11799 24809 -11696
rect 24927 -11799 25000 -11681
rect 21000 -11841 25000 -11799
rect 21000 -11959 21076 -11841
rect 21194 -11959 24809 -11841
rect 24927 -11959 25000 -11841
rect 21000 -12001 25000 -11959
rect 21000 -12119 21076 -12001
rect 21194 -12119 24809 -12001
rect 24927 -12119 25000 -12001
rect 21000 -12161 25000 -12119
rect 21000 -12279 21076 -12161
rect 21194 -12279 24809 -12161
rect 24927 -12279 25000 -12161
rect 21000 -12321 25000 -12279
rect 21000 -12439 21076 -12321
rect 21194 -12439 24809 -12321
rect 24927 -12439 25000 -12321
rect 21000 -12481 25000 -12439
rect 21000 -12599 21076 -12481
rect 21194 -12599 24809 -12481
rect 24927 -12599 25000 -12481
rect 21000 -12641 25000 -12599
rect 21000 -12759 21076 -12641
rect 21194 -12759 24809 -12641
rect 24927 -12759 25000 -12641
rect 21000 -12801 25000 -12759
rect 21000 -12919 21076 -12801
rect 21194 -12919 24809 -12801
rect 24927 -12919 25000 -12801
rect 21000 -12961 25000 -12919
rect 21000 -13079 21076 -12961
rect 21194 -13079 24809 -12961
rect 24927 -13079 25000 -12961
rect 21000 -13121 25000 -13079
rect 21000 -13239 21076 -13121
rect 21194 -13239 24809 -13121
rect 24927 -13239 25000 -13121
rect 21000 -13281 25000 -13239
rect 21000 -13399 21076 -13281
rect 21194 -13399 24809 -13281
rect 24927 -13399 25000 -13281
rect 21000 -13441 25000 -13399
rect 21000 -13559 21076 -13441
rect 21194 -13559 24809 -13441
rect 24927 -13559 25000 -13441
rect 21000 -13601 25000 -13559
rect 21000 -13719 21076 -13601
rect 21194 -13719 24809 -13601
rect 24927 -13719 25000 -13601
rect 21000 -13761 25000 -13719
rect 21000 -13879 21076 -13761
rect 21194 -13879 24809 -13761
rect 24927 -13879 25000 -13761
rect 21000 -13921 25000 -13879
rect 21000 -14039 21076 -13921
rect 21194 -14039 24809 -13921
rect 24927 -14039 25000 -13921
rect 21000 -14081 25000 -14039
rect 21000 -14199 21076 -14081
rect 21194 -14199 24809 -14081
rect 24927 -14199 25000 -14081
rect 21000 -14241 25000 -14199
rect 21000 -14359 21076 -14241
rect 21194 -14359 24809 -14241
rect 24927 -14359 25000 -14241
rect 21000 -14401 25000 -14359
rect 21000 -14519 21076 -14401
rect 21194 -14519 24809 -14401
rect 24927 -14519 25000 -14401
rect 21000 -14561 25000 -14519
rect 21000 -14679 21076 -14561
rect 21194 -14679 24809 -14561
rect 24927 -14679 25000 -14561
rect 21000 -14721 25000 -14679
rect 21000 -14839 21076 -14721
rect 21194 -14839 24809 -14721
rect 24927 -14839 25000 -14721
rect 21000 -14881 25000 -14839
rect 21000 -14999 21076 -14881
rect 21194 -14999 24809 -14881
rect 24927 -14999 25000 -14881
rect 21000 -15041 25000 -14999
rect 21000 -15159 21076 -15041
rect 21194 -15159 24809 -15041
rect 24927 -15159 25000 -15041
rect 21000 -15201 25000 -15159
rect 21000 -15319 21076 -15201
rect 21194 -15306 24809 -15201
rect 21194 -15319 21261 -15306
rect 21000 -15424 21261 -15319
rect 21379 -15424 21421 -15306
rect 21539 -15424 21581 -15306
rect 21699 -15424 21741 -15306
rect 21859 -15424 21901 -15306
rect 22019 -15424 22061 -15306
rect 22179 -15424 22221 -15306
rect 22339 -15424 22381 -15306
rect 22499 -15424 22541 -15306
rect 22659 -15424 22701 -15306
rect 22819 -15424 22861 -15306
rect 22979 -15424 23021 -15306
rect 23139 -15424 23181 -15306
rect 23299 -15424 23341 -15306
rect 23459 -15424 23501 -15306
rect 23619 -15424 23661 -15306
rect 23779 -15424 23821 -15306
rect 23939 -15424 23981 -15306
rect 24099 -15424 24141 -15306
rect 24259 -15424 24301 -15306
rect 24419 -15424 24461 -15306
rect 24579 -15424 24621 -15306
rect 24739 -15319 24809 -15306
rect 24927 -15319 25000 -15201
rect 24739 -15424 25000 -15319
rect 21000 -15500 25000 -15424
<< fillblock >>
rect 3000 -10000 4200 -9500
rect 9000 -10000 10200 -9500
rect 15000 -10000 16200 -9500
rect 21000 -10000 22200 -9500
rect 3000 -11500 3400 -10900
rect 9000 -11500 9400 -10910
rect 15000 -11500 16600 -11000
rect 21000 -11500 22200 -11000
<< comment >>
rect 900 -9500 1000 -5300
use cmota_gb_rp_gp  cmota_gb_rp_gp_1
timestamp 1671855392
transform 1 0 10100 0 1 -1250
box -3500 -3900 1401 300
use sky130hd_esd  sky130hd_esd_0
timestamp 1671850507
transform 0 -1 8680 -1 0 -5117
box 111 -30 333 290
use sky130hd_esd  sky130hd_esd_1
timestamp 1671850507
transform 1 0 11448 0 1 -3951
box 111 -30 333 290
use sky130hd_esd  sky130hd_esd_2
timestamp 1671850507
transform 1 0 11586 0 1 -3951
box 111 -30 333 290
<< labels >>
rlabel metal5 3600 -8800 6250 -6500 1 VHI
rlabel metal5 9750 -8700 12400 -6400 1 VLO
rlabel metal5 15650 -8700 18300 -6400 1 VIP
rlabel metal5 21650 -8700 24300 -6400 1 VOP
rlabel metal5 21650 -14600 24300 -12300 1 VIN
rlabel metal5 15650 -14650 18300 -12350 1 VREF
rlabel metal5 9700 -14650 12350 -12350 1 SBAR
rlabel metal5 3750 -14700 6400 -12400 1 S
<< end >>
