magic
tech sky130A
timestamp 1672031340
<< metal1 >>
rect -3 0 0 26
rect 26 0 29 26
<< via1 >>
rect 0 0 26 26
<< metal2 >>
rect -3 0 0 26
rect 26 0 29 26
<< end >>
