magic
tech sky130A
magscale 1 2
timestamp 1671378102
<< pwell >>
rect -53 637 369 767
rect -53 584 135 637
rect 189 584 369 637
rect -53 -53 369 584
<< nmos >>
rect 143 157 173 557
<< ndiff >>
rect 85 545 143 557
rect 85 169 97 545
rect 131 169 143 545
rect 85 157 143 169
rect 173 545 231 557
rect 173 169 185 545
rect 219 169 231 545
rect 173 157 231 169
<< ndiffc >>
rect 97 169 131 545
rect 185 169 219 545
<< psubdiff >>
rect -17 697 79 731
rect 237 697 333 731
rect -17 635 17 697
rect 299 635 333 697
rect -17 17 17 79
rect 299 17 333 79
rect -17 -17 79 17
rect 237 -17 333 17
<< psubdiffcont >>
rect 79 697 237 731
rect -17 79 17 635
rect 299 79 333 635
rect 79 -17 237 17
<< poly >>
rect 125 579 191 645
rect 143 557 173 579
rect 143 135 173 157
rect 125 119 191 135
rect 125 85 141 119
rect 175 85 191 119
rect 125 69 191 85
<< polycont >>
rect 141 85 175 119
<< locali >>
rect -51 697 79 731
rect 237 697 333 731
rect -51 635 17 697
rect -51 79 -17 635
rect 299 635 333 697
rect 97 545 131 561
rect 97 153 131 169
rect 185 545 219 561
rect 185 153 219 169
rect 125 85 141 119
rect 175 85 191 119
rect -51 17 17 79
rect 299 17 333 79
rect -51 -17 79 17
rect 237 -17 333 17
<< viali >>
rect -17 163 17 551
rect 97 169 131 545
rect 185 169 219 545
rect 141 85 175 119
<< metal1 >>
rect -51 551 137 557
rect -51 163 -17 551
rect 17 545 137 551
rect 17 533 97 545
rect 17 169 97 183
rect 131 169 137 545
rect 17 163 137 169
rect -51 157 137 163
rect 179 550 225 557
rect 179 545 340 550
rect 179 169 185 545
rect 219 540 340 545
rect 219 170 230 540
rect 330 170 340 540
rect 219 169 340 170
rect 179 160 340 169
rect 179 157 225 160
rect 45 119 191 125
rect 45 111 141 119
rect 45 59 59 111
rect 111 85 141 111
rect 175 85 191 119
rect 111 69 191 85
rect 111 59 125 69
rect 45 45 125 59
<< via1 >>
rect 7 183 17 533
rect 17 183 97 533
rect 97 183 117 533
rect 230 170 330 540
rect 59 59 111 111
<< metal2 >>
rect -3 533 127 543
rect -3 183 7 533
rect 117 183 127 533
rect -3 173 127 183
rect 220 540 340 550
rect 220 170 230 540
rect 330 170 340 540
rect 220 160 340 170
rect 45 120 125 125
rect 40 111 125 120
rect 40 59 59 111
rect 111 59 125 111
rect 40 50 125 59
rect 45 45 125 50
<< via2 >>
rect 7 183 107 533
rect 230 170 330 540
<< metal3 >>
rect -233 533 117 553
rect -233 413 7 533
rect -3 313 7 413
rect -233 183 7 313
rect 107 183 117 533
rect -233 173 117 183
rect 180 540 3780 560
rect 180 520 230 540
rect 330 520 3780 540
rect 180 200 220 520
rect 460 200 3780 520
rect 180 170 230 200
rect 330 170 3780 200
rect 180 166 3780 170
rect 220 160 340 166
<< via3 >>
rect 220 200 230 520
rect 230 200 330 520
rect 330 200 460 520
<< mimcap >>
rect 600 500 3740 520
rect 600 220 620 500
rect 3720 220 3740 500
rect 600 200 3740 220
<< mimcapcontact >>
rect 620 220 3720 500
<< metal4 >>
rect 180 520 500 560
rect 180 200 220 520
rect 460 200 500 520
rect 180 166 500 200
rect 560 550 3780 560
rect 560 500 3790 550
rect 560 220 620 500
rect 3720 220 3790 500
rect 560 170 3790 220
rect 560 166 3780 170
<< via4 >>
rect 220 200 460 520
<< mimcap2 >>
rect 600 500 3740 520
rect 600 220 620 500
rect 3720 220 3740 500
rect 600 200 3740 220
<< mimcap2contact >>
rect 620 220 3720 500
<< metal5 >>
rect 180 520 3780 560
rect 180 200 220 520
rect 460 500 3780 520
rect 460 220 620 500
rect 3720 220 3780 500
rect 460 200 3780 220
rect 180 166 3780 200
<< labels >>
rlabel metal1 -40 160 -20 550 1 VLO
rlabel metal2 40 50 50 120 1 S
rlabel metal4 3780 170 3790 550 7 C
<< end >>
