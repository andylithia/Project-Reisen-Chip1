magic
tech sky130A
magscale 1 2
timestamp 1671823942
<< locali >>
rect 250 300 400 310
rect 250 220 270 300
rect 380 220 400 300
rect 250 210 400 220
rect 440 300 590 310
rect 440 220 460 300
rect 570 220 590 300
rect 440 210 590 220
rect 635 261 687 277
rect 635 227 644 261
rect 678 227 687 261
rect 635 212 687 227
rect 779 261 831 277
rect 779 227 788 261
rect 822 227 831 261
rect 779 212 831 227
rect 982 261 1034 277
rect 982 227 991 261
rect 1025 227 1034 261
rect 982 212 1034 227
rect 1215 271 1267 287
rect 1215 237 1224 271
rect 1258 237 1267 271
rect 1215 222 1267 237
rect 1391 271 1443 287
rect 1391 237 1400 271
rect 1434 237 1443 271
rect 1391 222 1443 237
rect 1503 271 1555 287
rect 1503 237 1512 271
rect 1546 237 1555 271
rect 1503 222 1555 237
<< viali >>
rect 270 220 380 300
rect 460 220 570 300
rect 644 227 678 261
rect 788 227 822 261
rect 991 227 1025 261
rect 1224 237 1258 271
rect 1400 237 1434 271
rect 1512 237 1546 271
<< metal1 >>
rect 230 650 790 660
rect 230 580 240 650
rect 780 580 790 650
rect 230 570 790 580
rect 250 300 400 310
rect 250 220 260 300
rect 390 220 400 300
rect 250 210 400 220
rect 440 300 590 310
rect 440 220 450 300
rect 580 270 590 300
rect 1215 280 1267 287
rect 635 270 687 277
rect 580 220 635 270
rect 440 210 590 220
rect 635 212 687 218
rect 779 270 831 277
rect 779 212 831 218
rect 982 270 1034 277
rect 1215 222 1267 228
rect 1391 280 1443 287
rect 1391 222 1443 228
rect 1503 280 1555 287
rect 1503 222 1555 228
rect 982 212 1034 218
rect 1010 -10 1570 0
rect 1010 -80 1020 -10
rect 1560 -80 1570 -10
rect 1010 -90 1570 -80
<< via1 >>
rect 240 580 780 650
rect 260 220 270 300
rect 270 220 380 300
rect 380 220 390 300
rect 450 220 460 300
rect 460 220 570 300
rect 570 220 580 300
rect 635 261 687 270
rect 635 227 644 261
rect 644 227 678 261
rect 678 227 687 261
rect 635 218 687 227
rect 779 261 831 270
rect 779 227 788 261
rect 788 227 822 261
rect 822 227 831 261
rect 779 218 831 227
rect 982 261 1034 270
rect 982 227 991 261
rect 991 227 1025 261
rect 1025 227 1034 261
rect 982 218 1034 227
rect 1215 271 1267 280
rect 1215 237 1224 271
rect 1224 237 1258 271
rect 1258 237 1267 271
rect 1215 228 1267 237
rect 1391 271 1443 280
rect 1391 237 1400 271
rect 1400 237 1434 271
rect 1434 237 1443 271
rect 1391 228 1443 237
rect 1503 271 1555 280
rect 1503 237 1512 271
rect 1512 237 1546 271
rect 1546 237 1555 271
rect 1503 228 1555 237
rect 1020 -80 1560 -10
<< metal2 >>
rect 230 650 790 660
rect 230 580 240 650
rect 780 580 790 650
rect 230 570 790 580
rect 650 363 1255 393
rect 250 300 400 310
rect 250 220 260 300
rect 390 220 400 300
rect 250 210 400 220
rect 440 300 590 310
rect 440 220 450 300
rect 580 220 590 300
rect 650 277 680 363
rect 790 305 1135 335
rect 790 277 820 305
rect 440 210 590 220
rect 635 270 687 277
rect 635 212 687 218
rect 779 270 831 277
rect 779 212 831 218
rect 982 270 1034 277
rect 982 212 1034 218
rect 325 182 355 210
rect 790 182 820 212
rect 325 152 820 182
rect 1105 194 1135 305
rect 1225 287 1255 363
rect 1215 280 1267 287
rect 1215 222 1267 228
rect 1391 280 1443 287
rect 1391 222 1443 228
rect 1503 280 1555 287
rect 1503 222 1555 228
rect 1405 194 1435 222
rect 1105 164 1435 194
rect 1010 -10 1570 0
rect 1010 -80 1020 -10
rect 1560 -80 1570 -10
rect 1010 -90 1570 -80
<< via2 >>
rect 240 580 780 650
rect 260 220 370 300
rect 470 220 580 300
rect 1020 -80 1560 -10
<< metal3 >>
rect 230 650 790 660
rect 230 580 240 650
rect 780 580 790 650
rect 230 570 790 580
rect 250 300 380 310
rect 250 220 260 300
rect 370 220 380 300
rect 250 210 380 220
rect 460 300 590 310
rect 460 220 470 300
rect 580 220 590 300
rect 460 210 590 220
rect 1010 -10 1570 0
rect 1010 -80 1020 -10
rect 1560 -80 1570 -10
rect 1010 -90 1570 -80
use sky130_fd_sc_hs__and2_2  sky130_fd_sc_hs__and2_2_0 ~/openmpw/pdk_1/sky130A/libs.ref/sky130_fd_sc_hs/mag
timestamp 1670771148
transform 1 0 614 0 1 -48
box -38 -49 518 715
use sky130_fd_sc_hs__diode_2  sky130_fd_sc_hs__diode_2_0 ~/openmpw/pdk_1/sky130A/libs.ref/sky130_fd_sc_hs/mag
timestamp 1670771148
transform 1 0 230 0 1 -48
box -38 -49 230 715
use sky130_fd_sc_hs__diode_2  sky130_fd_sc_hs__diode_2_1
timestamp 1670771148
transform 1 0 422 0 1 -48
box -38 -49 230 715
use sky130_fd_sc_hs__nand2_2  sky130_fd_sc_hs__nand2_2_0 ~/openmpw/pdk_1/sky130A/libs.ref/sky130_fd_sc_hs/mag
timestamp 1670771148
transform 1 0 1094 0 1 -48
box -38 -49 518 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_0 ~/openmpw/pdk_1/sky130A/libs.ref/sky130_fd_sc_hs/mag
timestamp 1670771148
transform 1 0 1574 0 1 -48
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_1
timestamp 1670771148
transform 1 0 134 0 1 -48
box -38 -49 134 715
<< labels >>
rlabel locali 250 210 400 310 1 S1
rlabel locali 440 210 590 310 1 S2
rlabel metal2 982 212 1034 277 1 YAND
rlabel metal2 1503 222 1555 287 1 YNAND
rlabel metal3 230 570 790 660 1 VHI
rlabel metal3 1010 -90 1570 0 1 VLO
<< end >>
