magic
tech sky130A
timestamp 1671858438
<< pwell >>
rect -176 -282 176 282
<< psubdiff >>
rect -158 247 -110 264
rect 110 247 158 264
rect -158 216 -141 247
rect 141 216 158 247
rect -158 -247 -141 -216
rect 141 -247 158 -216
rect -158 -264 -110 -247
rect 110 -264 158 -247
<< psubdiffcont >>
rect -110 247 110 264
rect -158 -216 -141 216
rect 141 -216 158 216
rect -110 -264 110 -247
<< xpolycontact >>
rect -93 -199 -24 17
rect 24 -199 93 17
<< ppolyres >>
rect -93 130 93 199
rect -93 17 -24 130
rect 24 17 93 130
<< locali >>
rect -158 247 -110 264
rect 110 247 158 264
rect -158 216 -141 247
rect 141 216 158 247
rect -158 -247 -141 -216
rect 141 -247 158 -216
rect -158 -264 -110 -247
rect 110 -264 158 -247
<< properties >>
string FIXED_BBOX -149 -255 149 255
string gencell sky130_fd_pr__res_high_po_0p69
string library sky130
string parameters w 0.69 l 1.3 m 1 nx 2 wmin 0.690 lmin 0.50 rho 319.8 val 2.089k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 1 full_metal 1 wmax 0.690 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
