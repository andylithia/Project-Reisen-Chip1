magic
tech sky130A
magscale 1 2
timestamp 1671152619
<< error_p >>
rect -173 1072 -115 1078
rect 19 1072 77 1078
rect 211 1072 269 1078
rect -173 1038 -161 1072
rect 19 1038 31 1072
rect 211 1038 223 1072
rect -173 1032 -115 1038
rect 19 1032 77 1038
rect 211 1032 269 1038
rect -269 -1038 -211 -1032
rect -77 -1038 -19 -1032
rect 115 -1038 173 -1032
rect -269 -1072 -257 -1038
rect -77 -1072 -65 -1038
rect 115 -1072 127 -1038
rect -269 -1078 -211 -1072
rect -77 -1078 -19 -1072
rect 115 -1078 173 -1072
<< pwell >>
rect -455 -1210 455 1210
<< nmos >>
rect -255 -1000 -225 1000
rect -159 -1000 -129 1000
rect -63 -1000 -33 1000
rect 33 -1000 63 1000
rect 129 -1000 159 1000
rect 225 -1000 255 1000
<< ndiff >>
rect -317 988 -255 1000
rect -317 -988 -305 988
rect -271 -988 -255 988
rect -317 -1000 -255 -988
rect -225 988 -159 1000
rect -225 -988 -209 988
rect -175 -988 -159 988
rect -225 -1000 -159 -988
rect -129 988 -63 1000
rect -129 -988 -113 988
rect -79 -988 -63 988
rect -129 -1000 -63 -988
rect -33 988 33 1000
rect -33 -988 -17 988
rect 17 -988 33 988
rect -33 -1000 33 -988
rect 63 988 129 1000
rect 63 -988 79 988
rect 113 -988 129 988
rect 63 -1000 129 -988
rect 159 988 225 1000
rect 159 -988 175 988
rect 209 -988 225 988
rect 159 -1000 225 -988
rect 255 988 317 1000
rect 255 -988 271 988
rect 305 -988 317 988
rect 255 -1000 317 -988
<< ndiffc >>
rect -305 -988 -271 988
rect -209 -988 -175 988
rect -113 -988 -79 988
rect -17 -988 17 988
rect 79 -988 113 988
rect 175 -988 209 988
rect 271 -988 305 988
<< psubdiff >>
rect -419 1140 -323 1174
rect 323 1140 419 1174
rect -419 1078 -385 1140
rect 385 1078 419 1140
rect -419 -1140 -385 -1078
rect 385 -1140 419 -1078
rect -419 -1174 -323 -1140
rect 323 -1174 419 -1140
<< psubdiffcont >>
rect -323 1140 323 1174
rect -419 -1078 -385 1078
rect 385 -1078 419 1078
rect -323 -1174 323 -1140
<< poly >>
rect -177 1072 -111 1088
rect -177 1038 -161 1072
rect -127 1038 -111 1072
rect -255 1000 -225 1026
rect -177 1022 -111 1038
rect 15 1072 81 1088
rect 15 1038 31 1072
rect 65 1038 81 1072
rect -159 1000 -129 1022
rect -63 1000 -33 1026
rect 15 1022 81 1038
rect 207 1072 273 1088
rect 207 1038 223 1072
rect 257 1038 273 1072
rect 33 1000 63 1022
rect 129 1000 159 1026
rect 207 1022 273 1038
rect 225 1000 255 1022
rect -255 -1022 -225 -1000
rect -273 -1038 -207 -1022
rect -159 -1026 -129 -1000
rect -63 -1022 -33 -1000
rect -273 -1072 -257 -1038
rect -223 -1072 -207 -1038
rect -273 -1088 -207 -1072
rect -81 -1038 -15 -1022
rect 33 -1026 63 -1000
rect 129 -1022 159 -1000
rect -81 -1072 -65 -1038
rect -31 -1072 -15 -1038
rect -81 -1088 -15 -1072
rect 111 -1038 177 -1022
rect 225 -1026 255 -1000
rect 111 -1072 127 -1038
rect 161 -1072 177 -1038
rect 111 -1088 177 -1072
<< polycont >>
rect -161 1038 -127 1072
rect 31 1038 65 1072
rect 223 1038 257 1072
rect -257 -1072 -223 -1038
rect -65 -1072 -31 -1038
rect 127 -1072 161 -1038
<< locali >>
rect -419 1140 -323 1174
rect 323 1140 419 1174
rect -419 1078 -385 1140
rect 385 1078 419 1140
rect -177 1038 -161 1072
rect -127 1038 -111 1072
rect 15 1038 31 1072
rect 65 1038 81 1072
rect 207 1038 223 1072
rect 257 1038 273 1072
rect -305 988 -271 1004
rect -305 -1004 -271 -988
rect -209 988 -175 1004
rect -209 -1004 -175 -988
rect -113 988 -79 1004
rect -113 -1004 -79 -988
rect -17 988 17 1004
rect -17 -1004 17 -988
rect 79 988 113 1004
rect 79 -1004 113 -988
rect 175 988 209 1004
rect 175 -1004 209 -988
rect 271 988 305 1004
rect 271 -1004 305 -988
rect -273 -1072 -257 -1038
rect -223 -1072 -207 -1038
rect -81 -1072 -65 -1038
rect -31 -1072 -15 -1038
rect 111 -1072 127 -1038
rect 161 -1072 177 -1038
rect -419 -1140 -385 -1078
rect 385 -1140 419 -1078
rect -419 -1174 -323 -1140
rect 323 -1174 419 -1140
<< viali >>
rect -161 1038 -127 1072
rect 31 1038 65 1072
rect 223 1038 257 1072
rect -305 -988 -271 988
rect -209 -988 -175 988
rect -113 -988 -79 988
rect -17 -988 17 988
rect 79 -988 113 988
rect 175 -988 209 988
rect 271 -988 305 988
rect -257 -1072 -223 -1038
rect -65 -1072 -31 -1038
rect 127 -1072 161 -1038
<< metal1 >>
rect -173 1072 -115 1078
rect -173 1038 -161 1072
rect -127 1038 -115 1072
rect -173 1032 -115 1038
rect 19 1072 77 1078
rect 19 1038 31 1072
rect 65 1038 77 1072
rect 19 1032 77 1038
rect 211 1072 269 1078
rect 211 1038 223 1072
rect 257 1038 269 1072
rect 211 1032 269 1038
rect -311 988 -265 1000
rect -311 -988 -305 988
rect -271 -988 -265 988
rect -311 -1000 -265 -988
rect -215 988 -169 1000
rect -215 -988 -209 988
rect -175 -988 -169 988
rect -215 -1000 -169 -988
rect -119 988 -73 1000
rect -119 -988 -113 988
rect -79 -988 -73 988
rect -119 -1000 -73 -988
rect -23 988 23 1000
rect -23 -988 -17 988
rect 17 -988 23 988
rect -23 -1000 23 -988
rect 73 988 119 1000
rect 73 -988 79 988
rect 113 -988 119 988
rect 73 -1000 119 -988
rect 169 988 215 1000
rect 169 -988 175 988
rect 209 -988 215 988
rect 169 -1000 215 -988
rect 265 988 311 1000
rect 265 -988 271 988
rect 305 -988 311 988
rect 265 -1000 311 -988
rect -269 -1038 -211 -1032
rect -269 -1072 -257 -1038
rect -223 -1072 -211 -1038
rect -269 -1078 -211 -1072
rect -77 -1038 -19 -1032
rect -77 -1072 -65 -1038
rect -31 -1072 -19 -1038
rect -77 -1078 -19 -1072
rect 115 -1038 173 -1032
rect 115 -1072 127 -1038
rect 161 -1072 173 -1038
rect 115 -1078 173 -1072
<< properties >>
string FIXED_BBOX -402 -1157 402 1157
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 10 l 0.15 m 1 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
